library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_misc.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library UNISIM;
use UNISIM.vcomponents.all;

entity ram_master is
	port(clk             : in  std_logic;
        address_a       : in  std_logic_vector(31 downto 2);
        enable_a        : in  std_logic;
        wbe_a           : in  std_logic_vector(3 downto 0);
        data_write_a    : in  std_logic_vector(31 downto 0);
        data_read_a     : out std_logic_vector(31 downto 0);

        address_b       : in  std_logic_vector(31 downto 2);
        enable_b        : in  std_logic;
        wbe_b           : in  std_logic_vector(3 downto 0);
        data_write_b    : in  std_logic_vector(31 downto 0);
        data_read_b     : out std_logic_vector(31 downto 0));
end; --entity ram     

architecture ram_master of ram_master is
signal enable_a_lo       : std_logic;
signal wbe_a_lo          : std_logic_vector(3 downto 0);
signal data_write_a_lo   : std_logic_vector(31 downto 0);
signal data_read_a_lo    : std_logic_vector(31 downto 0);
signal enable_b_lo       : std_logic;
signal wbe_b_lo          : std_logic_vector(3 downto 0);
signal data_read_b_lo    : std_logic_vector(31 downto 0);
signal enable_a_hi       : std_logic;
signal wbe_a_hi          : std_logic_vector(3 downto 0);
signal data_read_a_hi   : std_logic_vector(31 downto 0);
signal enable_b_hi       : std_logic;
signal wbe_b_hi          : std_logic_vector(3 downto 0);
signal data_read_b_hi    : std_logic_vector(31 downto 0);
signal address_a_reg     : std_logic_vector(31 downto 2);
signal address_b_reg     : std_logic_vector(31 downto 2);
signal enable_a_lo_256       : std_logic;
signal wbe_a_lo_256          : std_logic_vector(3 downto 0);
signal data_write_a_lo_256   : std_logic_vector(31 downto 0);
signal data_read_a_lo_256    : std_logic_vector(31 downto 0);
signal enable_b_lo_256       : std_logic;
signal wbe_b_lo_256          : std_logic_vector(3 downto 0);
signal data_read_b_lo_256    : std_logic_vector(31 downto 0);
signal enable_a_hi_256       : std_logic;
signal wbe_a_hi_256          : std_logic_vector(3 downto 0);
signal data_read_a_hi_256   : std_logic_vector(31 downto 0);
signal enable_b_hi_256       : std_logic;
signal wbe_b_hi_256          : std_logic_vector(3 downto 0);
signal data_read_b_hi_256    : std_logic_vector(31 downto 0);
begin
process(clk)
begin
if rising_edge(clk) then
	address_a_reg <= address_a;
	address_b_reg <= address_b;
	end if;
end process;
data_read_a <= data_read_a_lo when (address_a_reg < x"0001000"&"00") else
data_read_a_hi when ((address_a_reg >= x"0001000"&"00") and (address_a_reg < x"0002000"&"00")) else 
data_read_a_lo_256 when ((address_a_reg >= x"0002000"&"00") and (address_a_reg < x"0003000"&"00")) else 
data_read_a_hi_256 when ((address_a_reg >= x"0003000"&"00") and (address_a_reg < x"0004000"&"00"));
data_read_b <= data_read_b_lo when (address_b_reg < x"0001000"&"00") else
data_read_b_hi when ((address_b_reg >= x"0001000"&"00") and (address_b_reg < x"0002000"&"00")) else
data_read_b_lo_256 when ((address_b_reg >= x"0002000"&"00") and (address_a_reg < x"0003000"&"00")) else 
data_read_b_hi_256 when ((address_b_reg >= x"0003000"&"00") and (address_b_reg< x"0004000"&"00"));
enable_a_lo <= enable_a when (address_a < x"0001000"&"00") else '0';
enable_b_lo <= enable_b when (address_b < x"0001000"&"00") else '0';
enable_a_hi <= enable_a when ((address_a >= x"0001000"&"00") and (address_a < x"0002000"&"00")) else '0';
enable_b_hi <= enable_b when ((address_b >= x"0001000"&"00") and (address_b < x"0002000"&"00")) else '0';
enable_a_lo_256 <= enable_a when ((address_a >= x"0002000"&"00") and (address_a < x"0003000"&"00")) else '0';
enable_b_lo_256 <= enable_b when ((address_b >= x"0002000"&"00") and (address_b < x"0003000"&"00")) else '0';
enable_a_hi_256 <= enable_a when ((address_a >= x"0003000"&"00") and (address_a < x"0004000"&"00")) else '0';
enable_b_hi_256 <= enable_b when ((address_b >= x"0003000"&"00") and (address_b < x"0004000"&"00")) else '0';
wbe_a_lo <= wbe_a when  enable_a_lo='1' else x"0";
wbe_a_hi <= wbe_a when  enable_a_hi='1' else x"0";
wbe_b_lo <= wbe_b when  enable_b_lo='1' else x"0";
wbe_b_hi <= wbe_b when  enable_b_hi='1' else x"0";
wbe_a_lo_256 <= wbe_a when  enable_a_lo_256='1' else x"0";
wbe_a_hi_256 <= wbe_a when  enable_a_hi_256='1' else x"0";
wbe_b_lo_256 <= wbe_b when  enable_b_lo_256='1' else x"0";
wbe_b_hi_256 <= wbe_b when  enable_b_hi_256='1' else x"0";



ram_bit_0_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"ED39BA795990D275FB4A6E96ACC4731DEA4598B0AFB54867F6EE4618C3749807",
INIT_01 => X"58A0047D8607944AC7DA180001ECA2544042106208408208C20022E9173734B3",
INIT_02 => X"9F775E7CB273E6CCA7DAAF00001000000478020113C9C38E09FB7CCCDD9F203E",
INIT_03 => X"441406267B4CB04443163C91110C58F24A31000B8028A810A3D0F8B169A01006",
INIT_04 => X"0005802424830120024121209088809DF81454ACA01E03501D0A3B91E00F0A00",
INIT_05 => X"C1E0039800112014C20B0232838F80D001C0100AEC83C008EF101A034C8CC300",
INIT_06 => X"8B0478B04A83405954592F9B9628000002C3F08754001B51881E007900060F01",
INIT_07 => X"39F36677EE1C387777622717EF711004A6818111086008E080FDC30594001017",
INIT_08 => X"160400195E83A3A0F61BC3929ECB622AABF5FF83860CEB164833F179B48CEE59",
INIT_09 => X"036D8004FDB47600000229410C61010016DC998C84B0128202C0DCB48F05D513",
INIT_0A => X"204122A033000182502440888420247041E876810099D35F900002DB00105C01",
INIT_0B => X"41C000947E16656074EA560F080544900960260144D201890018080D36191110",
INIT_0C => X"781EA781E2781EA781E2781EA781E2781C33C0613C0E00120800239450112ED4",
INIT_0D => X"872917095352BD2A90515A1CA44E7EA84B00001010043803120C3E04E03383E2",
INIT_0E => X"70C7E0B92800224008AE09B8942C48D1FC491204890244812250588601285432",
INIT_0F => X"B80C2038ABACB83C7E03EA5FF83C002783F103EA5FF83C002783F0120847A704",
INIT_10 => X"BD9870380230F2D7C103EACFF83C002783F103EACFF83C002783F310BBF7EFC2",
INIT_11 => X"1F10BBF7EFC61E01804E1E6EA1E3FA01FD97EFC4B80E008C7C2F678FF023FAF5",
INIT_12 => X"B801FCC8E8320C4DAC9220C6B2FF22EF72ADDE6F1A67C80600C2683E0EF8AE1F",
INIT_13 => X"4189B5C00FE651C6104C6D6400FFFB01FC0000FC07EE42FA7C07F22CE3082636",
INIT_14 => X"8BE9FC08FDF4195C0C2038A7C6CAFA7E289F9BA4570380131CAFB2003F9D190A",
INIT_15 => X"270AE9FE635BE11B7F0308D4A80092E0FC1FC662FA7E283FF68A8F0080AE1DDA",
INIT_16 => X"1204812058112C12411402056954AB0C280D000003350013024179498C2EC6B9",
INIT_17 => X"2048120481204812048120481204812048120481204812048120481204812048",
INIT_18 => X"0481204812048120481204812048120481204812048120481204812048120481",
INIT_19 => X"13043A85D4000000000000000001204812048120481204812048120481204812",
INIT_1A => X"82082082082082082218821390771C71C557CE263826D5B1D36AC59E0765D1CF",
INIT_1B => X"1F0F87C3E1F0F87C3E1F0F87C3E0820820820820820820820820820820820820",
INIT_1C => X"FFFFFFFE00000F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E",
INIT_1D => X"EF5D7BD7400000000000000000000000000000000000000000000061F007FFFF",
INIT_1E => X"A10A2D1574005D0428A10A2AAA8BEF552EBDFFF557BC01FF5D7BFFEBA5D55555",
INIT_1F => X"DEBAFFFFC2000AA8428AAAFFAAA8BFF00002AA10FF802ABEFA2D16AA00F7FBE8",
INIT_20 => X"975EFFF8002010002EAAAAAAAD1555FFFFAEA8B550051401450055575FF00517",
INIT_21 => X"4155FF0855575455D2AA8BFFA2D1575EF5D5555545FFFBE8A00087FC20BA5D2A",
INIT_22 => X"8028A00FFAE800AA082A820005D2E974BAA2D140145A2842AA00A284021FF5D0",
INIT_23 => X"2D17FFEF000017400FFD1555FF007FFFEBA55042AA00000017400FFAABFEBAFF",
INIT_24 => X"000000155F7D540000F7FBFFE105D7BE8ABAA284000105D0428BFFA2FBFDFFFA",
INIT_25 => X"75D7BFAEBA5551501D51C5FC7E00000000000000000000000000000000000000",
INIT_26 => X"28B6D16AA28EBF5EDA38AADE1543849557D492BF8E2DE00552EBFFC7552BC01D",
INIT_27 => X"000A85400E00E38A175FDE3F5C002DAAD42DAAAF784AFA82BC042DF47E3D1F80",
INIT_28 => X"AA150021C0092490E904BAFFD550A90FFA495FC7A05B555C257AAA8B45007540",
INIT_29 => X"2DA02402ABD4AD1D0E175D7140B455D516A1EAB45E2A000B4748717A095F571E",
INIT_2A => X"4004A8BC0ABFF7D03A17D1D5147540B454AA080038E9748542AE3D0051C7B6F0",
INIT_2B => X"FB6D4B8FC7BFFFD2168B68F57492F505FF5FA550490BFA482B420B8428A3DA85",
INIT_2C => X"0000000000000000000000016ABD554201543A1EDE9016D4AAB454AF400547AB",
INIT_2D => X"5D2EBDF55556BC35E7557FE8AB25D11415FD0151614000000000000000000000",
INIT_2E => X"9596CBEA41D7D3DECFAF7D43FABAAAD57DEBAAAFFD74AA04547EE18D680BE9A5",
INIT_2F => X"47D78228E5000EA422E10439C1FBCD282351BDAAF9C20AAAABCBEB1DFF803FC5",
INIT_30 => X"1E6284683ABBDD7DEAA100069C14B25495A00F38EBAC0E198B97605018053575",
INIT_31 => X"4408FE6A755ED8EFEFE41B2D17EAF02552BC0545556BD61E501001DF5DD3EBA3",
INIT_32 => X"556F922ACA8AB8283C8310FAB1588916D3861C0422C44082B52A81550A828141",
INIT_33 => X"A5FDBCD7D262E5AFAC4B6AADDD562AF57D7C369AF25495A23068A8301BA7FB95",
INIT_34 => X"003FE0000003FE0000003FE0000003FE0000003FE03D5789700282E9FEFB501E",
INIT_35 => X"0003FE0000003FE0000003FE0000003FE0000003FE0000003FE0000003FE0000",
INIT_36 => X"00000000000000000000000000000000000000000000000000000000003FE000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(0),        -- Port A data input
DOA(0)   => data_read_a_lo(0),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(0),        -- Port B data input
DOB(0)   => data_read_b_lo(0),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_1_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"212C001411984004084D000508C53810A03D1450E839B003342114428A000807",
INIT_01 => X"08000010400A0008010600000084004000400002000000000000000000140000",
INIT_02 => X"484DEBA0111800C004400D000000000028800001CC404E6008B4933336880010",
INIT_03 => X"650C00000848A0423183089008C604224200000100A200002C280810098C0001",
INIT_04 => X"00000004208B00200E010800006667BE7000102C00080000040012010000080C",
INIT_05 => X"0100000000002000600100208D04414000800000000200004800080000800200",
INIT_06 => X"010420104032C204071200000200000010104020000001000910000000040800",
INIT_07 => X"8C0060242183060CF118011281B00000220010400020002081A0008210000802",
INIT_08 => X"000400014812466427040098C000622AAAA43E3060C158AC97F0356BDBFBD008",
INIT_09 => X"026C000559102400200281400469000008B0800000901080004004308B434040",
INIT_0A => X"50502A2800800000400408200000201041000208000040020820034200005C00",
INIT_0B => X"13C051112A800008402002021128000081202205001000000028880004010500",
INIT_0C => X"191AC191A4191A4191AC191AC191A4191A00C8560C8D2940804060901210441E",
INIT_0D => X"C1C114417882F82C00181707044212080300001002081224002006406401918C",
INIT_0E => X"60C0C0B92C000000000400001004200044010200810040802040080200284401",
INIT_0F => X"380C200000043C2016000000F03C00280030000000F03C00280030000004860C",
INIT_10 => X"8D18703800000049C0000000F03C00280030000000F03C002800321080000BC2",
INIT_11 => X"0110800007861E0180000002A9001A00000007C4380E00000001E00230000000",
INIT_12 => X"688004C0C81200009480010280340000008082430A07C80600C0000009008610",
INIT_13 => X"4000134400241186100004A500007B00FC000000000E4A402C001208C3080002",
INIT_14 => X"A9002C0001E0181C0C200000025A400A200812A4070380000000B25000981902",
INIT_15 => X"0000804A0002410A170300C4A800800000020E22400A200096828F008000000A",
INIT_16 => X"020080200820040041002000010080000000000002340002004118010C228614",
INIT_17 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_18 => X"0080200802008020080200802008020080200802008020080200802008020080",
INIT_19 => X"2B5000A000000000000000000000200802008020080200802008020080200802",
INIT_1A => X"AA8A28A28A28A28AB2048634B03249249604CA291AEAFBF1528205C00020C745",
INIT_1B => X"974BA5D6EB75BADD6EB75BADD6EAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA",
INIT_1C => X"FFFFFFFF00000BA5D2E974BA5D2E974BA5D2E974BA5D2E974BA5D2E974BA5D2E",
INIT_1D => X"55AAAAAAA00000000000000000000000000000000000000000000181FFFFFFFF",
INIT_1E => X"BEF5D7BE8ABA5D557DFEFFFD17FEBA00042AAAAFFFFFFE00FF843DF45FFAE955",
INIT_1F => X"DFEF552A800AA5555575FFA2AE820BAFFAEBFF555500155EF552E975FFF7D168",
INIT_20 => X"6AA00A2FBEAABA5D55420AA00002AA00AAFBE8B55A280175455D002AA00A2AAB",
INIT_21 => X"BD75FFAA802AAAAFFAA801EF00517FFFFF7D56ABEF0004155550004154105D55",
INIT_22 => X"55575FF08557DEBAA2FBEAAAA552E955EF5D0415410A2AE97545A2AE954BAF7F",
INIT_23 => X"7D17DF55A2AEBDEAAFFFFC20AAFFFFFFFFFAAD5555FFFFAEAAB55A2D168B555D",
INIT_24 => X"0000000BAFFFBE8A00087FC20BA5D2A975EF5D0002010552E820AAFFD57FF55F",
INIT_25 => X"8FF8A38F45F7AA9217FA380AD400000000000000000000000000000000000000",
INIT_26 => X"D7552E975EFFFDF68BFF557BEAA925551785D7BFD5EFE3F08002FA92EBA5FDE2",
INIT_27 => X"43841017DE92BF8E3AA824924870BF5551555C7A28A821EFE3AABAE38005B575",
INIT_28 => X"0568005A1041055716DB7DB6FBEFEA81C55D0A0516802AA28BEF5EDB7DAA8A15",
INIT_29 => X"C7FEF1C043FE28E3FBD55FFAADE2DAAAE3A5C51C71C042DF45A3D1D00281E8A1",
INIT_2A => X"AA8B45B47F6FB55A95555E90F78E17F52FEF5EDA82FD249057F080417492AAAF",
INIT_2B => X"5FF8AAAA95B7AF45FF8F7DFEDFFAFF8E005FAE92A3AE3DBFF57FA2DF555D257A",
INIT_2C => X"000000000000000000000000A8F571EAA150021C0092490E905FFFD0550BD75C",
INIT_2D => X"00043DE00A2C57DE08FFAAA8B55F7EE801F7F2849EE000000000000000000000",
INIT_2E => X"6AAAE29F067155543A15D2E955EFFFFBEABEF557FEAA10595169BED83D1EBCA8",
INIT_2F => X"BAFFD57DEEAAA15976EB0444BFEB086808A8E3082C954BA5D7DD6145AAAA821A",
INIT_30 => X"B47FFD55D6107782001FF0812000A255D57FFBEF3B97EEAB2C40217B9778428A",
INIT_31 => X"35FF003F17418AEE817B540D11CA80BAAFA825EFAABEBCA18FE803755D08079E",
INIT_32 => X"8BDEBA2D757547D7862AF57ABFFCABE5553FD5FBEFE86353EFFFD03FE0275000",
INIT_33 => X"5A01F70C6AA04537957D6FB4807FFFB45F7EFFDA58FF2AA88A0F3C5014018AC2",
INIT_34 => X"00000000000000000000000000000000000000000B2DD7DEAA100069C14B2549",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(1),        -- Port A data input
DOA(0)   => data_read_a_lo(1),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(1),        -- Port B data input
DOB(0)   => data_read_b_lo(1),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_2_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10E006600180111284380310006289800480032283E000A34301002001A0816",
INIT_01 => X"0005A00810790848048044A54E404340404000720885800802000806EC910200",
INIT_02 => X"5C010802020408040C400850AA055254090541A111200A104A0000000908B510",
INIT_03 => X"0C1101100C00004401060A0010041028021560A0218808002440840008880550",
INIT_04 => X"8840C2802205140048281202180804040960986850688C99444090C10A124A69",
INIT_05 => X"910A21220A880010214000010340086856B141252252142242A068B090106372",
INIT_06 => X"4007A400E8A40086213090040001520500204088012121026050A54CE2154840",
INIT_07 => X"0204022420000004601120108108055200022025A83AA3008882004A001542CA",
INIT_08 => X"091C154429220A2824642010A010020282843E00000248000021100000884101",
INIT_09 => X"80442C1411D120828A2A116A24632885419244606001110AE11B202046439511",
INIT_0A => X"644022201204145003031012D40D718241108815384200904160AE42CE2818E2",
INIT_0B => X"1BF047118108829501009202A5A20068C003211551163A00E522B3000562082D",
INIT_0C => X"90D0490D2C90D0C90D2C90D0C90D2490D04486124868294032384890B8985534",
INIT_0D => X"184014960000008402028041005232001715A040820B11A401E2443243450D04",
INIT_0E => X"9306260000554015520481040100004504A08110000820440001009134000004",
INIT_0F => X"02000000001014000028052000400028040050052000400028040200501C8D38",
INIT_10 => X"4002000000000068005005200040002804002805200040002804000E00001000",
INIT_11 => X"0028400010008000000000102800009800601000040000000011820002140102",
INIT_12 => X"4022010110000000D00008310000801080102000A00004000000000009020000",
INIT_13 => X"00001A00C0082400000006802500008000000000080048000060041200000003",
INIT_14 => X"A000005400080600000000000850000014200411000000000010024440202200",
INIT_15 => X"0000000008840600002080200000000000021800000013000040000000000020",
INIT_16 => X"40902449022A800800002208090684819402120AA8001C800000000000100014",
INIT_17 => X"1902409024090240906419064190641902409024090240906419064190641902",
INIT_18 => X"9044190440900409004090041904419044190440900409004090641906419064",
INIT_19 => X"7D402A2953F81F81F83F03F03F04190441904419044090040900409004190441",
INIT_1A => X"4104104104104104609D21808205965965D65801004E35C300C2D50A22B1C50C",
INIT_1B => X"128944A25128944A25128944A250410410410410410410410410410410410410",
INIT_1C => X"FFFFFFFFE3F00944A25128944A25128944A25128944A25128944A25128944A25",
INIT_1D => X"100055400000000000000000000000000000000000000000000001E1F007FFFF",
INIT_1E => X"400FF843DF45FFAEBDF55082A82155082AAAA10F7FFEAB455500175FF5D2A800",
INIT_1F => X"ABEF082ABDF455D7BD5545F7D5574BAFFD16AAAAA28428ABA000428AAA5D7FD7",
INIT_20 => X"EAB455D7BEAABA5D2A97545552E975FFFFD168AAA5D7BE8BFF5D557FFEFFFD16",
INIT_21 => X"A955555555555FFA2AE820BAFFFFEAABA5555554BA5D0417545F7D56AAAAAAFB",
INIT_22 => X"002AA00AAAEBDFFF08042AABA087BD54BA08043DEAAFF843FF5508517FF55552",
INIT_23 => X"02A82010AAD1401FF002EBFF45A2FBFDFEF00042AA00AAFBEAB5500003FF5500",
INIT_24 => X"0000000BA0004155550004154105D556AA00A2FBEAABA085542145082A800BA0",
INIT_25 => X"D5500155FF552A87410007145400000000000000000000000000000000000000",
INIT_26 => X"9208002FABA4171D5400FF8A38F45F7AABA57D0000855FD1C2AAFA00EBA5E8B7",
INIT_27 => X"A92555178FD7BFD5FDFFA0020BFF78417BD5545F7F1554AAF7D16DABABFF57DE",
INIT_28 => X"756DFFDF6DAAAAAF1EFB6D417BEFA901C2E97F40552E975EFEBDF68ABA557BEA",
INIT_29 => X"2DB7DA3FBD21C7492E9256D555B555C7A2ABC20AAE3AABAE38005B574AA49041",
INIT_2A => X"5EDB7D1E803AF6D400028E02AB8A3A012540E2AABABC75D043A00003FE10E380",
INIT_2B => X"0EB8B7D0AAA800AA147085000FFDA001C7B47BFABC7BFFF7AB4714042AA38BEF",
INIT_2C => X"000000000000000000000000821E8A10568005A1041055716DA38B6FBEFFEF1C",
INIT_2D => X"5D2EBDE00AAC16ABEF5500155EF552A954000855544000000000000000000000",
INIT_2E => X"AF7D57DE0AFAD1EBEB400043DEAA085555400FFAAAAB55F7AEA8BF77004147EF",
INIT_2F => X"EFAAFBEABAF557FEA8515951E8B4D83D1EBDFF082CBDFEF005756145FFD5574A",
INIT_30 => X"E005951550100004155EFF7FFFDE08AA557FFFF083FFCEB95104210405D2E955",
INIT_31 => X"00AA002A3FE18AE803CBE7A3C014351082E951FF5D7FD6145AAAA820A2AAAD29",
INIT_32 => X"EAD45550028ABAFFD17FFED01001FFEF5542ABEB2AA848AAA2552EA8ABA75514",
INIT_33 => X"57FEBAF3F95EEE95C00B7CF12AAA800BA551417105FFFFC21555556EAB4CD6D5",
INIT_34 => X"00000000000000000000000000000000000000000187782001FF0812000A255D",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0400000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(2),        -- Port A data input
DOA(0)   => data_read_a_lo(2),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(2),        -- Port B data input
DOB(0)   => data_read_b_lo(2),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_3_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"210C00A20020000108430020001600B8156021104940741B3530400E02B92202",
INIT_01 => X"A00C9BC058B00968240402C992000B61404040028804A0080A000D16A8990A08",
INIT_02 => X"4809A902031800444445089866E331352180D468B8200E600C0081110B80ACD0",
INIT_03 => X"6D0A601008000142B1A30A040AC68428320006010A80881068A80D401C846330",
INIT_04 => X"482218076809C03B24841CD92CDD5A4402091278072948042640102107102D04",
INIT_05 => X"0B063006A6402109000104E40B04644B32A86D20014A0D204063296082000E34",
INIT_06 => X"01072010703402800606D0102800CAB31434442810B4858060D0500008C52828",
INIT_07 => X"8C00222420A14204E01C581091020CC8000E3226413990008D80001A00CCC4AA",
INIT_08 => X"0874732009120665255420184000220002843E14294258E805E0116002D95101",
INIT_09 => X"BA546AC411102029A61C974014EDBA1320B1046100C0B4034928002002211145",
INIT_0A => X"1052088250A1CC2041051913208CE802438000082040008000F399406BC07998",
INIT_0B => X"19E416590908884D00020242A500090801806801041358222302084204460020",
INIT_0C => X"1019010190101B0101B01019010198101B20805C080C880080506990125E0514",
INIT_0D => X"03400040A101C05C0088242D0000320013339310018011A044414400400101B0",
INIT_0E => X"6514CA601CCCC8B33204C0401104244000018380818040A07060090000280009",
INIT_0F => X"0000000000020000006000000000020000011000000000020000010072CC9251",
INIT_10 => X"0000000000010000014000000000020000013800000000020000010700000000",
INIT_11 => X"002C000000000000000000010000001A00000000000000000040000002440000",
INIT_12 => X"00B2000000000010002049910000011000500000000000000000008000000000",
INIT_13 => X"00020005500000000000800133000000000000000010000000C0000000000040",
INIT_14 => X"0000005300000000000000001000000110600000000000000000401540000000",
INIT_15 => X"8000000008200620000000000000000000400000000107000000000000000004",
INIT_16 => X"0280C0280C0205104100000A8D06C404440230B9980210020040000010010003",
INIT_17 => X"280C0280C0280C0280803808038080380803808038080380C0280C0280C0280C",
INIT_18 => X"80E0200C0280E0200C0280E030080380A030080380A030080380C0280C0280C0",
INIT_19 => X"291008A004D54AAB556AA9556AA830080380A030080380A030080380A0200C02",
INIT_1A => X"4904104104104104A20E85800004924924054C0F031E31C190A285040164C586",
INIT_1B => X"1A8D46A753A9D4EA753A9D4EA752492492492492492492492492492492492492",
INIT_1C => X"FFFFFFFEB6FECD46A351A8D46A351A8D46A351A8D46A351A8D46A351A8D46A35",
INIT_1D => X"00AA8400000000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"B455500175FF5D2AA8A10005540155087BEABFF552ABDF45A2D16AAAAF7D5400",
INIT_1F => X"201000556AB55552ABDE00AAD140010F7D17FF45A2AA82155082AAAA10F7FFEA",
INIT_20 => X"42155557FEAA10007FEAABA000428AAA557FD7400FF843DE00FFAEBFF55082A8",
INIT_21 => X"AA8A105D7BD5545F7D5574BAFF802AA00A2D168ABA085568BEFFFAE820000855",
INIT_22 => X"557FFEFF7D56ABEF557BD74BAFF8402145A2AEBFFEF552EAAABA5D0028BEF082",
INIT_23 => X"5043DEAAAAAA95410F7803FFFF55556AAAA552A975FFFFD16AAAA5D7BC01EF5D",
INIT_24 => X"0000000105D0417545F7D56AAAAAAFBEAB455D7BEAABA5D2A974005D55574005",
INIT_25 => X"5B6DF6FABAFFD547010AA8407400000000000000000000000000000000000000",
INIT_26 => X"6D1C2AAFA28EBF5E8B7D5500155FF552AAF0100071455451C75EABC74174BAF5",
INIT_27 => X"F45F7AABAF7D00009543D1C556AB6D4124BAE10BED542010FFD57AF55AAF5D75",
INIT_28 => X"ABFFEBA0870281C5F4716D5D7FEDA3A0955FF48208002FABA4171D5400FF8A38",
INIT_29 => X"B8EBA15203FFFF002AAFA384171D5545F7D0154AAF7D16DABABFF57DE92005F6",
INIT_2A => X"F68ABA417BC01D7555178FD7BFD5FDF571575D24BA438E021D5B6A4BAFFF5D2E",
INIT_2B => X"24BFE005D5B52428410E3AE92E3A490410EB843ABD71551FFE02552A975FFEBD",
INIT_2C => X"0000000000000000000000003849041756DFFDF6DAAAAAF1EFB6D417BEFBD71C",
INIT_2D => X"5D556AB45081028B55FFFFFFEBAFFD557400A280144000000000000000000000",
INIT_2E => X"0FFD56ABF5AAD15455F5D2EBDEAAA2D16ABEF5500175EF552ABDE00085554545",
INIT_2F => X"AA085555400FFAAAAB14F7AE28BF77004146BA557DEABEF00002BE10FFD54000",
INIT_30 => X"E0AF2D1EAEBA007FEABEFAA84174BA557FD55EF5D3BFEEB35055DEE1000043DE",
INIT_31 => X"0155FFAA28BF7592EABE0A0804ABFFB082EBDEAA005556145FFD5574AAF7D47D",
INIT_32 => X"EB8105D2E955EFAAFBE8AAA547FE21550853E8B4FABD5EBFF75D55420AA82AA8",
INIT_33 => X"57FFFF087FFCEF90104B780A557FC20AA082AAAE10AA8000000A2AC2ABFD2151",
INIT_34 => X"00000000000000000000000000000000000000000AA0004155EFF7FFFDE08AA5",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(3),        -- Port A data input
DOA(0)   => data_read_a_lo(3),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(3),        -- Port B data input
DOB(0)   => data_read_b_lo(3),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_4_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10804002061080A284201081034809800A002303500078B3432C82904204002",
INIT_01 => X"810398000008004C0420050E12100368403008418984014902030806A0910204",
INIT_02 => X"480108A000000000446448E01E80F00A41043118680402000800000009882390",
INIT_03 => X"065040108C0000408406080002101020260012E03000000030808902088000F0",
INIT_04 => X"9100EB8368155C1AE0B01CD60433B944028A90385AC0D438E02010E81C32E801",
INIT_05 => X"B81E4166DE080029204044C401041C4CF01C489433483C8042EAC190100074C4",
INIT_06 => X"400F0400688002A22010D4342045C50F0004028993B3A5260041E4500EB4C0E2",
INIT_07 => X"000000243020008461000812810003C300060064012E00048C82005800BC2888",
INIT_08 => X"08CC8F0109064220240410008000002202043E44001048000020114000881000",
INIT_09 => X"F0DC1EB5131020C7BE7D172251E53E80E891E5016041B4083945202002419104",
INIT_0A => X"7D6025AC2A0982500302003200872003FB108808280200204400786612CE2B08",
INIT_0B => X"11D0025980480A458100930201820964408268101000F022D8083B4044A0002C",
INIT_0C => X"90C3490C1490C3490C1490C1490C3490C104869A48618800B66305989ABA0434",
INIT_0D => X"220000000500021002100088004010001370F030808110204581043243050C54",
INIT_0E => X"06100C40903C1C30F20025440102200541204090600830045825050034010000",
INIT_0F => X"000000000012000000BC04000000020004018C040000000200040000721CD861",
INIT_10 => X"000000000001002001A40400000002000401DC04000000020004014D44001000",
INIT_11 => X"0065040010000000000000110000007600200000000000000050000005D40002",
INIT_12 => X"00DE00001000001040004A3B0000180088500000200000000000008000020000",
INIT_13 => X"0002080760000400000082024300008000000000081006000170000200000041",
INIT_14 => X"180002B200000200000000001806000192000010000000000010401F80000200",
INIT_15 => X"0814000114A00200000000200000000000401006000085C00040000000000024",
INIT_16 => X"40102459044481081044880A0986D4C1560636C7840A61803000820012113042",
INIT_17 => X"1900411064090041102409044110240900401064190040106409004110640904",
INIT_18 => X"9064090240100411044090241902401044110041902409064110241904401024",
INIT_19 => X"04048028064B261934D964C3269C090641100401044090641902401044010041",
INIT_1A => X"AA8A28A28A28A28A74C132343334514513028A2818E01F81400050E130106345",
INIT_1B => X"8341A0D46A351A8D46A351A8D46AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA",
INIT_1C => X"FFFFFFFE58C001A0D068341A0D068341A0D068341A0D068341A0D068341A0D06",
INIT_1D => X"10550015400000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"F45A2D16AAAAF7D568A00AA8400000AAFFC21FFF7D542000FFAE821FF552EAAA",
INIT_1F => X"0000AAAE820BA550015400087FD74BAFFD540000F7D155555087BEABFF552ABD",
INIT_20 => X"A8AAAF78015545FFD555555082AAAA10F7FFEAB455500175FF5D2AAAA1000554",
INIT_21 => X"56AB45552ABDE00AAD140010F7D17FF45A2FBC2000A2FFC21555551554005D2E",
INIT_22 => X"AEBFF55082E82145A280001EFF78402145A2AE801555D2E95555552E97410005",
INIT_23 => X"D517DF45557BD5410F7D555545F7AA97410000428AAA557FD5400FF843DE00FF",
INIT_24 => X"0000000AA085568BEFFFAE82000085542155557FEAA10007FEABEFAAD1400AA5",
INIT_25 => X"8EBAA801EF4920AFA10490A17000000000000000000000000000000000000000",
INIT_26 => X"451C75EABEF4124BAF55B6DF6FABAFFD56F010AA8407428A2F1C01FFF7D14202",
INIT_27 => X"5FF552AAFA10007155428A2AE850925D0010400087FD24AAE3DF47010E38E051",
INIT_28 => X"01555D51524004920ADA82EB8A12555EBFB4717D1C2AAFA28EBF5E8B7D550015",
INIT_29 => X"92555492A850381C5F6AB6D4124BAE10BED542010FFD57AF55AAF5D7410A2FBC",
INIT_2A => X"1D5400FF8A38E00F7AABAF7D0000955FDB684051D7F7840517DA2A4871554124",
INIT_2B => X"55D75EFBED5400825D557FF55007BD7410EBDB5017DE38E8708008002FAAA417",
INIT_2C => X"00000000000000000000000082005F6ABFFEBA0870281C5F4716D5D7FEDB7D09",
INIT_2D => X"AAD1401FFFFD5420BAA2AA821FF08043DE10002A964000000000000000000000",
INIT_2E => X"AA2FBD7410A2AE965555D556ABEF080028B55FFFFFDEBAFFD57FE00A280144BA",
INIT_2F => X"AAA2D16ABEF5500175EF552ABDE000855544AAAA82174105D0402000087FC00B",
INIT_30 => X"BF5AAD154400AAFBC015555554001008003FE00AAEA81154AAFFD65FF5D2EBDE",
INIT_31 => X"75EFA2AA155550004021E5582A964BE557FEABEF00002BE10FFD540000FFD56A",
INIT_32 => X"9661000043DEAA085555400FFAAAAA10F7AC28BF558001454DF78017555F7801",
INIT_33 => X"FD55EF5D7BFEEF35055487EFF7D1400105D517FF55087FD7410A2FBC01E7F2AE",
INIT_34 => X"0000000000000000000000000000000000000000010007FEABEFAA84174BA557",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0400000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(4),        -- Port A data input
DOA(0)   => data_read_a_lo(4),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(4),        -- Port B data input
DOB(0)   => data_read_b_lo(4),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_5_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50DF0A0791B3FC1694378283C81FD996A091A32152007AB36B20E03C040C006",
INIT_01 => X"081FBDC49830884C5C6A60000C34C24841280A00084000C8C212892EEA953231",
INIT_02 => X"C809AD5CB118E640A4F008F8011FF0002080000082CCC66609DB7DDDCB1F2036",
INIT_03 => X"25080626BE4C904210831C80084204720B20048A88800000B8E0F8102885500E",
INIT_04 => X"4005122024899100064520C01444429C7804103C0416C007198A3916E0551A04",
INIT_05 => X"46E1829941C9000944C8C022898FE2F20D7D7A104CB5C208E51417C054848912",
INIT_06 => X"CA075CA0E63342991612DF9A8205C0A0B030B20B10480900886E220801073711",
INIT_07 => X"8C732074B68D1A34E3180717FFD13FC72691924098712CE481FDC241D43C1ACD",
INIT_08 => X"16053F180A1286A4E51BD18840C320000075FE91A24458BA4DE0D57992D9BE58",
INIT_09 => X"0A4D8105BF3472304100930258E510601EDE1D8524309285FD416CB402259504",
INIT_0A => X"3110AC0D11C901B2112109204C28B67061E8928920CAD3CFC0140079065A4A65",
INIT_0B => X"C3404959321C284D356A964F8125CD7AC8632614005DFBAACFBC800024091128",
INIT_0C => X"380D6380B6380F638096380F6380B6380D51C04B1C07AD10C14020D233127AD5",
INIT_0D => X"992940513052F4CA8A0A0664A5023CA8470FF000908C383755AF1604E0538096",
INIT_0E => X"200040194FFC044FFA4B08BC85282C91F028D094284A34054A25508605135C01",
INIT_0F => X"BA0C2038ABACBC7C7806F94FF87C002F83F106F94FF87C002F83F2000A04C200",
INIT_10 => X"8D9A70380230F2DFC106F86FF87C002F83F106F86FF87C002F83F3601BFFEBC2",
INIT_11 => X"1F401BFFE7C69E01804E1E6EABE3F040FFD7C7C4BC0E008C7C2FE58FC0A9FFF5",
INIT_12 => X"F8BFDFC8C8120C4DBC802208B2EB2AE777ADFE6F0A47CC0600C2683E0FF8AE3F",
INIT_13 => X"4189B7C56DF47186104C6DE7037FFF00FC0000FC07EE4E7A7076FE28C3082636",
INIT_14 => X"B9E9F272FFFC181C0C2038A7C6DE7A7D909FBFA4070380131CAFB257FBD93902",
INIT_15 => X"2B34E9F56DFBEB1B7F2300C4A80092E0FC1FCE667A7C877FFE828F0080AE1DDA",
INIT_16 => X"51142511405EA00A1344612A898494801602081F87204A9452217159891640D4",
INIT_17 => X"0942511425014450940519425114650140519405194650146511405194050946",
INIT_18 => X"1465114250146501465194051944509445094051146501465014251140509445",
INIT_19 => X"7ED430A983124B2DA6924965B4D5014650142511425094450940519405094450",
INIT_1A => X"EFBEFBEFBEFBEFBE5FDFF3F7F773CF3CF7D796ED39FDEE76DFFCE9F84801B6DB",
INIT_1B => X"BDDEEF77BBDDEEF77BBDDEEF77BBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFB",
INIT_1C => X"FFFFFFFE433B5EEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77B",
INIT_1D => X"AAFFFBFFE00000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"000FFAE821FF552E820105500155555D2AA8A00AA843FFFFF78002155AAAE974",
INIT_1F => X"0000FFAE80000AAAE974BAFFAEAAB45AAAEBDEAAA2FFEAA00AAFFC21FFF7D542",
INIT_20 => X"7FE000055574BA557FFFF55087BEABFF552ABDF45A2D16AAAAF7D56AA00AA840",
INIT_21 => X"E820BA550015400087FD74BAFFD540000F780155555D7BE8B45085168BFFA2D1",
INIT_22 => X"2AAAA10005140145FFFBC01EFAAFFD75FF002E97555A2AABDEAAAAAAAAA00AAA",
INIT_23 => X"A84174BA5D043FF45AAAA974AAF7AEBFF55082AAAA10F7FFEAB455500175FF5D",
INIT_24 => X"000000000A2FFC21555551554005D2EA8AAAF78015545FFD555410552EA8BEFA",
INIT_25 => X"FFF8E0217DBEA4954AAE3FBFDE00000000000000000000000000000000000000",
INIT_26 => X"28A2F1C01D7F7D142028EBAA801EF492087A10490A171455D2EADA28B6803FFF",
INIT_27 => X"ABAFFD56FA10AA8417428E3AE87010A2A4974AAE3AEAFB6DAAA4BDEAAA2F1EDA",
INIT_28 => X"8B6D14516DBD7BEDB7DE381451554AA497FFFF451C75EABEF4124BAF55B6DF6F",
INIT_29 => X"BDEAAAAA0AFA28A2A4850925D0010400087FD24AAE3DF47010E38E0516D5D7BE",
INIT_2A => X"5E8B7D5500155FF552AAFA10007155545F7F1C21D7AAF1D55FF082A9057DA2AA",
INIT_2B => X"FB470384124ADBFFBE84174AA55043FF6DBEAE950AAEB8ABDF7D1C2AAFA28EBF",
INIT_2C => X"00000000000000000000000010A2FBC01555D51524004920ADA82EB8A12410EB",
INIT_2D => X"552EBFEBAF7843DFEFF7AE801EFF780174AAAAFBFEE000000000000000000000",
INIT_2E => X"FA2803FEBAAAD17CEAAAAD140155FFD5420BAA2AA821FF080415410002A96555",
INIT_2F => X"EF080028B55FFFFFDEBAFFD57FE00A280144AAA2AA97400A280174AAA2AEBDFE",
INIT_30 => X"410A2AE965FF557FE8BFF55557FF55FFFBFFEAA5D51554AA087BFEF555D556AB",
INIT_31 => X"55FF0004821FFAAAEBDEAAAA843CEAAAA80174105D0402000087FC00BAA2FBD7",
INIT_32 => X"BEFFF5D2EBDEAAA2D16ABEF5500175EF552ABDE00005554545F7D140145A2D55",
INIT_33 => X"03FE00AAAA81114AAFFD64BA00043FFFFFF80174AA55043DFFFFFAE974BAA2AE",
INIT_34 => X"0000000000000000000000000000000000000000000AAFBC0155555540010080",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"1800000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(5),        -- Port A data input
DOA(0)   => data_read_a_lo(5),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(5),        -- Port B data input
DOB(0)   => data_read_b_lo(5),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_6_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10844B0061A258A2840112C03002C18000402322520070B303301C0381A0086",
INIT_01 => X"0600404820094048008100000042026041000000090800090210080008510204",
INIT_02 => X"080108220C1000004440080000C008010000000001203240080080000988A050",
INIT_03 => X"040000000823404000020A600000002983800584488000103080040C08C00000",
INIT_04 => X"00101610A029B08400044800000000040000102A040810040400100500101800",
INIT_05 => X"05000000800C8300306420002900404400820000000A00804004084001200A00",
INIT_06 => X"64472644640C00808C10D00401823F0020204209101001002650020001052800",
INIT_07 => X"080000242000000461100050818080380900224000200008818028804883E10A",
INIT_08 => X"01FE80E0090242602C0020608000000000043E00000048800021140000881106",
INIT_09 => X"12447E041B102020208000424029006FE0B085013204D0200101006862119140",
INIT_0A => X"4D540B0D916BBE39059191200000200441040108000020006FC5FA6000816908",
INIT_0B => X"8BF05D11A20808454010834225A28962E40AA05510180022FFA6A8800402A06D",
INIT_0C => X"16C1416C5416C5416C3416C3416C7416C500B60A0B60AD04EB4104C093904535",
INIT_0D => X"59802817888180E80112A1660050900003400430CB4911B445A105B05B016C14",
INIT_0E => X"000000062003C90000442006439324280034E85A742D1A16CD2DA30046848048",
INIT_0F => X"00000000000157000600000000000028000C00000000000028000CE800048000",
INIT_10 => X"00000000000000483C00000000000028000C00000000000028000D1080000000",
INIT_11 => X"00108000000000000000000078000A00000000000000000000019A0030000000",
INIT_12 => X"4604000000000000934909080014000000000000000000000000000009005180",
INIT_13 => X"00001230B00000000000049B3C000000000000000001FA000C98000000000002",
INIT_14 => X"E8000E05000000000000000001720002A56000000000000000000FC080000000",
INIT_15 => X"0840000B000404A000000000000000000002099A0003B0000000000000000001",
INIT_16 => X"69DA5685A146D19D084488080904C0A1172240C0781400C81908000205208614",
INIT_17 => X"85A1695A769DA3685A169DA768DA1685A169DA7685A1685A769DA7685A168DA7",
INIT_18 => X"5A368DA1685A769DA168DA3695A569DA3685A169DA5695A368DA1695A569DA36",
INIT_19 => X"7F10800846638C31C71C718638E685A769DA5685A3685A569DA7685A168DA769",
INIT_1A => X"E38E38E38E38E38E76DDB3B7B377DF7DF7D7DE2F39FE3FC3D3EA55FF37F5F7CF",
INIT_1B => X"9FCFE7F3F9FCFE7F3F9FCFE7F3F8E38E38E38E38E38E38E38E38E38E38E38E38",
INIT_1C => X"FFFFFFFF61AC8FE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F",
INIT_1D => X"EFAAAABFE00000000000000000000000000000000000000000000181F007FFFF",
INIT_1E => X"FFFF78002155AAAE974AAFFFBFFE10F7FBE8BEF552E95555552EAABEF082E975",
INIT_1F => X"5410A2AAAAA10087FC01EF552EAAB45F7AE821550851555555D2AA8A00AA843F",
INIT_20 => X"2ABEFA2AEBDFFF552AAAA00AAFFC21FFF7D542000FFAE821FF552E8001055001",
INIT_21 => X"E80000AAAE974BAFFAEAAB45AAAEBDEAAA2FFEAB45552E800AA555568A105D00",
INIT_22 => X"D56AA00AA8400000007BC21FFAA803FFEF5551420105D5568B45FF8400000FFA",
INIT_23 => X"7FBC2155007FC20BAA2D5575FF087FFFF55087BEABFF552ABDF45A2D16AAAAF7",
INIT_24 => X"0000001555D7BE8B45085168BFFA2D17FE000055574BA557FFFE10F7AAA8A00F",
INIT_25 => X"D4924ADBD70820975FFA2A4BFE00000000000000000000000000000000000000",
INIT_26 => X"455D2EADA28B6803FFFFFF8E0217DBEA4954AAE3FBFDE38F7FFEABFF412A9056",
INIT_27 => X"1EF492087010490A07038B6A0AFA38007BC51EF4920AFB55EBA4851450855555",
INIT_28 => X"5082555F68A3855002FBC7BEA4BFFFF492EADA28A2F1C01D7F7D142028EBAA80",
INIT_29 => X"6DB45E38A07028E3AE87010A2A4974AAE3AEAFB6DAAA4BDEAAA2F1EDB55492A8",
INIT_2A => X"4BAF55B6DF6FABAFFD56FA10AA84174381C7FC01C7B68E3DFC75555400105D51",
INIT_2B => X"7FFFE38F7A0AFA38E3FFC21450071C2092A2D5571FF0851FDF451C75EABEF412",
INIT_2C => X"0000000000000000000000016D5D7BE8B6D14516DBD7BEDB7DE381451554AA49",
INIT_2D => X"F7FBEABEF002E801EF00003FF550800155FFA2803CE000000000000000000000",
INIT_2E => X"5A28417555085154555552EBFEBAF7843DFEFF7AE801EFF780174AAAAFBFEEAA",
INIT_2F => X"55FFD5420BAA2AA821FF080415410002A964AAFF803DEAA087FD55FF00043DF4",
INIT_30 => X"EBAAAD17CF55002E95410557BEAABA55043DF55F7803FFEF002ABEEAAAAD1401",
INIT_31 => X"DF455D51420105D517DF55AAAA964AAA2AA97400A280174AAA2AEBDFEFA2803F",
INIT_32 => X"7CF555D556ABEF080028B55FFFFFDEBAFFD57FE00A280144BA5D7FC2155FFAAB",
INIT_33 => X"BFFEAA5D51554AA087BFEEAAF7803DEAAAAFBC0155085540000A2D5575FF0851",
INIT_34 => X"00000000000000000000000000000000000000001FF557FE8BFF55557FF55FFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"1200000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(6),        -- Port A data input
DOA(0)   => data_read_a_lo(6),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(6),        -- Port B data input
DOB(0)   => data_read_b_lo(6),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_7_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10844B00482258A2842112C02450418800002300500030B303300C018180002",
INIT_01 => X"0200084020084048040080000201026040000000080000080200090000510204",
INIT_02 => X"4801082048100000444008040080000041000000000222400800000009000010",
INIT_03 => X"0401018108A144D0000208424000002103006480088000003080000408C10000",
INIT_04 => X"0000120022419000000C80000000000400201829040000050001940400301820",
INIT_05 => X"04000000800840092CC080214144004400000000000800065004004020220800",
INIT_06 => X"40870408600000808C10D4500080008020200008001001000240000061052002",
INIT_07 => X"08000024200000046010005281848001494020400031240C8C8238A06A000988",
INIT_08 => X"40050001090242602C0408408000000000243E00000048800020154000881024",
INIT_09 => X"024401041B132820000011424069004000B20403200891420101026A42210440",
INIT_0A => X"013800A0281400300C0010200008B20663970148004424006818026200004800",
INIT_0B => X"01C1103022881845421082C2C0082300401121810012004600001010040028A0",
INIT_0C => X"1200112001120011204112041120411206089010890100408040008012101414",
INIT_0D => X"09146817802988694902A02451109006230006E0808294008C02848148092001",
INIT_0E => X"000000042C00040002000004020020490020401020081004482501010C120948",
INIT_0F => X"0130C807144102420700052000003C00780B00052000003C007808450484C000",
INIT_10 => X"400002C0E00E0D003300052000003C00780B00052000003C0078099080001000",
INIT_11 => X"80908000100000661801E18042100E000060100000B038038380124038000102",
INIT_12 => X"053A010111848322020512000414400000002000A1001058300C0741C0054120",
INIT_13 => X"90644029D008240864231011BF00008000C3C003F00186040EE8041204321188",
INIT_14 => X"18100D770008060130C807182106040375600411004C2600E3400C2740202230",
INIT_15 => X"9094100A8CA406A0002C812240B0201F0380211604037740004010472041E201",
INIT_16 => X"40100401006E8118104428088904C4C414420080049450801000088444300601",
INIT_17 => X"0906409004010040104409024090240906401004010040102409024090240100",
INIT_18 => X"1024090241900401004090240902401004010040902409004010440100409024",
INIT_19 => X"004420A945841040002082080004110240902409004110040902409024110040",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFEDD9EC000000000000000000000000000000000000000000000000000",
INIT_1D => X"BA082AAAA00000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"555552EAABEF082E975EFAAAABFFEF002ABDF555D5157555F7FBC00AAAAD5400",
INIT_1F => X"FEAAAAAABDF55FFFBFDF55555568ABAAAD5401FF5D2AAAA10F7FBE8BEF552E95",
INIT_20 => X"400005D55554105D51401555D2AA8A00AA843FFFFF78002155AAAE974AAFFFBF",
INIT_21 => X"AAAA10087FC01EF552EAAB45F7AE821550851554AAF7FBFFEAA007BFFFEFF7D5",
INIT_22 => X"2E800105500155EF5D2EBFF450000020AA5D7BC0000F7D555545A28000010A2A",
INIT_23 => X"FAAA8A10FFD568ABAA2D56AAAAF7AABFE00AAFFC21FFF7D542000FFAE821FF55",
INIT_24 => X"000000145552E800AA555568A105D002ABEFA2AEBDFFF552AAAABAA2AE95555F",
INIT_25 => X"5E3F5C20BAAAD5420821C2EAAA00000000000000000000000000000000000000",
INIT_26 => X"38F7FFEABFF412A9056D4924ADBD70820975FFA2A4BFFFF1C2EB8F4555555054",
INIT_27 => X"17DBEA4954AAE3FBFDE82B6AEBAF55E3FFFAF55555F6FA92BED5421C75D20AAA",
INIT_28 => X"FE920075FDFD7F7D5400385D51504385D55401455D2EADA28B6803FFFFFF8E02",
INIT_29 => X"5057DB68E02038B6A0AFA38007BC51EF4920AFB55EBA485145085555492F7F5F",
INIT_2A => X"142028EBAA801EF492087010490A071EF4920B8F45140E07082417BC2000EBD5",
INIT_2B => X"2EADA92A2A09257DE3A4AAA10F7D16FAAABED56AE82F780BAE28A2F1C01D7F7D",
INIT_2C => X"00000000000000000000000155492A85082555F68A3855002FBC7BEA4BFFFF49",
INIT_2D => X"552EAAB455D5142155AAD1400AAA2D1420005D2EA9A000000000000000000000",
INIT_2E => X"0F7D1421555D042BAAAF7FBEABEF002E801EF00003FF550800155FFA2803CFFF",
INIT_2F => X"BAF7843DFEFF7AE801EFF780174AAAAFBFEE00F7AAAAB55AAFBEAB555D7BFDE0",
INIT_30 => X"555085154400FFD17FE1000517FF55FFD5420BA5D55400BA555543155552EBFE",
INIT_31 => X"5400087BC0000A2D5421EFF7AE810AAFF803DEAA087FD55FF00043DF45A28417",
INIT_32 => X"2BAAAAAD140155FFD5420BAA2AA821FF080415410002A965FF080428B45552A9",
INIT_33 => X"43DF55F7803FFEF002ABEE00A280001FFA28028A00FFD17DEAAF7D56AA10FF84",
INIT_34 => X"0000000000000000000000000000000000000000155002E95410557BEAABA550",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"01FFFFFFFFE00000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(7),        -- Port A data input
DOA(0)   => data_read_a_lo(7),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(7),        -- Port B data input
DOB(0)   => data_read_b_lo(7),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_8_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00000648E2840112C00000418000002700500030B3032000000000082",
INIT_01 => X"000009C21838284D1C2160000E12424840000000180800080200000040110204",
INIT_02 => X"080108000090000004400C040080000051000000000002400800000009000010",
INIT_03 => X"00000100043008D0000200024000000003800504488000103080880008800000",
INIT_04 => X"00009410A028A084000440000000000400001022040800150400808500321800",
INIT_05 => X"8500010080048A09302420202804400400800010200A00020204084011014A00",
INIT_06 => X"2447A244608800840490D0040007FE0021204288001000000050024001042800",
INIT_07 => X"4800002420000004201000D281040003182020400031241C0D80004041BFE88A",
INIT_08 => X"4005000108020220240000048000000000043E00000048800000010000881000",
INIT_09 => X"0204010519110020008111020069004008A28501120450220101214122509140",
INIT_0A => X"0528A52291490029019190200008B20E23008028000208804010024000004000",
INIT_0B => X"13C151312A8808454104824001280108A409A044001200020020989000000061",
INIT_0C => X"0000000000000000000000000000000000400020000229508040008012105400",
INIT_0D => X"48022817880508602102A1200810B2020340043248CA00240420000000400040",
INIT_0E => X"4100820020000C0000442142419120000014684A34251A12CD2CA30042840248",
INIT_0F => X"45F3D80000000001020404000783FC0000010404000783FC000000880284C010",
INIT_10 => X"02658FC7E0000000010404000783FC0000010404000783FC000001500000103D",
INIT_11 => X"40500000103961FE78000000000402400020003B43F1F8000000022010800002",
INIT_12 => X"0080001617CD800000080B000804080000020090659833F9F03C000000000000",
INIT_13 => X"B000000400018639EC000000000000FE03FFC00000000600840000C31CF60000",
INIT_14 => X"180204000001E2A3F3D80000000600802000401AA8FC7E00000000100002C2F5",
INIT_15 => X"005404020000104480DC372B47F060000000000600802000017570FF60000000",
INIT_16 => X"28CA328CA34650850A4C000009A494A015624080044440481908000220308640",
INIT_17 => X"8CA328CA328CA328CA3284A1284A1284A1284A1284A1284A328CA328CA328CA3",
INIT_18 => X"CA1284A1284A1284A128CA328CA328CA328CA3284A1284A1284A1284A128CA32",
INIT_19 => X"64108088440000000000000000028CA1284A1284A1284A128CA328CA328CA328",
INIT_1A => X"E79E79E79E79E79EDFC8F33637D6CB6CB2900A282950FAF15E8428917C51E75D",
INIT_1B => X"87D3E1F0F87C3E1F0F87C3E1F0F9E79E79E79E79E79E79E79E79E79E79E79E79",
INIT_1C => X"FFFFFFFECB0593E1F4F87D3E1F4F87D3E1F4F87D3E1F4F87D3E1F4F87D3E1F4F",
INIT_1D => X"10002ABFE00000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"555F7FBC00AAAAD5400BA082AAAA10000000010F7D5421EF007BC01FF5D7FFFE",
INIT_1F => X"FEAA5551554AAFF80021EF002A820BAFF8428A00A2AAAABEF002ABDF555D5157",
INIT_20 => X"E8BEFFFFFEAB55002ABFE10F7FBE8BEF552E95555552EAABEF082E975EFAAAAB",
INIT_21 => X"ABDF55FFFBFDF55555568ABAAAD5401FF5D2AAAB55FFD1400AA5D7FC01EFA2FF",
INIT_22 => X"AE974AAFFFBFFEAA08001555555516ABEFA280020AA5D043DF55557BEAAAAAAA",
INIT_23 => X"8042AB55005140145AAFFE8AAAF7D1401555D2AA8A00AA843FFFFF78002155AA",
INIT_24 => X"0000000AAF7FBFFEAA007BFFFEFF7D5400005D55554105D51400005551421EF0",
INIT_25 => X"71C7FC21EF5D75FFE10142EBAE00000000000000000000000000000000000000",
INIT_26 => X"FF1C2EB8F45555550545E3F5C20BAAAD5420821C2EAAA101C0005000E3D1401D",
INIT_27 => X"BD70820975FFA2A4BFE925D51554AAE384001FF142E800AAFF802AA28AAAEAFB",
INIT_28 => X"7092557BC21D7BEF5EDBC7FFF1EFB6D1420BAE38F7FFEABFF412A9056D4924AD",
INIT_29 => X"3AF55417BEDA82B6AEBAF55E3FFFAF55555F6FA92BED5421C75D20AAB45F7D14",
INIT_2A => X"03FFFFFF8E0217DBEA4954AAE3FBFDEAA1C001056D415F6ABEFA284020824904",
INIT_2B => X"55400385D51401EF00002FB45085F4016DAAF1EDAAAFFFB401455D2EADA28B68",
INIT_2C => X"00000000000000000000000092F7F5FFE920075FDFD7F7D5400385D51504385D",
INIT_2D => X"5D0417410AAD540155557FC01EF5D557DE105D2AA8A000000000000000000000",
INIT_2E => X"AF7842AABAA2AEBDFFF552EAAB455D5142155AAD1400AAA2D1420005D2EA9A10",
INIT_2F => X"EF002E801EF00003FF550800155FFA2803CE105D55574BAA280021EF5D2E820B",
INIT_30 => X"1555D042BB45FFD157410557FC0155F7D57FF55F7D57FFEF550028AAAF7FBEAB",
INIT_31 => X"8BFFAA8000000080428B55087FFFE00F7AAAAB55AAFBEAB555D7BFDE00F7D142",
INIT_32 => X"C2155552EBFEBAF7843DFEFF7AE801EFF780174AAAAFBFEEBA5D04021EF087BE",
INIT_33 => X"5420BA5D55400BA5555430BA5555421EF00043FF45007BC21FFA2D57FEBAF7FB",
INIT_34 => X"0000000000000000000000000000000000000000000FFD17FE1000517FF55FFD",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0800000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(8),        -- Port A data input
DOA(0)   => data_read_a_lo(8),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(8),        -- Port B data input
DOB(0)   => data_read_b_lo(8),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_9_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00018248A2840112C00002C18000002300500030B3032000000000006",
INIT_01 => X"000008000000004C0020000000100268413C0A61590001D90213C00000110204",
INIT_02 => X"680108200010000054400C040080000041000000010002400800800009082011",
INIT_03 => X"00040100000020D0000200124000000043800504488000103081880008800000",
INIT_04 => X"00001410A00AA084000400000200000400001020040010050020820400101880",
INIT_05 => X"0400040080048A09202420000C00410400000000000800020804004000000800",
INIT_06 => X"24478244640800840410D4144002008020200009301000000140000201042000",
INIT_07 => X"0800002C20000004301000128104000100002040003164040D80000040000888",
INIT_08 => X"40050003080202202400000080000000000C3E00000048800010230000881000",
INIT_09 => X"0024010411110420008010020021004000A204011200500001010000AA10C000",
INIT_0A => X"7945282804010009009090200008B20223800008020000004010024204000440",
INIT_0B => X"114100112208084540008240110001002400A000001000020008288000000420",
INIT_0C => X"010400100001040010000104001000010400080000820800000000801010100A",
INIT_0D => X"08403C16800100640182A0210010921003400412484202200400004004001040",
INIT_0E => X"410082002C000C000240004240932041401468CA34651A32CD28A22002840048",
INIT_0F => X"000000000000144002000420000000280001000420000000280000000284C010",
INIT_10 => X"4000000000000048010005000000002800010005000000002800001000001000",
INIT_11 => X"0010000010000000000000002A00020000201000000000000001820010000002",
INIT_12 => X"40BA00011000000090000B000004000000000000A00000000000000009000020",
INIT_13 => X"00001205D0080400000004803F0000800000000000004C0004E8001200000002",
INIT_14 => X"B000047700000600000000000054000135600011000000000000025740200200",
INIT_15 => X"001400020CA406A0000080200000000000020804000137400040000000000000",
INIT_16 => X"28CA328CA36651951A4CA8000984D4E557220080040440481908000001300614",
INIT_17 => X"84A1284A1284A1284A1284A1284A1284A1284A1284A1284A328CA328CA328CA3",
INIT_18 => X"4A1284A1284A1284A128CA328CA328CA328CA328CA328CA328CA328CA3284A12",
INIT_19 => X"2540A809010000000000000000028CA328CA328CA328CA3284A1284A1284A128",
INIT_1A => X"4534D34D34D34D344A2D840100E4920824055CD13333D2379A2A24018615C38E",
INIT_1B => X"268341A0D068341A0D068341A0D1451451451451451451451451451451451451",
INIT_1C => X"FFFFFFFE6DA90341A4D268341A0D069349A0D069349A0D068341A4D268341A4D",
INIT_1D => X"FFFFD557400000000000000000000000000000000000000000000001FFFFFFFF",
INIT_1E => X"1EF007BC01FF5D7FFFE10002ABFF55F7D168A00552E95555007BFFF55087BE8B",
INIT_1F => X"AA10F7FBC0145F7AE801EFF7FBFFF455D7BC0155F7D557410000000010F7D542",
INIT_20 => X"BDE00AA803FFEF5D55421EF002ABDF555D5157555F7FBC00AAAAD5400BA082AA",
INIT_21 => X"1554AAFF80021EF002A820BAFF8428A00A2AAAAAAAF7D17DE00FFFBD5555A2AA",
INIT_22 => X"2E975EFAAAABFFEF002A954BA5551421EF552E954105D00021455555420AA555",
INIT_23 => X"7D5575EFA2FFD75455D7BE8A005D5557410F7FBE8BEF552E95555552EAABEF08",
INIT_24 => X"000000155FFD1400AA5D7FC01EFA2FFE8BEFFFFFEAB55002ABFE10080028BFFF",
INIT_25 => X"D1C71F8F7D147BEFBEFEBD152400000000000000000000000000000000000000",
INIT_26 => X"101C0005000E3D1401D71C7FC21EF5D75FFE10142EBAF7DE3D16DA0041209056",
INIT_27 => X"0BAAAD5420821C2EAAA10E3FFC0145F7A0801FFEBFBF8F6D417BC716DEBD1524",
INIT_28 => X"DE28F7F5D0545B6AAB8E38B68A3AFFF5551471FF1C2EB8F45555550545E3F5C2",
INIT_29 => X"021455D5B470925D51554AAE384001FF142E800AAFF802AA28AAAEAFABAE3D17",
INIT_2A => X"A9056D4924ADBD70820975FFA2A4BFFFF082E974BA4155401C7552097428550E",
INIT_2B => X"20BAE0008002ABFFF7DB505FFAAFBD7555417FEFA00495B52438F7FFEABFF412",
INIT_2C => X"00000000000000000000000145F7D147092557BC21D7BEF5EDBC7FFF1EFB6D14",
INIT_2D => X"AAD17DE100804001EF55516ABFF557BFDFEFA2D5400000000000000000000000",
INIT_2E => X"F007FD55FFA2D5400105D0417410AAD540155557FC01EF5D557DE105D2AA8BEF",
INIT_2F => X"455D5142155AAD1400AAA2D1420005D2EA9A00A2FBC0145FF84001EFA2FFEABF",
INIT_30 => X"ABAA2AEBDEAAAAD17DEBAFFD142155FFAAAAABAFFAAAABFF5551555FF552EAAB",
INIT_31 => X"01555D00154AA552E801455D7BD54105D55574BAA280021EF5D2E820BAF7842A",
INIT_32 => X"C00AAF7FBEABEF002E801EF00003FF550800155FFA2803CFFF002E954BA00514",
INIT_33 => X"57FF55F7D57FFEF550028A10000428BEFF7FFC01FFA2FFD5545007BFDE10087F",
INIT_34 => X"0000000000000000000000000000000000000000145FFD157410557FC0155F7D",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"1000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(9),        -- Port A data input
DOA(0)   => data_read_a_lo(9),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(9),        -- Port B data input
DOB(0)   => data_read_b_lo(9),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_10_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000B0001800002840002C0000281800020030000000033122000400992006",
INIT_01 => X"A140098018300848180060000C00424040000000080000080200000000110200",
INIT_02 => X"0801080200100000046558000080000041000000002402400800000009008010",
INIT_03 => X"0001000084000040842242000210810803006400088000003080054288C10000",
INIT_04 => X"0000100022008000000C08000800000400A83A2044200C840000000400001820",
INIT_05 => X"0400000080000000248080210044000402000025000800000004203010100800",
INIT_06 => X"00078000600000040410D4102850008024240001981024A82000010461052000",
INIT_07 => X"0800002430204084281000128100000300002040003124040D80204040000888",
INIT_08 => X"0005000108020220240030008000000000043E0408104C800000010000881100",
INIT_09 => X"0004010511100020200000400021004008808060400111080000200002008400",
INIT_0A => X"0000000000010000060210200008B20223048808000200000010024000000000",
INIT_0B => X"03C0411009808245010002000028000080002105010000000020A34249020801",
INIT_0C => X"8004480044800048000480044800448000440002400221008840009012104400",
INIT_0D => X"0000540100000020088000000100100013000400000800040062400200440004",
INIT_0E => X"4100820020000400020000400200204900800000000000000000000100120800",
INIT_0F => X"0000000000101400020401000000002804010401000000002804000000048010",
INIT_10 => X"0000000000000068010400200000002804010400200000002804005000000000",
INIT_11 => X"0050000000000000000000102800024000400000000000000011820010800100",
INIT_12 => X"4000010000000000D00000080004080000002000000000000000000009020000",
INIT_13 => X"00001A000000200000000681000000000000000008004A000400040000000003",
INIT_14 => X"A800040000080000000000000852000020000400000000000010024000002000",
INIT_15 => X"0000000200000000002000000000000000021802000020000000000000000020",
INIT_16 => X"00000040002800100004200009048005C0000080000400000000000000200654",
INIT_17 => X"0802008020080200802008020080200802008020080200800000000000000000",
INIT_18 => X"0000000000000000000080200802008020080200802008020080200802008020",
INIT_19 => X"2054282101000000000000000000000000000000000000000000000000000000",
INIT_1A => X"A28A28A28A28A28A355950666151451453D51A242A503F834E5C49851D243555",
INIT_1B => X"994CA6532994CA6532994CA65328A28A28A28A28A28A28A28A28A28A28A28A28",
INIT_1C => X"FFFFFFFE8E31DCAE532994CA6532995CAE572B94CA6532994CA6572B95CAE532",
INIT_1D => X"AAFFFBC2000000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"555007BFFF55087BE8BFFFFD557400FF842ABEFA2AAA8B5500003DF55F7D568A",
INIT_1F => X"FE0008556ABFFA2D16AB550000021FFF7D17FFEF08042AB55F7D168A00552E95",
INIT_20 => X"3FF55A2D557400557BC2010000000010F7D5421EF007BC01FF5D7FFFE10002AB",
INIT_21 => X"BC0145F7AE801EFF7FBFFF455D7BC0155F7D557545FFAE820AA007BFDFEF5500",
INIT_22 => X"D5400BA082AAAA00FFAE820AAAAAABDFEFF78028BEF005140145A2842AA10F7F",
INIT_23 => X"AD56AB55A2D157400552EBFFEF5D7BD75EF002ABDF555D5157555F7FBC00AAAA",
INIT_24 => X"0000000AAF7D17DE00FFFBD5555A2AABDE00AA803FFEF5D55420BA08557FEBAA",
INIT_25 => X"51C0E3AF55F7DF68ABAE3F1C0000000000000000000000000000000000000000",
INIT_26 => X"7DE3D16DA0041209056D1C71F8F7D147BEFBEFEBD152400F7842FBD7B6AAAAB5",
INIT_27 => X"1EF5D75FFE10142EBAE0008556FBD7B6DB6AB7D1C0A001D7FFD178FC71C0E28B",
INIT_28 => X"2092147BFAFEF49043AF45A2DF504285D71C00101C0005000E3D1401D71C7FC2",
INIT_29 => X"4017DA28428A10E3FFC0145F7A0801FFEBFBF8F6D417BC716DEBD15256DF7AA8",
INIT_2A => X"550545E3F5C20BAAAD5420821C2EAAA00E3AA82092A2AABAFD7EB8A2ABC70855",
INIT_2B => X"51470821C557AE92A2DF6AB7DA2DF50410412ABDFC75D7BD55FF1C2EB8F45555",
INIT_2C => X"000000000000000000000000BAE3D17DE28F7F5D0545B6AAB8E38B68A3AFFF55",
INIT_2D => X"FF803DF45FFAEA8B555D2EAAB45F7FBE8ABAAAD5400000000000000000000000",
INIT_2E => X"5FFD168B55552AA8BEFAAD17DE100804001EF55516ABFF557BFDFEFA2D540010",
INIT_2F => X"10AAD540155557FC01EF5D557DE105D2AA8A0008557FF45FFFFE8BEF5D2E8015",
INIT_30 => X"5FFA2D5401FFF7AA800105D7FE8BEF08002AB45AAFFC00AA5D51400105D04174",
INIT_31 => X"AB55AAAEAAB450055421FFAA8428A00A2FBC0145FF84001EFA2FFEABFF007FD5",
INIT_32 => X"D55FF552EAAB455D5142155AAD1400AAA2D1420005D2EA9A10A2AA82010AAAEA",
INIT_33 => X"AAAABAFFAAAABFF555155400555568A10AAFBEABEFA2FFC0010082ABFF55557B",
INIT_34 => X"00000000000000000000000000000000000000000AAAAD17DEBAFFD142155FFA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"11FFFFFFFFE00000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(10),        -- Port A data input
DOA(0)   => data_read_a_lo(10),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(10),        -- Port B data input
DOB(0)   => data_read_b_lo(10),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_11_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10180B05A0010402840602C2D001019000000300000000330A20080EC180002",
INIT_01 => X"AB400984B83008481800E0000C26426040000000080000088200000802112220",
INIT_02 => X"8801081438106400A4F55800008000004100000040CCE24208005000C9060032",
INIT_03 => X"000406A492E6E440842254D002108153422004800880000030C0315688C00006",
INIT_04 => X"00001201200090001205400000000094108C322644240C840008030440111800",
INIT_05 => X"444000888008010028404002A002009402400025080880000C04223000170900",
INIT_06 => X"40871408620B00801410D94CAAD0018024242008A8102CA88A44010401042200",
INIT_07 => X"08320054B624408428100094ADD080011721A04000316C140CA1A8A1F9001889",
INIT_08 => X"140500090B02C2E0EC04D1C08000000000647E858A104C920C81A5011088A61C",
INIT_09 => X"002481041F165820000101024061004004800567603592A801014C4642601100",
INIT_0A => X"01002020000101B0070310200008B60A23A51B28020CE24E4010026004000440",
INIT_0B => X"03404110230CBA457670820140212100C0692644010001420038935269093161",
INIT_0C => X"2A0872A0C72A0872A0C72A0C72A0872A0C595043950421400800009010104280",
INIT_0D => X"8852141110244066C0820221480010AA73000420808CAC040464D280144050C7",
INIT_0E => X"410082022C000C0002020094030220C960A0409020481024482501A004014100",
INIT_0F => X"6DA02836090540355D86C046619A54052A5B86A0466196940631682800048010",
INIT_10 => X"8B68AA2C60289802AB86A046619A54052A5B86C04661969406316AC018B0E293",
INIT_11 => X"1FC09CB0E1076D4A200B2AC611A3D0405886C6EB211550815A8A2686EC81E2A4",
INIT_12 => X"9C0418CE0C5E8F650E48000892B37885620C1E1A06D7016A90A4626D82B10F1B",
INIT_13 => X"F1E164E02144D335546F28724001B030A56140A184483000C410A2699A2E32AC",
INIT_14 => X"415AAE8018A0A01B2990242E278056AAA203920E0BAE2012C08281808319C186",
INIT_15 => X"9B80D44F9051C049B18A12CB481042AD140C227002A0A02066954E7540CCDB58",
INIT_16 => X"4090240902468118104408000904C0C0964200800200108010003A02272400C1",
INIT_17 => X"0902409024090240902409024090240902409024090240902409024090240902",
INIT_18 => X"1004010040100401004090240902409024090240902409024090240902409024",
INIT_19 => X"2014002840000000000000000004010040100401004010040100401004010040",
INIT_1A => X"0020820820820820A069105251C00000015418982201060302C4281390042104",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFE0FC1C000000000000040200000000000000000001008000000000000",
INIT_1D => X"55000015400000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"B5500003DF55F7D568AAAFFFBC2010557BEAA10AAFBE8A00557BFFFEF007BC21",
INIT_1F => X"75455D7FE8BFF5D7FD540055003FFEFFFD142145000000000FF842ABEFA2AAA8",
INIT_20 => X"C0145557FC2010557FFDF55F7D168A00552E95555007BFFF55087BE8BFFFFD55",
INIT_21 => X"56ABFFA2D16AB550000021FFF7D17FFEF08042AB55A2AAAAB4508517FE00557B",
INIT_22 => X"7FFFE10002ABFE00AAFFE8AAAFF8402000550002145085555400F7FFE8A00085",
INIT_23 => X"8043FEBA002A975EFF7D17DFFFAA8000010000000010F7D5421EF007BC01FF5D",
INIT_24 => X"000000145FFAE820AA007BFDFEF55003FF55A2D557400557BC2145A2D1421450",
INIT_25 => X"8557BF8FEF1C7FC516D080E15400000000000000000000000000000000000000",
INIT_26 => X"00F7842FBD7B6AAAAB551C0E3AF55F7DF68ABAE3F1C00005D7BEDA00B6F1EFA2",
INIT_27 => X"F7D147BEFBEFEBD15257D5D7FEFBD7417BD5438550038FC7FFDF4216D080E070",
INIT_28 => X"DB4514517FE105575C216D5571C50104171FDF7DE3D16DA0041209056D1C71F8",
INIT_29 => X"52400FFF1EFA0008556FBD7B6DB6AB7D1C0A001D7FFD178FC71C0E28B6DA2AEA",
INIT_2A => X"1401D71C7FC21EF5D75FFE10142EBAE10A2FBEFA92F78A05028550E001451455",
INIT_2B => X"71C016DB6D54514500003FEBA1420905FFFFDF78FC7BE84050101C0005000E3D",
INIT_2C => X"0000000000000000000000016DF7AA82092147BFAFEF49043AF45A2DF504285D",
INIT_2D => X"5D7FFDE00F7D17FEBA557BEABEF557BD55EF082A974000000000000000000000",
INIT_2E => X"5F7FBC01FF082A97410FF803DF45FFAEA8B555D2EAAB45F7FBE8ABAAAD540010",
INIT_2F => X"100804001EF55516ABFF557BFDFEFA2D5401FF5D7FFDF55007BD74BA5D042AB4",
INIT_30 => X"B55552AA8BEFAAAABFF5555517FE005555401FF55515541000517FFEFAAD17DE",
INIT_31 => X"74BA5D2A801455D5140000FFD57FE0008557FF45FFFFE8BEF5D2E80155FFD168",
INIT_32 => X"174105D0417410AAD540155557FC01EF5D557DE105D2AA8A10AAFBFFE00F7AA9",
INIT_33 => X"02AB45AAFFC00AA5D51401FFFFD15555500003FEBA5D04001EFFFFFE8B55FF84",
INIT_34 => X"00000000000000000000000000000000000000001FFF7AA800105D7FE8BEF080",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"1000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(11),        -- Port A data input
DOA(0)   => data_read_a_lo(11),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(11),        -- Port B data input
DOB(0)   => data_read_b_lo(11),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_12_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50080B01BC002006940202C0DE041196A83183000000023322287E0FC000006",
INIT_01 => X"0E000C068000E04D40238000001702684000000008000008820009280A553231",
INIT_02 => X"2809AD0E7D180040945008040090000061800000C0E2F66009DA3D11CB148015",
INIT_03 => X"210D050012F6F8D2108216E24842005B8A20640008800000B8E0141C28851006",
INIT_04 => X"0080100022408000060DE0C00466630C70241837041000040800820480001AA4",
INIT_05 => X"04800018800000003C808003E0C8001401000000040900020904004000070800",
INIT_06 => X"00074000601300119E12D348438000803030800020100800AF08000261042400",
INIT_07 => X"8C53200CA4850224301807D1CB45900147E03040083124FC0CD0C8A1FF00198C",
INIT_08 => X"46050013081206A4A503A9E8C0812000001C7E11A24058B84D40E33992D98F7E",
INIT_09 => X"1004810491175C200000820018A5104010C01086003C13E000004EDF02040004",
INIT_0A => X"0000000000010000180018200408B27E234913E9004CFA09A818024800902109",
INIT_0B => X"014100580004304D267C06CCD0056600007827C00000008C00000000000219C0",
INIT_0C => X"2F0C32F0832F0832F0C32F0832F0832F0C197861978400040000208010120ACA",
INIT_0D => X"E0BF40403CFE7E03E8080382FD0018FE670004000006AE01180493C5BC1AF083",
INIT_0E => X"2000401EA0000440000800A0040028108000000000000000000000A74812DF00",
INIT_0F => X"C48DF8362F658A7E5F82CD23B6B0E403DBBE82C563B6A4E403DBB88C0E048200",
INIT_10 => X"454CFBE5403AB992F282C563B6B0E403DBBE82CD23B6A4E403DBBB1084E4B25A",
INIT_11 => X"851000E4B1D32BAB504BB74AD3F3FE04A8E0D0C319A7988B6F0C75CFD801A962",
INIT_12 => X"BEC4118D994B866E2E8C3808B6B63040328E7A33AF99B0AC20DE634D06C437BF",
INIT_13 => X"70CDC5F6214CA5991C6A7177402C49CA354D808D358A927EAD10A652CC8E3538",
INIT_14 => X"49F36E80083C3EAEB2003695430A7CDAA289553922990C11A4E494988231B325",
INIT_15 => X"3BC0FD5B304AD05A946D81616970A225658940BA7CDAA0A312666BD600E5550B",
INIT_16 => X"00000000001000000104200A89A4D0040000008003B81000000021CFEE02E280",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"8020080200802008020000000000000000000000000000000000000000000000",
INIT_19 => X"0544202101000000000000000000080200802008020080200802008020080200",
INIT_1A => X"4124924924924924481C040000B51451440146E518222204D82A5446021090CB",
INIT_1B => X"2C964B2190C86432190C86432190410410410410410410410410410410410410",
INIT_1C => X"FFFFFFFEF001D64B2592C964B2592C964B2592C964B2592C964B2592C964B259",
INIT_1D => X"00AAFBC2000000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"A00557BFFFEF007BC2155000015555087FC0010AAFBFFE100004020BAAAFFD54",
INIT_1F => X"2155AA8400000A2AABFF45550400000AAFBFFFEF550000010557BEAA10AAFBE8",
INIT_20 => X"C0010555155555FF8017400FF842ABEFA2AAA8B5500003DF55F7D568AAAFFFBC",
INIT_21 => X"FE8BFF5D7FD540055003FFEFFFD142145000000145A2AA821EFFFFFD7410007F",
INIT_22 => X"7BE8BFFFFD5574000051420BA557FC2145557FC20AAA2D57DEBAA2FBD55455D7",
INIT_23 => X"82EAAA00550415410AAFBFFFEF55042AB55F7D168A00552E95555007BFFF5508",
INIT_24 => X"000000155A2AAAAB4508517FE00557BC0145557FC2010557FFDE10AA84000000",
INIT_25 => X"0000A02092B6F5D2438A2FBC2000000000000000000000000000000000000000",
INIT_26 => X"005D7BEDA00B6F1EFA28557BF8FEF1C7FC516D080E1557D0075C7028B6F1FAE0",
INIT_27 => X"F55F7DF68ABAE3F1C017DAA8E07028B6A0BFF6D490E00000BEF5FAFEF4904070",
INIT_28 => X"51FFE3FBD0438007FC00385D555556DEB8410400F7842FBD7B6AAAAB551C0E3A",
INIT_29 => X"7DEBAA2FBD557D5D7FEFBD7417BD5438550038FC7FFDF4216D080E0716DAAA08",
INIT_2A => X"09056D1C71F8F7D147BEFBEFEBD152400005F450BA417BC51454971C20AAB6D1",
INIT_2B => X"71FDE10BE8E070280020AAA28410410400BEFBFAFEF49042AB7DE3D16DA00412",
INIT_2C => X"0000000000000000000000016DA2AEADB4514517FE105575C216D5571C501041",
INIT_2D => X"0055574BAFFD568A10002A82000FFD5400AAA2FBC00000000000000000000000",
INIT_2E => X"0FFD568BEF0004174105D7FFDE00F7D17FEBA557BEABEF557BD55EF082A975EF",
INIT_2F => X"45FFAEA8B555D2EAAB45F7FBE8ABAAAD5401EFA2AA974BAF7803FFFF002A8200",
INIT_30 => X"1FF082A975EFA280175FFAAFFC00BA087FC20AA5D55555FFA28000010FF803DF",
INIT_31 => X"75450851420BAFFD57DEAAAAFBD75FF5D7FFDF55007BD74BA5D042AB45F7FBC0",
INIT_32 => X"28BEFAAD17DE100804001EF55516ABFF557BFDFEFA2D540010007FD74AA007BD",
INIT_33 => X"5401FF55515541000517FE10F7AA954AA080428AAA000002010FFFFE8BEF0804",
INIT_34 => X"00000000000000000000000000000000000000001EFAAAABFF5555517FE00555",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"01FFFFFFFFE00000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(12),        -- Port A data input
DOA(0)   => data_read_a_lo(12),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(12),        -- Port B data input
DOB(0)   => data_read_b_lo(12),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_13_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10110A0441812402840402822007818000E00700000000330A3000000008042",
INIT_01 => X"A1400984B830C848180260000C0042404001000008220008A200100802110200",
INIT_02 => X"88010C02801040002475580400800000410000000064024608134C0CC9018034",
INIT_03 => X"00010100926220D084234212421085084300648A0880000630C0654288C10000",
INIT_04 => X"0004122122029100100C00001200009C40A83A2044360C84190BAC04E0101820",
INIT_05 => X"04E000008009050064C8C00104C10184034010250089C00EB004327064B60900",
INIT_06 => X"CA875CA8600000880410DA8C285001802424B008881024A8204E010461042700",
INIT_07 => X"08320014B02848A4A8100015C55500057801A04000712C040CB1F8806000088D",
INIT_08 => X"5005000908020220E40170008042000000557E048A144C800590010000882D00",
INIT_09 => X"00250104B5310020000100020821004016CC1C616401910801010100CA204000",
INIT_0A => X"0000000000010192072310200028B602234608080280074AC010025900100401",
INIT_0B => X"014100101118BA451000824150052110480121000140014200101352690BAC20",
INIT_0C => X"0000000040000000000000040000000000000020000000000000008010102A82",
INIT_0D => X"094040100000006C0802042501001C8017000C21908200028448400000000040",
INIT_0E => X"000000010C000C00081A08BC832A209AB0A85094284A14254A25510105130801",
INIT_0F => X"30BA901293C0F5012906A96DCD13042CE0C206E92DCD07042CE0C40D02048000",
INIT_10 => X"4CA4271CA2168ACB0E06E92DCD13042CE0C206A96DCD07042CE0C4408632C395",
INIT_11 => X"58408632C30D522CE80239CC2806AC44E954939AB299E000738F88296CA13B44",
INIT_12 => X"5145CD5306028F01990C080808494A64708B265CC4052B0F30302E060965EA00",
INIT_13 => X"51E0328A2CA9722094650CCAC0629112BA89C04A228568547B1654B9104A3286",
INIT_14 => X"A158BB80D4D8D48CB54012290470562EC29E44050B1DC60132282B68B9AA60C0",
INIT_15 => X"280000A5C11B9008FE2FA38F87804251CB0FAD40562EC0B426149D17E0044B10",
INIT_16 => X"509425094246A10A10441010090480C0964201800044109012001A000726E454",
INIT_17 => X"0942509425094250942509425094250942509425094250942509425094250942",
INIT_18 => X"9425094250942509425094250942509425094250942509425094250942509425",
INIT_19 => X"7E24502A80000000000000000005094250942509425094250942509425094250",
INIT_1A => X"AEBAEBAEBAEBAEBAFFD7F7F7F775555557DFBEEFBBFCFDF7DFFCF9F80089F7DF",
INIT_1B => X"BF5FAFD7EBF5FAFD7EBF5FAFD7EBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEB",
INIT_1C => X"FFFFFFFE0001DFAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7E",
INIT_1D => X"4500557DE00000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"E100004020BAAAFFD5400AAFBC2155AAAA97410FFFFEAAAAF7AA955EFF7803FF",
INIT_1F => X"5410F7AEBDE10FFFFFDEAAF7D568AAA5D002AB55005568B55087FC0010AAFBFF",
INIT_20 => X"555FF5D04154BAAAAEAAA10557BEAA10AAFBE8A00557BFFFEF007BC215500001",
INIT_21 => X"400000A2AABFF45550400000AAFBFFFEF550000155A28415410F7AEAABFFA2D1",
INIT_22 => X"D568AAAFFFBC21555D517FF45F7AEA8BFFA2AEAAA10A280021EF5D557FF55AA8",
INIT_23 => X"AAE974AAF7D142145082A975FF555568A00FF842ABEFA2AAA8B5500003DF55F7",
INIT_24 => X"000000145A2AA821EFFFFFD7410007FC0010555155555FF80174000055555EFA",
INIT_25 => X"2E3A0925C7E38E38F7D14557AE00000000000000000000000000000000000000",
INIT_26 => X"7D0075C7028B6F1FAE00000A02092B6F5D2438A2FBC2145B6A090428FFF5EAA9",
INIT_27 => X"FEF1C7FC516D080E15438E3A4BAE00FFF5FAE92F7D16AAAA41042FB7D145568B",
INIT_28 => X"2428FFA4AFBFFAAD1505FF490E174AABEA0ADA005D7BEDA00B6F1EFA28557BF8",
INIT_29 => X"001FF555F7FF7DAA8E07028B6A0BFF6D490E00000BEF5FAFEF490407155BE8E1",
INIT_2A => X"AAAB551C0E3AF55F7DF68ABAE3F1C0145415B78F45FFA4AFBC7BEA4AAA10A284",
INIT_2B => X"84104380055525FFBEAE90482E3D54216D0024975FF555F68A00F7842FBD7B6A",
INIT_2C => X"0000000000000000000000016DAAA0851FFE3FBD0438007FC00385D555556DEB",
INIT_2D => X"FF80020BAF7D16AA10A28402155A2AEA8BEF5D516AA000000000000000000000",
INIT_2E => X"A08003DFEF55516ABEF0055574BAFFD568A10002A82000FFD5400AAA2FBC0145",
INIT_2F => X"00F7D17FEBA557BEABEF557BD55EF082A974BAA28028A00F7D16AA10F7D56AAB",
INIT_30 => X"BEF000417545FFAA820BAFF843DFFFA2D5421FF002E954AAFF843DE105D7FFDE",
INIT_31 => X"DF55F7802AA10AA80001FF5D7FFDFEFA2AA974BAF7803FFFF002A82000FFD568",
INIT_32 => X"EAA10FF803DF45FFAEA8B555D2EAAB45F7FBE8ABAAAD540145007FE8B55FF843",
INIT_33 => X"FC20AA5D55555FFA280000BA0855401EFF7AA82010AAD1421FF0004155FF557F",
INIT_34 => X"00000000000000000000000000000000000000001EFA280175FFAAFFC00BA087",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"19FFFFFFFFE00000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(13),        -- Port A data input
DOA(0)   => data_read_a_lo(13),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(13),        -- Port B data input
DOB(0)   => data_read_b_lo(13),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_14_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10020A000180000284008280000281800000030000000033022000000580002",
INIT_01 => X"A140098018300848184860000C20C24040000000084000084200000000110200",
INIT_02 => X"88010C5A8010A600A4F558040080000041000000022C024008003CCCC9028030",
INIT_03 => X"000103A7A00904D0842242024210810803006480088000003081054288C10000",
INIT_04 => X"0000120122009000100C00000000000400A83A2044200C840000800400101820",
INIT_05 => X"040000008008010024C0C0010040000402000025000800020004207000100800",
INIT_06 => X"40870408600800800410D006A850018024240008881024A82040010461042000",
INIT_07 => X"08120054B42850B42A100010ED1500010001A040003164040CF5E20140000888",
INIT_08 => X"400500090A020220A40A7000800000000014FE8508144C924080C10000880140",
INIT_09 => X"0004010411110020000100020021004000800461600191080101000042200000",
INIT_0A => X"0000000000010190070310200008B202236D080802000002C010024000000000",
INIT_0B => X"0141001001088A45000082400000010040012100010000020000135249020820",
INIT_0C => X"0004000000000000004000000000000004000000000000000000008010100000",
INIT_0D => X"0840401000000044080200210100100017000420808200000440400000000040",
INIT_0E => X"0000000000000C00000000040302200800A04090204810244825010104130800",
INIT_0F => X"397468090008142014840100002C382800008401000038382800006402048000",
INIT_10 => X"83514072C000444C00840020002C38280000840020003838280002C09D010868",
INIT_11 => X"03C09D0104B01C57100440202900184414430534605E38048021800224804191",
INIT_12 => X"40049594C194000090450808802008830024F0E248C902AEF0024170CF180010",
INIT_13 => X"8000120020E5A08E6000048200196264BCF1C030C0604800001076C047300002",
INIT_14 => X"A00002003DEDE82C78900902A0D0000080019FAAA32D9602490302409292B832",
INIT_15 => X"2800D049100021171F6C34080240108AB292CA000000800AD1A19F6F000AA0C0",
INIT_16 => X"409024090246810810440000090480C096420080000010801001600001200454",
INIT_17 => X"0902409024090240902409024090240902409024090240902409024090240902",
INIT_18 => X"9024090240902409024090240902409024090240902409024090240902409024",
INIT_19 => X"6504002800000000000000000004090240902409024090240902409024090240",
INIT_1A => X"E79E79E79E79E79E7FDDF77777F3CF3CF7D55E6D39723FC3DEFA75D77B75F7DF",
INIT_1B => X"9FCFE7F3F9FCFE7F3F9FCFE7F3F9E79E79E79E79E79E79E79E79E79E79E79E79",
INIT_1C => X"FFFFFFFEFFFE0FE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F",
INIT_1D => X"55A28417400000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"AAAF7AA955EFF7803FF4500557DF45F7D16AB455D00001EFAAAAAAABA5555575",
INIT_1F => X"214555003FF450804001555D2AA8AAA002ABDE10082ABDF55AAAA97410FFFFEA",
INIT_20 => X"175EF5D5168A10082E80155087FC0010AAFBFFE100004020BAAAFFD5400AAFBC",
INIT_21 => X"EBDE10FFFFFDEAAF7D568AAA5D002AB55005568A00A2D5401455D00175FFFF84",
INIT_22 => X"7BC2155000015400AAD157545080402145087FD75FFF7AE82145A2D17FE10F7A",
INIT_23 => X"000000BAFFFBE8AAAA2FBFDE00087FD5410557BEAA10AAFBE8A00557BFFFEF00",
INIT_24 => X"000000155A28415410F7AEAABFFA2D1555FF5D04154BAAAAEAAA005D002AB450",
INIT_25 => X"7B6A0AAA82555157555B68012400000000000000000000000000000000000000",
INIT_26 => X"45B6A090428FFF5EAA92E3A0925C7E38E38F7D14557AF45FFDB6AB6D4100071C",
INIT_27 => X"092B6F5D2438A2FBC21455D0A3FF6D080407155552AAAA920020BFE10002EBAF",
INIT_28 => X"01454100175C7E380125D7555B6DA1014248217D0075C7028B6F1FAE00000A02",
INIT_29 => X"82145AAD178E38E3A4BAE00FFF5FAE92F7D16AAAA41042FB7D145568A38AADF4",
INIT_2A => X"1EFA28557BF8FEF1C7FC516D080E15400A2DB5754508040716D007BD05EFEBAA",
INIT_2B => X"A0ADA0055002AB6D0000020BAFFF1E8ABABEF1FAE001C7FD54005D7BEDA00B6F",
INIT_2C => X"00000000000000000000000155BE8E12428FFA4AFBFFAAD1505FF490E174AABE",
INIT_2D => X"F7FFEABFF080015555F78028A00555155555FF84000000000000000000000000",
INIT_2E => X"000003DE10082EAAB45FF80020BAF7D16AA10A28402155A2AEA8BEF5D516AB45",
INIT_2F => X"BAFFD568A10002A82000FFD5400AAA2FBC0145552ABFFFF000417555552EA8A1",
INIT_30 => X"FEF55516AABAAAFFC0145000417555A280001455D7FFDE105504021EF0055574",
INIT_31 => X"55FF007BC01FFAAAE80155AAD568ABAA28028A00F7D16AA10F7D56AABA08003D",
INIT_32 => X"D74105D7FFDE00F7D17FEBA557BEABEF557BD55EF082A97410AAFFD554508001",
INIT_33 => X"5421FF002E954AAFF843DE10550028BEF0004020BAF7D568AAAF7D168A105D7F",
INIT_34 => X"0000000000000000000000000000000000000000145FFAA820BAFF843DFFFA2D",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"01FFFFFFFFE00000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(14),        -- Port A data input
DOA(0)   => data_read_a_lo(14),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(14),        -- Port B data input
DOB(0)   => data_read_b_lo(14),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_15_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000A000000000284000280000001800020030000000033022000000180002",
INIT_01 => X"A140098018300848180060000C00424040000000080000080200000000110200",
INIT_02 => X"080108000010E60004E55800008000004100000000040240080000C009170016",
INIT_03 => X"0000000080000040842240000210810002000400888000003080014288C00000",
INIT_04 => X"0001100024A0800000440000000000040088322044200C840000011400151800",
INIT_05 => X"440002988000000020000000000B8094020000254C8800000514203000108800",
INIT_06 => X"00070000620040880410D00C285000802424000AA81024A80040010C01062001",
INIT_07 => X"086100043224489428100010811100010001A040003124040CAC600040000888",
INIT_08 => X"160500090A0282A06400100080C300000005BE0488104C800000010000880000",
INIT_09 => X"000581041110022000000002002100400080046140011008010100008A040000",
INIT_0A => X"0000000000010180060210200008B2022304080800000007C010024000000000",
INIT_0B => X"4140001001088A45000082000000010000002000010000020000034249000020",
INIT_0C => X"0004000040000400000000000000000004000020000200000000008010100000",
INIT_0D => X"094000100000004C000200250000188016000400000000000440400000000040",
INIT_0E => X"0000000108000C00000000000200200800800000000000004020000000000000",
INIT_0F => X"0000000000000000000404200000000000000404200000000000008C00048000",
INIT_10 => X"4000000000000000000405000000000000000405000000000000004000001000",
INIT_11 => X"0040000010000000000000000000004000201000000000000000000000800002",
INIT_12 => X"0004000110000000000C00080010180000000001A10240500000000000000000",
INIT_13 => X"0000000020080400000000020000008040020000000000000010001200000000",
INIT_14 => X"0000020000000611002800000000000080000011044220000000000080200200",
INIT_15 => X"8800000100000000009080E2E0A0000000000000000080000040000000000000",
INIT_16 => X"0000000000460000004400000904808094020080000010000000000000000041",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0004002800000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000004000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFE00000000000000000000000000000000000000000000000000000000",
INIT_1D => X"EF08517DE00000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"1EFAAAAAAABA555557555A284175FF000002010552A97400007BFDE10A2AA801",
INIT_1F => X"DFEF5D2AAAB45F7D17DF45087BC0155002A801FF08003DF45F7D16AB455D0000",
INIT_20 => X"C2145F7D568BEFAAD557555AAAA97410FFFFEAAAAF7AA955EFF7803FF4500557",
INIT_21 => X"03FF450804001555D2AA8AAA002ABDE10082ABDFFFF7D17FE10002E954AAF7FB",
INIT_22 => X"FFD5400AAFBC21EFA2AE95545A2D56ABFFAAD17DE10FFD1420AA007FC0145550",
INIT_23 => X"02A801550055401555D00174BA002AA8B55087FC0010AAFBFFE100004020BAAA",
INIT_24 => X"000000000A2D5401455D00175FFFF84175EF5D5168A10082E801FFFF8428A100",
INIT_25 => X"80871FAE00A2A0871EF145B7FE00000000000000000000000000000000000000",
INIT_26 => X"45FFDB6AB6D4100071C7B6A0AAA82555157555B680125C71C0E0500049209543",
INIT_27 => X"5C7E38E38F7D14557AFC75524AFB45FFD178F7D1C71C2145002E801C7140A3FF",
INIT_28 => X"AE000024954AAFFFBC2145F7DB6DBEFA2D557545B6A090428FFF5EAA92E3A092",
INIT_29 => X"470820071C71455D0A3FF6D080407155552AAAA920020BFE10002EBAFC7FFDF7",
INIT_2A => X"1FAE00000A02092B6F5D2438A2FBC21FFBEA090545B6D568BFFAADB7AE10F7D5",
INIT_2B => X"24821FFE3802FA2808208017D1C5142155410A104AA1420AFB7D0075C7028B6F",
INIT_2C => X"00000000000000000000000038AADF401454100175C7E380125D7555B6DA1014",
INIT_2D => X"552E954100004174AA00516AA10AA80155EF5D7BFDE000000000000000000000",
INIT_2E => X"5082E801555D2EBDF45F7FFEABFF080015555F78028A00555155555FF8400155",
INIT_2F => X"BAF7D16AA10A28402155A2AEA8BEF5D516AB555D043DF55F7D56ABEF55514015",
INIT_30 => X"E10082EAAB55FFFBE8A100804154AAF7FFC2145FFFFFDFEFAAD157545FF80020",
INIT_31 => X"ABEFA2FBE8A00FFD155410005555545552ABFFFF000417555552EA8A1000003D",
INIT_32 => X"3DFEF0055574BAFFD568A10002A82000FFD5400AAA2FBC01FFF78400155F7D16",
INIT_33 => X"0001455D7FFDE105504021FFAA843DEBA0000021EF555142155002E800AA5500",
INIT_34 => X"00000000000000000000000000000000000000000BAAAFFC0145000417555A28",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"1800000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(15),        -- Port A data input
DOA(0)   => data_read_a_lo(15),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(15),        -- Port B data input
DOB(0)   => data_read_b_lo(15),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_16_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"DA22C618B1000482B688B186588884862A400438255FC38381441205BA803003",
INIT_01 => X"8645A80028404C211203A952A90341080B173340412000E1005D628000820484",
INIT_02 => X"A101A9006DC1084833011850AAC55001349B10881802821808B4110007005E11",
INIT_03 => X"010108A802BB00080080006020020001A61036202800000D2410104200404550",
INIT_04 => X"8BFA58800005C40A46240252145148B38248030356415A4E62B6FC660F287240",
INIT_05 => X"1E0BD423CAC0000D610000000710296E542B6E3A825C15FB30A643695BFC2D56",
INIT_06 => X"000D0000C8008820CAE16020619156A5815006028179808C00A0D2152B90707A",
INIT_07 => X"F500240510A00205F0A407D0021A155378900002A002433A0AA00EE6E7956108",
INIT_08 => X"015995440C8327241440096A2800002828123D542910380004E0310362404076",
INIT_09 => X"10222D90409A05B2CB2CA400200209E5601044A24000000462A6001888010000",
INIT_0A => X"0000000000259200140001A15000017F0051D0F837248C005514AC40C0820500",
INIT_0B => X"01200848002912300200092BA80325A2000000000001514B5500030241C000CC",
INIT_0C => X"0001100011000110001100011000110001080008800080005202280801080395",
INIT_0D => X"17680002815014B90000205DA00880100095A64800008003561180063DB4F611",
INIT_0E => X"0280080922554515512174000000490009000000000000004010042A204A0C58",
INIT_0F => X"2DA0063EAA9C238B2D4C800632B266E828EE4C800632AAAB6830D0FC6B06C041",
INIT_10 => X"0839AA149339E8FB964C800632B266E82B2E4C800632AAAB683310872800EDA5",
INIT_11 => X"C087A800EB090D4AAC91268FFCBE81397826C4A20D2B6C510E8624792A4A30A4",
INIT_12 => X"3638E8849D5C532408DD6E004C90C06AC019D88B9795012CA96902C799912BC3",
INIT_13 => X"78706531C74485BD42A30906057FADAA456218FD8E3ED83B60E3A242DC0F1898",
INIT_14 => X"51727A06FB555793057C444CF45C5C9E89543B8BC6E80193DC36F6C71D1093A4",
INIT_15 => X"10DCD45DC02B331650CA8ACB4007E00D1C6A6A58395C917F7E74D936F650D69B",
INIT_16 => X"000000000012000081500008A422150884081ACAAC0542054004FC5884640508",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"3604000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"45145145145145147A7797E1E1A79E79E15634455131A436993071A616D4F68A",
INIT_1B => X"3E9F4FA7D1E9F47A7D1E9F47A7D3453453453453453453453453453453453453",
INIT_1C => X"FFFFFFFE00001F4FA7D3E9F4FA3D1E8F47A3D1E8F47A3D1E9F4FA7D3E9F4FA7D",
INIT_1D => X"00FF8015400000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"400007BFDE10A2AA801EF08517DE10FFFFFDFEFA2D16AB55A2FFFFEAA5D7FC00",
INIT_1F => X"74BA5D2EBDFEFAAD17FFFF002EBDE000800174AA55043FFFF000002010552A97",
INIT_20 => X"E8AAAAA80000105D557FF45F7D16AB455D00001EFAAAAAAABA555557555A2841",
INIT_21 => X"AAAB45F7D17DF45087BC0155002A801FF08003DE000004154BA002A800BA087F",
INIT_22 => X"803FF4500557DEAAF7D57DEBA082A82010FFAE975555D7FFDEAAFF80155EF5D2",
INIT_23 => X"2D57FFFF557FD55FF08003FE0055043FF55AAAA97410FFFFEAAAAF7AA955EFF7",
INIT_24 => X"0000001FFF7D17FE10002E954AAF7FBC2145F7D568BEFAAD557410552EA8BEFA",
INIT_25 => X"DB6FFFDEAA5571C7010FF8412400000000000000000000000000000000000000",
INIT_26 => X"C71C0E050004920954380871FAE00A2A0871EF145B7FE10E3F1F8FC7AAD56DB7",
INIT_27 => X"A82555157555B680124924124BDFEFA2D57FFC71C2EBDE280000174825D0E3FF",
INIT_28 => X"74821424800AA007FEDAAAA284020385D5F7AF45FFDB6AB6D4100071C7B6A0AA",
INIT_29 => X"F8EAAFF80175C75524AFB45FFD178F7D1C71C2145002E801C7140A3FE10080A1",
INIT_2A => X"5EAA92E3A0925C7E38E38F7D14557AE92EBDB78EAA1C2482010FFAE9556D557F",
INIT_2B => X"D557410492EADBEFA2D178FEF5575D55EF000A38E10490A3AF45B6A090428FFF",
INIT_2C => X"000000000000000000000001C7FFDF7AE000024954AAFFFBC2145F7DB6DBEFA2",
INIT_2D => X"A2D56AB45A2D57DFFFF7FBFFEAA555555400F780000000000000000000000000",
INIT_2E => X"A080415400552ABDF55552E954100004174AA00516AA10AA80155EF5D7BFDE10",
INIT_2F => X"FF080015555F78028A00555155555FF840000000043DFEFAAD17FF45552ABFEB",
INIT_30 => X"1555D2EBDE10002E974005D04020BA007BFDEBAA284000BA557FE8B45F7FFEAB",
INIT_31 => X"0000F7AE955EF5D7BE8ABAF784175555D043DF55F7D56ABEF555140155082E80",
INIT_32 => X"AAB45FF80020BAF7D16AA10A28402155A2AEA8BEF5D516AA00AAFBE8AAA55040",
INIT_33 => X"FC2145FFFFFDFEFAAD157410082ABFFEFAAD16ABFF5555575FF082AA8A00002A",
INIT_34 => X"0000000000000000000000000000000000000000155FFFBE8A100804154AAF7F",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0800000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(16),        -- Port A data input
DOA(0)   => data_read_a_lo(16),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(16),        -- Port B data input
DOB(0)   => data_read_b_lo(16),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_17_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"5284CE4FB7BD2C8994A13392DBD02E14006B82AC7E800D44D3DD2FD5F9B961C0",
INIT_01 => X"F8ACD01F7E03FC6793F2199B39FC233C11D93AE6F3BB92B32091DBC339B24542",
INIT_02 => X"8F333007FD6808092A2AFA6667033DB50853379C10BFF70F1BD011110F205F18",
INIT_03 => X"294ADB4AFFCBF0DAD63ABF836B58EAFE060478202022234B2E0303FDC9E18339",
INIT_04 => X"DB7A40806FE4040840EBC563A0150A0926146FECB04196482236FC2005282AE1",
INIT_05 => X"0807B4070670083DC68206D7E6D0250834336D1E81500FDB306045255BFC2076",
INIT_06 => X"00000000141C5AF3EA6AB187F7F8CE039786062C6CE092F5FE005236781C402A",
INIT_07 => X"1684248A38B022475DCA9BD00116E33CC3821774BB55F53BB42329AA3C0CEF60",
INIT_08 => X"60700CE0641527241060AD844E1C0088001223022D189A2800542219204903F8",
INIT_09 => X"D94C1C1C51DFF881861CBE0305A12A0321810217C01D34EDC98FFA1C8E000016",
INIT_0A => X"7E7D8F8FBDE40E001E000B3A5DAADAFDDA5DA79350DF70027CE86F047BEF19B6",
INIT_0B => X"814102F800633F1D0A7CC9AE74117FE0003A6AD055819D1F9984014B37BA5FFC",
INIT_0C => X"CF4FBCF4FBCF4FBCF4FBCF4FBCF4FBCF4FBE7A7DE7A7800617112E46F05D02DD",
INIT_0D => X"D7FE4A5A99FD6D3FEF4BEB5FF994F0FEFFCCF8430006CE8A3F06ABD73DBCF4FB",
INIT_0E => X"B29760593F33FA0CF170F40006001B1A05C0000000000000008004BA78428C7A",
INIT_0F => X"EDA57E46444357B3950A9BFBAC94CFA8581E0A9BFBAC8CCFA8580C7CAF51EF68",
INIT_10 => X"7DF76B5DB54A09003E0A9BFBAC94CFA8581E0A9BFBAC8CCFA8580E46FBFCB0CB",
INIT_11 => X"E7467BFCB1D5CFEB56A1A100D5345C1BFFE8FBDB892DB463034198E2881F3F78",
INIT_12 => X"4E0ADD39387F92B2935DFEAADDF38EBCFB9E3D636DCDF9B90F966BF92966D5D9",
INIT_13 => X"F256527055EB6D555CB294981B7FB5B2954CD3013013FDF5E82AF5B6AAAE594A",
INIT_14 => X"F7D7E835C67E655BAA868610117575EA1C34BD6975D48B44A0405FC15BA7270F",
INIT_15 => X"BD07F6CD2A47D0CBA96252756D7217E5E1C61DBDF5FA167F7AE5D3D21A414007",
INIT_16 => X"00000000005F08000179C16DECF67F08BC02F9067ED55805600545DFE45A80E7",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"F981800C00000000000000000000000000000000000000000000000000000000",
INIT_1A => X"A69A69A69A69A69A919261A1A6075D75D10DC800C027B731014BA4B864617114",
INIT_1B => X"8341A0D068351A8D068351A8D069A6BAE9A69A6BAE9A6BAE9A69A6BAE9A6BAE9",
INIT_1C => X"FFFFFFFE000011A8D46A351A8D46A351A8D46A351A8D46A341A0D068341A0D06",
INIT_1D => X"55AAFFD5400000000000000000000000000000000000000000000001FFFFFFFF",
INIT_1E => X"B55A2FFFFEAA5D7FC0000FF8015410FFFFFFFFFFFFFFDFEFF7D568A1008003DF",
INIT_1F => X"DF55A2D1400000804154BAF7D168A00A2803DE10FFAE95410FFFFFDFEFA2D16A",
INIT_20 => X"2AABAFFD56ABFF002EBDFFF000002010552A97400007BFDE10A2AA801EF08517",
INIT_21 => X"EBDFEFAAD17FFFF002EBDE000800174AA55043FEBA0004174AA5504000AA5504",
INIT_22 => X"5557555A284175FFFFFBE8B55A2FFFFF55F7803DEBA002AAAAAAF7FBD74BA5D2",
INIT_23 => X"D0417400FFD57DE00AAAAAAB45A2AA97545F7D16AB455D00001EFAAAAAAABA55",
INIT_24 => X"0000000000004154BA002A800BA087FE8AAAAA80000105D557FE00A2D5420AA5",
INIT_25 => X"7EBD16AA00000E3DF6DBEF5D2400000000000000000000000000000000000000",
INIT_26 => X"10E3F1F8FC7AAD56DB7DB6FFFDEAA5571C7010FF8412428FFFFFFFFFF7FBF8FD",
INIT_27 => X"E00A2A0871EF145B7FF7DA2D547038140E10492FFDF6DA28A28E3DE00F7A0924",
INIT_28 => X"2492550A020BA55002AA82F7DF6DBD71C2EBFFC71C0E050004920954380871FA",
INIT_29 => X"ADABAF7F5D74924124BDFEFA2D57FFC71C2EBDE280000174825D0E3FEAA14001",
INIT_2A => X"0071C7B6A0AAA82555157555B680125FFEBFFEDB55BEFFFAF6DE38E3DEAA002E",
INIT_2B => X"5F7AE28B6D545092490E10400FFDB7AE00A2AAADB45BEA092545FFDB6AB6D410",
INIT_2C => X"00000000000000000000000010080A174821424800AA007FEDAAAA284020385D",
INIT_2D => X"FFFBFDFEFF7FFEAB45A2D56AA00002EBDFFFF7D5400000000000000000000000",
INIT_2E => X"AA2AABDE10FF8400010A2D56AB45A2D57DFFFF7FBFFEAA555555400F780000AA",
INIT_2F => X"100004174AA00516AA10AA80155EF5D7BFDFEFAAD1554BA552E82000F7FFFFEA",
INIT_30 => X"400552ABDEBA5D0002000552A800BA55042AA10FFFFFDF55552EBDF55552E954",
INIT_31 => X"ABFFA2AEBFEAA082EBDEBAFFD55540000043DFEFAAD17FF45552ABFEBA080415",
INIT_32 => X"00145F7FFEABFF080015555F78028A00555155555FF84001FFAAFBFFF55FFFBE",
INIT_33 => X"BFDEBAA284000BA557FE8AAAFFD155400082A82000F7FFE8A00A2AABDF45F780",
INIT_34 => X"0000000000000000000000000000000000000000010002E974005D04020BA007",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"19FFFFFFFFE00000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(17),        -- Port A data input
DOA(0)   => data_read_a_lo(17),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(17),        -- Port B data input
DOB(0)   => data_read_b_lo(17),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_18_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"69844019080000A21A611406840014122A641074155FC28A2024001001801003",
INIT_01 => X"A643D920034004180005E9E3C90360C0041C0181002001602025800008440084",
INIT_02 => X"B7333980808408103F2000F81FC0FEDEAC2161B0B84D0002188011110C018041",
INIT_03 => X"0405D434003F2C020081587008020561E55116B0290000042B71240C800440F8",
INIT_04 => X"50805AC31007D6125724029216554A9847669903D640EC8E2001002604503004",
INIT_05 => X"0E010001C1CA11803850C800010022660C1C0065003C0404002646DC20A02D40",
INIT_06 => X"50AD050AC00000002A4F612449903FE080000000005889AC41E04508A9907020",
INIT_07 => X"5584280B10014003A8067400920810FF3C72024300A0030048221ACEE383E518",
INIT_08 => X"00C983E6041505253500F66E620428000B1804000152E52801A2020084090040",
INIT_09 => X"20500B90419005B0C309402030060860E01004A828408800440405E350294010",
INIT_0A => X"008010100007865421432121804021C20452880C2D200000045C18C0E0000A08",
INIT_0B => X"09700C04C44C92A88DC42215C882E82250811000000C1AE061861710A401A4E8",
INIT_0C => X"308003080030800308003080030800308001840018400400602A018809800371",
INIT_0D => X"0801010202021000780004200408C1002003F66CA1B13111C0D95C20C2030A00",
INIT_0E => X"02900806400FC503F08180050942E4200020C1B060D8306C182701404C197301",
INIT_0F => X"22AABABAF377DF1CA160820520EB3057E70E60820520F33057E72E9154159000",
INIT_10 => X"8A2AD5D48F37FAFEFE60820520EB3057E7CE60820520F33057E7EC658BF2DA78",
INIT_11 => X"32658BF2D4B2A80BF8FE39FD78EB0D882014A62C568FFAFC73FFDD9C2B30E046",
INIT_12 => X"C728C800DFC06F59F710107533C0C4E37619440FBFBAB2400AFC1600361D798F",
INIT_13 => X"0DEBBEB9454005BAA36DEFF894823A3D1A88A2FE29D5FC6DCAA2A002DD51B6E7",
INIT_14 => X"F3B7092A78606A28A5427AAB9FF4EDD251C7123E291660733EBF6FE519001BF4",
INIT_15 => X"82202AB58AFBFD5DE200A8EBE3A3EC110339E1DCEDC2590495BB2112E2BE4BF5",
INIT_16 => X"C1B06C1B06808348340000020301805002D008C1F92000A5F421B8000DB49103",
INIT_17 => X"1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06",
INIT_18 => X"B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C",
INIT_19 => X"16000000000000000000000000041B06C1B06C1B06C1B06C1B06C1B06C1B06C1",
INIT_1A => X"A28A28A28A28A28A244C16454170410412CA2EFB3AE03B85CF08C03F1A30F7DF",
INIT_1B => X"8944A25128954AA552A944A2512AAA8A28A28A2AAAAAA8A28A28A2AAAAAA8A28",
INIT_1C => X"FFFFFFFE000004A25128944A25128944A25128944A25128944A25128944A2512",
INIT_1D => X"105D2A80000000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"FEFF7D568A1008003DF55AAFFD5410FFFFFFFFFFFFFFFFFFFFFBFDEBA552E974",
INIT_1F => X"5410FFFFFFFFFF7FBE8B55AAD16AA1000516AA005D0400010FFFFFFFFFFFFFFD",
INIT_20 => X"FFE00087BC2155087BC0010FFFFFDFEFA2D16AB55A2FFFFEAA5D7FC0000FF801",
INIT_21 => X"1400000804154BAF7D168A00A2803DE10FFAE95555FFFBE8B45A2D56ABEFFFFF",
INIT_22 => X"AA801EF08517DF55000000010082A974AA08557DEBAFFAEBFF55AA8028B55A2D",
INIT_23 => X"52E800105D2AAAA10A2D1420AAFFAEA8BFF000002010552A97400007BFDE10A2",
INIT_24 => X"0000000BA0004174AA5504000AA55042AABAFFD56ABFF002EBDEBA0004020BA5",
INIT_25 => X"FF7FBFFEBA552A95410552485000000000000000000000000000000000000000",
INIT_26 => X"28FFFFFFFFFF7FBF8FD7EBD16AA00000E3DF6DBEF5D2438FFFFFFFFFFFFFFFFE",
INIT_27 => X"EAA5571C7010FF8412410FFFBF8FC7E3F5EAB45BEDB6FA3800556FA005504050",
INIT_28 => X"AB55BEDB6FBC7EBF5F8E10007BC516D1C71C5010E3F1F8FC7AAD56DB7DB6FFFD",
INIT_29 => X"BFF55BE8A2DB7DA2D547038140E10492FFDF6DA28A28E3DE00F7A09256DE3F1E",
INIT_2A => X"0954380871FAE00A2A0871EF145B7FF45080E070280820924AA145578E92F7A4",
INIT_2B => X"2EBFEBA1C0A00092412E850005D2AAFA38A2DF45082F7AAA8BC71C0E05000492",
INIT_2C => X"000000000000000000000000AA140012492550A020BA55002AA82F7DF6DBD71C",
INIT_2D => X"FFFFFFFFFFFFBFDFEFF7FFFDEAA5D2E954105504154000000000000000000000",
INIT_2E => X"A08557DE005500154AAFFFBFDFEFF7FFEAB45A2D56AA00002EBDFFFF7D5400AA",
INIT_2F => X"45A2D57DFFFF7FBFFEAA555555400F78000010F7FBE8B55AAD16AB55F7FBFDEA",
INIT_30 => X"E10FF84001FFAAD568B45FFFBFFF55A2D568A00087BD55FF5D5555410A2D56AB",
INIT_31 => X"00AA555168A10FF803DF45FFAABDFEFAAD1554BA552E82000F7FFFFEAAA2AABD",
INIT_32 => X"A8B55552E954100004174AA00516AA10AA80155EF5D7BFDF45002A974AA08000",
INIT_33 => X"42AA10FFFFFDF55552EBDEBA5D2E80010082A97410552EBDEBAA2FBD5400F7AA",
INIT_34 => X"00000000000000000000000000000000000000000BA5D0002000552A800BA550",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0800000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(18),        -- Port A data input
DOA(0)   => data_read_a_lo(18),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(18),        -- Port B data input
DOB(0)   => data_read_b_lo(18),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_19_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"042200000000000041088001001AA00000000000000000000000500802000003",
INIT_01 => X"200048000024000000000404000000000A22000800000800004A200000000001",
INIT_02 => X"032210008DEF00400060000001C008002489E0F0004037B00010101010000000",
INIT_03 => X"0000008128000000000000000000000024001620280000000000354200004008",
INIT_04 => X"000058800004C4024024001210001054B1C822009640000E2000002604003000",
INIT_05 => X"0E010001C0400000000000000000200604000000001C04000026400000002C40",
INIT_06 => X"000000000000000001800166A84004A080000000005884020020400009907020",
INIT_07 => X"E200201C00A14080082B26208008A00900120101402240440280040840802000",
INIT_08 => X"004180261C81210031000004340000200008105428020568040213003499C006",
INIT_09 => X"00000990000000B0C30800000000086020016000000000003838000000000000",
INIT_0A => X"000000000005860000000080A000206020408000000000000454080000000000",
INIT_0B => X"00000000000040002000044000000000000000000005E0003E00004049640004",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"00000000210001D8000000000000000020009640000000000000000000000000",
INIT_0E => X"040000000000C500300080000000000000000000000000000000000000000000",
INIT_0F => X"50500101088A37034E156600D740022800EC156600D740022800D01E0412D069",
INIT_10 => X"E61700224081044914156600D7400228002C156600D7400228001098F00D0FB7",
INIT_11 => X"CC98F00D0F2DD014010046037814EA63DBB31CE7605001008C41A061F0E7D693",
INIT_12 => X"361526D600000004089E12350C0E01FF23315422BABB46FEF5019146C0800380",
INIT_13 => X"00000130AA3592000000000629C03F3E60330C00C628908214551AC900000010",
INIT_14 => X"4208D65C006070845039014460088235ACC3123E2A29148841008482A4DAC000",
INIT_15 => X"6CD4953A66BE7A5040018D8A8AD9090A1EC20A188235AC509FB50C2D0500B409",
INIT_16 => X"00000000000000000000000000000000000008C0180027000006110008404608",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"9200000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"61861861861861861A2882313054D34D301C822EE8FC31C043198028002C7441",
INIT_1B => X"84C261349A4C26130984C261309861861861A69861861861861A698618618618",
INIT_1C => X"FFFFFFFE0000026130984C26130984C26130984C26130984C26130984C261309",
INIT_1D => X"00082E97400000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"FFFFFFBFDEBA552E974105D2A801EFFFFFFFFFFFFFFFFFFFFFFFFFEAA552E954",
INIT_1F => X"55EFFFFFFFFFFFFFFFFFEFF7FBFFEAA5D2E97545FFFFC2010FFFFFFFFFFFFFFF",
INIT_20 => X"6AA0008003DF555D5157410FFFFFFFFFFFFFFDFEFF7D568A1008003DF55AAFFD",
INIT_21 => X"FFFFFFF7FBE8B55AAD16AA1000516AA005D04001EFFFFFFFFFFFFFBFDF45AAD1",
INIT_22 => X"7FC0000FF80155EFFFFFFFFEFF7D16AB55A2D57DEBA557FEAA10080402010FFF",
INIT_23 => X"2D56AB45FFFBFDEBA5D7FC0155FFFFD7410FFFFFDFEFA2D16AB55A2FFFFEAA5D",
INIT_24 => X"000000155FFFBE8B45A2D56ABEFFFFFFFE00087BC2155087BC00AAFFFBFDF45A",
INIT_25 => X"FFFFFFDEAA552E95400002095400000000000000000000000000000000000000",
INIT_26 => X"38FFFFFFFFFFFFFFFFEFF7FBFFEBA552A954105524851C7FFFFFFFFFFFFFFFFF",
INIT_27 => X"A00000E3DF6DBEF5D25D7FFFFFFFFFFFFBFDFEFEBF5F8E92552E9556DEBF1C20",
INIT_28 => X"DFEFE3F1FAF55A2D568A0000003FF7D495155428FFFFFFFFFF7FBF8FD7EBD16A",
INIT_29 => X"EFA00000002010FFFBF8FC7E3F5EAB45BEDB6FA3800556FA005504051FFFFFFF",
INIT_2A => X"56DB7DB6FFFDEAA5571C7010FF84125EFF7F1F8FC7EBD568B6DBEDF7DEBA5571",
INIT_2B => X"71C5092E3F1F8F55AADB6DB7DEBF1FAE82557FC516DEBF1D0410E3F1F8FC7AAD",
INIT_2C => X"0000000000000000000000016DE3F1EAB55BEDB6FBC7EBF5F8E10007BC516D1C",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFBFDEAA5D2A954000800154000000000000000000000",
INIT_2E => X"0552A955EFAAD1400AAFFFFFFFFFFFFBFDFEFF7FFFDEAA5D2E95410550415545",
INIT_2F => X"EFF7FFEAB45A2D56AA00002EBDFFFF7D540145FFFFFFFEFF7FBFFFFFAAD16AA0",
INIT_30 => X"E005500155EFF7FBFDFEFAAD568B55AAD568A0008003DFFF0855554AAFFFBFDF",
INIT_31 => X"ABEFFFFFFFEAA55517DE10080400010F7FBE8B55AAD16AB55F7FBFDEAA08557D",
INIT_32 => X"40010A2D56AB45A2D57DFFFF7FBFFEAA555555400F780001FFF7D16AB55A2D16",
INIT_33 => X"568A00087BD55FF5D5555410AAD56AB45AAFFFFFEFAAD168A00557BD55FFA2D5",
INIT_34 => X"00000000000000000000000000000000000000001FFAAD568B45FFFBFFF55A2D",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"1000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(19),        -- Port A data input
DOA(0)   => data_read_a_lo(19),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(19),        -- Port B data input
DOB(0)   => data_read_b_lo(19),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_20_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000003",
INIT_01 => X"A75FF80000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"14088080800008400F655001FFCFF80018FA8044000000000000011000000007",
INIT_03 => X"0000000000000000000000000000000024001660380000000000000000004FF8",
INIT_04 => X"000079800014CC02C034001600000000000000101EC0012EE0C0026E1E80F000",
INIT_05 => X"3E1FE867DFC044003902100002203F2EFC040388137C3E20C8EEC00284033CC0",
INIT_06 => X"001F0001E0020002E80020000005FEAF91D10802ABFB80000021C8010FB0F0F4",
INIT_07 => X"00040007700000000000000001080FF900160000000200C00080001840BFE538",
INIT_08 => X"09FFBFE5181606000410A4000004202AA8043E0000000000000001209244C040",
INIT_09 => X"01227FB0000000F7DF78020004011FEFE0000000002003150200008388020000",
INIT_0A => X"000000000015BE0000004000000100000100506002008C2007D5FC8000002400",
INIT_0B => X"0000000000000000000000000000000400400520000000000000000400000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000020002",
INIT_0D => X"00010000000200000020000004000100203FF6C0000000000000000000000000",
INIT_0E => X"0000000600FFC53FF001800000002004080000000000000040900005C8485380",
INIT_0F => X"8000000009A9C300020080000800000003CC0080000800000003CC0200078000",
INIT_10 => X"00800000000012963C0080000800000003CC0080000800000003CC1008000000",
INIT_11 => X"00100800004000000000066C5000020020000000800000000C2E180010002000",
INIT_12 => X"96004000000000052B0200000014200040C2829000400000000000860F987980",
INIT_13 => X"0000A4B00400000000002958000240400000000007E1B0000402000000000014",
INIT_14 => X"400004004181800000000005C5A00000200C40808000000000AF0D8008000000",
INIT_15 => X"000800020141812737DC3020100400001C19C1D80000200400000000000015D1",
INIT_16 => X"0000004010080800801810100000000000093EDFF80200000000000010010010",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"4D20400200000000000000000000000000000000000000000000000000000000",
INIT_1A => X"CB0C30C30C30C30C8192608486879E79E681C000C00E08000402241560412010",
INIT_1B => X"2190C86432190C86432190C86432CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2",
INIT_1C => X"FFFFFFFE000010C86432190C86432190C86432190C86432190C86432190C8643",
INIT_1D => X"10080402000000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"FFFFFFFFFEAA552E95400082E975FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2A954",
INIT_1F => X"0000FFFFFFFFFFFFFFFFFFFFFFFDEAA5D2A954000800001EFFFFFFFFFFFFFFFF",
INIT_20 => X"FFEBA5D2A97400FF8017410FFFFFFFFFFFFFFFFFFFFFBFDEBA552E974105D2A8",
INIT_21 => X"FFFFFFFFFFFFFEFF7FBFFEAA5D2E97545FFFFC21FFFFFFFFFFFFFFFFFFFFF7FB",
INIT_22 => X"003DF55AAFFD5400FFFFFFFFFFFFFFDFEFF7FFEAA10000417555AAD5555EFFFF",
INIT_23 => X"FFBFDFEFAAD568A0000043DF45AAFBC2010FFFFFFFFFFFFFFDFEFF7D568A1008",
INIT_24 => X"0000001EFFFFFFFFFFFFFBFDF45AAD16AA0008003DF555D51574BAFFFFFFFFFF",
INIT_25 => X"FFFFFFFEBA5D2A95410000A00000000000000000000000000000000000000000",
INIT_26 => X"C7FFFFFFFFFFFFFFFFFFFFFFFDEAA552E954000020955FFFFFFFFFFFFFFFFFFF",
INIT_27 => X"EBA552A95410552485010FFFFFFFFFFFFFFFFFFF7FBFDEBA5D2E95400140E001",
INIT_28 => X"FFFFFFFFFDFEFF7FFFFEAA5D2E95400E38A17438FFFFFFFFFFFFFFFFEFF7FBFF",
INIT_29 => X"1557DBEDF575D7FFFFFFFFFFFFBFDFEFEBF5F8E92552E9556DEBF1C21C7FFFFF",
INIT_2A => X"BF8FD7EBD16AA00000E3DF6DBEF5D2438FFFFFFFFFF7FBFDFC7EBF1E8A00080A",
INIT_2B => X"5155492FFFFFFFEFF7F1F8FD7A2D168A1008043FF6DAAFBC5028FFFFFFFFFF7F",
INIT_2C => X"000000000000000000000001FFFFFFFDFEFE3F1FAF55A2D568A0000003FF7D49",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFEBA552A95410002E820000000000000000000000",
INIT_2E => X"A552E954005D2A82145FFFFFFFFFFFFFFFFFFFFFBFDEAA5D2A954000800155FF",
INIT_2F => X"FFFFFBFDFEFF7FFFDEAA5D2E95410550415410FFFFFFFFFFFFFFDFEFF7FBFFEB",
INIT_30 => X"5EFAAD140155FFFFFFFFFF7FBFDFFFFFFBFDEBA5D2A95400A2AA974AAFFFFFFF",
INIT_31 => X"FF55A2D568A10082E955FFFFFFD7545FFFFFFFEFF7FBFFFFFAAD16AA00552A95",
INIT_32 => X"D74AAFFFBFDFEFF7FFEAB45A2D56AA00002EBDFFFF7D5400BAFFFFFDFEFF7FBF",
INIT_33 => X"568A0008003DFFF085555410F7FBFDFEFFFD568B45AAD16AA1008003DFEFAAFB",
INIT_34 => X"00000000000000000000000000000000000000001EFF7FBFDFEFAAD568B55AAD",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"01FFFFFFFFE00000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(20),        -- Port A data input
DOA(0)   => data_read_a_lo(20),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(20),        -- Port B data input
DOB(0)   => data_read_b_lo(20),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_21_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"4A302428B824900A128C090A5C1800261500213C005FE812D10420054085A202",
INIT_01 => X"081FFE3440B609703B0427F801A40B8115BC4F655300340288A40D30040E4DD8",
INIT_02 => X"0109095C30C98809800000F9FFFFFFFF149FF1FCA4C0421B182E3490DF145FE4",
INIT_03 => X"084A76341244919000099486400026523C041660BA000100CC12701015007FF8",
INIT_04 => X"000079800014CC03C075161E001118653D2408041FC004AEF000816E1C11F541",
INIT_05 => X"7E1F00F7FFC000240100004683103E7FFE02482553FC3C0204EFC25010143CC0",
INIT_06 => X"801008011010421960E339A20205FEBF8140000203FFC806C8A1C1048FF0F0E0",
INIT_07 => X"750504800680102542AD800504530FF9061E8026998E9A00402CC25BD0FFF800",
INIT_08 => X"11FBFFE04691A5A00101818A6800088228000001A044C8168480D010F200AA08",
INIT_09 => X"E85A7FF080AC70FFDF78220010841EFFE7116E144071268DFD3E4C2404010000",
INIT_0A => X"54518A8A31B7FE00040009814C089202225412115428C03BC7D7FC15025B1AB6",
INIT_0B => X"88300E20806520398C682157A493896600E24E10100DFF22FF86002020ED110C",
INIT_0C => X"28D9228D9228D9228D9228D9228D9228D99146C9146C84006309044081A001B1",
INIT_0D => X"890000403000A01282088624001201A8C43FF7C0011529904595123203040D92",
INIT_0E => X"06102C4053FFD5BFF00A04A00200602CA5200110008800444021048034004001",
INIT_0F => X"2A00263009140094D81A5040605800B506901A30406054013605620272181965",
INIT_10 => X"890A202811209062801A3040605800B506901A50406054013605604350B81282",
INIT_11 => X"3F4350B811068C00049A0A5820A3C1725A8006C0A40404D058320496C2C9C600",
INIT_12 => X"98361AC808127C454402483153A3A895BB3C1E2E820704020381702C1AAA2C4B",
INIT_13 => X"4D910CC1B154510413CC2A200501B400A40018A00C80400040D8AA288209AA21",
INIT_14 => X"0048A0141AA00418080460678A4012288463B2050302019200B00206C3590102",
INIT_15 => X"233142440470C8A9310280C0180302A01427D060022011606E800E00169C19A0",
INIT_16 => X"4010040100448008004000000E07008010003EFFFE0373056024B01118011988",
INIT_17 => X"0100401004010040100401004010040100401004010040100401004010040100",
INIT_18 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_19 => X"7E00000000000000000000000004010040100401004010040100401004010040",
INIT_1A => X"EFBEFBEFBEFBEFBEFFFFF7F7FFF3CF3CFFFFBE7FBBFDFFF7DFFCFBF08103DFDF",
INIT_1B => X"FFFFFFF7FBFDFEFF7FBFDFEFF7FBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFB",
INIT_1C => X"FFFFFFFE00003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"00080002000000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"FFFFFFFFFEBA5D2A954100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_1F => X"75FFFFFFFFFFFFFFFFFFFFFFFFFFEBA552A97400082A975FFFFFFFFFFFFFFFFF",
INIT_20 => X"FDEAA5D2E974100800155EFFFFFFFFFFFFFFFFFFFFFFFFFEAA552E95400082E9",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFDEAA5D2A95400080000000FFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"2E974105D2A80000FFFFFFFFFFFFFFFFFFFFFBFDEBA5D2E974005D2E80000FFF",
INIT_23 => X"FFFFFFFFF7FBFDEBA552A954005D2E97410FFFFFFFFFFFFFFFFFFFFFBFDEBA55",
INIT_24 => X"0000001FFFFFFFFFFFFFFFFFFFFF7FBFFEBA5D2A97400FF80174BAFFFFFFFFFF",
INIT_25 => X"FFFFFFFEBA5D2E97400000400000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2A95410000A001FFFFFFFFFFFFFFFFFFF",
INIT_27 => X"EAA552E954000020955EFFFFFFFFFFFFFFFFFFFFFFFFFEAA552E97400002E955",
INIT_28 => X"FFFFFFFFFFFFFFFFBFDEAA5D2A974101400155C7FFFFFFFFFFFFFFFFFFFFFFFD",
INIT_29 => X"97400552A80010FFFFFFFFFFFFFFFFFFF7FBFDEBA5D2E95400140E00000FFFFF",
INIT_2A => X"FFFFEFF7FBFFEBA552A95410552485038FFFFFFFFFFFFFFFFFFF7FBFDEBA552E",
INIT_2B => X"8A174AAFFFFFFFFFFFFFFFFEFF7FBFFEAA5D2E97400412497438FFFFFFFFFFFF",
INIT_2C => X"000000000000000000000001C7FFFFFFFFFFFFFFDFEFF7FFFFEAA5D2E95400E3",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974000004000000000000000000000000",
INIT_2E => X"A552E97400002E975FFFFFFFFFFFFFFFFFFFFFFFFFFEBA552A95410002E821FF",
INIT_2F => X"FFFFFFFFFFFFFFBFDEAA5D2A954000800155EFFFFFFFFFFFFFFFFFFFFFFFFDEA",
INIT_30 => X"4005D2A82010FFFFFFFFFFFFFFFFEFF7FBFDEBA552A974105D0015545FFFFFFF",
INIT_31 => X"DFEFF7FFFFEAA5D2A974005D2E82010FFFFFFFFFFFFFFDFEFF7FBFFEBA552E95",
INIT_32 => X"154AAFFFFFFFFFFFFBFDFEFF7FFFDEAA5D2E954105504154AAFFFFFFFFFFFFFF",
INIT_33 => X"BFDEBA5D2A95400A2AA974BAFFFFFFFFFF7FBFDFEFFFFFFDEBA552E974000004",
INIT_34 => X"0000000000000000000000000000000000000000155FFFFFFFFFF7FBFDFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(21),        -- Port A data input
DOA(0)   => data_read_a_lo(21),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(21),        -- Port B data input
DOB(0)   => data_read_b_lo(21),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_22_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"5290F4CDE914905A14A43D33F488243E17122300F55FEB189B343A1140548380",
INIT_01 => X"A94007B259F6A975386262000C344BA9573C6FF57B18A5FB0ABFCD3C2C5F4F0C",
INIT_02 => X"877FE30EB378008D202551040030071869D0040180AC4B685F6E26FAA0810006",
INIT_03 => X"431965109E4481D6B5AAD6875AD6AB5A1815600802888808DEA83552954D3000",
INIT_04 => X"492C0020220001010E4916C884DCD607E5EC2A344103E48003D0800023D0072C",
INIT_05 => X"0020F8882001102D620A06D683018001023D37E5088043620101179092540112",
INIT_06 => X"0803008022385AAA447A3306AA50001035B41C0A88046CAEE8C23C08E040011C",
INIT_07 => X"1EC04ED017AB5497EB923F08182E20020689B735011FBFE7BC06260294401CA8",
INIT_08 => X"4A00401D4425ADA9035BE19C8F9442A8801200F4C9D7AC8093A051727B2AC349",
INIT_09 => X"50020040E48D50080002B00A0C00801014541E9504703680017F6CB405070015",
INIT_0A => X"54538A8A738041C23020131A80CFDFF3FE509A907C6AC050402204090090319A",
INIT_0B => X"40050220103D2A512C6A8C4F0011550008E06E000140009A000000424DE61920",
INIT_0C => X"A81C2A81C2A81C2A81C2A81C2A81C2A81C9540E1540E001400006100003202D0",
INIT_0D => X"8B2940D0E153941A8B1A262CA542A9A8D6C0010A101628013456520CA09281C2",
INIT_0E => X"80410089180008800143D83888281A2034A85014280A14050A01509E05085449",
INIT_0F => X"000C26706B3C189CD84ACD20B03001E387D04AC560B02401E387E1028AC04500",
INIT_10 => X"458870201570B036C04AC560B03001E387D04ACD20B02401E387E24708E7E242",
INIT_11 => X"044708E7E1C20A0106EA167C84EBF052A8E010C0180606E86C3F459DC08DA902",
INIT_12 => X"98225189980254CDEC22A98032A22C50EAC462030A01800407C2700C2ACA2C0F",
INIT_13 => X"4A99BCC1154C258012D86F601A2E49003400138C0DA2443A208AA612C0096C37",
INIT_14 => X"90E16025483C1E0C0006B085CEC03858958D15310201015504B512044A313300",
INIT_15 => X"6B0469512C6FC01A1421006028038720640310643858162712020B001AA415F2",
INIT_16 => X"11044110445E22022365034A8EA754008004C0200323001182122548881649D1",
INIT_17 => X"1044110441104411044110441104411044110441104411044110441104411044",
INIT_18 => X"0401004010040100401004010040100401004010040100401004411044110441",
INIT_19 => X"7D05122890000000003FFFFFFFF9004010040100401004010040100401004010",
INIT_1A => X"E79E79E79E79E79EFFDFF7F5F777DF7DF7DF7EFF7BFA3FC7DF7AF5BF7EFDF7DF",
INIT_1B => X"9FCFE7F3F9FCFE7F3F9FCFE7F3F9E79E79E79E79E79E79E79E79E79E79E79E79",
INIT_1C => X"FFFFFFFE00000FE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F",
INIT_1D => X"10000000000000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"FFFFFFFFFEBA5D2E974000800021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_1F => X"21FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E954000004001FFFFFFFFFFFFFFFFF",
INIT_20 => X"FFEBA552A97400002A801FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2A9541008040",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFEBA552A97400082A975FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"2E95400082E975FFFFFFFFFFFFFFFFFFFFFFFFFFEAA552E95410002A955FFFFF",
INIT_23 => X"FFFFFFFFFFFFFFEAA552E95400002E975EFFFFFFFFFFFFFFFFFFFFFFFFFEAA55",
INIT_24 => X"000000000FFFFFFFFFFFFFFFFFFFFFFFDEAA5D2E97410080015545FFFFFFFFFF",
INIT_25 => X"FFFFFFFEBA5D2E97410080002000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974000004001FFFFFFFFFFFFFFFFFFF",
INIT_27 => X"EBA5D2A95410000A001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2A954000804021",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFEBA552A97400082E821FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"95410082A975EFFFFFFFFFFFFFFFFFFFFFFFFFEAA552E97400002E955FFFFFFF",
INIT_2A => X"FFFFFFFFFFFDEAA552E954000020955C7FFFFFFFFFFFFFFFFFFFFFFFFEAA552E",
INIT_2B => X"0015545FFFFFFFFFFFFFFFFFFFFFFFDEAA5D2A974001C24975C7FFFFFFFFFFFF",
INIT_2C => X"00000000000000000000000000FFFFFFFFFFFFFFFFFFFFFBFDEAA5D2A9741014",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800020000000000000000000000",
INIT_2E => X"A5D2A954000800021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974000004001FF",
INIT_2F => X"FFFFFFFFFFFFFFFFFEBA552A95410002E821FFFFFFFFFFFFFFFFFFFFFFFFFFEB",
INIT_30 => X"400002E975EFFFFFFFFFFFFFFFFFFFFFFFFFEAA552A97400082A801FFFFFFFFF",
INIT_31 => X"FFFFFFFBFDEAA5D2E95410082E955EFFFFFFFFFFFFFFFFFFFFFFFFDEAA552E97",
INIT_32 => X"17545FFFFFFFFFFFFFFFFFFFFFBFDEAA5D2A95400080015545FFFFFFFFFFFFFF",
INIT_33 => X"BFDEBA552A974105D0015555FFFFFFFFFFFFFFFFFFF7FBFDEBA5D2A974005504",
INIT_34 => X"0000000000000000000000000000000000000000010FFFFFFFFFFFFFFFFEFF7F",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"01FFFFFFFFE00000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(22),        -- Port A data input
DOA(0)   => data_read_a_lo(22),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(22),        -- Port B data input
DOB(0)   => data_read_b_lo(22),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_23_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"EF20906D902424807BC8241BC81801B97D38AD3C0800103362A6741C80A12A02",
INIT_01 => X"001FFF8409F089003B4422000D80C80106804A7951C5B9D1C828043EA28838F9",
INIT_02 => X"073B8858218C2C50801000F9FFEFF8E72CA7F5FC2E048026496834D84721DFE0",
INIT_03 => X"2C4360101A4001001005080400401420350016E0BB222341C312000014006FF8",
INIT_04 => X"00017B810015DC03D034201E14000036486008101FC0002EE006297E1C05F561",
INIT_05 => X"7E1F02FFFFC80100004044800080BEFFFC0248005FFC3C18A5FFC2444484BCC0",
INIT_06 => X"4082040800000811224DE0A00005FFBF8000000003FF810640A1C0008FF2F0E1",
INIT_07 => X"D1D72040048D00388387D03D0E591FFD201F862691DFBE077C2BC45B40FFE458",
INIT_08 => X"1FFBFFEC440501A5604B31062356282AA84200D12342113EDC40000004582800",
INIT_09 => X"A890FFF0002023FFDF79000000000EFFE309606020008005FC00000040200000",
INIT_0A => X"000000000037FF50010103134CAFDF03BA18000F39A0106F87D7FA84024B0225",
INIT_0B => X"88300C48907120AC81083315A493886640030010540DFF20FF8610302409000C",
INIT_0C => X"10C1010C1010C1010C1010C1010C1010C10086080860840063090442A18001B1",
INIT_0D => X"0000280600020040030090000012A500003FF7E08181119A41C1443243050C10",
INIT_0E => X"06542C7043FFD5FFF00A04BC010A7724B1000080004000200004150030010004",
INIT_0F => X"B2080290C2909080A872BC4FC8500054840072FC0FC8440054840200705F9861",
INIT_10 => X"0C8220180F1082E00072FC0FC8500054840072BC4FC84400548402214A380380",
INIT_11 => X"19214A380344920080B21810240AB182EB37C380B40800707011001B43253EE5",
INIT_12 => X"0019CE4000026C00C00042BD4149067465910640A0050C060A0028063672A000",
INIT_13 => X"4D801800CCB050001344060211629580B80022480A444111706658280009A203",
INIT_14 => X"944CB232D6D0100C040250200845132C10BE200403018061101A220339C80000",
INIT_15 => X"402102A5493B8E287E03808480060E40C83C1405132C90742E408D0082140820",
INIT_16 => X"0080200802000100100000000000004002403EFFF8002385F034901019465001",
INIT_17 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_18 => X"8020080200802008020080200802008020080200802008020080200802008020",
INIT_19 => X"0000000000000000000000000000080200802008020080200802008020080200",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000004000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFE00000000000000000000000000000000000000000000000000000000",
INIT_1D => X"10080400000000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"FFFFFFFFFEBA5D2E974100000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_1F => X"21FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100004021FFFFFFFFFFFFFFFFF",
INIT_20 => X"FFEBA5D2E954000800001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9740008000",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E954000004001FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"2A954100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2A954100000021FFFFF",
INIT_23 => X"FFFFFFFFFFFFFFEBA5D2A954100800021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_24 => X"0000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA552A97400002A801FFFFFFFFFFFF",
INIT_25 => X"FFFFFFFEBA5D2E97410080400000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800021FFFFFFFFFFFFFFFFFFF",
INIT_27 => X"EBA5D2E974000004001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100004021",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFEBA5D2E954000800001FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"954100004021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2A954000804021FFFFFFF",
INIT_2A => X"FFFFFFFFFFFFEBA5D2A95410000A001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2A",
INIT_2B => X"2E821FFFFFFFFFFFFFFFFFFFFFFFFFFEBA552A97410080E001FFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA552A9740008",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804000000000000000000000000",
INIT_2E => X"A5D2E974100000021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800021FF",
INIT_2F => X"FFFFFFFFFFFFFFFFFEBA5D2E974000004001FFFFFFFFFFFFFFFFFFFFFFFFFFEB",
INIT_30 => X"4000800021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E954000804021FFFFFFFFF",
INIT_31 => X"FFFFFFFFFFEBA552A954100004001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2A95",
INIT_32 => X"821FFFFFFFFFFFFFFFFFFFFFFFFFFEBA552A95410002E821FFFFFFFFFFFFFFFF",
INIT_33 => X"FFFEAA552A97400082A801EFFFFFFFFFFFFFFFFFFFFFFFFFEAA552A97410002A",
INIT_34 => X"00000000000000000000000000000000000000001EFFFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"01FFFFFFFFE00000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(23),        -- Port A data input
DOA(0)   => data_read_a_lo(23),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(23),        -- Port B data input
DOB(0)   => data_read_b_lo(23),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_24_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100600007FFF000080108004000800020000840041000080808",
INIT_02 => X"172A00D000EF8210000000F9FFEFF8E7240FF1FC224087B1000639401D005FC0",
INIT_03 => X"00003A2E200811000000000400000000340016603A0000004860400014006FFF",
INIT_04 => X"000079800014CC03C034001E04010850300000101FC0002EE000006E1C00F500",
INIT_05 => X"3E1F0067FFC000000000000000003E2FFC024800137C3C0000EFC00000003CC0",
INIT_06 => X"000000000000001123820AA00005FEBF8000000003FF80000021C0000FF0F0E0",
INIT_07 => X"E600084002040A10812A000500590FF9001F95406A8000037230C01840FFE000",
INIT_08 => X"01FBFFEC4695A501604A000C7585080002C200408102F16C0184800026C92C10",
INIT_09 => X"A8107FF0000000FFDF78000000000EFFE001600000000005FC00000000000000",
INIT_0A => X"000000000037FF4000000AA0354000019C4000012800002387D7F804024B0224",
INIT_0B => X"88300C0081408000800001002482886600020010100DFA20FF8600000000000C",
INIT_0C => X"00C1000C1000C1000C1000C1000C1000C1000608006084006301044081800121",
INIT_0D => X"00000000900160000000000000000000003FF7C0010101904181003003000C10",
INIT_0E => X"16100C4043FFD5BFF00004100000000411000000000000000000040030000000",
INIT_0F => X"3A0421080012302010049400086C022004200494000878022004120270599965",
INIT_10 => X"C19240300081406100049400086C022004200494000878022004124819081840",
INIT_11 => X"2348190814C09C01010400132100106836001504240E01040051200200D06410",
INIT_12 => X"202CD680C0100010408240BD80008983596CD86EA84104060503C0B000020250",
INIT_13 => X"0002090164F40086000082062C1B6600BC000C300818044000B27A0043000041",
INIT_14 => X"110002577FE4080C08010842180C40018545BBA00301808A0810C0059AD01802",
INIT_15 => X"4820C04100852B931F00800010081980B042D2044001850ED8808F00050A002C",
INIT_16 => X"0000000000000000000000000000000000003EFFF80037046031E0110001100A",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"9900000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"EFBE7BE7BE7BE7BEC99E61848655D75D7FCB42BBABDB9F3044CB35CF612B4441",
INIT_1B => X"83C1E0F0783C1E0F0783C1E0F07BEFBEFBEF9E79E79E79E79E7BEFBEFBEFBEFB",
INIT_1C => X"FFFFFFFE000001E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F07",
INIT_1D => X"10080402000000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"FFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_1F => X"01FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800021FFFFFFFFFFFFFFFFF",
INIT_20 => X"FFEBA5D2E974100000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741000000",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974100004021FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"2E974000800021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974000004001FFFFF",
INIT_23 => X"FFFFFFFFFFFFFFEBA5D2E974000800001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_24 => X"0000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E954000800001FFFFFFFFFFFF",
INIT_25 => X"FFFFFFFEBA5D2E97410080402000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFF",
INIT_27 => X"EBA5D2E974100800021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800021",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFEBA5D2E974100000001FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974000004001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100004021FFFFFFF",
INIT_2A => X"FFFFFFFFFFFFEBA5D2E974000004001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E",
INIT_2B => X"00001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E954000800021FFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9540008",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804020000000000000000000000",
INIT_2E => X"A5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FF",
INIT_2F => X"FFFFFFFFFFFFFFFFFEBA5D2E974100800021FFFFFFFFFFFFFFFFFFFFFFFFFFEB",
INIT_30 => X"4100000021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100000001FFFFFFFFF",
INIT_31 => X"FFFFFFFFFFEBA5D2E974000004021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E97",
INIT_32 => X"021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974000004001FFFFFFFFFFFFFFFF",
INIT_33 => X"FFFEBA5D2E954000804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E954000004",
INIT_34 => X"00000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(24),        -- Port A data input
DOA(0)   => data_read_a_lo(24),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(24),        -- Port B data input
DOB(0)   => data_read_b_lo(24),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_25_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100200002000000080100004000000020000800041000080808",
INIT_02 => X"1000218000000800000000F9FFEFF8E738FFF1FC20400400000004455A375FE0",
INIT_03 => X"00002000000001000000000400000000340016623A0000004000000014006FFF",
INIT_04 => X"924279824C94CC1BE0B4001F20000000020380401FE0082EF000106E1C00F500",
INIT_05 => X"3E1F0067FFE048002582800100523E2FFE024820137C3C0040EFE02000003CE4",
INIT_06 => X"821B0821B8019819200020200005FEBF81C1002203FF80000021C1140FF8F0E0",
INIT_07 => X"00040000000000000000000500590FF9001F0000000000033020C01840FFFC78",
INIT_08 => X"01FBFFFD0004000100502000011400000282004001020000000001009015C000",
INIT_09 => X"B8DA7FF8004000FFDF7C062031863EFFF75D78004001010DFC00002005010000",
INIT_0A => X"000000000037FFC00602000000000001980400002800032387D7FE94FBEF2B2C",
INIT_0B => X"88300C0080400000800001002486887600020110100DFA20FF8603000000000C",
INIT_0C => X"00C1000C1000C1000C1000C1000C1000C10006080060840077330C4889CC2925",
INIT_0D => X"00000000000000000000000000002500003FF7C0010101904189003003000C10",
INIT_0E => X"06140C6043FFD5BFF00A04B80608003CB120C110608830445821140134120800",
INIT_0F => X"02000000000200200000900000400200000000900000400200000200701E1861",
INIT_10 => X"0002000000010000000090000040020000000090000040020000000008080000",
INIT_11 => X"0000080800008000000000010100000022000000040000000040000000002400",
INIT_12 => X"0000420000000010000040318020000041000001000244000000008008000010",
INIT_13 => X"0002000004100000000080000002040040000000001000400002080000000040",
INIT_14 => X"0100000042000010002000001000400000042000040200000000400008400000",
INIT_15 => X"0030800000010800000000C0A000000000400000400000040800000000000004",
INIT_16 => X"41104451044C82082068C0200000008014023EFFFC0063046020801000001000",
INIT_17 => X"1104411044110441104411044110441104411044110441104411044110441104",
INIT_18 => X"1044110441104411044110441104411044110441104411044110441104411044",
INIT_19 => X"A080800002FFFFFFFFFFFFFFFFFC110441104411044110441104411044110441",
INIT_1A => X"41041249041249042824014C48569A69AFEE8A252865AA3168A4CBDF860EC15D",
INIT_1B => X"58AC56231188C46231188C462312492492492492492492492490410410410410",
INIT_1C => X"FFFFFFFE00002C562B158AC562B158AC562B158AC562B158AC562B158AC562B1",
INIT_1D => X"10080400000000000000000000000000000000000000000000000001FFFFFFFF",
INIT_1E => X"FFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_1F => X"01FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFF",
INIT_20 => X"FFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008040",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800021FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"2E974100000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800001FFFFF",
INIT_23 => X"FFFFFFFFFFFFFFEBA5D2E974100000021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_24 => X"0000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100000001FFFFFFFFFFFF",
INIT_25 => X"FFFFFFFEBA5D2E97410080400000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFF",
INIT_27 => X"EBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974100800001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800021FFFFFFF",
INIT_2A => X"FFFFFFFFFFFFEBA5D2E974100800021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E",
INIT_2B => X"00001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100000021FFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741000",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804000000000000000000000000",
INIT_2E => X"A5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FF",
INIT_2F => X"FFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEB",
INIT_30 => X"4100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFF",
INIT_31 => X"FFFFFFFFFFEBA5D2E974100800001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E97",
INIT_32 => X"021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800021FFFFFFFFFFFFFFFF",
INIT_33 => X"FFFEBA5D2E974100000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800",
INIT_34 => X"00000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"01FFFFFFFFE00000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(25),        -- Port A data input
DOA(0)   => data_read_a_lo(25),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(25),        -- Port B data input
DOB(0)   => data_read_b_lo(25),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_26_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"E9264EAB20190CA3BA4997AA9002AE9C001006B0778015CFA17E0811039879C7",
INIT_01 => X"F1FFF9BB1F773C7F9BB07DFFFDD863FC5FFF3FEFFBBF9FFB22FFFBC7B9F30686",
INIT_02 => X"1B33188302E708180F6FFBFFFFCFFFFF9C7FF7FC24350B99082400001D00DFD8",
INIT_03 => X"4A53D958C50000DCE7366303739CD98C27C57EF57980014F271807E3C9E9CFF8",
INIT_04 => X"DBFAFBD7FB1CDEBEF1BE17F7AC88042787FBFFF8FEE9FF7EE6F4C0EE1FFAF869",
INIT_05 => X"BE1FFD67DFFEFFBDA7F7FED508707E2EFEBF6FFEB37C3FF302EEEDFF9B487CF6",
INIT_06 => X"75F7275F7CAC98E261EDF0253C7FFFEF87C74E8CCFFBB6FF70E1FE61FFBDF0FE",
INIT_07 => X"73840C07783060C72DF7D828912E6FFB80162776F3BFB7077E82255E40BFEEBA",
INIT_08 => X"69FFBFE43C872321367036163F1C0820A3063F460D1AEFC000060042648C4181",
INIT_09 => X"FB967FBD13D981F7DF7D7E6171AF3FEFE8A3E679FAC1FD1FFFBEB000763A8447",
INIT_0A => X"6AED1D1DAD7FBE7D67D7F3BB79CFFB83BF14EC1E7D7300B017F5FFE6FBEF73BE",
INIT_0B => X"99F51EDDCDEBCFF589807B70AD9A99EE7583F931109FFE33FF8E3FDFDAF64A3C",
INIT_0C => X"C0D78C0D78C0D78C0D78C0D78C0D78C0D7A606BC606B8C56F7730ECCDBDF1521",
INIT_0D => X"1D406B9EC20181CC1F73F87501DED3409BFFFEFFEBF341B867D3683A03A40F78",
INIT_0E => X"86D70CE04FFFFF3FF1F5F5475BD7F72E4D75EBFAF5FD7AFEFDFFAF59B6FF28FE",
INIT_0F => X"020007C040101480807D17B0004001F804007D17B0004001F8040212F35FFC6D",
INIT_10 => X"700200001DC00068007D17B0004001F804007D17B0004001F804006F60081400",
INIT_11 => X"206F60081800800007B000102C0801FB02683800040007700011801003DE050A",
INIT_12 => X"403E232130207080D012CEFF41008D188D502100B02004000F01900039020040",
INIT_13 => X"0E101A01F21A2C40039006823F80048100003F0008004D8100F90D162001C803",
INIT_14 => X"B604027F020A07400007C040085581019D602451500001EC00100247C4642608",
INIT_15 => X"CC3F02010EA40EA00020C830100F0D000022180581019F40084800001F100020",
INIT_16 => X"EBFAFEFFBFEFDFDDFE7DD87FEFF7FF796FFFFFDFFC017FEFFD7E841001D8197D",
INIT_17 => X"BFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAF",
INIT_18 => X"FAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFE",
INIT_19 => X"EDB5C88646FFFFFFFFFFFFFFFFFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEB",
INIT_1A => X"61861A69A6986186EBCAF55357E1C71C751D6C56F3D247859B3214FA76953F86",
INIT_1B => X"84C26130984C26130984C2613098618618618618618618618618618618618618",
INIT_1C => X"FFFFFFFE0000026130984C26130984C26130984C26130984C26130984C261309",
INIT_1D => X"10080400000000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"FFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_1F => X"21FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFF",
INIT_20 => X"FFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008040",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFF",
INIT_23 => X"FFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_24 => X"0000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFF",
INIT_25 => X"FFFFFFFEBA5D2E97410080400000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFF",
INIT_27 => X"EBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFF",
INIT_2A => X"FFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E",
INIT_2B => X"04021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804000000000000000000000000",
INIT_2E => X"A5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FF",
INIT_2F => X"FFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEB",
INIT_30 => X"4100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFF",
INIT_31 => X"FFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E97",
INIT_32 => X"001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFF",
INIT_33 => X"FFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804",
INIT_34 => X"00000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(26),        -- Port A data input
DOA(0)   => data_read_a_lo(26),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(26),        -- Port B data input
DOB(0)   => data_read_b_lo(26),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_27_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"00080A40000A41248002029000050A088000008242A0004404480002000A1155",
INIT_01 => X"F1FFF1C11F781C129C107DFFFE0860941E81258CA2B71C2220EC1B86E1A00002",
INIT_02 => X"4000002100000014400FF6FFFF0FFFFF8007F1FC211100014200800000887FC0",
INIT_03 => X"0842D85841000098C63061026318C18404C459757000015F00088BE3C0618FF8",
INIT_04 => X"DBEAE5D6D91C2EBCE1B21EA72C00000007FBE7C8F8E9EF79E6D440E91FDAE061",
INIT_05 => X"B91FF9671FE6B68984B5BCE408347E28FEBF6FEEB3723F7102E8EDBF8A4872F6",
INIT_06 => X"3573A357308418E40000D4113C7FFE4F86064C8DDFE3B6FF50D1FC61DE39C8FC",
INIT_07 => X"00000A20083060C00C81882A008C6FF880060424B39FB6037F00051C003FE04A",
INIT_08 => X"61FA3FE4010440410844060001040A00002200460D1A06000005040000001080",
INIT_09 => X"EB027E390A4881C7BEFC5F6171CE2F8FE823E778DAC16C1FFBBC900031589547",
INIT_0A => X"03813030213C3E2D62D6E21259CFDB039E806C024531008017C1F826FFEF41FE",
INIT_0B => X"9AB55F0DEFABC705488069302DBA98EAB582D835109FFC31FFAEAFCFDAF4423D",
INIT_0C => X"40C3440C3440C3440C3440C3440C3440C3C2061A2061AD46FF730E5CCBCD5521",
INIT_0D => X"0C407D1F820101441DA3A8310198C34089BFF8DD6B7941BC63F1683803C00E34",
INIT_0E => X"5710AE4047FFD23FF315D54358D593474955AB6AD5B56ADAB5FAAE58B2F628EA",
INIT_0F => X"020007C0400004C080791290004001D80001791290004001D8000210F1587971",
INIT_10 => X"300200001DC0000801791290004001D80001791290004001D800012F60080400",
INIT_11 => X"202F60080800800007B000000E0801BB020828000400077000008210035E0408",
INIT_12 => X"40BA2220202070801010C6F1410085188D500100102004000F01900031000060",
INIT_13 => X"0E100205D2120840039000813F80040100003F0000000F8100E909042001C800",
INIT_14 => X"3E04007F020201400007C040001781011D602040500001EC0000005744440408",
INIT_15 => X"C43F02000EA40EA000004810100F0D000020080781011F40080800001F100000",
INIT_16 => X"AB6ADAB6BDE75ED5EC71385FC2512E3565BBBF1FFC00636EED7E841000D81924",
INIT_17 => X"B6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6AD",
INIT_18 => X"6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADA",
INIT_19 => X"A471688747FFFFFFFFFFFFFFFFFAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB",
INIT_1A => X"0020800000000000780401CBC840000005243885A04012072A1810DA84002104",
INIT_1B => X"5028140201008040201008040200000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFE000028140A05028140A05028140A05028140A05028140A05028140A0",
INIT_1D => X"10080400000000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"FFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_1F => X"01FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFF",
INIT_20 => X"FFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008040",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFF",
INIT_23 => X"FFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_24 => X"0000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFF",
INIT_25 => X"FFFFFFFEBA5D2E97410080400000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFF",
INIT_27 => X"EBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFF",
INIT_2A => X"FFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E",
INIT_2B => X"04021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804000000000000000000000000",
INIT_2E => X"A5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FF",
INIT_2F => X"FFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEB",
INIT_30 => X"4100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFF",
INIT_31 => X"FFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E97",
INIT_32 => X"021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFF",
INIT_33 => X"FFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804",
INIT_34 => X"00000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"01FFFFFFFFE00000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(27),        -- Port A data input
DOA(0)   => data_read_a_lo(27),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(27),        -- Port B data input
DOB(0)   => data_read_b_lo(27),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_28_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"02200AA400180030808802A900002A08001280A08A801044104A1000001818C3",
INIT_01 => X"50A00011460214428114180000882214413D0A71592A01D92213D28005210202",
INIT_02 => X"1444428102100884000AA30200000000C1000401041108404400022220800000",
INIT_03 => X"461080404900000C6314A900318C52A40051081000888806108802A141288001",
INIT_04 => X"00800040110102000902002000888400081045A8A00003C00000500000080008",
INIT_05 => X"0000000000024CA0A0101800032000400000000B800000014000000B08180000",
INIT_06 => X"10280102802C0240041000011428004022220024440013511000013510000000",
INIT_07 => X"0804420009122448451020100020400080002041000000008000010400000880",
INIT_08 => X"2800000140200808021006108010422AAA800022448902849220114009224081",
INIT_09 => X"01C800004080A0000002480B04008100011000088800081002C19020150B0013",
INIT_0A => X"56D29A9A52800004004070208000000040006408001100105000020000001800",
INIT_0B => X"00040024440245400082D0220800008010001020458000010000040D96104210",
INIT_0C => X"50160501605016050160501605016050160280B0280B00120008430660210014",
INIT_0D => X"054001884200810C1631181500CA60400B4008072020500002002C0040010360",
INIT_0E => X"104420A00C000200005000010040A0020CC000200010000800920040804020A6",
INIT_0F => X"0000000000001400000102900000002800000102900000002800001001802104",
INIT_10 => X"3000000000000048000102900000002800000102900000002800000020000400",
INIT_11 => X"0000200008000000000000002800000100082800000000000001800000020008",
INIT_12 => X"4000202020200000901005480000000800000100102000000000000009000000",
INIT_13 => X"0000120002020840000004800080000100000000000048800001010420000002",
INIT_14 => X"A200000800020140000000000050800008000040500000000000024004040408",
INIT_15 => X"840A000002000000000048100000000000020800800008000008000000000000",
INIT_16 => X"8020080210810840861CD33548542A10209D4100000010200400000000880035",
INIT_17 => X"0200802008020080200802008020080200802008020080200802008020080200",
INIT_18 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_19 => X"40A0C22E10000000000000000000020080200802008020080200802008020080",
INIT_1A => X"08208208208208200360D4141D630C30C7788440B044280091A5CB03D01BD89A",
INIT_1B => X"582C16030180C06030180C060302082082082082082082082082082082082082",
INIT_1C => X"FFFFFFFE00002C160B0582C160B0582C160B0582C160B0582C160B0582C160B0",
INIT_1D => X"10080400000000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"FFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_1F => X"01FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFF",
INIT_20 => X"FFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008040",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFF",
INIT_23 => X"FFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_24 => X"0000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFF",
INIT_25 => X"FFFFFFFEBA5D2E97410080400000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFF",
INIT_27 => X"EBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFF",
INIT_2A => X"FFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E",
INIT_2B => X"04001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804000000000000000000000000",
INIT_2E => X"A5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FF",
INIT_2F => X"FFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEB",
INIT_30 => X"4100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFF",
INIT_31 => X"FFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E97",
INIT_32 => X"001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFF",
INIT_33 => X"FFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804",
INIT_34 => X"00000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"01FFFFFFFFE00000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(28),        -- Port A data input
DOA(0)   => data_read_a_lo(28),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(28),        -- Port B data input
DOB(0)   => data_read_b_lo(28),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_29_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"79964E4BA01DACAB9E659792D00AAE160002829C7FDFEFCEE97C2815039D70C3",
INIT_01 => X"50BFF9AB0775343F9AB01DF80D5821FC0FFF3FEFD1AF9FF1207FFBC7B9720586",
INIT_02 => X"0B33180300E700080F6AAA7BFFC007189C7FF2FC003503980A0000001D00DFD8",
INIT_03 => X"0401D940CD0000C8421A2B03210868AC23403E903900010E271006A148A0C000",
INIT_04 => X"49B87A417315D20A313E17F1800000058013DDF8BE21F36E02F0D06E03E8F800",
INIT_05 => X"3E00FC67C03A4D9C87525E5101603E6E023D27DA937C03E340EE25CB9B483C12",
INIT_06 => X"50B5050B540C004261EDE025142DFFE003C30E0447F877F930203E213F8CF01E",
INIT_07 => X"73800407781020476467D008910A4FFB80100332D1AE93059282215E40800678",
INIT_08 => X"21FF80003C832320342036063F08000001063F42050AEB4000221000248C0180",
INIT_09 => X"51547F8C1111A0F041056A0100A11FE000916249A800B915FE82B02052290002",
INIT_0A => X"2AAD1515AD5780540541619968C76980E914E4163D53002017F405C409A42A9A",
INIT_0B => X"014002D445624DB481806A6288100184500171200085FE030000157FDF124A10",
INIT_0C => X"D0068D0068D0068D0068D0068D0068D006A68034680300021410028450530014",
INIT_0D => X"15402B0E8201018C1561E855008C50401B7FFE27A0B2500806522C0A40A50268",
INIT_0E => X"928324400DFFFF0001F1F0050342D42A086040B02058102C48970541944B20FA",
INIT_0F => X"0000000000101480000507B00000002804000507B000000028040212034FAD28",
INIT_10 => X"7000000000000068000507B00000002804000507B00000002804004020001400",
INIT_11 => X"0040200018000000000000102C0000410068380000000000001180000082010A",
INIT_12 => X"4004212130200000D0120ED64000080800002100B02000000000000009020040",
INIT_13 => X"00001A00220A2C4000000682008000810000000008004D800011051620000003",
INIT_14 => X"B6000208000A0740000000000855800088000451500000000010024084242608",
INIT_15 => X"8C0F0001020000000020C8300000000000021805800088000048000000000020",
INIT_16 => X"C0B02C4B12C989489418D13FE7F3FFD8BADB7FC004012CA5141600000198087D",
INIT_17 => X"0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02",
INIT_18 => X"B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C",
INIT_19 => X"FEA0C00602FFFFFFFFFFFFFFFFFC0B02C0B02C0B02C0B02C0B02C0B02C0B02C0",
INIT_1A => X"FBAEBAEBAEBAEBAEFFFFF7E7EFBFFFFFFAEF3E7E5BB9FFF7DFF9E3F08843FFDF",
INIT_1B => X"FDFEFF7FBFDFEFF7FBFDFEFF7FBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBE",
INIT_1C => X"FFFFFFFE00003EFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FB",
INIT_1D => X"10080400000000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"FFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_1F => X"01FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFF",
INIT_20 => X"FFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008040",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFF",
INIT_23 => X"FFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_24 => X"0000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFF",
INIT_25 => X"FFFFFFFEBA5D2E97410080400000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFF",
INIT_27 => X"EBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFF",
INIT_2A => X"FFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E",
INIT_2B => X"04001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804000000000000000000000000",
INIT_2E => X"A5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FF",
INIT_2F => X"FFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEB",
INIT_30 => X"4100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFF",
INIT_31 => X"FFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E97",
INIT_32 => X"001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFF",
INIT_33 => X"FFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804",
INIT_34 => X"00000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(29),        -- Port A data input
DOA(0)   => data_read_a_lo(29),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(29),        -- Port B data input
DOB(0)   => data_read_b_lo(29),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_30_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"FD00000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"E79E79E79E79E79EEBFEF5D7D7F7DF7DFFDFFEFFFBFE7F87DFFEFFBF77BFFFDF",
INIT_1B => X"9FCFE7F3F9FCFE7F3F9FCFE7F3F9E79E79E79E79E79E79E79E79E79E79E79E79",
INIT_1C => X"FFFFFFFE00000FE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F",
INIT_1D => X"10080400000000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"FFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_1F => X"01FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFF",
INIT_20 => X"FFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008040",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFF",
INIT_23 => X"FFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_24 => X"0000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFF",
INIT_25 => X"FFFFFFFEBA5D2E97410080400000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFF",
INIT_27 => X"EBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFF",
INIT_2A => X"FFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E",
INIT_2B => X"04001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804000000000000000000000000",
INIT_2E => X"A5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FF",
INIT_2F => X"FFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEB",
INIT_30 => X"4100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFF",
INIT_31 => X"FFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E97",
INIT_32 => X"001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFF",
INIT_33 => X"FFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804",
INIT_34 => X"00000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(30),        -- Port A data input
DOA(0)   => data_read_a_lo(30),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(30),        -- Port B data input
DOB(0)   => data_read_b_lo(30),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_31_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"129000008004A00804A40000400800020000000C005FEA005800200400050100",
INIT_01 => X"A15FF18019700810180065FFFC0040801E80258CA2951C2200EC0906A0804140",
INIT_02 => X"0000000000000011000550FDFF0FFFFF0007F1FC200000011000000000205FC0",
INIT_03 => X"08425818000000908428C0024210A30004045060302223490002014280410FF8",
INIT_04 => X"DB6A618248140C18E0B016872400000007EBA24058E1ECA8E2D400681FD0E061",
INIT_05 => X"381FF8671FE01009048084C400103E28FE3F6FE513703F7000E8E5B4825030F6",
INIT_06 => X"00130001300018A00000D0002855FE0F84040C088BE3E4AE40C1FD04CE38C0FC",
INIT_07 => X"000008800020408008818838000C2FF800060424B39FB6037E000418003FE008",
INIT_08 => X"41FA3FE400040001004000000104088000020044091204000004000000000000",
INIT_09 => X"E8027E38004801C79E7C162231862E8FE00166704041240DF93D000000000004",
INIT_0A => X"0000000000343E002202021259CFDB039E0008024520000047C1F804FBEF01BE",
INIT_0B => X"88310E08812982050800A9102492986200824810110DFC30FF86036249E4002C",
INIT_0C => X"00C1000C1000C1000C1000C1000C1000C18006080060840477330C4889CC0121",
INIT_0D => X"08006816800100400902A0200110810080BFF0C80111019861D1403803800C10",
INIT_0E => X"06100C4043FFD03FF101D4000800130401808100408020401020041830120848",
INIT_0F => X"020007C04000008080781000004001D00000781000004001D0000200F0185861",
INIT_10 => X"000200001DC0000000781000004001D00000781000004001D000002F40080000",
INIT_11 => X"202F40080000800007B00000040801BA020000000400077000000010035C0400",
INIT_12 => X"003A0200000070800000C231410085108D500000000004000F01900030000040",
INIT_13 => X"0E100001D0100000039000003F00040000003F000000050100E808000001C800",
INIT_14 => X"14040077020000000007C0400005010115602000000001EC0000000740400000",
INIT_15 => X"403502000CA40EA000000000100F0D000020000501011740080000001F100000",
INIT_16 => X"01004010044602002061004A820104809402BE1FFC006304E036841000501900",
INIT_17 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_18 => X"0040100401004010040100401004010040100401004010040100401004010040",
INIT_19 => X"0001000802FFFFFFFFFFFFFFFFF8100401004010040100401004010040100401",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFE00000000000000000000000000000000000000000000000000000000",
INIT_1D => X"10080400000000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"FFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_1F => X"01FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFF",
INIT_20 => X"FFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008040",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFF",
INIT_23 => X"FFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_24 => X"0000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFF",
INIT_25 => X"FFFFFFFEBA5D2E97410080400000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFF",
INIT_27 => X"EBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFF",
INIT_2A => X"FFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E",
INIT_2B => X"04001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804000000000000000000000000",
INIT_2E => X"A5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FF",
INIT_2F => X"FFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEB",
INIT_30 => X"4100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFF",
INIT_31 => X"FFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E97",
INIT_32 => X"001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFF",
INIT_33 => X"FFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804",
INIT_34 => X"00000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(31),        -- Port A data input
DOA(0)   => data_read_a_lo(31),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(31),        -- Port B data input
DOB(0)   => data_read_b_lo(31),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_0_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"ED39BA795990D275FB4A6E96ACC4731DEA4598B0AFB54867F6EE4618C3749807",
INIT_01 => X"58A0047D8607944AC7DA180001ECA2544042106208408208C20022E9173734B3",
INIT_02 => X"9F775E7CB273E6CCA7DAAF00001000000478020113C9C38E09FB7CCCDD9F203E",
INIT_03 => X"441406267B4CB04443163C91110C58F24A31000B8028A810A3D0F8B169A01006",
INIT_04 => X"0005802424830120024121209088809DF81454ACA01E03501D0A3B91E00F0A00",
INIT_05 => X"C1E0039800112014C20B0232838F80D001C0100AEC83C008EF101A034C8CC300",
INIT_06 => X"8B0478B04A83405954592F9B9628000002C3F08754001B51881E007900060F01",
INIT_07 => X"39F36677EE1C387777622717EF711004A6818111086008E080FDC30594001017",
INIT_08 => X"160400195E83A3A0F61BC3929ECB622AABF5FF83860CEB164833F179B48CEE59",
INIT_09 => X"036D8004FDB47600000229410C61010016DC998C84B0128202C0DCB48F05D513",
INIT_0A => X"204122A033000182502440888420247041E876810099D35F900002DB00105C01",
INIT_0B => X"41C000947E16656074EA560F080544900960260144D201890018080D36191110",
INIT_0C => X"781EA781E2781EA781E2781EA781E2781C33C0613C0E00120800239450112ED4",
INIT_0D => X"872917095352BD2A90515A1CA44E7EA84B00001010043803120C3E04E03383E2",
INIT_0E => X"70C7E0B92800224008AE09B8942C48D1FC491204890244812250588601285432",
INIT_0F => X"B80C2038ABACB83C7E03EA5FF83C002783F103EA5FF83C002783F0120847A704",
INIT_10 => X"BD9870380230F2D7C103EACFF83C002783F103EACFF83C002783F310BBF7EFC2",
INIT_11 => X"1F10BBF7EFC61E01804E1E6EA1E3FA01FD97EFC4B80E008C7C2F678FF023FAF5",
INIT_12 => X"B801FCC8E8320C4DAC9220C6B2FF22EF72ADDE6F1A67C80600C2683E0EF8AE1F",
INIT_13 => X"4189B5C00FE651C6104C6D6400FFFB01FC0000FC07EE42FA7C07F22CE3082636",
INIT_14 => X"8BE9FC08FDF4195C0C2038A7C6CAFA7E289F9BA4570380131CAFB2003F9D190A",
INIT_15 => X"270AE9FE635BE11B7F0308D4A80092E0FC1FC662FA7E283FF68A8F0080AE1DDA",
INIT_16 => X"1204812058112C12411402056954AB0C280D000003350013024179498C2EC6B9",
INIT_17 => X"2048120481204812048120481204812048120481204812048120481204812048",
INIT_18 => X"0481204812048120481204812048120481204812048120481204812048120481",
INIT_19 => X"13043A85D4000000000000000001204812048120481204812048120481204812",
INIT_1A => X"82082082082082082218821390771C71C557CE263826D5B1D36AC59E0765D1CF",
INIT_1B => X"1F0F87C3E1F0F87C3E1F0F87C3E0820820820820820820820820820820820820",
INIT_1C => X"FFFFFFFE00000F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E",
INIT_1D => X"EF5D7BD7400000000000000000000000000000000000000000000061F007FFFF",
INIT_1E => X"A10A2D1574005D0428A10A2AAA8BEF552EBDFFF557BC01FF5D7BFFEBA5D55555",
INIT_1F => X"DEBAFFFFC2000AA8428AAAFFAAA8BFF00002AA10FF802ABEFA2D16AA00F7FBE8",
INIT_20 => X"975EFFF8002010002EAAAAAAAD1555FFFFAEA8B550051401450055575FF00517",
INIT_21 => X"4155FF0855575455D2AA8BFFA2D1575EF5D5555545FFFBE8A00087FC20BA5D2A",
INIT_22 => X"8028A00FFAE800AA082A820005D2E974BAA2D140145A2842AA00A284021FF5D0",
INIT_23 => X"2D17FFEF000017400FFD1555FF007FFFEBA55042AA00000017400FFAABFEBAFF",
INIT_24 => X"000000155F7D540000F7FBFFE105D7BE8ABAA284000105D0428BFFA2FBFDFFFA",
INIT_25 => X"75D7BFAEBA5551501D51C5FC7E00000000000000000000000000000000000000",
INIT_26 => X"28B6D16AA28EBF5EDA38AADE1543849557D492BF8E2DE00552EBFFC7552BC01D",
INIT_27 => X"000A85400E00E38A175FDE3F5C002DAAD42DAAAF784AFA82BC042DF47E3D1F80",
INIT_28 => X"AA150021C0092490E904BAFFD550A90FFA495FC7A05B555C257AAA8B45007540",
INIT_29 => X"2DA02402ABD4AD1D0E175D7140B455D516A1EAB45E2A000B4748717A095F571E",
INIT_2A => X"4004A8BC0ABFF7D03A17D1D5147540B454AA080038E9748542AE3D0051C7B6F0",
INIT_2B => X"FB6D4B8FC7BFFFD2168B68F57492F505FF5FA550490BFA482B420B8428A3DA85",
INIT_2C => X"0000000000000000000000016ABD554201543A1EDE9016D4AAB454AF400547AB",
INIT_2D => X"5D2EBDF55556BC35E7557FE8AB25D11415FD0151614000000000000000000000",
INIT_2E => X"9596CBEA41D7D3DECFAF7D43FABAAAD57DEBAAAFFD74AA04547EE18D680BE9A5",
INIT_2F => X"47D78228E5000EA422E10439C1FBCD282351BDAAF9C20AAAABCBEB1DFF803FC5",
INIT_30 => X"1E6284683ABBDD7DEAA100069C14B25495A00F38EBAC0E198B97605018053575",
INIT_31 => X"4408FE6A755ED8EFEFE41B2D17EAF02552BC0545556BD61E501001DF5DD3EBA3",
INIT_32 => X"556F922ACA8AB8283C8310FAB1588916D3861C0422C44082B52A81550A828141",
INIT_33 => X"A5FDBCD7D262E5AFAC4B6AADDD562AF57D7C369AF25495A23068A8301BA7FB95",
INIT_34 => X"003FE0000003FE0000003FE0000003FE0000003FE03D5789700282E9FEFB501E",
INIT_35 => X"0003FE0000003FE0000003FE0000003FE0000003FE0000003FE0000003FE0000",
INIT_36 => X"00000000000000000000000000000000000000000000000000000000003FE000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(0),        -- Port A data input
DOA(0)   => data_read_a_hi(0),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(0),        -- Port B data input
DOB(0)   => data_read_b_hi(0),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_1_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"212C001411984004084D000508C53810A03D1450E839B003342114428A000807",
INIT_01 => X"08000010400A0008010600000084004000400002000000000000000000140000",
INIT_02 => X"484DEBA0111800C004400D000000000028800001CC404E6008B4933336880010",
INIT_03 => X"650C00000848A0423183089008C604224200000100A200002C280810098C0001",
INIT_04 => X"00000004208B00200E010800006667BE7000102C00080000040012010000080C",
INIT_05 => X"0100000000002000600100208D04414000800000000200004800080000800200",
INIT_06 => X"010420104032C204071200000200000010104020000001000910000000040800",
INIT_07 => X"8C0060242183060CF118011281B00000220010400020002081A0008210000802",
INIT_08 => X"000400014812466427040098C000622AAAA43E3060C158AC97F0356BDBFBD008",
INIT_09 => X"026C000559102400200281400469000008B0800000901080004004308B434040",
INIT_0A => X"50502A2800800000400408200000201041000208000040020820034200005C00",
INIT_0B => X"13C051112A800008402002021128000081202205001000000028880004010500",
INIT_0C => X"191AC191A4191A4191AC191AC191A4191A00C8560C8D2940804060901210441E",
INIT_0D => X"C1C114417882F82C00181707044212080300001002081224002006406401918C",
INIT_0E => X"60C0C0B92C000000000400001004200044010200810040802040080200284401",
INIT_0F => X"380C200000043C2016000000F03C00280030000000F03C00280030000004860C",
INIT_10 => X"8D18703800000049C0000000F03C00280030000000F03C002800321080000BC2",
INIT_11 => X"0110800007861E0180000002A9001A00000007C4380E00000001E00230000000",
INIT_12 => X"688004C0C81200009480010280340000008082430A07C80600C0000009008610",
INIT_13 => X"4000134400241186100004A500007B00FC000000000E4A402C001208C3080002",
INIT_14 => X"A9002C0001E0181C0C200000025A400A200812A4070380000000B25000981902",
INIT_15 => X"0000804A0002410A170300C4A800800000020E22400A200096828F008000000A",
INIT_16 => X"020080200820040041002000010080000000000002340002004118010C228614",
INIT_17 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_18 => X"0080200802008020080200802008020080200802008020080200802008020080",
INIT_19 => X"2B5000A000000000000000000000200802008020080200802008020080200802",
INIT_1A => X"AA8A28A28A28A28AB2048634B03249249604CA291AEAFBF1528205C00020C745",
INIT_1B => X"974BA5D6EB75BADD6EB75BADD6EAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA",
INIT_1C => X"FFFFFFFF00000BA5D2E974BA5D2E974BA5D2E974BA5D2E974BA5D2E974BA5D2E",
INIT_1D => X"55AAAAAAA00000000000000000000000000000000000000000000181FFFFFFFF",
INIT_1E => X"BEF5D7BE8ABA5D557DFEFFFD17FEBA00042AAAAFFFFFFE00FF843DF45FFAE955",
INIT_1F => X"DFEF552A800AA5555575FFA2AE820BAFFAEBFF555500155EF552E975FFF7D168",
INIT_20 => X"6AA00A2FBEAABA5D55420AA00002AA00AAFBE8B55A280175455D002AA00A2AAB",
INIT_21 => X"BD75FFAA802AAAAFFAA801EF00517FFFFF7D56ABEF0004155550004154105D55",
INIT_22 => X"55575FF08557DEBAA2FBEAAAA552E955EF5D0415410A2AE97545A2AE954BAF7F",
INIT_23 => X"7D17DF55A2AEBDEAAFFFFC20AAFFFFFFFFFAAD5555FFFFAEAAB55A2D168B555D",
INIT_24 => X"0000000BAFFFBE8A00087FC20BA5D2A975EF5D0002010552E820AAFFD57FF55F",
INIT_25 => X"8FF8A38F45F7AA9217FA380AD400000000000000000000000000000000000000",
INIT_26 => X"D7552E975EFFFDF68BFF557BEAA925551785D7BFD5EFE3F08002FA92EBA5FDE2",
INIT_27 => X"43841017DE92BF8E3AA824924870BF5551555C7A28A821EFE3AABAE38005B575",
INIT_28 => X"0568005A1041055716DB7DB6FBEFEA81C55D0A0516802AA28BEF5EDB7DAA8A15",
INIT_29 => X"C7FEF1C043FE28E3FBD55FFAADE2DAAAE3A5C51C71C042DF45A3D1D00281E8A1",
INIT_2A => X"AA8B45B47F6FB55A95555E90F78E17F52FEF5EDA82FD249057F080417492AAAF",
INIT_2B => X"5FF8AAAA95B7AF45FF8F7DFEDFFAFF8E005FAE92A3AE3DBFF57FA2DF555D257A",
INIT_2C => X"000000000000000000000000A8F571EAA150021C0092490E905FFFD0550BD75C",
INIT_2D => X"00043DE00A2C57DE08FFAAA8B55F7EE801F7F2849EE000000000000000000000",
INIT_2E => X"6AAAE29F067155543A15D2E955EFFFFBEABEF557FEAA10595169BED83D1EBCA8",
INIT_2F => X"BAFFD57DEEAAA15976EB0444BFEB086808A8E3082C954BA5D7DD6145AAAA821A",
INIT_30 => X"B47FFD55D6107782001FF0812000A255D57FFBEF3B97EEAB2C40217B9778428A",
INIT_31 => X"35FF003F17418AEE817B540D11CA80BAAFA825EFAABEBCA18FE803755D08079E",
INIT_32 => X"8BDEBA2D757547D7862AF57ABFFCABE5553FD5FBEFE86353EFFFD03FE0275000",
INIT_33 => X"5A01F70C6AA04537957D6FB4807FFFB45F7EFFDA58FF2AA88A0F3C5014018AC2",
INIT_34 => X"00000000000000000000000000000000000000000B2DD7DEAA100069C14B2549",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(1),        -- Port A data input
DOA(0)   => data_read_a_hi(1),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(1),        -- Port B data input
DOB(0)   => data_read_b_hi(1),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_2_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10E006600180111284380310006289800480032283E000A34301002001A0816",
INIT_01 => X"0005A00810790848048044A54E404340404000720885800802000806EC910200",
INIT_02 => X"5C010802020408040C400850AA055254090541A111200A104A0000000908B510",
INIT_03 => X"0C1101100C00004401060A0010041028021560A0218808002440840008880550",
INIT_04 => X"8840C2802205140048281202180804040960986850688C99444090C10A124A69",
INIT_05 => X"910A21220A880010214000010340086856B141252252142242A068B090106372",
INIT_06 => X"4007A400E8A40086213090040001520500204088012121026050A54CE2154840",
INIT_07 => X"0204022420000004601120108108055200022025A83AA3008882004A001542CA",
INIT_08 => X"091C154429220A2824642010A010020282843E00000248000021100000884101",
INIT_09 => X"80442C1411D120828A2A116A24632885419244606001110AE11B202046439511",
INIT_0A => X"644022201204145003031012D40D718241108815384200904160AE42CE2818E2",
INIT_0B => X"1BF047118108829501009202A5A20068C003211551163A00E522B3000562082D",
INIT_0C => X"90D0490D2C90D0C90D2C90D0C90D2490D04486124868294032384890B8985534",
INIT_0D => X"184014960000008402028041005232001715A040820B11A401E2443243450D04",
INIT_0E => X"9306260000554015520481040100004504A08110000820440001009134000004",
INIT_0F => X"02000000001014000028052000400028040050052000400028040200501C8D38",
INIT_10 => X"4002000000000068005005200040002804002805200040002804000E00001000",
INIT_11 => X"0028400010008000000000102800009800601000040000000011820002140102",
INIT_12 => X"4022010110000000D00008310000801080102000A00004000000000009020000",
INIT_13 => X"00001A00C0082400000006802500008000000000080048000060041200000003",
INIT_14 => X"A000005400080600000000000850000014200411000000000010024440202200",
INIT_15 => X"0000000008840600002080200000000000021800000013000040000000000020",
INIT_16 => X"40902449022A800800002208090684819402120AA8001C800000000000100014",
INIT_17 => X"1902409024090240906419064190641902409024090240906419064190641902",
INIT_18 => X"9044190440900409004090041904419044190440900409004090641906419064",
INIT_19 => X"7D402A2953F81F81F83F03F03F04190441904419044090040900409004190441",
INIT_1A => X"4104104104104104609D21808205965965D65801004E35C300C2D50A22B1C50C",
INIT_1B => X"128944A25128944A25128944A250410410410410410410410410410410410410",
INIT_1C => X"FFFFFFFFE3F00944A25128944A25128944A25128944A25128944A25128944A25",
INIT_1D => X"100055400000000000000000000000000000000000000000000001E1F007FFFF",
INIT_1E => X"400FF843DF45FFAEBDF55082A82155082AAAA10F7FFEAB455500175FF5D2A800",
INIT_1F => X"ABEF082ABDF455D7BD5545F7D5574BAFFD16AAAAA28428ABA000428AAA5D7FD7",
INIT_20 => X"EAB455D7BEAABA5D2A97545552E975FFFFD168AAA5D7BE8BFF5D557FFEFFFD16",
INIT_21 => X"A955555555555FFA2AE820BAFFFFEAABA5555554BA5D0417545F7D56AAAAAAFB",
INIT_22 => X"002AA00AAAEBDFFF08042AABA087BD54BA08043DEAAFF843FF5508517FF55552",
INIT_23 => X"02A82010AAD1401FF002EBFF45A2FBFDFEF00042AA00AAFBEAB5500003FF5500",
INIT_24 => X"0000000BA0004155550004154105D556AA00A2FBEAABA085542145082A800BA0",
INIT_25 => X"D5500155FF552A87410007145400000000000000000000000000000000000000",
INIT_26 => X"9208002FABA4171D5400FF8A38F45F7AABA57D0000855FD1C2AAFA00EBA5E8B7",
INIT_27 => X"A92555178FD7BFD5FDFFA0020BFF78417BD5545F7F1554AAF7D16DABABFF57DE",
INIT_28 => X"756DFFDF6DAAAAAF1EFB6D417BEFA901C2E97F40552E975EFEBDF68ABA557BEA",
INIT_29 => X"2DB7DA3FBD21C7492E9256D555B555C7A2ABC20AAE3AABAE38005B574AA49041",
INIT_2A => X"5EDB7D1E803AF6D400028E02AB8A3A012540E2AABABC75D043A00003FE10E380",
INIT_2B => X"0EB8B7D0AAA800AA147085000FFDA001C7B47BFABC7BFFF7AB4714042AA38BEF",
INIT_2C => X"000000000000000000000000821E8A10568005A1041055716DA38B6FBEFFEF1C",
INIT_2D => X"5D2EBDE00AAC16ABEF5500155EF552A954000855544000000000000000000000",
INIT_2E => X"AF7D57DE0AFAD1EBEB400043DEAA085555400FFAAAAB55F7AEA8BF77004147EF",
INIT_2F => X"EFAAFBEABAF557FEA8515951E8B4D83D1EBDFF082CBDFEF005756145FFD5574A",
INIT_30 => X"E005951550100004155EFF7FFFDE08AA557FFFF083FFCEB95104210405D2E955",
INIT_31 => X"00AA002A3FE18AE803CBE7A3C014351082E951FF5D7FD6145AAAA820A2AAAD29",
INIT_32 => X"EAD45550028ABAFFD17FFED01001FFEF5542ABEB2AA848AAA2552EA8ABA75514",
INIT_33 => X"57FEBAF3F95EEE95C00B7CF12AAA800BA551417105FFFFC21555556EAB4CD6D5",
INIT_34 => X"00000000000000000000000000000000000000000187782001FF0812000A255D",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0400000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(2),        -- Port A data input
DOA(0)   => data_read_a_hi(2),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(2),        -- Port B data input
DOB(0)   => data_read_b_hi(2),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_3_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"210C00A20020000108430020001600B8156021104940741B3530400E02B92202",
INIT_01 => X"A00C9BC058B00968240402C992000B61404040028804A0080A000D16A8990A08",
INIT_02 => X"4809A902031800444445089866E331352180D468B8200E600C0081110B80ACD0",
INIT_03 => X"6D0A601008000142B1A30A040AC68428320006010A80881068A80D401C846330",
INIT_04 => X"482218076809C03B24841CD92CDD5A4402091278072948042640102107102D04",
INIT_05 => X"0B063006A6402109000104E40B04644B32A86D20014A0D204063296082000E34",
INIT_06 => X"01072010703402800606D0102800CAB31434442810B4858060D0500008C52828",
INIT_07 => X"8C00222420A14204E01C581091020CC8000E3226413990008D80001A00CCC4AA",
INIT_08 => X"0874732009120665255420184000220002843E14294258E805E0116002D95101",
INIT_09 => X"BA546AC411102029A61C974014EDBA1320B1046100C0B4034928002002211145",
INIT_0A => X"1052088250A1CC2041051913208CE802438000082040008000F399406BC07998",
INIT_0B => X"19E416590908884D00020242A500090801806801041358222302084204460020",
INIT_0C => X"1019010190101B0101B01019010198101B20805C080C880080506990125E0514",
INIT_0D => X"03400040A101C05C0088242D0000320013339310018011A044414400400101B0",
INIT_0E => X"6514CA601CCCC8B33204C0401104244000018380818040A07060090000280009",
INIT_0F => X"0000000000020000006000000000020000011000000000020000010072CC9251",
INIT_10 => X"0000000000010000014000000000020000013800000000020000010700000000",
INIT_11 => X"002C000000000000000000010000001A00000000000000000040000002440000",
INIT_12 => X"00B2000000000010002049910000011000500000000000000000008000000000",
INIT_13 => X"00020005500000000000800133000000000000000010000000C0000000000040",
INIT_14 => X"0000005300000000000000001000000110600000000000000000401540000000",
INIT_15 => X"8000000008200620000000000000000000400000000107000000000000000004",
INIT_16 => X"0280C0280C0205104100000A8D06C404440230B9980210020040000010010003",
INIT_17 => X"280C0280C0280C0280803808038080380803808038080380C0280C0280C0280C",
INIT_18 => X"80E0200C0280E0200C0280E030080380A030080380A030080380C0280C0280C0",
INIT_19 => X"291008A004D54AAB556AA9556AA830080380A030080380A030080380A0200C02",
INIT_1A => X"4904104104104104A20E85800004924924054C0F031E31C190A285040164C586",
INIT_1B => X"1A8D46A753A9D4EA753A9D4EA752492492492492492492492492492492492492",
INIT_1C => X"FFFFFFFEB6FECD46A351A8D46A351A8D46A351A8D46A351A8D46A351A8D46A35",
INIT_1D => X"00AA8400000000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"B455500175FF5D2AA8A10005540155087BEABFF552ABDF45A2D16AAAAF7D5400",
INIT_1F => X"201000556AB55552ABDE00AAD140010F7D17FF45A2AA82155082AAAA10F7FFEA",
INIT_20 => X"42155557FEAA10007FEAABA000428AAA557FD7400FF843DE00FFAEBFF55082A8",
INIT_21 => X"AA8A105D7BD5545F7D5574BAFF802AA00A2D168ABA085568BEFFFAE820000855",
INIT_22 => X"557FFEFF7D56ABEF557BD74BAFF8402145A2AEBFFEF552EAAABA5D0028BEF082",
INIT_23 => X"5043DEAAAAAA95410F7803FFFF55556AAAA552A975FFFFD16AAAA5D7BC01EF5D",
INIT_24 => X"0000000105D0417545F7D56AAAAAAFBEAB455D7BEAABA5D2A974005D55574005",
INIT_25 => X"5B6DF6FABAFFD547010AA8407400000000000000000000000000000000000000",
INIT_26 => X"6D1C2AAFA28EBF5E8B7D5500155FF552AAF0100071455451C75EABC74174BAF5",
INIT_27 => X"F45F7AABAF7D00009543D1C556AB6D4124BAE10BED542010FFD57AF55AAF5D75",
INIT_28 => X"ABFFEBA0870281C5F4716D5D7FEDA3A0955FF48208002FABA4171D5400FF8A38",
INIT_29 => X"B8EBA15203FFFF002AAFA384171D5545F7D0154AAF7D16DABABFF57DE92005F6",
INIT_2A => X"F68ABA417BC01D7555178FD7BFD5FDF571575D24BA438E021D5B6A4BAFFF5D2E",
INIT_2B => X"24BFE005D5B52428410E3AE92E3A490410EB843ABD71551FFE02552A975FFEBD",
INIT_2C => X"0000000000000000000000003849041756DFFDF6DAAAAAF1EFB6D417BEFBD71C",
INIT_2D => X"5D556AB45081028B55FFFFFFEBAFFD557400A280144000000000000000000000",
INIT_2E => X"0FFD56ABF5AAD15455F5D2EBDEAAA2D16ABEF5500175EF552ABDE00085554545",
INIT_2F => X"AA085555400FFAAAAB14F7AE28BF77004146BA557DEABEF00002BE10FFD54000",
INIT_30 => X"E0AF2D1EAEBA007FEABEFAA84174BA557FD55EF5D3BFEEB35055DEE1000043DE",
INIT_31 => X"0155FFAA28BF7592EABE0A0804ABFFB082EBDEAA005556145FFD5574AAF7D47D",
INIT_32 => X"EB8105D2E955EFAAFBE8AAA547FE21550853E8B4FABD5EBFF75D55420AA82AA8",
INIT_33 => X"57FFFF087FFCEF90104B780A557FC20AA082AAAE10AA8000000A2AC2ABFD2151",
INIT_34 => X"00000000000000000000000000000000000000000AA0004155EFF7FFFDE08AA5",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(3),        -- Port A data input
DOA(0)   => data_read_a_hi(3),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(3),        -- Port B data input
DOB(0)   => data_read_b_hi(3),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_4_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10804002061080A284201081034809800A002303500078B3432C82904204002",
INIT_01 => X"810398000008004C0420050E12100368403008418984014902030806A0910204",
INIT_02 => X"480108A000000000446448E01E80F00A41043118680402000800000009882390",
INIT_03 => X"065040108C0000408406080002101020260012E03000000030808902088000F0",
INIT_04 => X"9100EB8368155C1AE0B01CD60433B944028A90385AC0D438E02010E81C32E801",
INIT_05 => X"B81E4166DE080029204044C401041C4CF01C489433483C8042EAC190100074C4",
INIT_06 => X"400F0400688002A22010D4342045C50F0004028993B3A5260041E4500EB4C0E2",
INIT_07 => X"000000243020008461000812810003C300060064012E00048C82005800BC2888",
INIT_08 => X"08CC8F0109064220240410008000002202043E44001048000020114000881000",
INIT_09 => X"F0DC1EB5131020C7BE7D172251E53E80E891E5016041B4083945202002419104",
INIT_0A => X"7D6025AC2A0982500302003200872003FB108808280200204400786612CE2B08",
INIT_0B => X"11D0025980480A458100930201820964408268101000F022D8083B4044A0002C",
INIT_0C => X"90C3490C1490C3490C1490C1490C3490C104869A48618800B66305989ABA0434",
INIT_0D => X"220000000500021002100088004010001370F030808110204581043243050C54",
INIT_0E => X"06100C40903C1C30F20025440102200541204090600830045825050034010000",
INIT_0F => X"000000000012000000BC04000000020004018C040000000200040000721CD861",
INIT_10 => X"000000000001002001A40400000002000401DC04000000020004014D44001000",
INIT_11 => X"0065040010000000000000110000007600200000000000000050000005D40002",
INIT_12 => X"00DE00001000001040004A3B0000180088500000200000000000008000020000",
INIT_13 => X"0002080760000400000082024300008000000000081006000170000200000041",
INIT_14 => X"180002B200000200000000001806000192000010000000000010401F80000200",
INIT_15 => X"0814000114A00200000000200000000000401006000085C00040000000000024",
INIT_16 => X"40102459044481081044880A0986D4C1560636C7840A61803000820012113042",
INIT_17 => X"1900411064090041102409044110240900401064190040106409004110640904",
INIT_18 => X"9064090240100411044090241902401044110041902409064110241904401024",
INIT_19 => X"04048028064B261934D964C3269C090641100401044090641902401044010041",
INIT_1A => X"AA8A28A28A28A28A74C132343334514513028A2818E01F81400050E130106345",
INIT_1B => X"8341A0D46A351A8D46A351A8D46AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA",
INIT_1C => X"FFFFFFFE58C001A0D068341A0D068341A0D068341A0D068341A0D068341A0D06",
INIT_1D => X"10550015400000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"F45A2D16AAAAF7D568A00AA8400000AAFFC21FFF7D542000FFAE821FF552EAAA",
INIT_1F => X"0000AAAE820BA550015400087FD74BAFFD540000F7D155555087BEABFF552ABD",
INIT_20 => X"A8AAAF78015545FFD555555082AAAA10F7FFEAB455500175FF5D2AAAA1000554",
INIT_21 => X"56AB45552ABDE00AAD140010F7D17FF45A2FBC2000A2FFC21555551554005D2E",
INIT_22 => X"AEBFF55082E82145A280001EFF78402145A2AE801555D2E95555552E97410005",
INIT_23 => X"D517DF45557BD5410F7D555545F7AA97410000428AAA557FD5400FF843DE00FF",
INIT_24 => X"0000000AA085568BEFFFAE82000085542155557FEAA10007FEABEFAAD1400AA5",
INIT_25 => X"8EBAA801EF4920AFA10490A17000000000000000000000000000000000000000",
INIT_26 => X"451C75EABEF4124BAF55B6DF6FABAFFD56F010AA8407428A2F1C01FFF7D14202",
INIT_27 => X"5FF552AAFA10007155428A2AE850925D0010400087FD24AAE3DF47010E38E051",
INIT_28 => X"01555D51524004920ADA82EB8A12555EBFB4717D1C2AAFA28EBF5E8B7D550015",
INIT_29 => X"92555492A850381C5F6AB6D4124BAE10BED542010FFD57AF55AAF5D7410A2FBC",
INIT_2A => X"1D5400FF8A38E00F7AABAF7D0000955FDB684051D7F7840517DA2A4871554124",
INIT_2B => X"55D75EFBED5400825D557FF55007BD7410EBDB5017DE38E8708008002FAAA417",
INIT_2C => X"00000000000000000000000082005F6ABFFEBA0870281C5F4716D5D7FEDB7D09",
INIT_2D => X"AAD1401FFFFD5420BAA2AA821FF08043DE10002A964000000000000000000000",
INIT_2E => X"AA2FBD7410A2AE965555D556ABEF080028B55FFFFFDEBAFFD57FE00A280144BA",
INIT_2F => X"AAA2D16ABEF5500175EF552ABDE000855544AAAA82174105D0402000087FC00B",
INIT_30 => X"BF5AAD154400AAFBC015555554001008003FE00AAEA81154AAFFD65FF5D2EBDE",
INIT_31 => X"75EFA2AA155550004021E5582A964BE557FEABEF00002BE10FFD540000FFD56A",
INIT_32 => X"9661000043DEAA085555400FFAAAAA10F7AC28BF558001454DF78017555F7801",
INIT_33 => X"FD55EF5D7BFEEF35055487EFF7D1400105D517FF55087FD7410A2FBC01E7F2AE",
INIT_34 => X"0000000000000000000000000000000000000000010007FEABEFAA84174BA557",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0400000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(4),        -- Port A data input
DOA(0)   => data_read_a_hi(4),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(4),        -- Port B data input
DOB(0)   => data_read_b_hi(4),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_5_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50DF0A0791B3FC1694378283C81FD996A091A32152007AB36B20E03C040C006",
INIT_01 => X"081FBDC49830884C5C6A60000C34C24841280A00084000C8C212892EEA953231",
INIT_02 => X"C809AD5CB118E640A4F008F8011FF0002080000082CCC66609DB7DDDCB1F2036",
INIT_03 => X"25080626BE4C904210831C80084204720B20048A88800000B8E0F8102885500E",
INIT_04 => X"4005122024899100064520C01444429C7804103C0416C007198A3916E0551A04",
INIT_05 => X"46E1829941C9000944C8C022898FE2F20D7D7A104CB5C208E51417C054848912",
INIT_06 => X"CA075CA0E63342991612DF9A8205C0A0B030B20B10480900886E220801073711",
INIT_07 => X"8C732074B68D1A34E3180717FFD13FC72691924098712CE481FDC241D43C1ACD",
INIT_08 => X"16053F180A1286A4E51BD18840C320000075FE91A24458BA4DE0D57992D9BE58",
INIT_09 => X"0A4D8105BF3472304100930258E510601EDE1D8524309285FD416CB402259504",
INIT_0A => X"3110AC0D11C901B2112109204C28B67061E8928920CAD3CFC0140079065A4A65",
INIT_0B => X"C3404959321C284D356A964F8125CD7AC8632614005DFBAACFBC800024091128",
INIT_0C => X"380D6380B6380F638096380F6380B6380D51C04B1C07AD10C14020D233127AD5",
INIT_0D => X"992940513052F4CA8A0A0664A5023CA8470FF000908C383755AF1604E0538096",
INIT_0E => X"200040194FFC044FFA4B08BC85282C91F028D094284A34054A25508605135C01",
INIT_0F => X"BA0C2038ABACBC7C7806F94FF87C002F83F106F94FF87C002F83F2000A04C200",
INIT_10 => X"8D9A70380230F2DFC106F86FF87C002F83F106F86FF87C002F83F3601BFFEBC2",
INIT_11 => X"1F401BFFE7C69E01804E1E6EABE3F040FFD7C7C4BC0E008C7C2FE58FC0A9FFF5",
INIT_12 => X"F8BFDFC8C8120C4DBC802208B2EB2AE777ADFE6F0A47CC0600C2683E0FF8AE3F",
INIT_13 => X"4189B7C56DF47186104C6DE7037FFF00FC0000FC07EE4E7A7076FE28C3082636",
INIT_14 => X"B9E9F272FFFC181C0C2038A7C6DE7A7D909FBFA4070380131CAFB257FBD93902",
INIT_15 => X"2B34E9F56DFBEB1B7F2300C4A80092E0FC1FCE667A7C877FFE828F0080AE1DDA",
INIT_16 => X"51142511405EA00A1344612A898494801602081F87204A9452217159891640D4",
INIT_17 => X"0942511425014450940519425114650140519405194650146511405194050946",
INIT_18 => X"1465114250146501465194051944509445094051146501465014251140509445",
INIT_19 => X"7ED430A983124B2DA6924965B4D5014650142511425094450940519405094450",
INIT_1A => X"EFBEFBEFBEFBEFBE5FDFF3F7F773CF3CF7D796ED39FDEE76DFFCE9F84801B6DB",
INIT_1B => X"BDDEEF77BBDDEEF77BBDDEEF77BBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFB",
INIT_1C => X"FFFFFFFE433B5EEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77B",
INIT_1D => X"AAFFFBFFE00000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"000FFAE821FF552E820105500155555D2AA8A00AA843FFFFF78002155AAAE974",
INIT_1F => X"0000FFAE80000AAAE974BAFFAEAAB45AAAEBDEAAA2FFEAA00AAFFC21FFF7D542",
INIT_20 => X"7FE000055574BA557FFFF55087BEABFF552ABDF45A2D16AAAAF7D56AA00AA840",
INIT_21 => X"E820BA550015400087FD74BAFFD540000F780155555D7BE8B45085168BFFA2D1",
INIT_22 => X"2AAAA10005140145FFFBC01EFAAFFD75FF002E97555A2AABDEAAAAAAAAA00AAA",
INIT_23 => X"A84174BA5D043FF45AAAA974AAF7AEBFF55082AAAA10F7FFEAB455500175FF5D",
INIT_24 => X"000000000A2FFC21555551554005D2EA8AAAF78015545FFD555410552EA8BEFA",
INIT_25 => X"FFF8E0217DBEA4954AAE3FBFDE00000000000000000000000000000000000000",
INIT_26 => X"28A2F1C01D7F7D142028EBAA801EF492087A10490A171455D2EADA28B6803FFF",
INIT_27 => X"ABAFFD56FA10AA8417428E3AE87010A2A4974AAE3AEAFB6DAAA4BDEAAA2F1EDA",
INIT_28 => X"8B6D14516DBD7BEDB7DE381451554AA497FFFF451C75EABEF4124BAF55B6DF6F",
INIT_29 => X"BDEAAAAA0AFA28A2A4850925D0010400087FD24AAE3DF47010E38E0516D5D7BE",
INIT_2A => X"5E8B7D5500155FF552AAFA10007155545F7F1C21D7AAF1D55FF082A9057DA2AA",
INIT_2B => X"FB470384124ADBFFBE84174AA55043FF6DBEAE950AAEB8ABDF7D1C2AAFA28EBF",
INIT_2C => X"00000000000000000000000010A2FBC01555D51524004920ADA82EB8A12410EB",
INIT_2D => X"552EBFEBAF7843DFEFF7AE801EFF780174AAAAFBFEE000000000000000000000",
INIT_2E => X"FA2803FEBAAAD17CEAAAAD140155FFD5420BAA2AA821FF080415410002A96555",
INIT_2F => X"EF080028B55FFFFFDEBAFFD57FE00A280144AAA2AA97400A280174AAA2AEBDFE",
INIT_30 => X"410A2AE965FF557FE8BFF55557FF55FFFBFFEAA5D51554AA087BFEF555D556AB",
INIT_31 => X"55FF0004821FFAAAEBDEAAAA843CEAAAA80174105D0402000087FC00BAA2FBD7",
INIT_32 => X"BEFFF5D2EBDEAAA2D16ABEF5500175EF552ABDE00005554545F7D140145A2D55",
INIT_33 => X"03FE00AAAA81114AAFFD64BA00043FFFFFF80174AA55043DFFFFFAE974BAA2AE",
INIT_34 => X"0000000000000000000000000000000000000000000AAFBC0155555540010080",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"1800000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(5),        -- Port A data input
DOA(0)   => data_read_a_hi(5),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(5),        -- Port B data input
DOB(0)   => data_read_b_hi(5),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_6_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10844B0061A258A2840112C03002C18000402322520070B303301C0381A0086",
INIT_01 => X"0600404820094048008100000042026041000000090800090210080008510204",
INIT_02 => X"080108220C1000004440080000C008010000000001203240080080000988A050",
INIT_03 => X"040000000823404000020A600000002983800584488000103080040C08C00000",
INIT_04 => X"00101610A029B08400044800000000040000102A040810040400100500101800",
INIT_05 => X"05000000800C8300306420002900404400820000000A00804004084001200A00",
INIT_06 => X"64472644640C00808C10D00401823F0020204209101001002650020001052800",
INIT_07 => X"080000242000000461100050818080380900224000200008818028804883E10A",
INIT_08 => X"01FE80E0090242602C0020608000000000043E00000048800021140000881106",
INIT_09 => X"12447E041B102020208000424029006FE0B085013204D0200101006862119140",
INIT_0A => X"4D540B0D916BBE39059191200000200441040108000020006FC5FA6000816908",
INIT_0B => X"8BF05D11A20808454010834225A28962E40AA05510180022FFA6A8800402A06D",
INIT_0C => X"16C1416C5416C5416C3416C3416C7416C500B60A0B60AD04EB4104C093904535",
INIT_0D => X"59802817888180E80112A1660050900003400430CB4911B445A105B05B016C14",
INIT_0E => X"000000062003C90000442006439324280034E85A742D1A16CD2DA30046848048",
INIT_0F => X"00000000000157000600000000000028000C00000000000028000CE800048000",
INIT_10 => X"00000000000000483C00000000000028000C00000000000028000D1080000000",
INIT_11 => X"00108000000000000000000078000A00000000000000000000019A0030000000",
INIT_12 => X"4604000000000000934909080014000000000000000000000000000009005180",
INIT_13 => X"00001230B00000000000049B3C000000000000000001FA000C98000000000002",
INIT_14 => X"E8000E05000000000000000001720002A56000000000000000000FC080000000",
INIT_15 => X"0840000B000404A000000000000000000002099A0003B0000000000000000001",
INIT_16 => X"69DA5685A146D19D084488080904C0A1172240C0781400C81908000205208614",
INIT_17 => X"85A1695A769DA3685A169DA768DA1685A169DA7685A1685A769DA7685A168DA7",
INIT_18 => X"5A368DA1685A769DA168DA3695A569DA3685A169DA5695A368DA1695A569DA36",
INIT_19 => X"7F10800846638C31C71C718638E685A769DA5685A3685A569DA7685A168DA769",
INIT_1A => X"E38E38E38E38E38E76DDB3B7B377DF7DF7D7DE2F39FE3FC3D3EA55FF37F5F7CF",
INIT_1B => X"9FCFE7F3F9FCFE7F3F9FCFE7F3F8E38E38E38E38E38E38E38E38E38E38E38E38",
INIT_1C => X"FFFFFFFF61AC8FE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F",
INIT_1D => X"EFAAAABFE00000000000000000000000000000000000000000000181F007FFFF",
INIT_1E => X"FFFF78002155AAAE974AAFFFBFFE10F7FBE8BEF552E95555552EAABEF082E975",
INIT_1F => X"5410A2AAAAA10087FC01EF552EAAB45F7AE821550851555555D2AA8A00AA843F",
INIT_20 => X"2ABEFA2AEBDFFF552AAAA00AAFFC21FFF7D542000FFAE821FF552E8001055001",
INIT_21 => X"E80000AAAE974BAFFAEAAB45AAAEBDEAAA2FFEAB45552E800AA555568A105D00",
INIT_22 => X"D56AA00AA8400000007BC21FFAA803FFEF5551420105D5568B45FF8400000FFA",
INIT_23 => X"7FBC2155007FC20BAA2D5575FF087FFFF55087BEABFF552ABDF45A2D16AAAAF7",
INIT_24 => X"0000001555D7BE8B45085168BFFA2D17FE000055574BA557FFFE10F7AAA8A00F",
INIT_25 => X"D4924ADBD70820975FFA2A4BFE00000000000000000000000000000000000000",
INIT_26 => X"455D2EADA28B6803FFFFFF8E0217DBEA4954AAE3FBFDE38F7FFEABFF412A9056",
INIT_27 => X"1EF492087010490A07038B6A0AFA38007BC51EF4920AFB55EBA4851450855555",
INIT_28 => X"5082555F68A3855002FBC7BEA4BFFFF492EADA28A2F1C01D7F7D142028EBAA80",
INIT_29 => X"6DB45E38A07028E3AE87010A2A4974AAE3AEAFB6DAAA4BDEAAA2F1EDB55492A8",
INIT_2A => X"4BAF55B6DF6FABAFFD56FA10AA84174381C7FC01C7B68E3DFC75555400105D51",
INIT_2B => X"7FFFE38F7A0AFA38E3FFC21450071C2092A2D5571FF0851FDF451C75EABEF412",
INIT_2C => X"0000000000000000000000016D5D7BE8B6D14516DBD7BEDB7DE381451554AA49",
INIT_2D => X"F7FBEABEF002E801EF00003FF550800155FFA2803CE000000000000000000000",
INIT_2E => X"5A28417555085154555552EBFEBAF7843DFEFF7AE801EFF780174AAAAFBFEEAA",
INIT_2F => X"55FFD5420BAA2AA821FF080415410002A964AAFF803DEAA087FD55FF00043DF4",
INIT_30 => X"EBAAAD17CF55002E95410557BEAABA55043DF55F7803FFEF002ABEEAAAAD1401",
INIT_31 => X"DF455D51420105D517DF55AAAA964AAA2AA97400A280174AAA2AEBDFEFA2803F",
INIT_32 => X"7CF555D556ABEF080028B55FFFFFDEBAFFD57FE00A280144BA5D7FC2155FFAAB",
INIT_33 => X"BFFEAA5D51554AA087BFEEAAF7803DEAAAAFBC0155085540000A2D5575FF0851",
INIT_34 => X"00000000000000000000000000000000000000001FF557FE8BFF55557FF55FFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"1200000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(6),        -- Port A data input
DOA(0)   => data_read_a_hi(6),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(6),        -- Port B data input
DOB(0)   => data_read_b_hi(6),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_7_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10844B00482258A2842112C02450418800002300500030B303300C018180002",
INIT_01 => X"0200084020084048040080000201026040000000080000080200090000510204",
INIT_02 => X"4801082048100000444008040080000041000000000222400800000009000010",
INIT_03 => X"0401018108A144D0000208424000002103006480088000003080000408C10000",
INIT_04 => X"0000120022419000000C80000000000400201829040000050001940400301820",
INIT_05 => X"04000000800840092CC080214144004400000000000800065004004020220800",
INIT_06 => X"40870408600000808C10D4500080008020200008001001000240000061052002",
INIT_07 => X"08000024200000046010005281848001494020400031240C8C8238A06A000988",
INIT_08 => X"40050001090242602C0408408000000000243E00000048800020154000881024",
INIT_09 => X"024401041B132820000011424069004000B20403200891420101026A42210440",
INIT_0A => X"013800A0281400300C0010200008B20663970148004424006818026200004800",
INIT_0B => X"01C1103022881845421082C2C0082300401121810012004600001010040028A0",
INIT_0C => X"1200112001120011204112041120411206089010890100408040008012101414",
INIT_0D => X"09146817802988694902A02451109006230006E0808294008C02848148092001",
INIT_0E => X"000000042C00040002000004020020490020401020081004482501010C120948",
INIT_0F => X"0130C807144102420700052000003C00780B00052000003C007808450484C000",
INIT_10 => X"400002C0E00E0D003300052000003C00780B00052000003C0078099080001000",
INIT_11 => X"80908000100000661801E18042100E000060100000B038038380124038000102",
INIT_12 => X"053A010111848322020512000414400000002000A1001058300C0741C0054120",
INIT_13 => X"90644029D008240864231011BF00008000C3C003F00186040EE8041204321188",
INIT_14 => X"18100D770008060130C807182106040375600411004C2600E3400C2740202230",
INIT_15 => X"9094100A8CA406A0002C812240B0201F0380211604037740004010472041E201",
INIT_16 => X"40100401006E8118104428088904C4C414420080049450801000088444300601",
INIT_17 => X"0906409004010040104409024090240906401004010040102409024090240100",
INIT_18 => X"1024090241900401004090240902401004010040902409004010440100409024",
INIT_19 => X"004420A945841040002082080004110240902409004110040902409024110040",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFEDD9EC000000000000000000000000000000000000000000000000000",
INIT_1D => X"BA082AAAA00000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"555552EAABEF082E975EFAAAABFFEF002ABDF555D5157555F7FBC00AAAAD5400",
INIT_1F => X"FEAAAAAABDF55FFFBFDF55555568ABAAAD5401FF5D2AAAA10F7FBE8BEF552E95",
INIT_20 => X"400005D55554105D51401555D2AA8A00AA843FFFFF78002155AAAE974AAFFFBF",
INIT_21 => X"AAAA10087FC01EF552EAAB45F7AE821550851554AAF7FBFFEAA007BFFFEFF7D5",
INIT_22 => X"2E800105500155EF5D2EBFF450000020AA5D7BC0000F7D555545A28000010A2A",
INIT_23 => X"FAAA8A10FFD568ABAA2D56AAAAF7AABFE00AAFFC21FFF7D542000FFAE821FF55",
INIT_24 => X"000000145552E800AA555568A105D002ABEFA2AEBDFFF552AAAABAA2AE95555F",
INIT_25 => X"5E3F5C20BAAAD5420821C2EAAA00000000000000000000000000000000000000",
INIT_26 => X"38F7FFEABFF412A9056D4924ADBD70820975FFA2A4BFFFF1C2EB8F4555555054",
INIT_27 => X"17DBEA4954AAE3FBFDE82B6AEBAF55E3FFFAF55555F6FA92BED5421C75D20AAA",
INIT_28 => X"FE920075FDFD7F7D5400385D51504385D55401455D2EADA28B6803FFFFFF8E02",
INIT_29 => X"5057DB68E02038B6A0AFA38007BC51EF4920AFB55EBA485145085555492F7F5F",
INIT_2A => X"142028EBAA801EF492087010490A071EF4920B8F45140E07082417BC2000EBD5",
INIT_2B => X"2EADA92A2A09257DE3A4AAA10F7D16FAAABED56AE82F780BAE28A2F1C01D7F7D",
INIT_2C => X"00000000000000000000000155492A85082555F68A3855002FBC7BEA4BFFFF49",
INIT_2D => X"552EAAB455D5142155AAD1400AAA2D1420005D2EA9A000000000000000000000",
INIT_2E => X"0F7D1421555D042BAAAF7FBEABEF002E801EF00003FF550800155FFA2803CFFF",
INIT_2F => X"BAF7843DFEFF7AE801EFF780174AAAAFBFEE00F7AAAAB55AAFBEAB555D7BFDE0",
INIT_30 => X"555085154400FFD17FE1000517FF55FFD5420BA5D55400BA555543155552EBFE",
INIT_31 => X"5400087BC0000A2D5421EFF7AE810AAFF803DEAA087FD55FF00043DF45A28417",
INIT_32 => X"2BAAAAAD140155FFD5420BAA2AA821FF080415410002A965FF080428B45552A9",
INIT_33 => X"43DF55F7803FFEF002ABEE00A280001FFA28028A00FFD17DEAAF7D56AA10FF84",
INIT_34 => X"0000000000000000000000000000000000000000155002E95410557BEAABA550",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"01FFFFFFFFE00000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(7),        -- Port A data input
DOA(0)   => data_read_a_hi(7),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(7),        -- Port B data input
DOB(0)   => data_read_b_hi(7),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_8_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00000648E2840112C00000418000002700500030B3032000000000082",
INIT_01 => X"000009C21838284D1C2160000E12424840000000180800080200000040110204",
INIT_02 => X"080108000090000004400C040080000051000000000002400800000009000010",
INIT_03 => X"00000100043008D0000200024000000003800504488000103080880008800000",
INIT_04 => X"00009410A028A084000440000000000400001022040800150400808500321800",
INIT_05 => X"8500010080048A09302420202804400400800010200A00020204084011014A00",
INIT_06 => X"2447A244608800840490D0040007FE0021204288001000000050024001042800",
INIT_07 => X"4800002420000004201000D281040003182020400031241C0D80004041BFE88A",
INIT_08 => X"4005000108020220240000048000000000043E00000048800000010000881000",
INIT_09 => X"0204010519110020008111020069004008A28501120450220101214122509140",
INIT_0A => X"0528A52291490029019190200008B20E23008028000208804010024000004000",
INIT_0B => X"13C151312A8808454104824001280108A409A044001200020020989000000061",
INIT_0C => X"0000000000000000000000000000000000400020000229508040008012105400",
INIT_0D => X"48022817880508602102A1200810B2020340043248CA00240420000000400040",
INIT_0E => X"4100820020000C0000442142419120000014684A34251A12CD2CA30042840248",
INIT_0F => X"45F3D80000000001020404000783FC0000010404000783FC000000880284C010",
INIT_10 => X"02658FC7E0000000010404000783FC0000010404000783FC000001500000103D",
INIT_11 => X"40500000103961FE78000000000402400020003B43F1F8000000022010800002",
INIT_12 => X"0080001617CD800000080B000804080000020090659833F9F03C000000000000",
INIT_13 => X"B000000400018639EC000000000000FE03FFC00000000600840000C31CF60000",
INIT_14 => X"180204000001E2A3F3D80000000600802000401AA8FC7E00000000100002C2F5",
INIT_15 => X"005404020000104480DC372B47F060000000000600802000017570FF60000000",
INIT_16 => X"28CA328CA34650850A4C000009A494A015624080044440481908000220308640",
INIT_17 => X"8CA328CA328CA328CA3284A1284A1284A1284A1284A1284A328CA328CA328CA3",
INIT_18 => X"CA1284A1284A1284A128CA328CA328CA328CA3284A1284A1284A1284A128CA32",
INIT_19 => X"64108088440000000000000000028CA1284A1284A1284A128CA328CA328CA328",
INIT_1A => X"E79E79E79E79E79EDFC8F33637D6CB6CB2900A282950FAF15E8428917C51E75D",
INIT_1B => X"87D3E1F0F87C3E1F0F87C3E1F0F9E79E79E79E79E79E79E79E79E79E79E79E79",
INIT_1C => X"FFFFFFFECB0593E1F4F87D3E1F4F87D3E1F4F87D3E1F4F87D3E1F4F87D3E1F4F",
INIT_1D => X"10002ABFE00000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"555F7FBC00AAAAD5400BA082AAAA10000000010F7D5421EF007BC01FF5D7FFFE",
INIT_1F => X"FEAA5551554AAFF80021EF002A820BAFF8428A00A2AAAABEF002ABDF555D5157",
INIT_20 => X"E8BEFFFFFEAB55002ABFE10F7FBE8BEF552E95555552EAABEF082E975EFAAAAB",
INIT_21 => X"ABDF55FFFBFDF55555568ABAAAD5401FF5D2AAAB55FFD1400AA5D7FC01EFA2FF",
INIT_22 => X"AE974AAFFFBFFEAA08001555555516ABEFA280020AA5D043DF55557BEAAAAAAA",
INIT_23 => X"8042AB55005140145AAFFE8AAAF7D1401555D2AA8A00AA843FFFFF78002155AA",
INIT_24 => X"0000000AAF7FBFFEAA007BFFFEFF7D5400005D55554105D51400005551421EF0",
INIT_25 => X"71C7FC21EF5D75FFE10142EBAE00000000000000000000000000000000000000",
INIT_26 => X"FF1C2EB8F45555550545E3F5C20BAAAD5420821C2EAAA101C0005000E3D1401D",
INIT_27 => X"BD70820975FFA2A4BFE925D51554AAE384001FF142E800AAFF802AA28AAAEAFB",
INIT_28 => X"7092557BC21D7BEF5EDBC7FFF1EFB6D1420BAE38F7FFEABFF412A9056D4924AD",
INIT_29 => X"3AF55417BEDA82B6AEBAF55E3FFFAF55555F6FA92BED5421C75D20AAB45F7D14",
INIT_2A => X"03FFFFFF8E0217DBEA4954AAE3FBFDEAA1C001056D415F6ABEFA284020824904",
INIT_2B => X"55400385D51401EF00002FB45085F4016DAAF1EDAAAFFFB401455D2EADA28B68",
INIT_2C => X"00000000000000000000000092F7F5FFE920075FDFD7F7D5400385D51504385D",
INIT_2D => X"5D0417410AAD540155557FC01EF5D557DE105D2AA8A000000000000000000000",
INIT_2E => X"AF7842AABAA2AEBDFFF552EAAB455D5142155AAD1400AAA2D1420005D2EA9A10",
INIT_2F => X"EF002E801EF00003FF550800155FFA2803CE105D55574BAA280021EF5D2E820B",
INIT_30 => X"1555D042BB45FFD157410557FC0155F7D57FF55F7D57FFEF550028AAAF7FBEAB",
INIT_31 => X"8BFFAA8000000080428B55087FFFE00F7AAAAB55AAFBEAB555D7BFDE00F7D142",
INIT_32 => X"C2155552EBFEBAF7843DFEFF7AE801EFF780174AAAAFBFEEBA5D04021EF087BE",
INIT_33 => X"5420BA5D55400BA5555430BA5555421EF00043FF45007BC21FFA2D57FEBAF7FB",
INIT_34 => X"0000000000000000000000000000000000000000000FFD17FE1000517FF55FFD",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0800000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(8),        -- Port A data input
DOA(0)   => data_read_a_hi(8),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(8),        -- Port B data input
DOB(0)   => data_read_b_hi(8),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_9_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00018248A2840112C00002C18000002300500030B3032000000000006",
INIT_01 => X"000008000000004C0020000000100268413C0A61590001D90213C00000110204",
INIT_02 => X"680108200010000054400C040080000041000000010002400800800009082011",
INIT_03 => X"00040100000020D0000200124000000043800504488000103081880008800000",
INIT_04 => X"00001410A00AA084000400000200000400001020040010050020820400101880",
INIT_05 => X"0400040080048A09202420000C00410400000000000800020804004000000800",
INIT_06 => X"24478244640800840410D4144002008020200009301000000140000201042000",
INIT_07 => X"0800002C20000004301000128104000100002040003164040D80000040000888",
INIT_08 => X"40050003080202202400000080000000000C3E00000048800010230000881000",
INIT_09 => X"0024010411110420008010020021004000A204011200500001010000AA10C000",
INIT_0A => X"7945282804010009009090200008B20223800008020000004010024204000440",
INIT_0B => X"114100112208084540008240110001002400A000001000020008288000000420",
INIT_0C => X"010400100001040010000104001000010400080000820800000000801010100A",
INIT_0D => X"08403C16800100640182A0210010921003400412484202200400004004001040",
INIT_0E => X"410082002C000C000240004240932041401468CA34651A32CD28A22002840048",
INIT_0F => X"000000000000144002000420000000280001000420000000280000000284C010",
INIT_10 => X"4000000000000048010005000000002800010005000000002800001000001000",
INIT_11 => X"0010000010000000000000002A00020000201000000000000001820010000002",
INIT_12 => X"40BA00011000000090000B000004000000000000A00000000000000009000020",
INIT_13 => X"00001205D0080400000004803F0000800000000000004C0004E8001200000002",
INIT_14 => X"B000047700000600000000000054000135600011000000000000025740200200",
INIT_15 => X"001400020CA406A0000080200000000000020804000137400040000000000000",
INIT_16 => X"28CA328CA36651951A4CA8000984D4E557220080040440481908000001300614",
INIT_17 => X"84A1284A1284A1284A1284A1284A1284A1284A1284A1284A328CA328CA328CA3",
INIT_18 => X"4A1284A1284A1284A128CA328CA328CA328CA328CA328CA328CA328CA3284A12",
INIT_19 => X"2540A809010000000000000000028CA328CA328CA328CA3284A1284A1284A128",
INIT_1A => X"4534D34D34D34D344A2D840100E4920824055CD13333D2379A2A24018615C38E",
INIT_1B => X"268341A0D068341A0D068341A0D1451451451451451451451451451451451451",
INIT_1C => X"FFFFFFFE6DA90341A4D268341A0D069349A0D069349A0D068341A4D268341A4D",
INIT_1D => X"FFFFD557400000000000000000000000000000000000000000000001FFFFFFFF",
INIT_1E => X"1EF007BC01FF5D7FFFE10002ABFF55F7D168A00552E95555007BFFF55087BE8B",
INIT_1F => X"AA10F7FBC0145F7AE801EFF7FBFFF455D7BC0155F7D557410000000010F7D542",
INIT_20 => X"BDE00AA803FFEF5D55421EF002ABDF555D5157555F7FBC00AAAAD5400BA082AA",
INIT_21 => X"1554AAFF80021EF002A820BAFF8428A00A2AAAAAAAF7D17DE00FFFBD5555A2AA",
INIT_22 => X"2E975EFAAAABFFEF002A954BA5551421EF552E954105D00021455555420AA555",
INIT_23 => X"7D5575EFA2FFD75455D7BE8A005D5557410F7FBE8BEF552E95555552EAABEF08",
INIT_24 => X"000000155FFD1400AA5D7FC01EFA2FFE8BEFFFFFEAB55002ABFE10080028BFFF",
INIT_25 => X"D1C71F8F7D147BEFBEFEBD152400000000000000000000000000000000000000",
INIT_26 => X"101C0005000E3D1401D71C7FC21EF5D75FFE10142EBAF7DE3D16DA0041209056",
INIT_27 => X"0BAAAD5420821C2EAAA10E3FFC0145F7A0801FFEBFBF8F6D417BC716DEBD1524",
INIT_28 => X"DE28F7F5D0545B6AAB8E38B68A3AFFF5551471FF1C2EB8F45555550545E3F5C2",
INIT_29 => X"021455D5B470925D51554AAE384001FF142E800AAFF802AA28AAAEAFABAE3D17",
INIT_2A => X"A9056D4924ADBD70820975FFA2A4BFFFF082E974BA4155401C7552097428550E",
INIT_2B => X"20BAE0008002ABFFF7DB505FFAAFBD7555417FEFA00495B52438F7FFEABFF412",
INIT_2C => X"00000000000000000000000145F7D147092557BC21D7BEF5EDBC7FFF1EFB6D14",
INIT_2D => X"AAD17DE100804001EF55516ABFF557BFDFEFA2D5400000000000000000000000",
INIT_2E => X"F007FD55FFA2D5400105D0417410AAD540155557FC01EF5D557DE105D2AA8BEF",
INIT_2F => X"455D5142155AAD1400AAA2D1420005D2EA9A00A2FBC0145FF84001EFA2FFEABF",
INIT_30 => X"ABAA2AEBDEAAAAD17DEBAFFD142155FFAAAAABAFFAAAABFF5551555FF552EAAB",
INIT_31 => X"01555D00154AA552E801455D7BD54105D55574BAA280021EF5D2E820BAF7842A",
INIT_32 => X"C00AAF7FBEABEF002E801EF00003FF550800155FFA2803CFFF002E954BA00514",
INIT_33 => X"57FF55F7D57FFEF550028A10000428BEFF7FFC01FFA2FFD5545007BFDE10087F",
INIT_34 => X"0000000000000000000000000000000000000000145FFD157410557FC0155F7D",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"1000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(9),        -- Port A data input
DOA(0)   => data_read_a_hi(9),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(9),        -- Port B data input
DOB(0)   => data_read_b_hi(9),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_10_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000B0001800002840002C0000281800020030000000033122000400992006",
INIT_01 => X"A140098018300848180060000C00424040000000080000080200000000110200",
INIT_02 => X"0801080200100000046558000080000041000000002402400800000009008010",
INIT_03 => X"0001000084000040842242000210810803006400088000003080054288C10000",
INIT_04 => X"0000100022008000000C08000800000400A83A2044200C840000000400001820",
INIT_05 => X"0400000080000000248080210044000402000025000800000004203010100800",
INIT_06 => X"00078000600000040410D4102850008024240001981024A82000010461052000",
INIT_07 => X"0800002430204084281000128100000300002040003124040D80204040000888",
INIT_08 => X"0005000108020220240030008000000000043E0408104C800000010000881100",
INIT_09 => X"0004010511100020200000400021004008808060400111080000200002008400",
INIT_0A => X"0000000000010000060210200008B20223048808000200000010024000000000",
INIT_0B => X"03C0411009808245010002000028000080002105010000000020A34249020801",
INIT_0C => X"8004480044800048000480044800448000440002400221008840009012104400",
INIT_0D => X"0000540100000020088000000100100013000400000800040062400200440004",
INIT_0E => X"4100820020000400020000400200204900800000000000000000000100120800",
INIT_0F => X"0000000000101400020401000000002804010401000000002804000000048010",
INIT_10 => X"0000000000000068010400200000002804010400200000002804005000000000",
INIT_11 => X"0050000000000000000000102800024000400000000000000011820010800100",
INIT_12 => X"4000010000000000D00000080004080000002000000000000000000009020000",
INIT_13 => X"00001A000000200000000681000000000000000008004A000400040000000003",
INIT_14 => X"A800040000080000000000000852000020000400000000000010024000002000",
INIT_15 => X"0000000200000000002000000000000000021802000020000000000000000020",
INIT_16 => X"00000040002800100004200009048005C0000080000400000000000000200654",
INIT_17 => X"0802008020080200802008020080200802008020080200800000000000000000",
INIT_18 => X"0000000000000000000080200802008020080200802008020080200802008020",
INIT_19 => X"2054282101000000000000000000000000000000000000000000000000000000",
INIT_1A => X"A28A28A28A28A28A355950666151451453D51A242A503F834E5C49851D243555",
INIT_1B => X"994CA6532994CA6532994CA65328A28A28A28A28A28A28A28A28A28A28A28A28",
INIT_1C => X"FFFFFFFE8E31DCAE532994CA6532995CAE572B94CA6532994CA6572B95CAE532",
INIT_1D => X"AAFFFBC2000000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"555007BFFF55087BE8BFFFFD557400FF842ABEFA2AAA8B5500003DF55F7D568A",
INIT_1F => X"FE0008556ABFFA2D16AB550000021FFF7D17FFEF08042AB55F7D168A00552E95",
INIT_20 => X"3FF55A2D557400557BC2010000000010F7D5421EF007BC01FF5D7FFFE10002AB",
INIT_21 => X"BC0145F7AE801EFF7FBFFF455D7BC0155F7D557545FFAE820AA007BFDFEF5500",
INIT_22 => X"D5400BA082AAAA00FFAE820AAAAAABDFEFF78028BEF005140145A2842AA10F7F",
INIT_23 => X"AD56AB55A2D157400552EBFFEF5D7BD75EF002ABDF555D5157555F7FBC00AAAA",
INIT_24 => X"0000000AAF7D17DE00FFFBD5555A2AABDE00AA803FFEF5D55420BA08557FEBAA",
INIT_25 => X"51C0E3AF55F7DF68ABAE3F1C0000000000000000000000000000000000000000",
INIT_26 => X"7DE3D16DA0041209056D1C71F8F7D147BEFBEFEBD152400F7842FBD7B6AAAAB5",
INIT_27 => X"1EF5D75FFE10142EBAE0008556FBD7B6DB6AB7D1C0A001D7FFD178FC71C0E28B",
INIT_28 => X"2092147BFAFEF49043AF45A2DF504285D71C00101C0005000E3D1401D71C7FC2",
INIT_29 => X"4017DA28428A10E3FFC0145F7A0801FFEBFBF8F6D417BC716DEBD15256DF7AA8",
INIT_2A => X"550545E3F5C20BAAAD5420821C2EAAA00E3AA82092A2AABAFD7EB8A2ABC70855",
INIT_2B => X"51470821C557AE92A2DF6AB7DA2DF50410412ABDFC75D7BD55FF1C2EB8F45555",
INIT_2C => X"000000000000000000000000BAE3D17DE28F7F5D0545B6AAB8E38B68A3AFFF55",
INIT_2D => X"FF803DF45FFAEA8B555D2EAAB45F7FBE8ABAAAD5400000000000000000000000",
INIT_2E => X"5FFD168B55552AA8BEFAAD17DE100804001EF55516ABFF557BFDFEFA2D540010",
INIT_2F => X"10AAD540155557FC01EF5D557DE105D2AA8A0008557FF45FFFFE8BEF5D2E8015",
INIT_30 => X"5FFA2D5401FFF7AA800105D7FE8BEF08002AB45AAFFC00AA5D51400105D04174",
INIT_31 => X"AB55AAAEAAB450055421FFAA8428A00A2FBC0145FF84001EFA2FFEABFF007FD5",
INIT_32 => X"D55FF552EAAB455D5142155AAD1400AAA2D1420005D2EA9A10A2AA82010AAAEA",
INIT_33 => X"AAAABAFFAAAABFF555155400555568A10AAFBEABEFA2FFC0010082ABFF55557B",
INIT_34 => X"00000000000000000000000000000000000000000AAAAD17DEBAFFD142155FFA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"11FFFFFFFFE00000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(10),        -- Port A data input
DOA(0)   => data_read_a_hi(10),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(10),        -- Port B data input
DOB(0)   => data_read_b_hi(10),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_11_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10180B05A0010402840602C2D001019000000300000000330A20080EC180002",
INIT_01 => X"AB400984B83008481800E0000C26426040000000080000088200000802112220",
INIT_02 => X"8801081438106400A4F55800008000004100000040CCE24208005000C9060032",
INIT_03 => X"000406A492E6E440842254D002108153422004800880000030C0315688C00006",
INIT_04 => X"00001201200090001205400000000094108C322644240C840008030440111800",
INIT_05 => X"444000888008010028404002A002009402400025080880000C04223000170900",
INIT_06 => X"40871408620B00801410D94CAAD0018024242008A8102CA88A44010401042200",
INIT_07 => X"08320054B624408428100094ADD080011721A04000316C140CA1A8A1F9001889",
INIT_08 => X"140500090B02C2E0EC04D1C08000000000647E858A104C920C81A5011088A61C",
INIT_09 => X"002481041F165820000101024061004004800567603592A801014C4642601100",
INIT_0A => X"01002020000101B0070310200008B60A23A51B28020CE24E4010026004000440",
INIT_0B => X"03404110230CBA457670820140212100C0692644010001420038935269093161",
INIT_0C => X"2A0872A0C72A0872A0C72A0C72A0872A0C595043950421400800009010104280",
INIT_0D => X"8852141110244066C0820221480010AA73000420808CAC040464D280144050C7",
INIT_0E => X"410082022C000C0002020094030220C960A0409020481024482501A004014100",
INIT_0F => X"6DA02836090540355D86C046619A54052A5B86A0466196940631682800048010",
INIT_10 => X"8B68AA2C60289802AB86A046619A54052A5B86C04661969406316AC018B0E293",
INIT_11 => X"1FC09CB0E1076D4A200B2AC611A3D0405886C6EB211550815A8A2686EC81E2A4",
INIT_12 => X"9C0418CE0C5E8F650E48000892B37885620C1E1A06D7016A90A4626D82B10F1B",
INIT_13 => X"F1E164E02144D335546F28724001B030A56140A184483000C410A2699A2E32AC",
INIT_14 => X"415AAE8018A0A01B2990242E278056AAA203920E0BAE2012C08281808319C186",
INIT_15 => X"9B80D44F9051C049B18A12CB481042AD140C227002A0A02066954E7540CCDB58",
INIT_16 => X"4090240902468118104408000904C0C0964200800200108010003A02272400C1",
INIT_17 => X"0902409024090240902409024090240902409024090240902409024090240902",
INIT_18 => X"1004010040100401004090240902409024090240902409024090240902409024",
INIT_19 => X"2014002840000000000000000004010040100401004010040100401004010040",
INIT_1A => X"0020820820820820A069105251C00000015418982201060302C4281390042104",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFE0FC1C000000000000040200000000000000000001008000000000000",
INIT_1D => X"55000015400000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"B5500003DF55F7D568AAAFFFBC2010557BEAA10AAFBE8A00557BFFFEF007BC21",
INIT_1F => X"75455D7FE8BFF5D7FD540055003FFEFFFD142145000000000FF842ABEFA2AAA8",
INIT_20 => X"C0145557FC2010557FFDF55F7D168A00552E95555007BFFF55087BE8BFFFFD55",
INIT_21 => X"56ABFFA2D16AB550000021FFF7D17FFEF08042AB55A2AAAAB4508517FE00557B",
INIT_22 => X"7FFFE10002ABFE00AAFFE8AAAFF8402000550002145085555400F7FFE8A00085",
INIT_23 => X"8043FEBA002A975EFF7D17DFFFAA8000010000000010F7D5421EF007BC01FF5D",
INIT_24 => X"000000145FFAE820AA007BFDFEF55003FF55A2D557400557BC2145A2D1421450",
INIT_25 => X"8557BF8FEF1C7FC516D080E15400000000000000000000000000000000000000",
INIT_26 => X"00F7842FBD7B6AAAAB551C0E3AF55F7DF68ABAE3F1C00005D7BEDA00B6F1EFA2",
INIT_27 => X"F7D147BEFBEFEBD15257D5D7FEFBD7417BD5438550038FC7FFDF4216D080E070",
INIT_28 => X"DB4514517FE105575C216D5571C50104171FDF7DE3D16DA0041209056D1C71F8",
INIT_29 => X"52400FFF1EFA0008556FBD7B6DB6AB7D1C0A001D7FFD178FC71C0E28B6DA2AEA",
INIT_2A => X"1401D71C7FC21EF5D75FFE10142EBAE10A2FBEFA92F78A05028550E001451455",
INIT_2B => X"71C016DB6D54514500003FEBA1420905FFFFDF78FC7BE84050101C0005000E3D",
INIT_2C => X"0000000000000000000000016DF7AA82092147BFAFEF49043AF45A2DF504285D",
INIT_2D => X"5D7FFDE00F7D17FEBA557BEABEF557BD55EF082A974000000000000000000000",
INIT_2E => X"5F7FBC01FF082A97410FF803DF45FFAEA8B555D2EAAB45F7FBE8ABAAAD540010",
INIT_2F => X"100804001EF55516ABFF557BFDFEFA2D5401FF5D7FFDF55007BD74BA5D042AB4",
INIT_30 => X"B55552AA8BEFAAAABFF5555517FE005555401FF55515541000517FFEFAAD17DE",
INIT_31 => X"74BA5D2A801455D5140000FFD57FE0008557FF45FFFFE8BEF5D2E80155FFD168",
INIT_32 => X"174105D0417410AAD540155557FC01EF5D557DE105D2AA8A10AAFBFFE00F7AA9",
INIT_33 => X"02AB45AAFFC00AA5D51401FFFFD15555500003FEBA5D04001EFFFFFE8B55FF84",
INIT_34 => X"00000000000000000000000000000000000000001FFF7AA800105D7FE8BEF080",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"1000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(11),        -- Port A data input
DOA(0)   => data_read_a_hi(11),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(11),        -- Port B data input
DOB(0)   => data_read_b_hi(11),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_12_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50080B01BC002006940202C0DE041196A83183000000023322287E0FC000006",
INIT_01 => X"0E000C068000E04D40238000001702684000000008000008820009280A553231",
INIT_02 => X"2809AD0E7D180040945008040090000061800000C0E2F66009DA3D11CB148015",
INIT_03 => X"210D050012F6F8D2108216E24842005B8A20640008800000B8E0141C28851006",
INIT_04 => X"0080100022408000060DE0C00466630C70241837041000040800820480001AA4",
INIT_05 => X"04800018800000003C808003E0C8001401000000040900020904004000070800",
INIT_06 => X"00074000601300119E12D348438000803030800020100800AF08000261042400",
INIT_07 => X"8C53200CA4850224301807D1CB45900147E03040083124FC0CD0C8A1FF00198C",
INIT_08 => X"46050013081206A4A503A9E8C0812000001C7E11A24058B84D40E33992D98F7E",
INIT_09 => X"1004810491175C200000820018A5104010C01086003C13E000004EDF02040004",
INIT_0A => X"0000000000010000180018200408B27E234913E9004CFA09A818024800902109",
INIT_0B => X"014100580004304D267C06CCD0056600007827C00000008C00000000000219C0",
INIT_0C => X"2F0C32F0832F0832F0C32F0832F0832F0C197861978400040000208010120ACA",
INIT_0D => X"E0BF40403CFE7E03E8080382FD0018FE670004000006AE01180493C5BC1AF083",
INIT_0E => X"2000401EA0000440000800A0040028108000000000000000000000A74812DF00",
INIT_0F => X"C48DF8362F658A7E5F82CD23B6B0E403DBBE82C563B6A4E403DBB88C0E048200",
INIT_10 => X"454CFBE5403AB992F282C563B6B0E403DBBE82CD23B6A4E403DBBB1084E4B25A",
INIT_11 => X"851000E4B1D32BAB504BB74AD3F3FE04A8E0D0C319A7988B6F0C75CFD801A962",
INIT_12 => X"BEC4118D994B866E2E8C3808B6B63040328E7A33AF99B0AC20DE634D06C437BF",
INIT_13 => X"70CDC5F6214CA5991C6A7177402C49CA354D808D358A927EAD10A652CC8E3538",
INIT_14 => X"49F36E80083C3EAEB2003695430A7CDAA289553922990C11A4E494988231B325",
INIT_15 => X"3BC0FD5B304AD05A946D81616970A225658940BA7CDAA0A312666BD600E5550B",
INIT_16 => X"00000000001000000104200A89A4D0040000008003B81000000021CFEE02E280",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"8020080200802008020000000000000000000000000000000000000000000000",
INIT_19 => X"0544202101000000000000000000080200802008020080200802008020080200",
INIT_1A => X"4124924924924924481C040000B51451440146E518222204D82A5446021090CB",
INIT_1B => X"2C964B2190C86432190C86432190410410410410410410410410410410410410",
INIT_1C => X"FFFFFFFEF001D64B2592C964B2592C964B2592C964B2592C964B2592C964B259",
INIT_1D => X"00AAFBC2000000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"A00557BFFFEF007BC2155000015555087FC0010AAFBFFE100004020BAAAFFD54",
INIT_1F => X"2155AA8400000A2AABFF45550400000AAFBFFFEF550000010557BEAA10AAFBE8",
INIT_20 => X"C0010555155555FF8017400FF842ABEFA2AAA8B5500003DF55F7D568AAAFFFBC",
INIT_21 => X"FE8BFF5D7FD540055003FFEFFFD142145000000145A2AA821EFFFFFD7410007F",
INIT_22 => X"7BE8BFFFFD5574000051420BA557FC2145557FC20AAA2D57DEBAA2FBD55455D7",
INIT_23 => X"82EAAA00550415410AAFBFFFEF55042AB55F7D168A00552E95555007BFFF5508",
INIT_24 => X"000000155A2AAAAB4508517FE00557BC0145557FC2010557FFDE10AA84000000",
INIT_25 => X"0000A02092B6F5D2438A2FBC2000000000000000000000000000000000000000",
INIT_26 => X"005D7BEDA00B6F1EFA28557BF8FEF1C7FC516D080E1557D0075C7028B6F1FAE0",
INIT_27 => X"F55F7DF68ABAE3F1C017DAA8E07028B6A0BFF6D490E00000BEF5FAFEF4904070",
INIT_28 => X"51FFE3FBD0438007FC00385D555556DEB8410400F7842FBD7B6AAAAB551C0E3A",
INIT_29 => X"7DEBAA2FBD557D5D7FEFBD7417BD5438550038FC7FFDF4216D080E0716DAAA08",
INIT_2A => X"09056D1C71F8F7D147BEFBEFEBD152400005F450BA417BC51454971C20AAB6D1",
INIT_2B => X"71FDE10BE8E070280020AAA28410410400BEFBFAFEF49042AB7DE3D16DA00412",
INIT_2C => X"0000000000000000000000016DA2AEADB4514517FE105575C216D5571C501041",
INIT_2D => X"0055574BAFFD568A10002A82000FFD5400AAA2FBC00000000000000000000000",
INIT_2E => X"0FFD568BEF0004174105D7FFDE00F7D17FEBA557BEABEF557BD55EF082A975EF",
INIT_2F => X"45FFAEA8B555D2EAAB45F7FBE8ABAAAD5401EFA2AA974BAF7803FFFF002A8200",
INIT_30 => X"1FF082A975EFA280175FFAAFFC00BA087FC20AA5D55555FFA28000010FF803DF",
INIT_31 => X"75450851420BAFFD57DEAAAAFBD75FF5D7FFDF55007BD74BA5D042AB45F7FBC0",
INIT_32 => X"28BEFAAD17DE100804001EF55516ABFF557BFDFEFA2D540010007FD74AA007BD",
INIT_33 => X"5401FF55515541000517FE10F7AA954AA080428AAA000002010FFFFE8BEF0804",
INIT_34 => X"00000000000000000000000000000000000000001EFAAAABFF5555517FE00555",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"01FFFFFFFFE00000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(12),        -- Port A data input
DOA(0)   => data_read_a_hi(12),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(12),        -- Port B data input
DOB(0)   => data_read_b_hi(12),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_13_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10110A0441812402840402822007818000E00700000000330A3000000008042",
INIT_01 => X"A1400984B830C848180260000C0042404001000008220008A200100802110200",
INIT_02 => X"88010C02801040002475580400800000410000000064024608134C0CC9018034",
INIT_03 => X"00010100926220D084234212421085084300648A0880000630C0654288C10000",
INIT_04 => X"0004122122029100100C00001200009C40A83A2044360C84190BAC04E0101820",
INIT_05 => X"04E000008009050064C8C00104C10184034010250089C00EB004327064B60900",
INIT_06 => X"CA875CA8600000880410DA8C285001802424B008881024A8204E010461042700",
INIT_07 => X"08320014B02848A4A8100015C55500057801A04000712C040CB1F8806000088D",
INIT_08 => X"5005000908020220E40170008042000000557E048A144C800590010000882D00",
INIT_09 => X"00250104B5310020000100020821004016CC1C616401910801010100CA204000",
INIT_0A => X"0000000000010192072310200028B602234608080280074AC010025900100401",
INIT_0B => X"014100101118BA451000824150052110480121000140014200101352690BAC20",
INIT_0C => X"0000000040000000000000040000000000000020000000000000008010102A82",
INIT_0D => X"094040100000006C0802042501001C8017000C21908200028448400000000040",
INIT_0E => X"000000010C000C00081A08BC832A209AB0A85094284A14254A25510105130801",
INIT_0F => X"30BA901293C0F5012906A96DCD13042CE0C206E92DCD07042CE0C40D02048000",
INIT_10 => X"4CA4271CA2168ACB0E06E92DCD13042CE0C206A96DCD07042CE0C4408632C395",
INIT_11 => X"58408632C30D522CE80239CC2806AC44E954939AB299E000738F88296CA13B44",
INIT_12 => X"5145CD5306028F01990C080808494A64708B265CC4052B0F30302E060965EA00",
INIT_13 => X"51E0328A2CA9722094650CCAC0629112BA89C04A228568547B1654B9104A3286",
INIT_14 => X"A158BB80D4D8D48CB54012290470562EC29E44050B1DC60132282B68B9AA60C0",
INIT_15 => X"280000A5C11B9008FE2FA38F87804251CB0FAD40562EC0B426149D17E0044B10",
INIT_16 => X"509425094246A10A10441010090480C0964201800044109012001A000726E454",
INIT_17 => X"0942509425094250942509425094250942509425094250942509425094250942",
INIT_18 => X"9425094250942509425094250942509425094250942509425094250942509425",
INIT_19 => X"7E24502A80000000000000000005094250942509425094250942509425094250",
INIT_1A => X"AEBAEBAEBAEBAEBAFFD7F7F7F775555557DFBEEFBBFCFDF7DFFCF9F80089F7DF",
INIT_1B => X"BF5FAFD7EBF5FAFD7EBF5FAFD7EBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEB",
INIT_1C => X"FFFFFFFE0001DFAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7E",
INIT_1D => X"4500557DE00000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"E100004020BAAAFFD5400AAFBC2155AAAA97410FFFFEAAAAF7AA955EFF7803FF",
INIT_1F => X"5410F7AEBDE10FFFFFDEAAF7D568AAA5D002AB55005568B55087FC0010AAFBFF",
INIT_20 => X"555FF5D04154BAAAAEAAA10557BEAA10AAFBE8A00557BFFFEF007BC215500001",
INIT_21 => X"400000A2AABFF45550400000AAFBFFFEF550000155A28415410F7AEAABFFA2D1",
INIT_22 => X"D568AAAFFFBC21555D517FF45F7AEA8BFFA2AEAAA10A280021EF5D557FF55AA8",
INIT_23 => X"AAE974AAF7D142145082A975FF555568A00FF842ABEFA2AAA8B5500003DF55F7",
INIT_24 => X"000000145A2AA821EFFFFFD7410007FC0010555155555FF80174000055555EFA",
INIT_25 => X"2E3A0925C7E38E38F7D14557AE00000000000000000000000000000000000000",
INIT_26 => X"7D0075C7028B6F1FAE00000A02092B6F5D2438A2FBC2145B6A090428FFF5EAA9",
INIT_27 => X"FEF1C7FC516D080E15438E3A4BAE00FFF5FAE92F7D16AAAA41042FB7D145568B",
INIT_28 => X"2428FFA4AFBFFAAD1505FF490E174AABEA0ADA005D7BEDA00B6F1EFA28557BF8",
INIT_29 => X"001FF555F7FF7DAA8E07028B6A0BFF6D490E00000BEF5FAFEF490407155BE8E1",
INIT_2A => X"AAAB551C0E3AF55F7DF68ABAE3F1C0145415B78F45FFA4AFBC7BEA4AAA10A284",
INIT_2B => X"84104380055525FFBEAE90482E3D54216D0024975FF555F68A00F7842FBD7B6A",
INIT_2C => X"0000000000000000000000016DAAA0851FFE3FBD0438007FC00385D555556DEB",
INIT_2D => X"FF80020BAF7D16AA10A28402155A2AEA8BEF5D516AA000000000000000000000",
INIT_2E => X"A08003DFEF55516ABEF0055574BAFFD568A10002A82000FFD5400AAA2FBC0145",
INIT_2F => X"00F7D17FEBA557BEABEF557BD55EF082A974BAA28028A00F7D16AA10F7D56AAB",
INIT_30 => X"BEF000417545FFAA820BAFF843DFFFA2D5421FF002E954AAFF843DE105D7FFDE",
INIT_31 => X"DF55F7802AA10AA80001FF5D7FFDFEFA2AA974BAF7803FFFF002A82000FFD568",
INIT_32 => X"EAA10FF803DF45FFAEA8B555D2EAAB45F7FBE8ABAAAD540145007FE8B55FF843",
INIT_33 => X"FC20AA5D55555FFA280000BA0855401EFF7AA82010AAD1421FF0004155FF557F",
INIT_34 => X"00000000000000000000000000000000000000001EFA280175FFAAFFC00BA087",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"19FFFFFFFFE00000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(13),        -- Port A data input
DOA(0)   => data_read_a_hi(13),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(13),        -- Port B data input
DOB(0)   => data_read_b_hi(13),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_14_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10020A000180000284008280000281800000030000000033022000000580002",
INIT_01 => X"A140098018300848184860000C20C24040000000084000084200000000110200",
INIT_02 => X"88010C5A8010A600A4F558040080000041000000022C024008003CCCC9028030",
INIT_03 => X"000103A7A00904D0842242024210810803006480088000003081054288C10000",
INIT_04 => X"0000120122009000100C00000000000400A83A2044200C840000800400101820",
INIT_05 => X"040000008008010024C0C0010040000402000025000800020004207000100800",
INIT_06 => X"40870408600800800410D006A850018024240008881024A82040010461042000",
INIT_07 => X"08120054B42850B42A100010ED1500010001A040003164040CF5E20140000888",
INIT_08 => X"400500090A020220A40A7000800000000014FE8508144C924080C10000880140",
INIT_09 => X"0004010411110020000100020021004000800461600191080101000042200000",
INIT_0A => X"0000000000010190070310200008B202236D080802000002C010024000000000",
INIT_0B => X"0141001001088A45000082400000010040012100010000020000135249020820",
INIT_0C => X"0004000000000000004000000000000004000000000000000000008010100000",
INIT_0D => X"0840401000000044080200210100100017000420808200000440400000000040",
INIT_0E => X"0000000000000C00000000040302200800A04090204810244825010104130800",
INIT_0F => X"397468090008142014840100002C382800008401000038382800006402048000",
INIT_10 => X"83514072C000444C00840020002C38280000840020003838280002C09D010868",
INIT_11 => X"03C09D0104B01C57100440202900184414430534605E38048021800224804191",
INIT_12 => X"40049594C194000090450808802008830024F0E248C902AEF0024170CF180010",
INIT_13 => X"8000120020E5A08E6000048200196264BCF1C030C0604800001076C047300002",
INIT_14 => X"A00002003DEDE82C78900902A0D0000080019FAAA32D9602490302409292B832",
INIT_15 => X"2800D049100021171F6C34080240108AB292CA000000800AD1A19F6F000AA0C0",
INIT_16 => X"409024090246810810440000090480C096420080000010801001600001200454",
INIT_17 => X"0902409024090240902409024090240902409024090240902409024090240902",
INIT_18 => X"9024090240902409024090240902409024090240902409024090240902409024",
INIT_19 => X"6504002800000000000000000004090240902409024090240902409024090240",
INIT_1A => X"E79E79E79E79E79E7FDDF77777F3CF3CF7D55E6D39723FC3DEFA75D77B75F7DF",
INIT_1B => X"9FCFE7F3F9FCFE7F3F9FCFE7F3F9E79E79E79E79E79E79E79E79E79E79E79E79",
INIT_1C => X"FFFFFFFEFFFE0FE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F",
INIT_1D => X"55A28417400000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"AAAF7AA955EFF7803FF4500557DF45F7D16AB455D00001EFAAAAAAABA5555575",
INIT_1F => X"214555003FF450804001555D2AA8AAA002ABDE10082ABDF55AAAA97410FFFFEA",
INIT_20 => X"175EF5D5168A10082E80155087FC0010AAFBFFE100004020BAAAFFD5400AAFBC",
INIT_21 => X"EBDE10FFFFFDEAAF7D568AAA5D002AB55005568A00A2D5401455D00175FFFF84",
INIT_22 => X"7BC2155000015400AAD157545080402145087FD75FFF7AE82145A2D17FE10F7A",
INIT_23 => X"000000BAFFFBE8AAAA2FBFDE00087FD5410557BEAA10AAFBE8A00557BFFFEF00",
INIT_24 => X"000000155A28415410F7AEAABFFA2D1555FF5D04154BAAAAEAAA005D002AB450",
INIT_25 => X"7B6A0AAA82555157555B68012400000000000000000000000000000000000000",
INIT_26 => X"45B6A090428FFF5EAA92E3A0925C7E38E38F7D14557AF45FFDB6AB6D4100071C",
INIT_27 => X"092B6F5D2438A2FBC21455D0A3FF6D080407155552AAAA920020BFE10002EBAF",
INIT_28 => X"01454100175C7E380125D7555B6DA1014248217D0075C7028B6F1FAE00000A02",
INIT_29 => X"82145AAD178E38E3A4BAE00FFF5FAE92F7D16AAAA41042FB7D145568A38AADF4",
INIT_2A => X"1EFA28557BF8FEF1C7FC516D080E15400A2DB5754508040716D007BD05EFEBAA",
INIT_2B => X"A0ADA0055002AB6D0000020BAFFF1E8ABABEF1FAE001C7FD54005D7BEDA00B6F",
INIT_2C => X"00000000000000000000000155BE8E12428FFA4AFBFFAAD1505FF490E174AABE",
INIT_2D => X"F7FFEABFF080015555F78028A00555155555FF84000000000000000000000000",
INIT_2E => X"000003DE10082EAAB45FF80020BAF7D16AA10A28402155A2AEA8BEF5D516AB45",
INIT_2F => X"BAFFD568A10002A82000FFD5400AAA2FBC0145552ABFFFF000417555552EA8A1",
INIT_30 => X"FEF55516AABAAAFFC0145000417555A280001455D7FFDE105504021EF0055574",
INIT_31 => X"55FF007BC01FFAAAE80155AAD568ABAA28028A00F7D16AA10F7D56AABA08003D",
INIT_32 => X"D74105D7FFDE00F7D17FEBA557BEABEF557BD55EF082A97410AAFFD554508001",
INIT_33 => X"5421FF002E954AAFF843DE10550028BEF0004020BAF7D568AAAF7D168A105D7F",
INIT_34 => X"0000000000000000000000000000000000000000145FFAA820BAFF843DFFFA2D",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"01FFFFFFFFE00000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(14),        -- Port A data input
DOA(0)   => data_read_a_hi(14),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(14),        -- Port B data input
DOB(0)   => data_read_b_hi(14),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_15_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000A000000000284000280000001800020030000000033022000000180002",
INIT_01 => X"A140098018300848180060000C00424040000000080000080200000000110200",
INIT_02 => X"080108000010E60004E55800008000004100000000040240080000C009170016",
INIT_03 => X"0000000080000040842240000210810002000400888000003080014288C00000",
INIT_04 => X"0001100024A0800000440000000000040088322044200C840000011400151800",
INIT_05 => X"440002988000000020000000000B8094020000254C8800000514203000108800",
INIT_06 => X"00070000620040880410D00C285000802424000AA81024A80040010C01062001",
INIT_07 => X"086100043224489428100010811100010001A040003124040CAC600040000888",
INIT_08 => X"160500090A0282A06400100080C300000005BE0488104C800000010000880000",
INIT_09 => X"000581041110022000000002002100400080046140011008010100008A040000",
INIT_0A => X"0000000000010180060210200008B2022304080800000007C010024000000000",
INIT_0B => X"4140001001088A45000082000000010000002000010000020000034249000020",
INIT_0C => X"0004000040000400000000000000000004000020000200000000008010100000",
INIT_0D => X"094000100000004C000200250000188016000400000000000440400000000040",
INIT_0E => X"0000000108000C00000000000200200800800000000000004020000000000000",
INIT_0F => X"0000000000000000000404200000000000000404200000000000008C00048000",
INIT_10 => X"4000000000000000000405000000000000000405000000000000004000001000",
INIT_11 => X"0040000010000000000000000000004000201000000000000000000000800002",
INIT_12 => X"0004000110000000000C00080010180000000001A10240500000000000000000",
INIT_13 => X"0000000020080400000000020000008040020000000000000010001200000000",
INIT_14 => X"0000020000000611002800000000000080000011044220000000000080200200",
INIT_15 => X"8800000100000000009080E2E0A0000000000000000080000040000000000000",
INIT_16 => X"0000000000460000004400000904808094020080000010000000000000000041",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0004002800000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000004000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFE00000000000000000000000000000000000000000000000000000000",
INIT_1D => X"EF08517DE00000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"1EFAAAAAAABA555557555A284175FF000002010552A97400007BFDE10A2AA801",
INIT_1F => X"DFEF5D2AAAB45F7D17DF45087BC0155002A801FF08003DF45F7D16AB455D0000",
INIT_20 => X"C2145F7D568BEFAAD557555AAAA97410FFFFEAAAAF7AA955EFF7803FF4500557",
INIT_21 => X"03FF450804001555D2AA8AAA002ABDE10082ABDFFFF7D17FE10002E954AAF7FB",
INIT_22 => X"FFD5400AAFBC21EFA2AE95545A2D56ABFFAAD17DE10FFD1420AA007FC0145550",
INIT_23 => X"02A801550055401555D00174BA002AA8B55087FC0010AAFBFFE100004020BAAA",
INIT_24 => X"000000000A2D5401455D00175FFFF84175EF5D5168A10082E801FFFF8428A100",
INIT_25 => X"80871FAE00A2A0871EF145B7FE00000000000000000000000000000000000000",
INIT_26 => X"45FFDB6AB6D4100071C7B6A0AAA82555157555B680125C71C0E0500049209543",
INIT_27 => X"5C7E38E38F7D14557AFC75524AFB45FFD178F7D1C71C2145002E801C7140A3FF",
INIT_28 => X"AE000024954AAFFFBC2145F7DB6DBEFA2D557545B6A090428FFF5EAA92E3A092",
INIT_29 => X"470820071C71455D0A3FF6D080407155552AAAA920020BFE10002EBAFC7FFDF7",
INIT_2A => X"1FAE00000A02092B6F5D2438A2FBC21FFBEA090545B6D568BFFAADB7AE10F7D5",
INIT_2B => X"24821FFE3802FA2808208017D1C5142155410A104AA1420AFB7D0075C7028B6F",
INIT_2C => X"00000000000000000000000038AADF401454100175C7E380125D7555B6DA1014",
INIT_2D => X"552E954100004174AA00516AA10AA80155EF5D7BFDE000000000000000000000",
INIT_2E => X"5082E801555D2EBDF45F7FFEABFF080015555F78028A00555155555FF8400155",
INIT_2F => X"BAF7D16AA10A28402155A2AEA8BEF5D516AB555D043DF55F7D56ABEF55514015",
INIT_30 => X"E10082EAAB55FFFBE8A100804154AAF7FFC2145FFFFFDFEFAAD157545FF80020",
INIT_31 => X"ABEFA2FBE8A00FFD155410005555545552ABFFFF000417555552EA8A1000003D",
INIT_32 => X"3DFEF0055574BAFFD568A10002A82000FFD5400AAA2FBC01FFF78400155F7D16",
INIT_33 => X"0001455D7FFDE105504021FFAA843DEBA0000021EF555142155002E800AA5500",
INIT_34 => X"00000000000000000000000000000000000000000BAAAFFC0145000417555A28",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"1800000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(15),        -- Port A data input
DOA(0)   => data_read_a_hi(15),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(15),        -- Port B data input
DOB(0)   => data_read_b_hi(15),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_16_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"DA22C618B1000482B688B186588884862A400438255FC38381441205BA803003",
INIT_01 => X"8645A80028404C211203A952A90341080B173340412000E1005D628000820484",
INIT_02 => X"A101A9006DC1084833011850AAC55001349B10881802821808B4110007005E11",
INIT_03 => X"010108A802BB00080080006020020001A61036202800000D2410104200404550",
INIT_04 => X"8BFA58800005C40A46240252145148B38248030356415A4E62B6FC660F287240",
INIT_05 => X"1E0BD423CAC0000D610000000710296E542B6E3A825C15FB30A643695BFC2D56",
INIT_06 => X"000D0000C8008820CAE16020619156A5815006028179808C00A0D2152B90707A",
INIT_07 => X"F500240510A00205F0A407D0021A155378900002A002433A0AA00EE6E7956108",
INIT_08 => X"015995440C8327241440096A2800002828123D542910380004E0310362404076",
INIT_09 => X"10222D90409A05B2CB2CA400200209E5601044A24000000462A6001888010000",
INIT_0A => X"0000000000259200140001A15000017F0051D0F837248C005514AC40C0820500",
INIT_0B => X"01200848002912300200092BA80325A2000000000001514B5500030241C000CC",
INIT_0C => X"0001100011000110001100011000110001080008800080005202280801080395",
INIT_0D => X"17680002815014B90000205DA00880100095A64800008003561180063DB4F611",
INIT_0E => X"0280080922554515512174000000490009000000000000004010042A204A0C58",
INIT_0F => X"2DA0063EAA9C238B2D4C800632B266E828EE4C800632AAAB6830D0FC6B06C041",
INIT_10 => X"0839AA149339E8FB964C800632B266E82B2E4C800632AAAB683310872800EDA5",
INIT_11 => X"C087A800EB090D4AAC91268FFCBE81397826C4A20D2B6C510E8624792A4A30A4",
INIT_12 => X"3638E8849D5C532408DD6E004C90C06AC019D88B9795012CA96902C799912BC3",
INIT_13 => X"78706531C74485BD42A30906057FADAA456218FD8E3ED83B60E3A242DC0F1898",
INIT_14 => X"51727A06FB555793057C444CF45C5C9E89543B8BC6E80193DC36F6C71D1093A4",
INIT_15 => X"10DCD45DC02B331650CA8ACB4007E00D1C6A6A58395C917F7E74D936F650D69B",
INIT_16 => X"000000000012000081500008A422150884081ACAAC0542054004FC5884640508",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"3604000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"45145145145145147A7797E1E1A79E79E15634455131A436993071A616D4F68A",
INIT_1B => X"3E9F4FA7D1E9F47A7D1E9F47A7D3453453453453453453453453453453453453",
INIT_1C => X"FFFFFFFE00001F4FA7D3E9F4FA3D1E8F47A3D1E8F47A3D1E9F4FA7D3E9F4FA7D",
INIT_1D => X"00FF8015400000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"400007BFDE10A2AA801EF08517DE10FFFFFDFEFA2D16AB55A2FFFFEAA5D7FC00",
INIT_1F => X"74BA5D2EBDFEFAAD17FFFF002EBDE000800174AA55043FFFF000002010552A97",
INIT_20 => X"E8AAAAA80000105D557FF45F7D16AB455D00001EFAAAAAAABA555557555A2841",
INIT_21 => X"AAAB45F7D17DF45087BC0155002A801FF08003DE000004154BA002A800BA087F",
INIT_22 => X"803FF4500557DEAAF7D57DEBA082A82010FFAE975555D7FFDEAAFF80155EF5D2",
INIT_23 => X"2D57FFFF557FD55FF08003FE0055043FF55AAAA97410FFFFEAAAAF7AA955EFF7",
INIT_24 => X"0000001FFF7D17FE10002E954AAF7FBC2145F7D568BEFAAD557410552EA8BEFA",
INIT_25 => X"DB6FFFDEAA5571C7010FF8412400000000000000000000000000000000000000",
INIT_26 => X"C71C0E050004920954380871FAE00A2A0871EF145B7FE10E3F1F8FC7AAD56DB7",
INIT_27 => X"A82555157555B680124924124BDFEFA2D57FFC71C2EBDE280000174825D0E3FF",
INIT_28 => X"74821424800AA007FEDAAAA284020385D5F7AF45FFDB6AB6D4100071C7B6A0AA",
INIT_29 => X"F8EAAFF80175C75524AFB45FFD178F7D1C71C2145002E801C7140A3FE10080A1",
INIT_2A => X"5EAA92E3A0925C7E38E38F7D14557AE92EBDB78EAA1C2482010FFAE9556D557F",
INIT_2B => X"D557410492EADBEFA2D178FEF5575D55EF000A38E10490A3AF45B6A090428FFF",
INIT_2C => X"000000000000000000000001C7FFDF7AE000024954AAFFFBC2145F7DB6DBEFA2",
INIT_2D => X"A2D56AB45A2D57DFFFF7FBFFEAA555555400F780000000000000000000000000",
INIT_2E => X"A080415400552ABDF55552E954100004174AA00516AA10AA80155EF5D7BFDE10",
INIT_2F => X"FF080015555F78028A00555155555FF840000000043DFEFAAD17FF45552ABFEB",
INIT_30 => X"1555D2EBDE10002E974005D04020BA007BFDEBAA284000BA557FE8B45F7FFEAB",
INIT_31 => X"0000F7AE955EF5D7BE8ABAF784175555D043DF55F7D56ABEF555140155082E80",
INIT_32 => X"AAB45FF80020BAF7D16AA10A28402155A2AEA8BEF5D516AA00AAFBE8AAA55040",
INIT_33 => X"FC2145FFFFFDFEFAAD157410082ABFFEFAAD16ABFF5555575FF082AA8A00002A",
INIT_34 => X"0000000000000000000000000000000000000000155FFFBE8A100804154AAF7F",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0800000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(16),        -- Port A data input
DOA(0)   => data_read_a_hi(16),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(16),        -- Port B data input
DOB(0)   => data_read_b_hi(16),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_17_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"5284CE4FB7BD2C8994A13392DBD02E14006B82AC7E800D44D3DD2FD5F9B961C0",
INIT_01 => X"F8ACD01F7E03FC6793F2199B39FC233C11D93AE6F3BB92B32091DBC339B24542",
INIT_02 => X"8F333007FD6808092A2AFA6667033DB50853379C10BFF70F1BD011110F205F18",
INIT_03 => X"294ADB4AFFCBF0DAD63ABF836B58EAFE060478202022234B2E0303FDC9E18339",
INIT_04 => X"DB7A40806FE4040840EBC563A0150A0926146FECB04196482236FC2005282AE1",
INIT_05 => X"0807B4070670083DC68206D7E6D0250834336D1E81500FDB306045255BFC2076",
INIT_06 => X"00000000141C5AF3EA6AB187F7F8CE039786062C6CE092F5FE005236781C402A",
INIT_07 => X"1684248A38B022475DCA9BD00116E33CC3821774BB55F53BB42329AA3C0CEF60",
INIT_08 => X"60700CE0641527241060AD844E1C0088001223022D189A2800542219204903F8",
INIT_09 => X"D94C1C1C51DFF881861CBE0305A12A0321810217C01D34EDC98FFA1C8E000016",
INIT_0A => X"7E7D8F8FBDE40E001E000B3A5DAADAFDDA5DA79350DF70027CE86F047BEF19B6",
INIT_0B => X"814102F800633F1D0A7CC9AE74117FE0003A6AD055819D1F9984014B37BA5FFC",
INIT_0C => X"CF4FBCF4FBCF4FBCF4FBCF4FBCF4FBCF4FBE7A7DE7A7800617112E46F05D02DD",
INIT_0D => X"D7FE4A5A99FD6D3FEF4BEB5FF994F0FEFFCCF8430006CE8A3F06ABD73DBCF4FB",
INIT_0E => X"B29760593F33FA0CF170F40006001B1A05C0000000000000008004BA78428C7A",
INIT_0F => X"EDA57E46444357B3950A9BFBAC94CFA8581E0A9BFBAC8CCFA8580C7CAF51EF68",
INIT_10 => X"7DF76B5DB54A09003E0A9BFBAC94CFA8581E0A9BFBAC8CCFA8580E46FBFCB0CB",
INIT_11 => X"E7467BFCB1D5CFEB56A1A100D5345C1BFFE8FBDB892DB463034198E2881F3F78",
INIT_12 => X"4E0ADD39387F92B2935DFEAADDF38EBCFB9E3D636DCDF9B90F966BF92966D5D9",
INIT_13 => X"F256527055EB6D555CB294981B7FB5B2954CD3013013FDF5E82AF5B6AAAE594A",
INIT_14 => X"F7D7E835C67E655BAA868610117575EA1C34BD6975D48B44A0405FC15BA7270F",
INIT_15 => X"BD07F6CD2A47D0CBA96252756D7217E5E1C61DBDF5FA167F7AE5D3D21A414007",
INIT_16 => X"00000000005F08000179C16DECF67F08BC02F9067ED55805600545DFE45A80E7",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"F981800C00000000000000000000000000000000000000000000000000000000",
INIT_1A => X"A69A69A69A69A69A919261A1A6075D75D10DC800C027B731014BA4B864617114",
INIT_1B => X"8341A0D068351A8D068351A8D069A6BAE9A69A6BAE9A6BAE9A69A6BAE9A6BAE9",
INIT_1C => X"FFFFFFFE000011A8D46A351A8D46A351A8D46A351A8D46A341A0D068341A0D06",
INIT_1D => X"55AAFFD5400000000000000000000000000000000000000000000001FFFFFFFF",
INIT_1E => X"B55A2FFFFEAA5D7FC0000FF8015410FFFFFFFFFFFFFFDFEFF7D568A1008003DF",
INIT_1F => X"DF55A2D1400000804154BAF7D168A00A2803DE10FFAE95410FFFFFDFEFA2D16A",
INIT_20 => X"2AABAFFD56ABFF002EBDFFF000002010552A97400007BFDE10A2AA801EF08517",
INIT_21 => X"EBDFEFAAD17FFFF002EBDE000800174AA55043FEBA0004174AA5504000AA5504",
INIT_22 => X"5557555A284175FFFFFBE8B55A2FFFFF55F7803DEBA002AAAAAAF7FBD74BA5D2",
INIT_23 => X"D0417400FFD57DE00AAAAAAB45A2AA97545F7D16AB455D00001EFAAAAAAABA55",
INIT_24 => X"0000000000004154BA002A800BA087FE8AAAAA80000105D557FE00A2D5420AA5",
INIT_25 => X"7EBD16AA00000E3DF6DBEF5D2400000000000000000000000000000000000000",
INIT_26 => X"10E3F1F8FC7AAD56DB7DB6FFFDEAA5571C7010FF8412428FFFFFFFFFF7FBF8FD",
INIT_27 => X"E00A2A0871EF145B7FF7DA2D547038140E10492FFDF6DA28A28E3DE00F7A0924",
INIT_28 => X"2492550A020BA55002AA82F7DF6DBD71C2EBFFC71C0E050004920954380871FA",
INIT_29 => X"ADABAF7F5D74924124BDFEFA2D57FFC71C2EBDE280000174825D0E3FEAA14001",
INIT_2A => X"0071C7B6A0AAA82555157555B680125FFEBFFEDB55BEFFFAF6DE38E3DEAA002E",
INIT_2B => X"5F7AE28B6D545092490E10400FFDB7AE00A2AAADB45BEA092545FFDB6AB6D410",
INIT_2C => X"00000000000000000000000010080A174821424800AA007FEDAAAA284020385D",
INIT_2D => X"FFFBFDFEFF7FFEAB45A2D56AA00002EBDFFFF7D5400000000000000000000000",
INIT_2E => X"AA2AABDE10FF8400010A2D56AB45A2D57DFFFF7FBFFEAA555555400F780000AA",
INIT_2F => X"100004174AA00516AA10AA80155EF5D7BFDFEFAAD1554BA552E82000F7FFFFEA",
INIT_30 => X"400552ABDEBA5D0002000552A800BA55042AA10FFFFFDF55552EBDF55552E954",
INIT_31 => X"ABFFA2AEBFEAA082EBDEBAFFD55540000043DFEFAAD17FF45552ABFEBA080415",
INIT_32 => X"00145F7FFEABFF080015555F78028A00555155555FF84001FFAAFBFFF55FFFBE",
INIT_33 => X"BFDEBAA284000BA557FE8AAAFFD155400082A82000F7FFE8A00A2AABDF45F780",
INIT_34 => X"0000000000000000000000000000000000000000010002E974005D04020BA007",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"19FFFFFFFFE00000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(17),        -- Port A data input
DOA(0)   => data_read_a_hi(17),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(17),        -- Port B data input
DOB(0)   => data_read_b_hi(17),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_18_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"69844019080000A21A611406840014122A641074155FC28A2024001001801003",
INIT_01 => X"A643D920034004180005E9E3C90360C0041C0181002001602025800008440084",
INIT_02 => X"B7333980808408103F2000F81FC0FEDEAC2161B0B84D0002188011110C018041",
INIT_03 => X"0405D434003F2C020081587008020561E55116B0290000042B71240C800440F8",
INIT_04 => X"50805AC31007D6125724029216554A9847669903D640EC8E2001002604503004",
INIT_05 => X"0E010001C1CA11803850C800010022660C1C0065003C0404002646DC20A02D40",
INIT_06 => X"50AD050AC00000002A4F612449903FE080000000005889AC41E04508A9907020",
INIT_07 => X"5584280B10014003A8067400920810FF3C72024300A0030048221ACEE383E518",
INIT_08 => X"00C983E6041505253500F66E620428000B1804000152E52801A2020084090040",
INIT_09 => X"20500B90419005B0C309402030060860E01004A828408800440405E350294010",
INIT_0A => X"008010100007865421432121804021C20452880C2D200000045C18C0E0000A08",
INIT_0B => X"09700C04C44C92A88DC42215C882E82250811000000C1AE061861710A401A4E8",
INIT_0C => X"308003080030800308003080030800308001840018400400602A018809800371",
INIT_0D => X"0801010202021000780004200408C1002003F66CA1B13111C0D95C20C2030A00",
INIT_0E => X"02900806400FC503F08180050942E4200020C1B060D8306C182701404C197301",
INIT_0F => X"22AABABAF377DF1CA160820520EB3057E70E60820520F33057E72E9154159000",
INIT_10 => X"8A2AD5D48F37FAFEFE60820520EB3057E7CE60820520F33057E7EC658BF2DA78",
INIT_11 => X"32658BF2D4B2A80BF8FE39FD78EB0D882014A62C568FFAFC73FFDD9C2B30E046",
INIT_12 => X"C728C800DFC06F59F710107533C0C4E37619440FBFBAB2400AFC1600361D798F",
INIT_13 => X"0DEBBEB9454005BAA36DEFF894823A3D1A88A2FE29D5FC6DCAA2A002DD51B6E7",
INIT_14 => X"F3B7092A78606A28A5427AAB9FF4EDD251C7123E291660733EBF6FE519001BF4",
INIT_15 => X"82202AB58AFBFD5DE200A8EBE3A3EC110339E1DCEDC2590495BB2112E2BE4BF5",
INIT_16 => X"C1B06C1B06808348340000020301805002D008C1F92000A5F421B8000DB49103",
INIT_17 => X"1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06",
INIT_18 => X"B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C",
INIT_19 => X"16000000000000000000000000041B06C1B06C1B06C1B06C1B06C1B06C1B06C1",
INIT_1A => X"A28A28A28A28A28A244C16454170410412CA2EFB3AE03B85CF08C03F1A30F7DF",
INIT_1B => X"8944A25128954AA552A944A2512AAA8A28A28A2AAAAAA8A28A28A2AAAAAA8A28",
INIT_1C => X"FFFFFFFE000004A25128944A25128944A25128944A25128944A25128944A2512",
INIT_1D => X"105D2A80000000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"FEFF7D568A1008003DF55AAFFD5410FFFFFFFFFFFFFFFFFFFFFBFDEBA552E974",
INIT_1F => X"5410FFFFFFFFFF7FBE8B55AAD16AA1000516AA005D0400010FFFFFFFFFFFFFFD",
INIT_20 => X"FFE00087BC2155087BC0010FFFFFDFEFA2D16AB55A2FFFFEAA5D7FC0000FF801",
INIT_21 => X"1400000804154BAF7D168A00A2803DE10FFAE95555FFFBE8B45A2D56ABEFFFFF",
INIT_22 => X"AA801EF08517DF55000000010082A974AA08557DEBAFFAEBFF55AA8028B55A2D",
INIT_23 => X"52E800105D2AAAA10A2D1420AAFFAEA8BFF000002010552A97400007BFDE10A2",
INIT_24 => X"0000000BA0004174AA5504000AA55042AABAFFD56ABFF002EBDEBA0004020BA5",
INIT_25 => X"FF7FBFFEBA552A95410552485000000000000000000000000000000000000000",
INIT_26 => X"28FFFFFFFFFF7FBF8FD7EBD16AA00000E3DF6DBEF5D2438FFFFFFFFFFFFFFFFE",
INIT_27 => X"EAA5571C7010FF8412410FFFBF8FC7E3F5EAB45BEDB6FA3800556FA005504050",
INIT_28 => X"AB55BEDB6FBC7EBF5F8E10007BC516D1C71C5010E3F1F8FC7AAD56DB7DB6FFFD",
INIT_29 => X"BFF55BE8A2DB7DA2D547038140E10492FFDF6DA28A28E3DE00F7A09256DE3F1E",
INIT_2A => X"0954380871FAE00A2A0871EF145B7FF45080E070280820924AA145578E92F7A4",
INIT_2B => X"2EBFEBA1C0A00092412E850005D2AAFA38A2DF45082F7AAA8BC71C0E05000492",
INIT_2C => X"000000000000000000000000AA140012492550A020BA55002AA82F7DF6DBD71C",
INIT_2D => X"FFFFFFFFFFFFBFDFEFF7FFFDEAA5D2E954105504154000000000000000000000",
INIT_2E => X"A08557DE005500154AAFFFBFDFEFF7FFEAB45A2D56AA00002EBDFFFF7D5400AA",
INIT_2F => X"45A2D57DFFFF7FBFFEAA555555400F78000010F7FBE8B55AAD16AB55F7FBFDEA",
INIT_30 => X"E10FF84001FFAAD568B45FFFBFFF55A2D568A00087BD55FF5D5555410A2D56AB",
INIT_31 => X"00AA555168A10FF803DF45FFAABDFEFAAD1554BA552E82000F7FFFFEAAA2AABD",
INIT_32 => X"A8B55552E954100004174AA00516AA10AA80155EF5D7BFDF45002A974AA08000",
INIT_33 => X"42AA10FFFFFDF55552EBDEBA5D2E80010082A97410552EBDEBAA2FBD5400F7AA",
INIT_34 => X"00000000000000000000000000000000000000000BA5D0002000552A800BA550",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0800000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(18),        -- Port A data input
DOA(0)   => data_read_a_hi(18),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(18),        -- Port B data input
DOB(0)   => data_read_b_hi(18),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_19_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"042200000000000041088001001AA00000000000000000000000500802000003",
INIT_01 => X"200048000024000000000404000000000A22000800000800004A200000000001",
INIT_02 => X"032210008DEF00400060000001C008002489E0F0004037B00010101010000000",
INIT_03 => X"0000008128000000000000000000000024001620280000000000354200004008",
INIT_04 => X"000058800004C4024024001210001054B1C822009640000E2000002604003000",
INIT_05 => X"0E010001C0400000000000000000200604000000001C04000026400000002C40",
INIT_06 => X"000000000000000001800166A84004A080000000005884020020400009907020",
INIT_07 => X"E200201C00A14080082B26208008A00900120101402240440280040840802000",
INIT_08 => X"004180261C81210031000004340000200008105428020568040213003499C006",
INIT_09 => X"00000990000000B0C30800000000086020016000000000003838000000000000",
INIT_0A => X"000000000005860000000080A000206020408000000000000454080000000000",
INIT_0B => X"00000000000040002000044000000000000000000005E0003E00004049640004",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"00000000210001D8000000000000000020009640000000000000000000000000",
INIT_0E => X"040000000000C500300080000000000000000000000000000000000000000000",
INIT_0F => X"50500101088A37034E156600D740022800EC156600D740022800D01E0412D069",
INIT_10 => X"E61700224081044914156600D7400228002C156600D7400228001098F00D0FB7",
INIT_11 => X"CC98F00D0F2DD014010046037814EA63DBB31CE7605001008C41A061F0E7D693",
INIT_12 => X"361526D600000004089E12350C0E01FF23315422BABB46FEF5019146C0800380",
INIT_13 => X"00000130AA3592000000000629C03F3E60330C00C628908214551AC900000010",
INIT_14 => X"4208D65C006070845039014460088235ACC3123E2A29148841008482A4DAC000",
INIT_15 => X"6CD4953A66BE7A5040018D8A8AD9090A1EC20A188235AC509FB50C2D0500B409",
INIT_16 => X"00000000000000000000000000000000000008C0180027000006110008404608",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"9200000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"61861861861861861A2882313054D34D301C822EE8FC31C043198028002C7441",
INIT_1B => X"84C261349A4C26130984C261309861861861A69861861861861A698618618618",
INIT_1C => X"FFFFFFFE0000026130984C26130984C26130984C26130984C26130984C261309",
INIT_1D => X"00082E97400000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"FFFFFFBFDEBA552E974105D2A801EFFFFFFFFFFFFFFFFFFFFFFFFFEAA552E954",
INIT_1F => X"55EFFFFFFFFFFFFFFFFFEFF7FBFFEAA5D2E97545FFFFC2010FFFFFFFFFFFFFFF",
INIT_20 => X"6AA0008003DF555D5157410FFFFFFFFFFFFFFDFEFF7D568A1008003DF55AAFFD",
INIT_21 => X"FFFFFFF7FBE8B55AAD16AA1000516AA005D04001EFFFFFFFFFFFFFBFDF45AAD1",
INIT_22 => X"7FC0000FF80155EFFFFFFFFEFF7D16AB55A2D57DEBA557FEAA10080402010FFF",
INIT_23 => X"2D56AB45FFFBFDEBA5D7FC0155FFFFD7410FFFFFDFEFA2D16AB55A2FFFFEAA5D",
INIT_24 => X"000000155FFFBE8B45A2D56ABEFFFFFFFE00087BC2155087BC00AAFFFBFDF45A",
INIT_25 => X"FFFFFFDEAA552E95400002095400000000000000000000000000000000000000",
INIT_26 => X"38FFFFFFFFFFFFFFFFEFF7FBFFEBA552A954105524851C7FFFFFFFFFFFFFFFFF",
INIT_27 => X"A00000E3DF6DBEF5D25D7FFFFFFFFFFFFBFDFEFEBF5F8E92552E9556DEBF1C20",
INIT_28 => X"DFEFE3F1FAF55A2D568A0000003FF7D495155428FFFFFFFFFF7FBF8FD7EBD16A",
INIT_29 => X"EFA00000002010FFFBF8FC7E3F5EAB45BEDB6FA3800556FA005504051FFFFFFF",
INIT_2A => X"56DB7DB6FFFDEAA5571C7010FF84125EFF7F1F8FC7EBD568B6DBEDF7DEBA5571",
INIT_2B => X"71C5092E3F1F8F55AADB6DB7DEBF1FAE82557FC516DEBF1D0410E3F1F8FC7AAD",
INIT_2C => X"0000000000000000000000016DE3F1EAB55BEDB6FBC7EBF5F8E10007BC516D1C",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFBFDEAA5D2A954000800154000000000000000000000",
INIT_2E => X"0552A955EFAAD1400AAFFFFFFFFFFFFBFDFEFF7FFFDEAA5D2E95410550415545",
INIT_2F => X"EFF7FFEAB45A2D56AA00002EBDFFFF7D540145FFFFFFFEFF7FBFFFFFAAD16AA0",
INIT_30 => X"E005500155EFF7FBFDFEFAAD568B55AAD568A0008003DFFF0855554AAFFFBFDF",
INIT_31 => X"ABEFFFFFFFEAA55517DE10080400010F7FBE8B55AAD16AB55F7FBFDEAA08557D",
INIT_32 => X"40010A2D56AB45A2D57DFFFF7FBFFEAA555555400F780001FFF7D16AB55A2D16",
INIT_33 => X"568A00087BD55FF5D5555410AAD56AB45AAFFFFFEFAAD168A00557BD55FFA2D5",
INIT_34 => X"00000000000000000000000000000000000000001FFAAD568B45FFFBFFF55A2D",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"1000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(19),        -- Port A data input
DOA(0)   => data_read_a_hi(19),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(19),        -- Port B data input
DOB(0)   => data_read_b_hi(19),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_20_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000003",
INIT_01 => X"A75FF80000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"14088080800008400F655001FFCFF80018FA8044000000000000011000000007",
INIT_03 => X"0000000000000000000000000000000024001660380000000000000000004FF8",
INIT_04 => X"000079800014CC02C034001600000000000000101EC0012EE0C0026E1E80F000",
INIT_05 => X"3E1FE867DFC044003902100002203F2EFC040388137C3E20C8EEC00284033CC0",
INIT_06 => X"001F0001E0020002E80020000005FEAF91D10802ABFB80000021C8010FB0F0F4",
INIT_07 => X"00040007700000000000000001080FF900160000000200C00080001840BFE538",
INIT_08 => X"09FFBFE5181606000410A4000004202AA8043E0000000000000001209244C040",
INIT_09 => X"01227FB0000000F7DF78020004011FEFE0000000002003150200008388020000",
INIT_0A => X"000000000015BE0000004000000100000100506002008C2007D5FC8000002400",
INIT_0B => X"0000000000000000000000000000000400400520000000000000000400000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000020002",
INIT_0D => X"00010000000200000020000004000100203FF6C0000000000000000000000000",
INIT_0E => X"0000000600FFC53FF001800000002004080000000000000040900005C8485380",
INIT_0F => X"8000000009A9C300020080000800000003CC0080000800000003CC0200078000",
INIT_10 => X"00800000000012963C0080000800000003CC0080000800000003CC1008000000",
INIT_11 => X"00100800004000000000066C5000020020000000800000000C2E180010002000",
INIT_12 => X"96004000000000052B0200000014200040C2829000400000000000860F987980",
INIT_13 => X"0000A4B00400000000002958000240400000000007E1B0000402000000000014",
INIT_14 => X"400004004181800000000005C5A00000200C40808000000000AF0D8008000000",
INIT_15 => X"000800020141812737DC3020100400001C19C1D80000200400000000000015D1",
INIT_16 => X"0000004010080800801810100000000000093EDFF80200000000000010010010",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"4D20400200000000000000000000000000000000000000000000000000000000",
INIT_1A => X"CB0C30C30C30C30C8192608486879E79E681C000C00E08000402241560412010",
INIT_1B => X"2190C86432190C86432190C86432CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2",
INIT_1C => X"FFFFFFFE000010C86432190C86432190C86432190C86432190C86432190C8643",
INIT_1D => X"10080402000000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"FFFFFFFFFEAA552E95400082E975FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2A954",
INIT_1F => X"0000FFFFFFFFFFFFFFFFFFFFFFFDEAA5D2A954000800001EFFFFFFFFFFFFFFFF",
INIT_20 => X"FFEBA5D2A97400FF8017410FFFFFFFFFFFFFFFFFFFFFBFDEBA552E974105D2A8",
INIT_21 => X"FFFFFFFFFFFFFEFF7FBFFEAA5D2E97545FFFFC21FFFFFFFFFFFFFFFFFFFFF7FB",
INIT_22 => X"003DF55AAFFD5400FFFFFFFFFFFFFFDFEFF7FFEAA10000417555AAD5555EFFFF",
INIT_23 => X"FFBFDFEFAAD568A0000043DF45AAFBC2010FFFFFFFFFFFFFFDFEFF7D568A1008",
INIT_24 => X"0000001EFFFFFFFFFFFFFBFDF45AAD16AA0008003DF555D51574BAFFFFFFFFFF",
INIT_25 => X"FFFFFFFEBA5D2A95410000A00000000000000000000000000000000000000000",
INIT_26 => X"C7FFFFFFFFFFFFFFFFFFFFFFFDEAA552E954000020955FFFFFFFFFFFFFFFFFFF",
INIT_27 => X"EBA552A95410552485010FFFFFFFFFFFFFFFFFFF7FBFDEBA5D2E95400140E001",
INIT_28 => X"FFFFFFFFFDFEFF7FFFFEAA5D2E95400E38A17438FFFFFFFFFFFFFFFFEFF7FBFF",
INIT_29 => X"1557DBEDF575D7FFFFFFFFFFFFBFDFEFEBF5F8E92552E9556DEBF1C21C7FFFFF",
INIT_2A => X"BF8FD7EBD16AA00000E3DF6DBEF5D2438FFFFFFFFFF7FBFDFC7EBF1E8A00080A",
INIT_2B => X"5155492FFFFFFFEFF7F1F8FD7A2D168A1008043FF6DAAFBC5028FFFFFFFFFF7F",
INIT_2C => X"000000000000000000000001FFFFFFFDFEFE3F1FAF55A2D568A0000003FF7D49",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFEBA552A95410002E820000000000000000000000",
INIT_2E => X"A552E954005D2A82145FFFFFFFFFFFFFFFFFFFFFBFDEAA5D2A954000800155FF",
INIT_2F => X"FFFFFBFDFEFF7FFFDEAA5D2E95410550415410FFFFFFFFFFFFFFDFEFF7FBFFEB",
INIT_30 => X"5EFAAD140155FFFFFFFFFF7FBFDFFFFFFBFDEBA5D2A95400A2AA974AAFFFFFFF",
INIT_31 => X"FF55A2D568A10082E955FFFFFFD7545FFFFFFFEFF7FBFFFFFAAD16AA00552A95",
INIT_32 => X"D74AAFFFBFDFEFF7FFEAB45A2D56AA00002EBDFFFF7D5400BAFFFFFDFEFF7FBF",
INIT_33 => X"568A0008003DFFF085555410F7FBFDFEFFFD568B45AAD16AA1008003DFEFAAFB",
INIT_34 => X"00000000000000000000000000000000000000001EFF7FBFDFEFAAD568B55AAD",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"01FFFFFFFFE00000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(20),        -- Port A data input
DOA(0)   => data_read_a_hi(20),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(20),        -- Port B data input
DOB(0)   => data_read_b_hi(20),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_21_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"4A302428B824900A128C090A5C1800261500213C005FE812D10420054085A202",
INIT_01 => X"081FFE3440B609703B0427F801A40B8115BC4F655300340288A40D30040E4DD8",
INIT_02 => X"0109095C30C98809800000F9FFFFFFFF149FF1FCA4C0421B182E3490DF145FE4",
INIT_03 => X"084A76341244919000099486400026523C041660BA000100CC12701015007FF8",
INIT_04 => X"000079800014CC03C075161E001118653D2408041FC004AEF000816E1C11F541",
INIT_05 => X"7E1F00F7FFC000240100004683103E7FFE02482553FC3C0204EFC25010143CC0",
INIT_06 => X"801008011010421960E339A20205FEBF8140000203FFC806C8A1C1048FF0F0E0",
INIT_07 => X"750504800680102542AD800504530FF9061E8026998E9A00402CC25BD0FFF800",
INIT_08 => X"11FBFFE04691A5A00101818A6800088228000001A044C8168480D010F200AA08",
INIT_09 => X"E85A7FF080AC70FFDF78220010841EFFE7116E144071268DFD3E4C2404010000",
INIT_0A => X"54518A8A31B7FE00040009814C089202225412115428C03BC7D7FC15025B1AB6",
INIT_0B => X"88300E20806520398C682157A493896600E24E10100DFF22FF86002020ED110C",
INIT_0C => X"28D9228D9228D9228D9228D9228D9228D99146C9146C84006309044081A001B1",
INIT_0D => X"890000403000A01282088624001201A8C43FF7C0011529904595123203040D92",
INIT_0E => X"06102C4053FFD5BFF00A04A00200602CA5200110008800444021048034004001",
INIT_0F => X"2A00263009140094D81A5040605800B506901A30406054013605620272181965",
INIT_10 => X"890A202811209062801A3040605800B506901A50406054013605604350B81282",
INIT_11 => X"3F4350B811068C00049A0A5820A3C1725A8006C0A40404D058320496C2C9C600",
INIT_12 => X"98361AC808127C454402483153A3A895BB3C1E2E820704020381702C1AAA2C4B",
INIT_13 => X"4D910CC1B154510413CC2A200501B400A40018A00C80400040D8AA288209AA21",
INIT_14 => X"0048A0141AA00418080460678A4012288463B2050302019200B00206C3590102",
INIT_15 => X"233142440470C8A9310280C0180302A01427D060022011606E800E00169C19A0",
INIT_16 => X"4010040100448008004000000E07008010003EFFFE0373056024B01118011988",
INIT_17 => X"0100401004010040100401004010040100401004010040100401004010040100",
INIT_18 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_19 => X"7E00000000000000000000000004010040100401004010040100401004010040",
INIT_1A => X"EFBEFBEFBEFBEFBEFFFFF7F7FFF3CF3CFFFFBE7FBBFDFFF7DFFCFBF08103DFDF",
INIT_1B => X"FFFFFFF7FBFDFEFF7FBFDFEFF7FBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFB",
INIT_1C => X"FFFFFFFE00003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"00080002000000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"FFFFFFFFFEBA5D2A954100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_1F => X"75FFFFFFFFFFFFFFFFFFFFFFFFFFEBA552A97400082A975FFFFFFFFFFFFFFFFF",
INIT_20 => X"FDEAA5D2E974100800155EFFFFFFFFFFFFFFFFFFFFFFFFFEAA552E95400082E9",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFDEAA5D2A95400080000000FFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"2E974105D2A80000FFFFFFFFFFFFFFFFFFFFFBFDEBA5D2E974005D2E80000FFF",
INIT_23 => X"FFFFFFFFF7FBFDEBA552A954005D2E97410FFFFFFFFFFFFFFFFFFFFFBFDEBA55",
INIT_24 => X"0000001FFFFFFFFFFFFFFFFFFFFF7FBFFEBA5D2A97400FF80174BAFFFFFFFFFF",
INIT_25 => X"FFFFFFFEBA5D2E97400000400000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2A95410000A001FFFFFFFFFFFFFFFFFFF",
INIT_27 => X"EAA552E954000020955EFFFFFFFFFFFFFFFFFFFFFFFFFEAA552E97400002E955",
INIT_28 => X"FFFFFFFFFFFFFFFFBFDEAA5D2A974101400155C7FFFFFFFFFFFFFFFFFFFFFFFD",
INIT_29 => X"97400552A80010FFFFFFFFFFFFFFFFFFF7FBFDEBA5D2E95400140E00000FFFFF",
INIT_2A => X"FFFFEFF7FBFFEBA552A95410552485038FFFFFFFFFFFFFFFFFFF7FBFDEBA552E",
INIT_2B => X"8A174AAFFFFFFFFFFFFFFFFEFF7FBFFEAA5D2E97400412497438FFFFFFFFFFFF",
INIT_2C => X"000000000000000000000001C7FFFFFFFFFFFFFFDFEFF7FFFFEAA5D2E95400E3",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974000004000000000000000000000000",
INIT_2E => X"A552E97400002E975FFFFFFFFFFFFFFFFFFFFFFFFFFEBA552A95410002E821FF",
INIT_2F => X"FFFFFFFFFFFFFFBFDEAA5D2A954000800155EFFFFFFFFFFFFFFFFFFFFFFFFDEA",
INIT_30 => X"4005D2A82010FFFFFFFFFFFFFFFFEFF7FBFDEBA552A974105D0015545FFFFFFF",
INIT_31 => X"DFEFF7FFFFEAA5D2A974005D2E82010FFFFFFFFFFFFFFDFEFF7FBFFEBA552E95",
INIT_32 => X"154AAFFFFFFFFFFFFBFDFEFF7FFFDEAA5D2E954105504154AAFFFFFFFFFFFFFF",
INIT_33 => X"BFDEBA5D2A95400A2AA974BAFFFFFFFFFF7FBFDFEFFFFFFDEBA552E974000004",
INIT_34 => X"0000000000000000000000000000000000000000155FFFFFFFFFF7FBFDFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(21),        -- Port A data input
DOA(0)   => data_read_a_hi(21),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(21),        -- Port B data input
DOB(0)   => data_read_b_hi(21),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_22_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"5290F4CDE914905A14A43D33F488243E17122300F55FEB189B343A1140548380",
INIT_01 => X"A94007B259F6A975386262000C344BA9573C6FF57B18A5FB0ABFCD3C2C5F4F0C",
INIT_02 => X"877FE30EB378008D202551040030071869D0040180AC4B685F6E26FAA0810006",
INIT_03 => X"431965109E4481D6B5AAD6875AD6AB5A1815600802888808DEA83552954D3000",
INIT_04 => X"492C0020220001010E4916C884DCD607E5EC2A344103E48003D0800023D0072C",
INIT_05 => X"0020F8882001102D620A06D683018001023D37E5088043620101179092540112",
INIT_06 => X"0803008022385AAA447A3306AA50001035B41C0A88046CAEE8C23C08E040011C",
INIT_07 => X"1EC04ED017AB5497EB923F08182E20020689B735011FBFE7BC06260294401CA8",
INIT_08 => X"4A00401D4425ADA9035BE19C8F9442A8801200F4C9D7AC8093A051727B2AC349",
INIT_09 => X"50020040E48D50080002B00A0C00801014541E9504703680017F6CB405070015",
INIT_0A => X"54538A8A738041C23020131A80CFDFF3FE509A907C6AC050402204090090319A",
INIT_0B => X"40050220103D2A512C6A8C4F0011550008E06E000140009A000000424DE61920",
INIT_0C => X"A81C2A81C2A81C2A81C2A81C2A81C2A81C9540E1540E001400006100003202D0",
INIT_0D => X"8B2940D0E153941A8B1A262CA542A9A8D6C0010A101628013456520CA09281C2",
INIT_0E => X"80410089180008800143D83888281A2034A85014280A14050A01509E05085449",
INIT_0F => X"000C26706B3C189CD84ACD20B03001E387D04AC560B02401E387E1028AC04500",
INIT_10 => X"458870201570B036C04AC560B03001E387D04ACD20B02401E387E24708E7E242",
INIT_11 => X"044708E7E1C20A0106EA167C84EBF052A8E010C0180606E86C3F459DC08DA902",
INIT_12 => X"98225189980254CDEC22A98032A22C50EAC462030A01800407C2700C2ACA2C0F",
INIT_13 => X"4A99BCC1154C258012D86F601A2E49003400138C0DA2443A208AA612C0096C37",
INIT_14 => X"90E16025483C1E0C0006B085CEC03858958D15310201015504B512044A313300",
INIT_15 => X"6B0469512C6FC01A1421006028038720640310643858162712020B001AA415F2",
INIT_16 => X"11044110445E22022365034A8EA754008004C0200323001182122548881649D1",
INIT_17 => X"1044110441104411044110441104411044110441104411044110441104411044",
INIT_18 => X"0401004010040100401004010040100401004010040100401004411044110441",
INIT_19 => X"7D05122890000000003FFFFFFFF9004010040100401004010040100401004010",
INIT_1A => X"E79E79E79E79E79EFFDFF7F5F777DF7DF7DF7EFF7BFA3FC7DF7AF5BF7EFDF7DF",
INIT_1B => X"9FCFE7F3F9FCFE7F3F9FCFE7F3F9E79E79E79E79E79E79E79E79E79E79E79E79",
INIT_1C => X"FFFFFFFE00000FE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F",
INIT_1D => X"10000000000000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"FFFFFFFFFEBA5D2E974000800021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_1F => X"21FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E954000004001FFFFFFFFFFFFFFFFF",
INIT_20 => X"FFEBA552A97400002A801FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2A9541008040",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFEBA552A97400082A975FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"2E95400082E975FFFFFFFFFFFFFFFFFFFFFFFFFFEAA552E95410002A955FFFFF",
INIT_23 => X"FFFFFFFFFFFFFFEAA552E95400002E975EFFFFFFFFFFFFFFFFFFFFFFFFFEAA55",
INIT_24 => X"000000000FFFFFFFFFFFFFFFFFFFFFFFDEAA5D2E97410080015545FFFFFFFFFF",
INIT_25 => X"FFFFFFFEBA5D2E97410080002000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974000004001FFFFFFFFFFFFFFFFFFF",
INIT_27 => X"EBA5D2A95410000A001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2A954000804021",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFEBA552A97400082E821FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"95410082A975EFFFFFFFFFFFFFFFFFFFFFFFFFEAA552E97400002E955FFFFFFF",
INIT_2A => X"FFFFFFFFFFFDEAA552E954000020955C7FFFFFFFFFFFFFFFFFFFFFFFFEAA552E",
INIT_2B => X"0015545FFFFFFFFFFFFFFFFFFFFFFFDEAA5D2A974001C24975C7FFFFFFFFFFFF",
INIT_2C => X"00000000000000000000000000FFFFFFFFFFFFFFFFFFFFFBFDEAA5D2A9741014",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800020000000000000000000000",
INIT_2E => X"A5D2A954000800021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974000004001FF",
INIT_2F => X"FFFFFFFFFFFFFFFFFEBA552A95410002E821FFFFFFFFFFFFFFFFFFFFFFFFFFEB",
INIT_30 => X"400002E975EFFFFFFFFFFFFFFFFFFFFFFFFFEAA552A97400082A801FFFFFFFFF",
INIT_31 => X"FFFFFFFBFDEAA5D2E95410082E955EFFFFFFFFFFFFFFFFFFFFFFFFDEAA552E97",
INIT_32 => X"17545FFFFFFFFFFFFFFFFFFFFFBFDEAA5D2A95400080015545FFFFFFFFFFFFFF",
INIT_33 => X"BFDEBA552A974105D0015555FFFFFFFFFFFFFFFFFFF7FBFDEBA5D2A974005504",
INIT_34 => X"0000000000000000000000000000000000000000010FFFFFFFFFFFFFFFFEFF7F",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"01FFFFFFFFE00000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(22),        -- Port A data input
DOA(0)   => data_read_a_hi(22),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(22),        -- Port B data input
DOB(0)   => data_read_b_hi(22),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_23_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"EF20906D902424807BC8241BC81801B97D38AD3C0800103362A6741C80A12A02",
INIT_01 => X"001FFF8409F089003B4422000D80C80106804A7951C5B9D1C828043EA28838F9",
INIT_02 => X"073B8858218C2C50801000F9FFEFF8E72CA7F5FC2E048026496834D84721DFE0",
INIT_03 => X"2C4360101A4001001005080400401420350016E0BB222341C312000014006FF8",
INIT_04 => X"00017B810015DC03D034201E14000036486008101FC0002EE006297E1C05F561",
INIT_05 => X"7E1F02FFFFC80100004044800080BEFFFC0248005FFC3C18A5FFC2444484BCC0",
INIT_06 => X"4082040800000811224DE0A00005FFBF8000000003FF810640A1C0008FF2F0E1",
INIT_07 => X"D1D72040048D00388387D03D0E591FFD201F862691DFBE077C2BC45B40FFE458",
INIT_08 => X"1FFBFFEC440501A5604B31062356282AA84200D12342113EDC40000004582800",
INIT_09 => X"A890FFF0002023FFDF79000000000EFFE309606020008005FC00000040200000",
INIT_0A => X"000000000037FF50010103134CAFDF03BA18000F39A0106F87D7FA84024B0225",
INIT_0B => X"88300C48907120AC81083315A493886640030010540DFF20FF8610302409000C",
INIT_0C => X"10C1010C1010C1010C1010C1010C1010C10086080860840063090442A18001B1",
INIT_0D => X"0000280600020040030090000012A500003FF7E08181119A41C1443243050C10",
INIT_0E => X"06542C7043FFD5FFF00A04BC010A7724B1000080004000200004150030010004",
INIT_0F => X"B2080290C2909080A872BC4FC8500054840072FC0FC8440054840200705F9861",
INIT_10 => X"0C8220180F1082E00072FC0FC8500054840072BC4FC84400548402214A380380",
INIT_11 => X"19214A380344920080B21810240AB182EB37C380B40800707011001B43253EE5",
INIT_12 => X"0019CE4000026C00C00042BD4149067465910640A0050C060A0028063672A000",
INIT_13 => X"4D801800CCB050001344060211629580B80022480A444111706658280009A203",
INIT_14 => X"944CB232D6D0100C040250200845132C10BE200403018061101A220339C80000",
INIT_15 => X"402102A5493B8E287E03808480060E40C83C1405132C90742E408D0082140820",
INIT_16 => X"0080200802000100100000000000004002403EFFF8002385F034901019465001",
INIT_17 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_18 => X"8020080200802008020080200802008020080200802008020080200802008020",
INIT_19 => X"0000000000000000000000000000080200802008020080200802008020080200",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000004000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFE00000000000000000000000000000000000000000000000000000000",
INIT_1D => X"10080400000000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"FFFFFFFFFEBA5D2E974100000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_1F => X"21FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100004021FFFFFFFFFFFFFFFFF",
INIT_20 => X"FFEBA5D2E954000800001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9740008000",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E954000004001FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"2A954100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2A954100000021FFFFF",
INIT_23 => X"FFFFFFFFFFFFFFEBA5D2A954100800021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_24 => X"0000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA552A97400002A801FFFFFFFFFFFF",
INIT_25 => X"FFFFFFFEBA5D2E97410080400000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800021FFFFFFFFFFFFFFFFFFF",
INIT_27 => X"EBA5D2E974000004001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100004021",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFEBA5D2E954000800001FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"954100004021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2A954000804021FFFFFFF",
INIT_2A => X"FFFFFFFFFFFFEBA5D2A95410000A001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2A",
INIT_2B => X"2E821FFFFFFFFFFFFFFFFFFFFFFFFFFEBA552A97410080E001FFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA552A9740008",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804000000000000000000000000",
INIT_2E => X"A5D2E974100000021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800021FF",
INIT_2F => X"FFFFFFFFFFFFFFFFFEBA5D2E974000004001FFFFFFFFFFFFFFFFFFFFFFFFFFEB",
INIT_30 => X"4000800021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E954000804021FFFFFFFFF",
INIT_31 => X"FFFFFFFFFFEBA552A954100004001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2A95",
INIT_32 => X"821FFFFFFFFFFFFFFFFFFFFFFFFFFEBA552A95410002E821FFFFFFFFFFFFFFFF",
INIT_33 => X"FFFEAA552A97400082A801EFFFFFFFFFFFFFFFFFFFFFFFFFEAA552A97410002A",
INIT_34 => X"00000000000000000000000000000000000000001EFFFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"01FFFFFFFFE00000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(23),        -- Port A data input
DOA(0)   => data_read_a_hi(23),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(23),        -- Port B data input
DOB(0)   => data_read_b_hi(23),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_24_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100600007FFF000080108004000800020000840041000080808",
INIT_02 => X"172A00D000EF8210000000F9FFEFF8E7240FF1FC224087B1000639401D005FC0",
INIT_03 => X"00003A2E200811000000000400000000340016603A0000004860400014006FFF",
INIT_04 => X"000079800014CC03C034001E04010850300000101FC0002EE000006E1C00F500",
INIT_05 => X"3E1F0067FFC000000000000000003E2FFC024800137C3C0000EFC00000003CC0",
INIT_06 => X"000000000000001123820AA00005FEBF8000000003FF80000021C0000FF0F0E0",
INIT_07 => X"E600084002040A10812A000500590FF9001F95406A8000037230C01840FFE000",
INIT_08 => X"01FBFFEC4695A501604A000C7585080002C200408102F16C0184800026C92C10",
INIT_09 => X"A8107FF0000000FFDF78000000000EFFE001600000000005FC00000000000000",
INIT_0A => X"000000000037FF4000000AA0354000019C4000012800002387D7F804024B0224",
INIT_0B => X"88300C0081408000800001002482886600020010100DFA20FF8600000000000C",
INIT_0C => X"00C1000C1000C1000C1000C1000C1000C1000608006084006301044081800121",
INIT_0D => X"00000000900160000000000000000000003FF7C0010101904181003003000C10",
INIT_0E => X"16100C4043FFD5BFF00004100000000411000000000000000000040030000000",
INIT_0F => X"3A0421080012302010049400086C022004200494000878022004120270599965",
INIT_10 => X"C19240300081406100049400086C022004200494000878022004124819081840",
INIT_11 => X"2348190814C09C01010400132100106836001504240E01040051200200D06410",
INIT_12 => X"202CD680C0100010408240BD80008983596CD86EA84104060503C0B000020250",
INIT_13 => X"0002090164F40086000082062C1B6600BC000C300818044000B27A0043000041",
INIT_14 => X"110002577FE4080C08010842180C40018545BBA00301808A0810C0059AD01802",
INIT_15 => X"4820C04100852B931F00800010081980B042D2044001850ED8808F00050A002C",
INIT_16 => X"0000000000000000000000000000000000003EFFF80037046031E0110001100A",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"9900000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"EFBE7BE7BE7BE7BEC99E61848655D75D7FCB42BBABDB9F3044CB35CF612B4441",
INIT_1B => X"83C1E0F0783C1E0F0783C1E0F07BEFBEFBEF9E79E79E79E79E7BEFBEFBEFBEFB",
INIT_1C => X"FFFFFFFE000001E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F07",
INIT_1D => X"10080402000000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"FFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_1F => X"01FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800021FFFFFFFFFFFFFFFFF",
INIT_20 => X"FFEBA5D2E974100000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741000000",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974100004021FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"2E974000800021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974000004001FFFFF",
INIT_23 => X"FFFFFFFFFFFFFFEBA5D2E974000800001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_24 => X"0000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E954000800001FFFFFFFFFFFF",
INIT_25 => X"FFFFFFFEBA5D2E97410080402000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFF",
INIT_27 => X"EBA5D2E974100800021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800021",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFEBA5D2E974100000001FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974000004001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100004021FFFFFFF",
INIT_2A => X"FFFFFFFFFFFFEBA5D2E974000004001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E",
INIT_2B => X"00001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E954000800021FFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9540008",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804020000000000000000000000",
INIT_2E => X"A5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FF",
INIT_2F => X"FFFFFFFFFFFFFFFFFEBA5D2E974100800021FFFFFFFFFFFFFFFFFFFFFFFFFFEB",
INIT_30 => X"4100000021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100000001FFFFFFFFF",
INIT_31 => X"FFFFFFFFFFEBA5D2E974000004021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E97",
INIT_32 => X"021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974000004001FFFFFFFFFFFFFFFF",
INIT_33 => X"FFFEBA5D2E954000804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E954000004",
INIT_34 => X"00000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(24),        -- Port A data input
DOA(0)   => data_read_a_hi(24),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(24),        -- Port B data input
DOB(0)   => data_read_b_hi(24),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_25_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100200002000000080100004000000020000800041000080808",
INIT_02 => X"1000218000000800000000F9FFEFF8E738FFF1FC20400400000004455A375FE0",
INIT_03 => X"00002000000001000000000400000000340016623A0000004000000014006FFF",
INIT_04 => X"924279824C94CC1BE0B4001F20000000020380401FE0082EF000106E1C00F500",
INIT_05 => X"3E1F0067FFE048002582800100523E2FFE024820137C3C0040EFE02000003CE4",
INIT_06 => X"821B0821B8019819200020200005FEBF81C1002203FF80000021C1140FF8F0E0",
INIT_07 => X"00040000000000000000000500590FF9001F0000000000033020C01840FFFC78",
INIT_08 => X"01FBFFFD0004000100502000011400000282004001020000000001009015C000",
INIT_09 => X"B8DA7FF8004000FFDF7C062031863EFFF75D78004001010DFC00002005010000",
INIT_0A => X"000000000037FFC00602000000000001980400002800032387D7FE94FBEF2B2C",
INIT_0B => X"88300C0080400000800001002486887600020110100DFA20FF8603000000000C",
INIT_0C => X"00C1000C1000C1000C1000C1000C1000C10006080060840077330C4889CC2925",
INIT_0D => X"00000000000000000000000000002500003FF7C0010101904189003003000C10",
INIT_0E => X"06140C6043FFD5BFF00A04B80608003CB120C110608830445821140134120800",
INIT_0F => X"02000000000200200000900000400200000000900000400200000200701E1861",
INIT_10 => X"0002000000010000000090000040020000000090000040020000000008080000",
INIT_11 => X"0000080800008000000000010100000022000000040000000040000000002400",
INIT_12 => X"0000420000000010000040318020000041000001000244000000008008000010",
INIT_13 => X"0002000004100000000080000002040040000000001000400002080000000040",
INIT_14 => X"0100000042000010002000001000400000042000040200000000400008400000",
INIT_15 => X"0030800000010800000000C0A000000000400000400000040800000000000004",
INIT_16 => X"41104451044C82082068C0200000008014023EFFFC0063046020801000001000",
INIT_17 => X"1104411044110441104411044110441104411044110441104411044110441104",
INIT_18 => X"1044110441104411044110441104411044110441104411044110441104411044",
INIT_19 => X"A080800002FFFFFFFFFFFFFFFFFC110441104411044110441104411044110441",
INIT_1A => X"41041249041249042824014C48569A69AFEE8A252865AA3168A4CBDF860EC15D",
INIT_1B => X"58AC56231188C46231188C462312492492492492492492492490410410410410",
INIT_1C => X"FFFFFFFE00002C562B158AC562B158AC562B158AC562B158AC562B158AC562B1",
INIT_1D => X"10080400000000000000000000000000000000000000000000000001FFFFFFFF",
INIT_1E => X"FFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_1F => X"01FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFF",
INIT_20 => X"FFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008040",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800021FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"2E974100000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800001FFFFF",
INIT_23 => X"FFFFFFFFFFFFFFEBA5D2E974100000021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_24 => X"0000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100000001FFFFFFFFFFFF",
INIT_25 => X"FFFFFFFEBA5D2E97410080400000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFF",
INIT_27 => X"EBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974100800001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800021FFFFFFF",
INIT_2A => X"FFFFFFFFFFFFEBA5D2E974100800021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E",
INIT_2B => X"00001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100000021FFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741000",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804000000000000000000000000",
INIT_2E => X"A5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FF",
INIT_2F => X"FFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEB",
INIT_30 => X"4100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFF",
INIT_31 => X"FFFFFFFFFFEBA5D2E974100800001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E97",
INIT_32 => X"021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800021FFFFFFFFFFFFFFFF",
INIT_33 => X"FFFEBA5D2E974100000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800",
INIT_34 => X"00000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"01FFFFFFFFE00000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(25),        -- Port A data input
DOA(0)   => data_read_a_hi(25),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(25),        -- Port B data input
DOB(0)   => data_read_b_hi(25),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_26_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"E9264EAB20190CA3BA4997AA9002AE9C001006B0778015CFA17E0811039879C7",
INIT_01 => X"F1FFF9BB1F773C7F9BB07DFFFDD863FC5FFF3FEFFBBF9FFB22FFFBC7B9F30686",
INIT_02 => X"1B33188302E708180F6FFBFFFFCFFFFF9C7FF7FC24350B99082400001D00DFD8",
INIT_03 => X"4A53D958C50000DCE7366303739CD98C27C57EF57980014F271807E3C9E9CFF8",
INIT_04 => X"DBFAFBD7FB1CDEBEF1BE17F7AC88042787FBFFF8FEE9FF7EE6F4C0EE1FFAF869",
INIT_05 => X"BE1FFD67DFFEFFBDA7F7FED508707E2EFEBF6FFEB37C3FF302EEEDFF9B487CF6",
INIT_06 => X"75F7275F7CAC98E261EDF0253C7FFFEF87C74E8CCFFBB6FF70E1FE61FFBDF0FE",
INIT_07 => X"73840C07783060C72DF7D828912E6FFB80162776F3BFB7077E82255E40BFEEBA",
INIT_08 => X"69FFBFE43C872321367036163F1C0820A3063F460D1AEFC000060042648C4181",
INIT_09 => X"FB967FBD13D981F7DF7D7E6171AF3FEFE8A3E679FAC1FD1FFFBEB000763A8447",
INIT_0A => X"6AED1D1DAD7FBE7D67D7F3BB79CFFB83BF14EC1E7D7300B017F5FFE6FBEF73BE",
INIT_0B => X"99F51EDDCDEBCFF589807B70AD9A99EE7583F931109FFE33FF8E3FDFDAF64A3C",
INIT_0C => X"C0D78C0D78C0D78C0D78C0D78C0D78C0D7A606BC606B8C56F7730ECCDBDF1521",
INIT_0D => X"1D406B9EC20181CC1F73F87501DED3409BFFFEFFEBF341B867D3683A03A40F78",
INIT_0E => X"86D70CE04FFFFF3FF1F5F5475BD7F72E4D75EBFAF5FD7AFEFDFFAF59B6FF28FE",
INIT_0F => X"020007C040101480807D17B0004001F804007D17B0004001F8040212F35FFC6D",
INIT_10 => X"700200001DC00068007D17B0004001F804007D17B0004001F804006F60081400",
INIT_11 => X"206F60081800800007B000102C0801FB02683800040007700011801003DE050A",
INIT_12 => X"403E232130207080D012CEFF41008D188D502100B02004000F01900039020040",
INIT_13 => X"0E101A01F21A2C40039006823F80048100003F0008004D8100F90D162001C803",
INIT_14 => X"B604027F020A07400007C040085581019D602451500001EC00100247C4642608",
INIT_15 => X"CC3F02010EA40EA00020C830100F0D000022180581019F40084800001F100020",
INIT_16 => X"EBFAFEFFBFEFDFDDFE7DD87FEFF7FF796FFFFFDFFC017FEFFD7E841001D8197D",
INIT_17 => X"BFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAF",
INIT_18 => X"FAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFE",
INIT_19 => X"EDB5C88646FFFFFFFFFFFFFFFFFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEB",
INIT_1A => X"61861A69A6986186EBCAF55357E1C71C751D6C56F3D247859B3214FA76953F86",
INIT_1B => X"84C26130984C26130984C2613098618618618618618618618618618618618618",
INIT_1C => X"FFFFFFFE0000026130984C26130984C26130984C26130984C26130984C261309",
INIT_1D => X"10080400000000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"FFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_1F => X"21FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFF",
INIT_20 => X"FFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008040",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFF",
INIT_23 => X"FFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_24 => X"0000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFF",
INIT_25 => X"FFFFFFFEBA5D2E97410080400000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFF",
INIT_27 => X"EBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFF",
INIT_2A => X"FFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E",
INIT_2B => X"04021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804000000000000000000000000",
INIT_2E => X"A5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FF",
INIT_2F => X"FFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEB",
INIT_30 => X"4100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFF",
INIT_31 => X"FFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E97",
INIT_32 => X"001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFF",
INIT_33 => X"FFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804",
INIT_34 => X"00000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(26),        -- Port A data input
DOA(0)   => data_read_a_hi(26),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(26),        -- Port B data input
DOB(0)   => data_read_b_hi(26),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_27_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"00080A40000A41248002029000050A088000008242A0004404480002000A1155",
INIT_01 => X"F1FFF1C11F781C129C107DFFFE0860941E81258CA2B71C2220EC1B86E1A00002",
INIT_02 => X"4000002100000014400FF6FFFF0FFFFF8007F1FC211100014200800000887FC0",
INIT_03 => X"0842D85841000098C63061026318C18404C459757000015F00088BE3C0618FF8",
INIT_04 => X"DBEAE5D6D91C2EBCE1B21EA72C00000007FBE7C8F8E9EF79E6D440E91FDAE061",
INIT_05 => X"B91FF9671FE6B68984B5BCE408347E28FEBF6FEEB3723F7102E8EDBF8A4872F6",
INIT_06 => X"3573A357308418E40000D4113C7FFE4F86064C8DDFE3B6FF50D1FC61DE39C8FC",
INIT_07 => X"00000A20083060C00C81882A008C6FF880060424B39FB6037F00051C003FE04A",
INIT_08 => X"61FA3FE4010440410844060001040A00002200460D1A06000005040000001080",
INIT_09 => X"EB027E390A4881C7BEFC5F6171CE2F8FE823E778DAC16C1FFBBC900031589547",
INIT_0A => X"03813030213C3E2D62D6E21259CFDB039E806C024531008017C1F826FFEF41FE",
INIT_0B => X"9AB55F0DEFABC705488069302DBA98EAB582D835109FFC31FFAEAFCFDAF4423D",
INIT_0C => X"40C3440C3440C3440C3440C3440C3440C3C2061A2061AD46FF730E5CCBCD5521",
INIT_0D => X"0C407D1F820101441DA3A8310198C34089BFF8DD6B7941BC63F1683803C00E34",
INIT_0E => X"5710AE4047FFD23FF315D54358D593474955AB6AD5B56ADAB5FAAE58B2F628EA",
INIT_0F => X"020007C0400004C080791290004001D80001791290004001D8000210F1587971",
INIT_10 => X"300200001DC0000801791290004001D80001791290004001D800012F60080400",
INIT_11 => X"202F60080800800007B000000E0801BB020828000400077000008210035E0408",
INIT_12 => X"40BA2220202070801010C6F1410085188D500100102004000F01900031000060",
INIT_13 => X"0E100205D2120840039000813F80040100003F0000000F8100E909042001C800",
INIT_14 => X"3E04007F020201400007C040001781011D602040500001EC0000005744440408",
INIT_15 => X"C43F02000EA40EA000004810100F0D000020080781011F40080800001F100000",
INIT_16 => X"AB6ADAB6BDE75ED5EC71385FC2512E3565BBBF1FFC00636EED7E841000D81924",
INIT_17 => X"B6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6AD",
INIT_18 => X"6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADA",
INIT_19 => X"A471688747FFFFFFFFFFFFFFFFFAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB",
INIT_1A => X"0020800000000000780401CBC840000005243885A04012072A1810DA84002104",
INIT_1B => X"5028140201008040201008040200000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFE000028140A05028140A05028140A05028140A05028140A05028140A0",
INIT_1D => X"10080400000000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"FFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_1F => X"01FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFF",
INIT_20 => X"FFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008040",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFF",
INIT_23 => X"FFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_24 => X"0000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFF",
INIT_25 => X"FFFFFFFEBA5D2E97410080400000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFF",
INIT_27 => X"EBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFF",
INIT_2A => X"FFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E",
INIT_2B => X"04021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804000000000000000000000000",
INIT_2E => X"A5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FF",
INIT_2F => X"FFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEB",
INIT_30 => X"4100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFF",
INIT_31 => X"FFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E97",
INIT_32 => X"021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFF",
INIT_33 => X"FFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804",
INIT_34 => X"00000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"01FFFFFFFFE00000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(27),        -- Port A data input
DOA(0)   => data_read_a_hi(27),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(27),        -- Port B data input
DOB(0)   => data_read_b_hi(27),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_28_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"02200AA400180030808802A900002A08001280A08A801044104A1000001818C3",
INIT_01 => X"50A00011460214428114180000882214413D0A71592A01D92213D28005210202",
INIT_02 => X"1444428102100884000AA30200000000C1000401041108404400022220800000",
INIT_03 => X"461080404900000C6314A900318C52A40051081000888806108802A141288001",
INIT_04 => X"00800040110102000902002000888400081045A8A00003C00000500000080008",
INIT_05 => X"0000000000024CA0A0101800032000400000000B800000014000000B08180000",
INIT_06 => X"10280102802C0240041000011428004022220024440013511000013510000000",
INIT_07 => X"0804420009122448451020100020400080002041000000008000010400000880",
INIT_08 => X"2800000140200808021006108010422AAA800022448902849220114009224081",
INIT_09 => X"01C800004080A0000002480B04008100011000088800081002C19020150B0013",
INIT_0A => X"56D29A9A52800004004070208000000040006408001100105000020000001800",
INIT_0B => X"00040024440245400082D0220800008010001020458000010000040D96104210",
INIT_0C => X"50160501605016050160501605016050160280B0280B00120008430660210014",
INIT_0D => X"054001884200810C1631181500CA60400B4008072020500002002C0040010360",
INIT_0E => X"104420A00C000200005000010040A0020CC000200010000800920040804020A6",
INIT_0F => X"0000000000001400000102900000002800000102900000002800001001802104",
INIT_10 => X"3000000000000048000102900000002800000102900000002800000020000400",
INIT_11 => X"0000200008000000000000002800000100082800000000000001800000020008",
INIT_12 => X"4000202020200000901005480000000800000100102000000000000009000000",
INIT_13 => X"0000120002020840000004800080000100000000000048800001010420000002",
INIT_14 => X"A200000800020140000000000050800008000040500000000000024004040408",
INIT_15 => X"840A000002000000000048100000000000020800800008000008000000000000",
INIT_16 => X"8020080210810840861CD33548542A10209D4100000010200400000000880035",
INIT_17 => X"0200802008020080200802008020080200802008020080200802008020080200",
INIT_18 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_19 => X"40A0C22E10000000000000000000020080200802008020080200802008020080",
INIT_1A => X"08208208208208200360D4141D630C30C7788440B044280091A5CB03D01BD89A",
INIT_1B => X"582C16030180C06030180C060302082082082082082082082082082082082082",
INIT_1C => X"FFFFFFFE00002C160B0582C160B0582C160B0582C160B0582C160B0582C160B0",
INIT_1D => X"10080400000000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"FFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_1F => X"01FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFF",
INIT_20 => X"FFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008040",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFF",
INIT_23 => X"FFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_24 => X"0000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFF",
INIT_25 => X"FFFFFFFEBA5D2E97410080400000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFF",
INIT_27 => X"EBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFF",
INIT_2A => X"FFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E",
INIT_2B => X"04001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804000000000000000000000000",
INIT_2E => X"A5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FF",
INIT_2F => X"FFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEB",
INIT_30 => X"4100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFF",
INIT_31 => X"FFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E97",
INIT_32 => X"001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFF",
INIT_33 => X"FFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804",
INIT_34 => X"00000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"01FFFFFFFFE00000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(28),        -- Port A data input
DOA(0)   => data_read_a_hi(28),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(28),        -- Port B data input
DOB(0)   => data_read_b_hi(28),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_29_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"79964E4BA01DACAB9E659792D00AAE160002829C7FDFEFCEE97C2815039D70C3",
INIT_01 => X"50BFF9AB0775343F9AB01DF80D5821FC0FFF3FEFD1AF9FF1207FFBC7B9720586",
INIT_02 => X"0B33180300E700080F6AAA7BFFC007189C7FF2FC003503980A0000001D00DFD8",
INIT_03 => X"0401D940CD0000C8421A2B03210868AC23403E903900010E271006A148A0C000",
INIT_04 => X"49B87A417315D20A313E17F1800000058013DDF8BE21F36E02F0D06E03E8F800",
INIT_05 => X"3E00FC67C03A4D9C87525E5101603E6E023D27DA937C03E340EE25CB9B483C12",
INIT_06 => X"50B5050B540C004261EDE025142DFFE003C30E0447F877F930203E213F8CF01E",
INIT_07 => X"73800407781020476467D008910A4FFB80100332D1AE93059282215E40800678",
INIT_08 => X"21FF80003C832320342036063F08000001063F42050AEB4000221000248C0180",
INIT_09 => X"51547F8C1111A0F041056A0100A11FE000916249A800B915FE82B02052290002",
INIT_0A => X"2AAD1515AD5780540541619968C76980E914E4163D53002017F405C409A42A9A",
INIT_0B => X"014002D445624DB481806A6288100184500171200085FE030000157FDF124A10",
INIT_0C => X"D0068D0068D0068D0068D0068D0068D006A68034680300021410028450530014",
INIT_0D => X"15402B0E8201018C1561E855008C50401B7FFE27A0B2500806522C0A40A50268",
INIT_0E => X"928324400DFFFF0001F1F0050342D42A086040B02058102C48970541944B20FA",
INIT_0F => X"0000000000101480000507B00000002804000507B000000028040212034FAD28",
INIT_10 => X"7000000000000068000507B00000002804000507B00000002804004020001400",
INIT_11 => X"0040200018000000000000102C0000410068380000000000001180000082010A",
INIT_12 => X"4004212130200000D0120ED64000080800002100B02000000000000009020040",
INIT_13 => X"00001A00220A2C4000000682008000810000000008004D800011051620000003",
INIT_14 => X"B6000208000A0740000000000855800088000451500000000010024084242608",
INIT_15 => X"8C0F0001020000000020C8300000000000021805800088000048000000000020",
INIT_16 => X"C0B02C4B12C989489418D13FE7F3FFD8BADB7FC004012CA5141600000198087D",
INIT_17 => X"0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02",
INIT_18 => X"B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C",
INIT_19 => X"FEA0C00602FFFFFFFFFFFFFFFFFC0B02C0B02C0B02C0B02C0B02C0B02C0B02C0",
INIT_1A => X"FBAEBAEBAEBAEBAEFFFFF7E7EFBFFFFFFAEF3E7E5BB9FFF7DFF9E3F08843FFDF",
INIT_1B => X"FDFEFF7FBFDFEFF7FBFDFEFF7FBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBE",
INIT_1C => X"FFFFFFFE00003EFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FB",
INIT_1D => X"10080400000000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"FFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_1F => X"01FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFF",
INIT_20 => X"FFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008040",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFF",
INIT_23 => X"FFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_24 => X"0000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFF",
INIT_25 => X"FFFFFFFEBA5D2E97410080400000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFF",
INIT_27 => X"EBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFF",
INIT_2A => X"FFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E",
INIT_2B => X"04001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804000000000000000000000000",
INIT_2E => X"A5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FF",
INIT_2F => X"FFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEB",
INIT_30 => X"4100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFF",
INIT_31 => X"FFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E97",
INIT_32 => X"001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFF",
INIT_33 => X"FFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804",
INIT_34 => X"00000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(29),        -- Port A data input
DOA(0)   => data_read_a_hi(29),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(29),        -- Port B data input
DOB(0)   => data_read_b_hi(29),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_30_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"FD00000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"E79E79E79E79E79EEBFEF5D7D7F7DF7DFFDFFEFFFBFE7F87DFFEFFBF77BFFFDF",
INIT_1B => X"9FCFE7F3F9FCFE7F3F9FCFE7F3F9E79E79E79E79E79E79E79E79E79E79E79E79",
INIT_1C => X"FFFFFFFE00000FE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F",
INIT_1D => X"10080400000000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"FFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_1F => X"01FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFF",
INIT_20 => X"FFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008040",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFF",
INIT_23 => X"FFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_24 => X"0000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFF",
INIT_25 => X"FFFFFFFEBA5D2E97410080400000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFF",
INIT_27 => X"EBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFF",
INIT_2A => X"FFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E",
INIT_2B => X"04001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804000000000000000000000000",
INIT_2E => X"A5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FF",
INIT_2F => X"FFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEB",
INIT_30 => X"4100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFF",
INIT_31 => X"FFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E97",
INIT_32 => X"001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFF",
INIT_33 => X"FFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804",
INIT_34 => X"00000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(30),        -- Port A data input
DOA(0)   => data_read_a_hi(30),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(30),        -- Port B data input
DOB(0)   => data_read_b_hi(30),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_31_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"129000008004A00804A40000400800020000000C005FEA005800200400050100",
INIT_01 => X"A15FF18019700810180065FFFC0040801E80258CA2951C2200EC0906A0804140",
INIT_02 => X"0000000000000011000550FDFF0FFFFF0007F1FC200000011000000000205FC0",
INIT_03 => X"08425818000000908428C0024210A30004045060302223490002014280410FF8",
INIT_04 => X"DB6A618248140C18E0B016872400000007EBA24058E1ECA8E2D400681FD0E061",
INIT_05 => X"381FF8671FE01009048084C400103E28FE3F6FE513703F7000E8E5B4825030F6",
INIT_06 => X"00130001300018A00000D0002855FE0F84040C088BE3E4AE40C1FD04CE38C0FC",
INIT_07 => X"000008800020408008818838000C2FF800060424B39FB6037E000418003FE008",
INIT_08 => X"41FA3FE400040001004000000104088000020044091204000004000000000000",
INIT_09 => X"E8027E38004801C79E7C162231862E8FE00166704041240DF93D000000000004",
INIT_0A => X"0000000000343E002202021259CFDB039E0008024520000047C1F804FBEF01BE",
INIT_0B => X"88310E08812982050800A9102492986200824810110DFC30FF86036249E4002C",
INIT_0C => X"00C1000C1000C1000C1000C1000C1000C18006080060840477330C4889CC0121",
INIT_0D => X"08006816800100400902A0200110810080BFF0C80111019861D1403803800C10",
INIT_0E => X"06100C4043FFD03FF101D4000800130401808100408020401020041830120848",
INIT_0F => X"020007C04000008080781000004001D00000781000004001D0000200F0185861",
INIT_10 => X"000200001DC0000000781000004001D00000781000004001D000002F40080000",
INIT_11 => X"202F40080000800007B00000040801BA020000000400077000000010035C0400",
INIT_12 => X"003A0200000070800000C231410085108D500000000004000F01900030000040",
INIT_13 => X"0E100001D0100000039000003F00040000003F000000050100E808000001C800",
INIT_14 => X"14040077020000000007C0400005010115602000000001EC0000000740400000",
INIT_15 => X"403502000CA40EA000000000100F0D000020000501011740080000001F100000",
INIT_16 => X"01004010044602002061004A820104809402BE1FFC006304E036841000501900",
INIT_17 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_18 => X"0040100401004010040100401004010040100401004010040100401004010040",
INIT_19 => X"0001000802FFFFFFFFFFFFFFFFF8100401004010040100401004010040100401",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFE00000000000000000000000000000000000000000000000000000000",
INIT_1D => X"10080400000000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"FFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_1F => X"01FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFF",
INIT_20 => X"FFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008040",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFF",
INIT_23 => X"FFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_24 => X"0000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFF",
INIT_25 => X"FFFFFFFEBA5D2E97410080400000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFF",
INIT_27 => X"EBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFF",
INIT_2A => X"FFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E",
INIT_2B => X"04001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804000000000000000000000000",
INIT_2E => X"A5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FF",
INIT_2F => X"FFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEB",
INIT_30 => X"4100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFF",
INIT_31 => X"FFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E97",
INIT_32 => X"001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFF",
INIT_33 => X"FFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804",
INIT_34 => X"00000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(31),        -- Port A data input
DOA(0)   => data_read_a_hi(31),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(31),        -- Port B data input
DOB(0)   => data_read_b_hi(31),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_0_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"ED39BA795990D275FB4A6E96ACC4731DEA4598B0AFB54867F6EE4618C3749807",
INIT_01 => X"58A0047D8607944AC7DA180001ECA2544042106208408208C20022E9173734B3",
INIT_02 => X"9F775E7CB273E6CCA7DAAF00001000000478020113C9C38E09FB7CCCDD9F203E",
INIT_03 => X"441406267B4CB04443163C91110C58F24A31000B8028A810A3D0F8B169A01006",
INIT_04 => X"0005802424830120024121209088809DF81454ACA01E03501D0A3B91E00F0A00",
INIT_05 => X"C1E0039800112014C20B0232838F80D001C0100AEC83C008EF101A034C8CC300",
INIT_06 => X"8B0478B04A83405954592F9B9628000002C3F08754001B51881E007900060F01",
INIT_07 => X"39F36677EE1C387777622717EF711004A6818111086008E080FDC30594001017",
INIT_08 => X"160400195E83A3A0F61BC3929ECB622AABF5FF83860CEB164833F179B48CEE59",
INIT_09 => X"036D8004FDB47600000229410C61010016DC998C84B0128202C0DCB48F05D513",
INIT_0A => X"204122A033000182502440888420247041E876810099D35F900002DB00105C01",
INIT_0B => X"41C000947E16656074EA560F080544900960260144D201890018080D36191110",
INIT_0C => X"781EA781E2781EA781E2781EA781E2781C33C0613C0E00120800239450112ED4",
INIT_0D => X"872917095352BD2A90515A1CA44E7EA84B00001010043803120C3E04E03383E2",
INIT_0E => X"70C7E0B92800224008AE09B8942C48D1FC491204890244812250588601285432",
INIT_0F => X"B80C2038ABACB83C7E03EA5FF83C002783F103EA5FF83C002783F0120847A704",
INIT_10 => X"BD9870380230F2D7C103EACFF83C002783F103EACFF83C002783F310BBF7EFC2",
INIT_11 => X"1F10BBF7EFC61E01804E1E6EA1E3FA01FD97EFC4B80E008C7C2F678FF023FAF5",
INIT_12 => X"B801FCC8E8320C4DAC9220C6B2FF22EF72ADDE6F1A67C80600C2683E0EF8AE1F",
INIT_13 => X"4189B5C00FE651C6104C6D6400FFFB01FC0000FC07EE42FA7C07F22CE3082636",
INIT_14 => X"8BE9FC08FDF4195C0C2038A7C6CAFA7E289F9BA4570380131CAFB2003F9D190A",
INIT_15 => X"270AE9FE635BE11B7F0308D4A80092E0FC1FC662FA7E283FF68A8F0080AE1DDA",
INIT_16 => X"1204812058112C12411402056954AB0C280D000003350013024179498C2EC6B9",
INIT_17 => X"2048120481204812048120481204812048120481204812048120481204812048",
INIT_18 => X"0481204812048120481204812048120481204812048120481204812048120481",
INIT_19 => X"13043A85D4000000000000000001204812048120481204812048120481204812",
INIT_1A => X"82082082082082082218821390771C71C557CE263826D5B1D36AC59E0765D1CF",
INIT_1B => X"1F0F87C3E1F0F87C3E1F0F87C3E0820820820820820820820820820820820820",
INIT_1C => X"FFFFFFFE00000F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E",
INIT_1D => X"EF5D7BD7400000000000000000000000000000000000000000000061F007FFFF",
INIT_1E => X"A10A2D1574005D0428A10A2AAA8BEF552EBDFFF557BC01FF5D7BFFEBA5D55555",
INIT_1F => X"DEBAFFFFC2000AA8428AAAFFAAA8BFF00002AA10FF802ABEFA2D16AA00F7FBE8",
INIT_20 => X"975EFFF8002010002EAAAAAAAD1555FFFFAEA8B550051401450055575FF00517",
INIT_21 => X"4155FF0855575455D2AA8BFFA2D1575EF5D5555545FFFBE8A00087FC20BA5D2A",
INIT_22 => X"8028A00FFAE800AA082A820005D2E974BAA2D140145A2842AA00A284021FF5D0",
INIT_23 => X"2D17FFEF000017400FFD1555FF007FFFEBA55042AA00000017400FFAABFEBAFF",
INIT_24 => X"000000155F7D540000F7FBFFE105D7BE8ABAA284000105D0428BFFA2FBFDFFFA",
INIT_25 => X"75D7BFAEBA5551501D51C5FC7E00000000000000000000000000000000000000",
INIT_26 => X"28B6D16AA28EBF5EDA38AADE1543849557D492BF8E2DE00552EBFFC7552BC01D",
INIT_27 => X"000A85400E00E38A175FDE3F5C002DAAD42DAAAF784AFA82BC042DF47E3D1F80",
INIT_28 => X"AA150021C0092490E904BAFFD550A90FFA495FC7A05B555C257AAA8B45007540",
INIT_29 => X"2DA02402ABD4AD1D0E175D7140B455D516A1EAB45E2A000B4748717A095F571E",
INIT_2A => X"4004A8BC0ABFF7D03A17D1D5147540B454AA080038E9748542AE3D0051C7B6F0",
INIT_2B => X"FB6D4B8FC7BFFFD2168B68F57492F505FF5FA550490BFA482B420B8428A3DA85",
INIT_2C => X"0000000000000000000000016ABD554201543A1EDE9016D4AAB454AF400547AB",
INIT_2D => X"5D2EBDF55556BC35E7557FE8AB25D11415FD0151614000000000000000000000",
INIT_2E => X"9596CBEA41D7D3DECFAF7D43FABAAAD57DEBAAAFFD74AA04547EE18D680BE9A5",
INIT_2F => X"47D78228E5000EA422E10439C1FBCD282351BDAAF9C20AAAABCBEB1DFF803FC5",
INIT_30 => X"1E6284683ABBDD7DEAA100069C14B25495A00F38EBAC0E198B97605018053575",
INIT_31 => X"4408FE6A755ED8EFEFE41B2D17EAF02552BC0545556BD61E501001DF5DD3EBA3",
INIT_32 => X"556F922ACA8AB8283C8310FAB1588916D3861C0422C44082B52A81550A828141",
INIT_33 => X"A5FDBCD7D262E5AFAC4B6AADDD562AF57D7C369AF25495A23068A8301BA7FB95",
INIT_34 => X"003FE0000003FE0000003FE0000003FE0000003FE03D5789700282E9FEFB501E",
INIT_35 => X"0003FE0000003FE0000003FE0000003FE0000003FE0000003FE0000003FE0000",
INIT_36 => X"00000000000000000000000000000000000000000000000000000000003FE000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(0),        -- Port A data input
DOA(0)   => data_read_a_lo_256(0),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(0),        -- Port B data input
DOB(0)   => data_read_b_lo_256(0),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_1_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"212C001411984004084D000508C53810A03D1450E839B003342114428A000807",
INIT_01 => X"08000010400A0008010600000084004000400002000000000000000000140000",
INIT_02 => X"484DEBA0111800C004400D000000000028800001CC404E6008B4933336880010",
INIT_03 => X"650C00000848A0423183089008C604224200000100A200002C280810098C0001",
INIT_04 => X"00000004208B00200E010800006667BE7000102C00080000040012010000080C",
INIT_05 => X"0100000000002000600100208D04414000800000000200004800080000800200",
INIT_06 => X"010420104032C204071200000200000010104020000001000910000000040800",
INIT_07 => X"8C0060242183060CF118011281B00000220010400020002081A0008210000802",
INIT_08 => X"000400014812466427040098C000622AAAA43E3060C158AC97F0356BDBFBD008",
INIT_09 => X"026C000559102400200281400469000008B0800000901080004004308B434040",
INIT_0A => X"50502A2800800000400408200000201041000208000040020820034200005C00",
INIT_0B => X"13C051112A800008402002021128000081202205001000000028880004010500",
INIT_0C => X"191AC191A4191A4191AC191AC191A4191A00C8560C8D2940804060901210441E",
INIT_0D => X"C1C114417882F82C00181707044212080300001002081224002006406401918C",
INIT_0E => X"60C0C0B92C000000000400001004200044010200810040802040080200284401",
INIT_0F => X"380C200000043C2016000000F03C00280030000000F03C00280030000004860C",
INIT_10 => X"8D18703800000049C0000000F03C00280030000000F03C002800321080000BC2",
INIT_11 => X"0110800007861E0180000002A9001A00000007C4380E00000001E00230000000",
INIT_12 => X"688004C0C81200009480010280340000008082430A07C80600C0000009008610",
INIT_13 => X"4000134400241186100004A500007B00FC000000000E4A402C001208C3080002",
INIT_14 => X"A9002C0001E0181C0C200000025A400A200812A4070380000000B25000981902",
INIT_15 => X"0000804A0002410A170300C4A800800000020E22400A200096828F008000000A",
INIT_16 => X"020080200820040041002000010080000000000002340002004118010C228614",
INIT_17 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_18 => X"0080200802008020080200802008020080200802008020080200802008020080",
INIT_19 => X"2B5000A000000000000000000000200802008020080200802008020080200802",
INIT_1A => X"AA8A28A28A28A28AB2048634B03249249604CA291AEAFBF1528205C00020C745",
INIT_1B => X"974BA5D6EB75BADD6EB75BADD6EAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA",
INIT_1C => X"FFFFFFFF00000BA5D2E974BA5D2E974BA5D2E974BA5D2E974BA5D2E974BA5D2E",
INIT_1D => X"55AAAAAAA00000000000000000000000000000000000000000000181FFFFFFFF",
INIT_1E => X"BEF5D7BE8ABA5D557DFEFFFD17FEBA00042AAAAFFFFFFE00FF843DF45FFAE955",
INIT_1F => X"DFEF552A800AA5555575FFA2AE820BAFFAEBFF555500155EF552E975FFF7D168",
INIT_20 => X"6AA00A2FBEAABA5D55420AA00002AA00AAFBE8B55A280175455D002AA00A2AAB",
INIT_21 => X"BD75FFAA802AAAAFFAA801EF00517FFFFF7D56ABEF0004155550004154105D55",
INIT_22 => X"55575FF08557DEBAA2FBEAAAA552E955EF5D0415410A2AE97545A2AE954BAF7F",
INIT_23 => X"7D17DF55A2AEBDEAAFFFFC20AAFFFFFFFFFAAD5555FFFFAEAAB55A2D168B555D",
INIT_24 => X"0000000BAFFFBE8A00087FC20BA5D2A975EF5D0002010552E820AAFFD57FF55F",
INIT_25 => X"8FF8A38F45F7AA9217FA380AD400000000000000000000000000000000000000",
INIT_26 => X"D7552E975EFFFDF68BFF557BEAA925551785D7BFD5EFE3F08002FA92EBA5FDE2",
INIT_27 => X"43841017DE92BF8E3AA824924870BF5551555C7A28A821EFE3AABAE38005B575",
INIT_28 => X"0568005A1041055716DB7DB6FBEFEA81C55D0A0516802AA28BEF5EDB7DAA8A15",
INIT_29 => X"C7FEF1C043FE28E3FBD55FFAADE2DAAAE3A5C51C71C042DF45A3D1D00281E8A1",
INIT_2A => X"AA8B45B47F6FB55A95555E90F78E17F52FEF5EDA82FD249057F080417492AAAF",
INIT_2B => X"5FF8AAAA95B7AF45FF8F7DFEDFFAFF8E005FAE92A3AE3DBFF57FA2DF555D257A",
INIT_2C => X"000000000000000000000000A8F571EAA150021C0092490E905FFFD0550BD75C",
INIT_2D => X"00043DE00A2C57DE08FFAAA8B55F7EE801F7F2849EE000000000000000000000",
INIT_2E => X"6AAAE29F067155543A15D2E955EFFFFBEABEF557FEAA10595169BED83D1EBCA8",
INIT_2F => X"BAFFD57DEEAAA15976EB0444BFEB086808A8E3082C954BA5D7DD6145AAAA821A",
INIT_30 => X"B47FFD55D6107782001FF0812000A255D57FFBEF3B97EEAB2C40217B9778428A",
INIT_31 => X"35FF003F17418AEE817B540D11CA80BAAFA825EFAABEBCA18FE803755D08079E",
INIT_32 => X"8BDEBA2D757547D7862AF57ABFFCABE5553FD5FBEFE86353EFFFD03FE0275000",
INIT_33 => X"5A01F70C6AA04537957D6FB4807FFFB45F7EFFDA58FF2AA88A0F3C5014018AC2",
INIT_34 => X"00000000000000000000000000000000000000000B2DD7DEAA100069C14B2549",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(1),        -- Port A data input
DOA(0)   => data_read_a_lo_256(1),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(1),        -- Port B data input
DOB(0)   => data_read_b_lo_256(1),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_2_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10E006600180111284380310006289800480032283E000A34301002001A0816",
INIT_01 => X"0005A00810790848048044A54E404340404000720885800802000806EC910200",
INIT_02 => X"5C010802020408040C400850AA055254090541A111200A104A0000000908B510",
INIT_03 => X"0C1101100C00004401060A0010041028021560A0218808002440840008880550",
INIT_04 => X"8840C2802205140048281202180804040960986850688C99444090C10A124A69",
INIT_05 => X"910A21220A880010214000010340086856B141252252142242A068B090106372",
INIT_06 => X"4007A400E8A40086213090040001520500204088012121026050A54CE2154840",
INIT_07 => X"0204022420000004601120108108055200022025A83AA3008882004A001542CA",
INIT_08 => X"091C154429220A2824642010A010020282843E00000248000021100000884101",
INIT_09 => X"80442C1411D120828A2A116A24632885419244606001110AE11B202046439511",
INIT_0A => X"644022201204145003031012D40D718241108815384200904160AE42CE2818E2",
INIT_0B => X"1BF047118108829501009202A5A20068C003211551163A00E522B3000562082D",
INIT_0C => X"90D0490D2C90D0C90D2C90D0C90D2490D04486124868294032384890B8985534",
INIT_0D => X"184014960000008402028041005232001715A040820B11A401E2443243450D04",
INIT_0E => X"9306260000554015520481040100004504A08110000820440001009134000004",
INIT_0F => X"02000000001014000028052000400028040050052000400028040200501C8D38",
INIT_10 => X"4002000000000068005005200040002804002805200040002804000E00001000",
INIT_11 => X"0028400010008000000000102800009800601000040000000011820002140102",
INIT_12 => X"4022010110000000D00008310000801080102000A00004000000000009020000",
INIT_13 => X"00001A00C0082400000006802500008000000000080048000060041200000003",
INIT_14 => X"A000005400080600000000000850000014200411000000000010024440202200",
INIT_15 => X"0000000008840600002080200000000000021800000013000040000000000020",
INIT_16 => X"40902449022A800800002208090684819402120AA8001C800000000000100014",
INIT_17 => X"1902409024090240906419064190641902409024090240906419064190641902",
INIT_18 => X"9044190440900409004090041904419044190440900409004090641906419064",
INIT_19 => X"7D402A2953F81F81F83F03F03F04190441904419044090040900409004190441",
INIT_1A => X"4104104104104104609D21808205965965D65801004E35C300C2D50A22B1C50C",
INIT_1B => X"128944A25128944A25128944A250410410410410410410410410410410410410",
INIT_1C => X"FFFFFFFFE3F00944A25128944A25128944A25128944A25128944A25128944A25",
INIT_1D => X"100055400000000000000000000000000000000000000000000001E1F007FFFF",
INIT_1E => X"400FF843DF45FFAEBDF55082A82155082AAAA10F7FFEAB455500175FF5D2A800",
INIT_1F => X"ABEF082ABDF455D7BD5545F7D5574BAFFD16AAAAA28428ABA000428AAA5D7FD7",
INIT_20 => X"EAB455D7BEAABA5D2A97545552E975FFFFD168AAA5D7BE8BFF5D557FFEFFFD16",
INIT_21 => X"A955555555555FFA2AE820BAFFFFEAABA5555554BA5D0417545F7D56AAAAAAFB",
INIT_22 => X"002AA00AAAEBDFFF08042AABA087BD54BA08043DEAAFF843FF5508517FF55552",
INIT_23 => X"02A82010AAD1401FF002EBFF45A2FBFDFEF00042AA00AAFBEAB5500003FF5500",
INIT_24 => X"0000000BA0004155550004154105D556AA00A2FBEAABA085542145082A800BA0",
INIT_25 => X"D5500155FF552A87410007145400000000000000000000000000000000000000",
INIT_26 => X"9208002FABA4171D5400FF8A38F45F7AABA57D0000855FD1C2AAFA00EBA5E8B7",
INIT_27 => X"A92555178FD7BFD5FDFFA0020BFF78417BD5545F7F1554AAF7D16DABABFF57DE",
INIT_28 => X"756DFFDF6DAAAAAF1EFB6D417BEFA901C2E97F40552E975EFEBDF68ABA557BEA",
INIT_29 => X"2DB7DA3FBD21C7492E9256D555B555C7A2ABC20AAE3AABAE38005B574AA49041",
INIT_2A => X"5EDB7D1E803AF6D400028E02AB8A3A012540E2AABABC75D043A00003FE10E380",
INIT_2B => X"0EB8B7D0AAA800AA147085000FFDA001C7B47BFABC7BFFF7AB4714042AA38BEF",
INIT_2C => X"000000000000000000000000821E8A10568005A1041055716DA38B6FBEFFEF1C",
INIT_2D => X"5D2EBDE00AAC16ABEF5500155EF552A954000855544000000000000000000000",
INIT_2E => X"AF7D57DE0AFAD1EBEB400043DEAA085555400FFAAAAB55F7AEA8BF77004147EF",
INIT_2F => X"EFAAFBEABAF557FEA8515951E8B4D83D1EBDFF082CBDFEF005756145FFD5574A",
INIT_30 => X"E005951550100004155EFF7FFFDE08AA557FFFF083FFCEB95104210405D2E955",
INIT_31 => X"00AA002A3FE18AE803CBE7A3C014351082E951FF5D7FD6145AAAA820A2AAAD29",
INIT_32 => X"EAD45550028ABAFFD17FFED01001FFEF5542ABEB2AA848AAA2552EA8ABA75514",
INIT_33 => X"57FEBAF3F95EEE95C00B7CF12AAA800BA551417105FFFFC21555556EAB4CD6D5",
INIT_34 => X"00000000000000000000000000000000000000000187782001FF0812000A255D",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0400000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(2),        -- Port A data input
DOA(0)   => data_read_a_lo_256(2),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(2),        -- Port B data input
DOB(0)   => data_read_b_lo_256(2),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_3_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"210C00A20020000108430020001600B8156021104940741B3530400E02B92202",
INIT_01 => X"A00C9BC058B00968240402C992000B61404040028804A0080A000D16A8990A08",
INIT_02 => X"4809A902031800444445089866E331352180D468B8200E600C0081110B80ACD0",
INIT_03 => X"6D0A601008000142B1A30A040AC68428320006010A80881068A80D401C846330",
INIT_04 => X"482218076809C03B24841CD92CDD5A4402091278072948042640102107102D04",
INIT_05 => X"0B063006A6402109000104E40B04644B32A86D20014A0D204063296082000E34",
INIT_06 => X"01072010703402800606D0102800CAB31434442810B4858060D0500008C52828",
INIT_07 => X"8C00222420A14204E01C581091020CC8000E3226413990008D80001A00CCC4AA",
INIT_08 => X"0874732009120665255420184000220002843E14294258E805E0116002D95101",
INIT_09 => X"BA546AC411102029A61C974014EDBA1320B1046100C0B4034928002002211145",
INIT_0A => X"1052088250A1CC2041051913208CE802438000082040008000F399406BC07998",
INIT_0B => X"19E416590908884D00020242A500090801806801041358222302084204460020",
INIT_0C => X"1019010190101B0101B01019010198101B20805C080C880080506990125E0514",
INIT_0D => X"03400040A101C05C0088242D0000320013339310018011A044414400400101B0",
INIT_0E => X"6514CA601CCCC8B33204C0401104244000018380818040A07060090000280009",
INIT_0F => X"0000000000020000006000000000020000011000000000020000010072CC9251",
INIT_10 => X"0000000000010000014000000000020000013800000000020000010700000000",
INIT_11 => X"002C000000000000000000010000001A00000000000000000040000002440000",
INIT_12 => X"00B2000000000010002049910000011000500000000000000000008000000000",
INIT_13 => X"00020005500000000000800133000000000000000010000000C0000000000040",
INIT_14 => X"0000005300000000000000001000000110600000000000000000401540000000",
INIT_15 => X"8000000008200620000000000000000000400000000107000000000000000004",
INIT_16 => X"0280C0280C0205104100000A8D06C404440230B9980210020040000010010003",
INIT_17 => X"280C0280C0280C0280803808038080380803808038080380C0280C0280C0280C",
INIT_18 => X"80E0200C0280E0200C0280E030080380A030080380A030080380C0280C0280C0",
INIT_19 => X"291008A004D54AAB556AA9556AA830080380A030080380A030080380A0200C02",
INIT_1A => X"4904104104104104A20E85800004924924054C0F031E31C190A285040164C586",
INIT_1B => X"1A8D46A753A9D4EA753A9D4EA752492492492492492492492492492492492492",
INIT_1C => X"FFFFFFFEB6FECD46A351A8D46A351A8D46A351A8D46A351A8D46A351A8D46A35",
INIT_1D => X"00AA8400000000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"B455500175FF5D2AA8A10005540155087BEABFF552ABDF45A2D16AAAAF7D5400",
INIT_1F => X"201000556AB55552ABDE00AAD140010F7D17FF45A2AA82155082AAAA10F7FFEA",
INIT_20 => X"42155557FEAA10007FEAABA000428AAA557FD7400FF843DE00FFAEBFF55082A8",
INIT_21 => X"AA8A105D7BD5545F7D5574BAFF802AA00A2D168ABA085568BEFFFAE820000855",
INIT_22 => X"557FFEFF7D56ABEF557BD74BAFF8402145A2AEBFFEF552EAAABA5D0028BEF082",
INIT_23 => X"5043DEAAAAAA95410F7803FFFF55556AAAA552A975FFFFD16AAAA5D7BC01EF5D",
INIT_24 => X"0000000105D0417545F7D56AAAAAAFBEAB455D7BEAABA5D2A974005D55574005",
INIT_25 => X"5B6DF6FABAFFD547010AA8407400000000000000000000000000000000000000",
INIT_26 => X"6D1C2AAFA28EBF5E8B7D5500155FF552AAF0100071455451C75EABC74174BAF5",
INIT_27 => X"F45F7AABAF7D00009543D1C556AB6D4124BAE10BED542010FFD57AF55AAF5D75",
INIT_28 => X"ABFFEBA0870281C5F4716D5D7FEDA3A0955FF48208002FABA4171D5400FF8A38",
INIT_29 => X"B8EBA15203FFFF002AAFA384171D5545F7D0154AAF7D16DABABFF57DE92005F6",
INIT_2A => X"F68ABA417BC01D7555178FD7BFD5FDF571575D24BA438E021D5B6A4BAFFF5D2E",
INIT_2B => X"24BFE005D5B52428410E3AE92E3A490410EB843ABD71551FFE02552A975FFEBD",
INIT_2C => X"0000000000000000000000003849041756DFFDF6DAAAAAF1EFB6D417BEFBD71C",
INIT_2D => X"5D556AB45081028B55FFFFFFEBAFFD557400A280144000000000000000000000",
INIT_2E => X"0FFD56ABF5AAD15455F5D2EBDEAAA2D16ABEF5500175EF552ABDE00085554545",
INIT_2F => X"AA085555400FFAAAAB14F7AE28BF77004146BA557DEABEF00002BE10FFD54000",
INIT_30 => X"E0AF2D1EAEBA007FEABEFAA84174BA557FD55EF5D3BFEEB35055DEE1000043DE",
INIT_31 => X"0155FFAA28BF7592EABE0A0804ABFFB082EBDEAA005556145FFD5574AAF7D47D",
INIT_32 => X"EB8105D2E955EFAAFBE8AAA547FE21550853E8B4FABD5EBFF75D55420AA82AA8",
INIT_33 => X"57FFFF087FFCEF90104B780A557FC20AA082AAAE10AA8000000A2AC2ABFD2151",
INIT_34 => X"00000000000000000000000000000000000000000AA0004155EFF7FFFDE08AA5",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(3),        -- Port A data input
DOA(0)   => data_read_a_lo_256(3),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(3),        -- Port B data input
DOB(0)   => data_read_b_lo_256(3),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_4_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10804002061080A284201081034809800A002303500078B3432C82904204002",
INIT_01 => X"810398000008004C0420050E12100368403008418984014902030806A0910204",
INIT_02 => X"480108A000000000446448E01E80F00A41043118680402000800000009882390",
INIT_03 => X"065040108C0000408406080002101020260012E03000000030808902088000F0",
INIT_04 => X"9100EB8368155C1AE0B01CD60433B944028A90385AC0D438E02010E81C32E801",
INIT_05 => X"B81E4166DE080029204044C401041C4CF01C489433483C8042EAC190100074C4",
INIT_06 => X"400F0400688002A22010D4342045C50F0004028993B3A5260041E4500EB4C0E2",
INIT_07 => X"000000243020008461000812810003C300060064012E00048C82005800BC2888",
INIT_08 => X"08CC8F0109064220240410008000002202043E44001048000020114000881000",
INIT_09 => X"F0DC1EB5131020C7BE7D172251E53E80E891E5016041B4083945202002419104",
INIT_0A => X"7D6025AC2A0982500302003200872003FB108808280200204400786612CE2B08",
INIT_0B => X"11D0025980480A458100930201820964408268101000F022D8083B4044A0002C",
INIT_0C => X"90C3490C1490C3490C1490C1490C3490C104869A48618800B66305989ABA0434",
INIT_0D => X"220000000500021002100088004010001370F030808110204581043243050C54",
INIT_0E => X"06100C40903C1C30F20025440102200541204090600830045825050034010000",
INIT_0F => X"000000000012000000BC04000000020004018C040000000200040000721CD861",
INIT_10 => X"000000000001002001A40400000002000401DC04000000020004014D44001000",
INIT_11 => X"0065040010000000000000110000007600200000000000000050000005D40002",
INIT_12 => X"00DE00001000001040004A3B0000180088500000200000000000008000020000",
INIT_13 => X"0002080760000400000082024300008000000000081006000170000200000041",
INIT_14 => X"180002B200000200000000001806000192000010000000000010401F80000200",
INIT_15 => X"0814000114A00200000000200000000000401006000085C00040000000000024",
INIT_16 => X"40102459044481081044880A0986D4C1560636C7840A61803000820012113042",
INIT_17 => X"1900411064090041102409044110240900401064190040106409004110640904",
INIT_18 => X"9064090240100411044090241902401044110041902409064110241904401024",
INIT_19 => X"04048028064B261934D964C3269C090641100401044090641902401044010041",
INIT_1A => X"AA8A28A28A28A28A74C132343334514513028A2818E01F81400050E130106345",
INIT_1B => X"8341A0D46A351A8D46A351A8D46AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA",
INIT_1C => X"FFFFFFFE58C001A0D068341A0D068341A0D068341A0D068341A0D068341A0D06",
INIT_1D => X"10550015400000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"F45A2D16AAAAF7D568A00AA8400000AAFFC21FFF7D542000FFAE821FF552EAAA",
INIT_1F => X"0000AAAE820BA550015400087FD74BAFFD540000F7D155555087BEABFF552ABD",
INIT_20 => X"A8AAAF78015545FFD555555082AAAA10F7FFEAB455500175FF5D2AAAA1000554",
INIT_21 => X"56AB45552ABDE00AAD140010F7D17FF45A2FBC2000A2FFC21555551554005D2E",
INIT_22 => X"AEBFF55082E82145A280001EFF78402145A2AE801555D2E95555552E97410005",
INIT_23 => X"D517DF45557BD5410F7D555545F7AA97410000428AAA557FD5400FF843DE00FF",
INIT_24 => X"0000000AA085568BEFFFAE82000085542155557FEAA10007FEABEFAAD1400AA5",
INIT_25 => X"8EBAA801EF4920AFA10490A17000000000000000000000000000000000000000",
INIT_26 => X"451C75EABEF4124BAF55B6DF6FABAFFD56F010AA8407428A2F1C01FFF7D14202",
INIT_27 => X"5FF552AAFA10007155428A2AE850925D0010400087FD24AAE3DF47010E38E051",
INIT_28 => X"01555D51524004920ADA82EB8A12555EBFB4717D1C2AAFA28EBF5E8B7D550015",
INIT_29 => X"92555492A850381C5F6AB6D4124BAE10BED542010FFD57AF55AAF5D7410A2FBC",
INIT_2A => X"1D5400FF8A38E00F7AABAF7D0000955FDB684051D7F7840517DA2A4871554124",
INIT_2B => X"55D75EFBED5400825D557FF55007BD7410EBDB5017DE38E8708008002FAAA417",
INIT_2C => X"00000000000000000000000082005F6ABFFEBA0870281C5F4716D5D7FEDB7D09",
INIT_2D => X"AAD1401FFFFD5420BAA2AA821FF08043DE10002A964000000000000000000000",
INIT_2E => X"AA2FBD7410A2AE965555D556ABEF080028B55FFFFFDEBAFFD57FE00A280144BA",
INIT_2F => X"AAA2D16ABEF5500175EF552ABDE000855544AAAA82174105D0402000087FC00B",
INIT_30 => X"BF5AAD154400AAFBC015555554001008003FE00AAEA81154AAFFD65FF5D2EBDE",
INIT_31 => X"75EFA2AA155550004021E5582A964BE557FEABEF00002BE10FFD540000FFD56A",
INIT_32 => X"9661000043DEAA085555400FFAAAAA10F7AC28BF558001454DF78017555F7801",
INIT_33 => X"FD55EF5D7BFEEF35055487EFF7D1400105D517FF55087FD7410A2FBC01E7F2AE",
INIT_34 => X"0000000000000000000000000000000000000000010007FEABEFAA84174BA557",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0400000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(4),        -- Port A data input
DOA(0)   => data_read_a_lo_256(4),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(4),        -- Port B data input
DOB(0)   => data_read_b_lo_256(4),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_5_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50DF0A0791B3FC1694378283C81FD996A091A32152007AB36B20E03C040C006",
INIT_01 => X"081FBDC49830884C5C6A60000C34C24841280A00084000C8C212892EEA953231",
INIT_02 => X"C809AD5CB118E640A4F008F8011FF0002080000082CCC66609DB7DDDCB1F2036",
INIT_03 => X"25080626BE4C904210831C80084204720B20048A88800000B8E0F8102885500E",
INIT_04 => X"4005122024899100064520C01444429C7804103C0416C007198A3916E0551A04",
INIT_05 => X"46E1829941C9000944C8C022898FE2F20D7D7A104CB5C208E51417C054848912",
INIT_06 => X"CA075CA0E63342991612DF9A8205C0A0B030B20B10480900886E220801073711",
INIT_07 => X"8C732074B68D1A34E3180717FFD13FC72691924098712CE481FDC241D43C1ACD",
INIT_08 => X"16053F180A1286A4E51BD18840C320000075FE91A24458BA4DE0D57992D9BE58",
INIT_09 => X"0A4D8105BF3472304100930258E510601EDE1D8524309285FD416CB402259504",
INIT_0A => X"3110AC0D11C901B2112109204C28B67061E8928920CAD3CFC0140079065A4A65",
INIT_0B => X"C3404959321C284D356A964F8125CD7AC8632614005DFBAACFBC800024091128",
INIT_0C => X"380D6380B6380F638096380F6380B6380D51C04B1C07AD10C14020D233127AD5",
INIT_0D => X"992940513052F4CA8A0A0664A5023CA8470FF000908C383755AF1604E0538096",
INIT_0E => X"200040194FFC044FFA4B08BC85282C91F028D094284A34054A25508605135C01",
INIT_0F => X"BA0C2038ABACBC7C7806F94FF87C002F83F106F94FF87C002F83F2000A04C200",
INIT_10 => X"8D9A70380230F2DFC106F86FF87C002F83F106F86FF87C002F83F3601BFFEBC2",
INIT_11 => X"1F401BFFE7C69E01804E1E6EABE3F040FFD7C7C4BC0E008C7C2FE58FC0A9FFF5",
INIT_12 => X"F8BFDFC8C8120C4DBC802208B2EB2AE777ADFE6F0A47CC0600C2683E0FF8AE3F",
INIT_13 => X"4189B7C56DF47186104C6DE7037FFF00FC0000FC07EE4E7A7076FE28C3082636",
INIT_14 => X"B9E9F272FFFC181C0C2038A7C6DE7A7D909FBFA4070380131CAFB257FBD93902",
INIT_15 => X"2B34E9F56DFBEB1B7F2300C4A80092E0FC1FCE667A7C877FFE828F0080AE1DDA",
INIT_16 => X"51142511405EA00A1344612A898494801602081F87204A9452217159891640D4",
INIT_17 => X"0942511425014450940519425114650140519405194650146511405194050946",
INIT_18 => X"1465114250146501465194051944509445094051146501465014251140509445",
INIT_19 => X"7ED430A983124B2DA6924965B4D5014650142511425094450940519405094450",
INIT_1A => X"EFBEFBEFBEFBEFBE5FDFF3F7F773CF3CF7D796ED39FDEE76DFFCE9F84801B6DB",
INIT_1B => X"BDDEEF77BBDDEEF77BBDDEEF77BBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFB",
INIT_1C => X"FFFFFFFE433B5EEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77B",
INIT_1D => X"AAFFFBFFE00000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"000FFAE821FF552E820105500155555D2AA8A00AA843FFFFF78002155AAAE974",
INIT_1F => X"0000FFAE80000AAAE974BAFFAEAAB45AAAEBDEAAA2FFEAA00AAFFC21FFF7D542",
INIT_20 => X"7FE000055574BA557FFFF55087BEABFF552ABDF45A2D16AAAAF7D56AA00AA840",
INIT_21 => X"E820BA550015400087FD74BAFFD540000F780155555D7BE8B45085168BFFA2D1",
INIT_22 => X"2AAAA10005140145FFFBC01EFAAFFD75FF002E97555A2AABDEAAAAAAAAA00AAA",
INIT_23 => X"A84174BA5D043FF45AAAA974AAF7AEBFF55082AAAA10F7FFEAB455500175FF5D",
INIT_24 => X"000000000A2FFC21555551554005D2EA8AAAF78015545FFD555410552EA8BEFA",
INIT_25 => X"FFF8E0217DBEA4954AAE3FBFDE00000000000000000000000000000000000000",
INIT_26 => X"28A2F1C01D7F7D142028EBAA801EF492087A10490A171455D2EADA28B6803FFF",
INIT_27 => X"ABAFFD56FA10AA8417428E3AE87010A2A4974AAE3AEAFB6DAAA4BDEAAA2F1EDA",
INIT_28 => X"8B6D14516DBD7BEDB7DE381451554AA497FFFF451C75EABEF4124BAF55B6DF6F",
INIT_29 => X"BDEAAAAA0AFA28A2A4850925D0010400087FD24AAE3DF47010E38E0516D5D7BE",
INIT_2A => X"5E8B7D5500155FF552AAFA10007155545F7F1C21D7AAF1D55FF082A9057DA2AA",
INIT_2B => X"FB470384124ADBFFBE84174AA55043FF6DBEAE950AAEB8ABDF7D1C2AAFA28EBF",
INIT_2C => X"00000000000000000000000010A2FBC01555D51524004920ADA82EB8A12410EB",
INIT_2D => X"552EBFEBAF7843DFEFF7AE801EFF780174AAAAFBFEE000000000000000000000",
INIT_2E => X"FA2803FEBAAAD17CEAAAAD140155FFD5420BAA2AA821FF080415410002A96555",
INIT_2F => X"EF080028B55FFFFFDEBAFFD57FE00A280144AAA2AA97400A280174AAA2AEBDFE",
INIT_30 => X"410A2AE965FF557FE8BFF55557FF55FFFBFFEAA5D51554AA087BFEF555D556AB",
INIT_31 => X"55FF0004821FFAAAEBDEAAAA843CEAAAA80174105D0402000087FC00BAA2FBD7",
INIT_32 => X"BEFFF5D2EBDEAAA2D16ABEF5500175EF552ABDE00005554545F7D140145A2D55",
INIT_33 => X"03FE00AAAA81114AAFFD64BA00043FFFFFF80174AA55043DFFFFFAE974BAA2AE",
INIT_34 => X"0000000000000000000000000000000000000000000AAFBC0155555540010080",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"1800000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(5),        -- Port A data input
DOA(0)   => data_read_a_lo_256(5),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(5),        -- Port B data input
DOB(0)   => data_read_b_lo_256(5),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_6_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10844B0061A258A2840112C03002C18000402322520070B303301C0381A0086",
INIT_01 => X"0600404820094048008100000042026041000000090800090210080008510204",
INIT_02 => X"080108220C1000004440080000C008010000000001203240080080000988A050",
INIT_03 => X"040000000823404000020A600000002983800584488000103080040C08C00000",
INIT_04 => X"00101610A029B08400044800000000040000102A040810040400100500101800",
INIT_05 => X"05000000800C8300306420002900404400820000000A00804004084001200A00",
INIT_06 => X"64472644640C00808C10D00401823F0020204209101001002650020001052800",
INIT_07 => X"080000242000000461100050818080380900224000200008818028804883E10A",
INIT_08 => X"01FE80E0090242602C0020608000000000043E00000048800021140000881106",
INIT_09 => X"12447E041B102020208000424029006FE0B085013204D0200101006862119140",
INIT_0A => X"4D540B0D916BBE39059191200000200441040108000020006FC5FA6000816908",
INIT_0B => X"8BF05D11A20808454010834225A28962E40AA05510180022FFA6A8800402A06D",
INIT_0C => X"16C1416C5416C5416C3416C3416C7416C500B60A0B60AD04EB4104C093904535",
INIT_0D => X"59802817888180E80112A1660050900003400430CB4911B445A105B05B016C14",
INIT_0E => X"000000062003C90000442006439324280034E85A742D1A16CD2DA30046848048",
INIT_0F => X"00000000000157000600000000000028000C00000000000028000CE800048000",
INIT_10 => X"00000000000000483C00000000000028000C00000000000028000D1080000000",
INIT_11 => X"00108000000000000000000078000A00000000000000000000019A0030000000",
INIT_12 => X"4604000000000000934909080014000000000000000000000000000009005180",
INIT_13 => X"00001230B00000000000049B3C000000000000000001FA000C98000000000002",
INIT_14 => X"E8000E05000000000000000001720002A56000000000000000000FC080000000",
INIT_15 => X"0840000B000404A000000000000000000002099A0003B0000000000000000001",
INIT_16 => X"69DA5685A146D19D084488080904C0A1172240C0781400C81908000205208614",
INIT_17 => X"85A1695A769DA3685A169DA768DA1685A169DA7685A1685A769DA7685A168DA7",
INIT_18 => X"5A368DA1685A769DA168DA3695A569DA3685A169DA5695A368DA1695A569DA36",
INIT_19 => X"7F10800846638C31C71C718638E685A769DA5685A3685A569DA7685A168DA769",
INIT_1A => X"E38E38E38E38E38E76DDB3B7B377DF7DF7D7DE2F39FE3FC3D3EA55FF37F5F7CF",
INIT_1B => X"9FCFE7F3F9FCFE7F3F9FCFE7F3F8E38E38E38E38E38E38E38E38E38E38E38E38",
INIT_1C => X"FFFFFFFF61AC8FE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F",
INIT_1D => X"EFAAAABFE00000000000000000000000000000000000000000000181F007FFFF",
INIT_1E => X"FFFF78002155AAAE974AAFFFBFFE10F7FBE8BEF552E95555552EAABEF082E975",
INIT_1F => X"5410A2AAAAA10087FC01EF552EAAB45F7AE821550851555555D2AA8A00AA843F",
INIT_20 => X"2ABEFA2AEBDFFF552AAAA00AAFFC21FFF7D542000FFAE821FF552E8001055001",
INIT_21 => X"E80000AAAE974BAFFAEAAB45AAAEBDEAAA2FFEAB45552E800AA555568A105D00",
INIT_22 => X"D56AA00AA8400000007BC21FFAA803FFEF5551420105D5568B45FF8400000FFA",
INIT_23 => X"7FBC2155007FC20BAA2D5575FF087FFFF55087BEABFF552ABDF45A2D16AAAAF7",
INIT_24 => X"0000001555D7BE8B45085168BFFA2D17FE000055574BA557FFFE10F7AAA8A00F",
INIT_25 => X"D4924ADBD70820975FFA2A4BFE00000000000000000000000000000000000000",
INIT_26 => X"455D2EADA28B6803FFFFFF8E0217DBEA4954AAE3FBFDE38F7FFEABFF412A9056",
INIT_27 => X"1EF492087010490A07038B6A0AFA38007BC51EF4920AFB55EBA4851450855555",
INIT_28 => X"5082555F68A3855002FBC7BEA4BFFFF492EADA28A2F1C01D7F7D142028EBAA80",
INIT_29 => X"6DB45E38A07028E3AE87010A2A4974AAE3AEAFB6DAAA4BDEAAA2F1EDB55492A8",
INIT_2A => X"4BAF55B6DF6FABAFFD56FA10AA84174381C7FC01C7B68E3DFC75555400105D51",
INIT_2B => X"7FFFE38F7A0AFA38E3FFC21450071C2092A2D5571FF0851FDF451C75EABEF412",
INIT_2C => X"0000000000000000000000016D5D7BE8B6D14516DBD7BEDB7DE381451554AA49",
INIT_2D => X"F7FBEABEF002E801EF00003FF550800155FFA2803CE000000000000000000000",
INIT_2E => X"5A28417555085154555552EBFEBAF7843DFEFF7AE801EFF780174AAAAFBFEEAA",
INIT_2F => X"55FFD5420BAA2AA821FF080415410002A964AAFF803DEAA087FD55FF00043DF4",
INIT_30 => X"EBAAAD17CF55002E95410557BEAABA55043DF55F7803FFEF002ABEEAAAAD1401",
INIT_31 => X"DF455D51420105D517DF55AAAA964AAA2AA97400A280174AAA2AEBDFEFA2803F",
INIT_32 => X"7CF555D556ABEF080028B55FFFFFDEBAFFD57FE00A280144BA5D7FC2155FFAAB",
INIT_33 => X"BFFEAA5D51554AA087BFEEAAF7803DEAAAAFBC0155085540000A2D5575FF0851",
INIT_34 => X"00000000000000000000000000000000000000001FF557FE8BFF55557FF55FFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"1200000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(6),        -- Port A data input
DOA(0)   => data_read_a_lo_256(6),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(6),        -- Port B data input
DOB(0)   => data_read_b_lo_256(6),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_7_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10844B00482258A2842112C02450418800002300500030B303300C018180002",
INIT_01 => X"0200084020084048040080000201026040000000080000080200090000510204",
INIT_02 => X"4801082048100000444008040080000041000000000222400800000009000010",
INIT_03 => X"0401018108A144D0000208424000002103006480088000003080000408C10000",
INIT_04 => X"0000120022419000000C80000000000400201829040000050001940400301820",
INIT_05 => X"04000000800840092CC080214144004400000000000800065004004020220800",
INIT_06 => X"40870408600000808C10D4500080008020200008001001000240000061052002",
INIT_07 => X"08000024200000046010005281848001494020400031240C8C8238A06A000988",
INIT_08 => X"40050001090242602C0408408000000000243E00000048800020154000881024",
INIT_09 => X"024401041B132820000011424069004000B20403200891420101026A42210440",
INIT_0A => X"013800A0281400300C0010200008B20663970148004424006818026200004800",
INIT_0B => X"01C1103022881845421082C2C0082300401121810012004600001010040028A0",
INIT_0C => X"1200112001120011204112041120411206089010890100408040008012101414",
INIT_0D => X"09146817802988694902A02451109006230006E0808294008C02848148092001",
INIT_0E => X"000000042C00040002000004020020490020401020081004482501010C120948",
INIT_0F => X"0130C807144102420700052000003C00780B00052000003C007808450484C000",
INIT_10 => X"400002C0E00E0D003300052000003C00780B00052000003C0078099080001000",
INIT_11 => X"80908000100000661801E18042100E000060100000B038038380124038000102",
INIT_12 => X"053A010111848322020512000414400000002000A1001058300C0741C0054120",
INIT_13 => X"90644029D008240864231011BF00008000C3C003F00186040EE8041204321188",
INIT_14 => X"18100D770008060130C807182106040375600411004C2600E3400C2740202230",
INIT_15 => X"9094100A8CA406A0002C812240B0201F0380211604037740004010472041E201",
INIT_16 => X"40100401006E8118104428088904C4C414420080049450801000088444300601",
INIT_17 => X"0906409004010040104409024090240906401004010040102409024090240100",
INIT_18 => X"1024090241900401004090240902401004010040902409004010440100409024",
INIT_19 => X"004420A945841040002082080004110240902409004110040902409024110040",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFEDD9EC000000000000000000000000000000000000000000000000000",
INIT_1D => X"BA082AAAA00000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"555552EAABEF082E975EFAAAABFFEF002ABDF555D5157555F7FBC00AAAAD5400",
INIT_1F => X"FEAAAAAABDF55FFFBFDF55555568ABAAAD5401FF5D2AAAA10F7FBE8BEF552E95",
INIT_20 => X"400005D55554105D51401555D2AA8A00AA843FFFFF78002155AAAE974AAFFFBF",
INIT_21 => X"AAAA10087FC01EF552EAAB45F7AE821550851554AAF7FBFFEAA007BFFFEFF7D5",
INIT_22 => X"2E800105500155EF5D2EBFF450000020AA5D7BC0000F7D555545A28000010A2A",
INIT_23 => X"FAAA8A10FFD568ABAA2D56AAAAF7AABFE00AAFFC21FFF7D542000FFAE821FF55",
INIT_24 => X"000000145552E800AA555568A105D002ABEFA2AEBDFFF552AAAABAA2AE95555F",
INIT_25 => X"5E3F5C20BAAAD5420821C2EAAA00000000000000000000000000000000000000",
INIT_26 => X"38F7FFEABFF412A9056D4924ADBD70820975FFA2A4BFFFF1C2EB8F4555555054",
INIT_27 => X"17DBEA4954AAE3FBFDE82B6AEBAF55E3FFFAF55555F6FA92BED5421C75D20AAA",
INIT_28 => X"FE920075FDFD7F7D5400385D51504385D55401455D2EADA28B6803FFFFFF8E02",
INIT_29 => X"5057DB68E02038B6A0AFA38007BC51EF4920AFB55EBA485145085555492F7F5F",
INIT_2A => X"142028EBAA801EF492087010490A071EF4920B8F45140E07082417BC2000EBD5",
INIT_2B => X"2EADA92A2A09257DE3A4AAA10F7D16FAAABED56AE82F780BAE28A2F1C01D7F7D",
INIT_2C => X"00000000000000000000000155492A85082555F68A3855002FBC7BEA4BFFFF49",
INIT_2D => X"552EAAB455D5142155AAD1400AAA2D1420005D2EA9A000000000000000000000",
INIT_2E => X"0F7D1421555D042BAAAF7FBEABEF002E801EF00003FF550800155FFA2803CFFF",
INIT_2F => X"BAF7843DFEFF7AE801EFF780174AAAAFBFEE00F7AAAAB55AAFBEAB555D7BFDE0",
INIT_30 => X"555085154400FFD17FE1000517FF55FFD5420BA5D55400BA555543155552EBFE",
INIT_31 => X"5400087BC0000A2D5421EFF7AE810AAFF803DEAA087FD55FF00043DF45A28417",
INIT_32 => X"2BAAAAAD140155FFD5420BAA2AA821FF080415410002A965FF080428B45552A9",
INIT_33 => X"43DF55F7803FFEF002ABEE00A280001FFA28028A00FFD17DEAAF7D56AA10FF84",
INIT_34 => X"0000000000000000000000000000000000000000155002E95410557BEAABA550",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"01FFFFFFFFE00000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(7),        -- Port A data input
DOA(0)   => data_read_a_lo_256(7),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(7),        -- Port B data input
DOB(0)   => data_read_b_lo_256(7),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_8_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00000648E2840112C00000418000002700500030B3032000000000082",
INIT_01 => X"000009C21838284D1C2160000E12424840000000180800080200000040110204",
INIT_02 => X"080108000090000004400C040080000051000000000002400800000009000010",
INIT_03 => X"00000100043008D0000200024000000003800504488000103080880008800000",
INIT_04 => X"00009410A028A084000440000000000400001022040800150400808500321800",
INIT_05 => X"8500010080048A09302420202804400400800010200A00020204084011014A00",
INIT_06 => X"2447A244608800840490D0040007FE0021204288001000000050024001042800",
INIT_07 => X"4800002420000004201000D281040003182020400031241C0D80004041BFE88A",
INIT_08 => X"4005000108020220240000048000000000043E00000048800000010000881000",
INIT_09 => X"0204010519110020008111020069004008A28501120450220101214122509140",
INIT_0A => X"0528A52291490029019190200008B20E23008028000208804010024000004000",
INIT_0B => X"13C151312A8808454104824001280108A409A044001200020020989000000061",
INIT_0C => X"0000000000000000000000000000000000400020000229508040008012105400",
INIT_0D => X"48022817880508602102A1200810B2020340043248CA00240420000000400040",
INIT_0E => X"4100820020000C0000442142419120000014684A34251A12CD2CA30042840248",
INIT_0F => X"45F3D80000000001020404000783FC0000010404000783FC000000880284C010",
INIT_10 => X"02658FC7E0000000010404000783FC0000010404000783FC000001500000103D",
INIT_11 => X"40500000103961FE78000000000402400020003B43F1F8000000022010800002",
INIT_12 => X"0080001617CD800000080B000804080000020090659833F9F03C000000000000",
INIT_13 => X"B000000400018639EC000000000000FE03FFC00000000600840000C31CF60000",
INIT_14 => X"180204000001E2A3F3D80000000600802000401AA8FC7E00000000100002C2F5",
INIT_15 => X"005404020000104480DC372B47F060000000000600802000017570FF60000000",
INIT_16 => X"28CA328CA34650850A4C000009A494A015624080044440481908000220308640",
INIT_17 => X"8CA328CA328CA328CA3284A1284A1284A1284A1284A1284A328CA328CA328CA3",
INIT_18 => X"CA1284A1284A1284A128CA328CA328CA328CA3284A1284A1284A1284A128CA32",
INIT_19 => X"64108088440000000000000000028CA1284A1284A1284A128CA328CA328CA328",
INIT_1A => X"E79E79E79E79E79EDFC8F33637D6CB6CB2900A282950FAF15E8428917C51E75D",
INIT_1B => X"87D3E1F0F87C3E1F0F87C3E1F0F9E79E79E79E79E79E79E79E79E79E79E79E79",
INIT_1C => X"FFFFFFFECB0593E1F4F87D3E1F4F87D3E1F4F87D3E1F4F87D3E1F4F87D3E1F4F",
INIT_1D => X"10002ABFE00000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"555F7FBC00AAAAD5400BA082AAAA10000000010F7D5421EF007BC01FF5D7FFFE",
INIT_1F => X"FEAA5551554AAFF80021EF002A820BAFF8428A00A2AAAABEF002ABDF555D5157",
INIT_20 => X"E8BEFFFFFEAB55002ABFE10F7FBE8BEF552E95555552EAABEF082E975EFAAAAB",
INIT_21 => X"ABDF55FFFBFDF55555568ABAAAD5401FF5D2AAAB55FFD1400AA5D7FC01EFA2FF",
INIT_22 => X"AE974AAFFFBFFEAA08001555555516ABEFA280020AA5D043DF55557BEAAAAAAA",
INIT_23 => X"8042AB55005140145AAFFE8AAAF7D1401555D2AA8A00AA843FFFFF78002155AA",
INIT_24 => X"0000000AAF7FBFFEAA007BFFFEFF7D5400005D55554105D51400005551421EF0",
INIT_25 => X"71C7FC21EF5D75FFE10142EBAE00000000000000000000000000000000000000",
INIT_26 => X"FF1C2EB8F45555550545E3F5C20BAAAD5420821C2EAAA101C0005000E3D1401D",
INIT_27 => X"BD70820975FFA2A4BFE925D51554AAE384001FF142E800AAFF802AA28AAAEAFB",
INIT_28 => X"7092557BC21D7BEF5EDBC7FFF1EFB6D1420BAE38F7FFEABFF412A9056D4924AD",
INIT_29 => X"3AF55417BEDA82B6AEBAF55E3FFFAF55555F6FA92BED5421C75D20AAB45F7D14",
INIT_2A => X"03FFFFFF8E0217DBEA4954AAE3FBFDEAA1C001056D415F6ABEFA284020824904",
INIT_2B => X"55400385D51401EF00002FB45085F4016DAAF1EDAAAFFFB401455D2EADA28B68",
INIT_2C => X"00000000000000000000000092F7F5FFE920075FDFD7F7D5400385D51504385D",
INIT_2D => X"5D0417410AAD540155557FC01EF5D557DE105D2AA8A000000000000000000000",
INIT_2E => X"AF7842AABAA2AEBDFFF552EAAB455D5142155AAD1400AAA2D1420005D2EA9A10",
INIT_2F => X"EF002E801EF00003FF550800155FFA2803CE105D55574BAA280021EF5D2E820B",
INIT_30 => X"1555D042BB45FFD157410557FC0155F7D57FF55F7D57FFEF550028AAAF7FBEAB",
INIT_31 => X"8BFFAA8000000080428B55087FFFE00F7AAAAB55AAFBEAB555D7BFDE00F7D142",
INIT_32 => X"C2155552EBFEBAF7843DFEFF7AE801EFF780174AAAAFBFEEBA5D04021EF087BE",
INIT_33 => X"5420BA5D55400BA5555430BA5555421EF00043FF45007BC21FFA2D57FEBAF7FB",
INIT_34 => X"0000000000000000000000000000000000000000000FFD17FE1000517FF55FFD",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0800000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(8),        -- Port A data input
DOA(0)   => data_read_a_lo_256(8),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(8),        -- Port B data input
DOB(0)   => data_read_b_lo_256(8),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_9_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00018248A2840112C00002C18000002300500030B3032000000000006",
INIT_01 => X"000008000000004C0020000000100268413C0A61590001D90213C00000110204",
INIT_02 => X"680108200010000054400C040080000041000000010002400800800009082011",
INIT_03 => X"00040100000020D0000200124000000043800504488000103081880008800000",
INIT_04 => X"00001410A00AA084000400000200000400001020040010050020820400101880",
INIT_05 => X"0400040080048A09202420000C00410400000000000800020804004000000800",
INIT_06 => X"24478244640800840410D4144002008020200009301000000140000201042000",
INIT_07 => X"0800002C20000004301000128104000100002040003164040D80000040000888",
INIT_08 => X"40050003080202202400000080000000000C3E00000048800010230000881000",
INIT_09 => X"0024010411110420008010020021004000A204011200500001010000AA10C000",
INIT_0A => X"7945282804010009009090200008B20223800008020000004010024204000440",
INIT_0B => X"114100112208084540008240110001002400A000001000020008288000000420",
INIT_0C => X"010400100001040010000104001000010400080000820800000000801010100A",
INIT_0D => X"08403C16800100640182A0210010921003400412484202200400004004001040",
INIT_0E => X"410082002C000C000240004240932041401468CA34651A32CD28A22002840048",
INIT_0F => X"000000000000144002000420000000280001000420000000280000000284C010",
INIT_10 => X"4000000000000048010005000000002800010005000000002800001000001000",
INIT_11 => X"0010000010000000000000002A00020000201000000000000001820010000002",
INIT_12 => X"40BA00011000000090000B000004000000000000A00000000000000009000020",
INIT_13 => X"00001205D0080400000004803F0000800000000000004C0004E8001200000002",
INIT_14 => X"B000047700000600000000000054000135600011000000000000025740200200",
INIT_15 => X"001400020CA406A0000080200000000000020804000137400040000000000000",
INIT_16 => X"28CA328CA36651951A4CA8000984D4E557220080040440481908000001300614",
INIT_17 => X"84A1284A1284A1284A1284A1284A1284A1284A1284A1284A328CA328CA328CA3",
INIT_18 => X"4A1284A1284A1284A128CA328CA328CA328CA328CA328CA328CA328CA3284A12",
INIT_19 => X"2540A809010000000000000000028CA328CA328CA328CA3284A1284A1284A128",
INIT_1A => X"4534D34D34D34D344A2D840100E4920824055CD13333D2379A2A24018615C38E",
INIT_1B => X"268341A0D068341A0D068341A0D1451451451451451451451451451451451451",
INIT_1C => X"FFFFFFFE6DA90341A4D268341A0D069349A0D069349A0D068341A4D268341A4D",
INIT_1D => X"FFFFD557400000000000000000000000000000000000000000000001FFFFFFFF",
INIT_1E => X"1EF007BC01FF5D7FFFE10002ABFF55F7D168A00552E95555007BFFF55087BE8B",
INIT_1F => X"AA10F7FBC0145F7AE801EFF7FBFFF455D7BC0155F7D557410000000010F7D542",
INIT_20 => X"BDE00AA803FFEF5D55421EF002ABDF555D5157555F7FBC00AAAAD5400BA082AA",
INIT_21 => X"1554AAFF80021EF002A820BAFF8428A00A2AAAAAAAF7D17DE00FFFBD5555A2AA",
INIT_22 => X"2E975EFAAAABFFEF002A954BA5551421EF552E954105D00021455555420AA555",
INIT_23 => X"7D5575EFA2FFD75455D7BE8A005D5557410F7FBE8BEF552E95555552EAABEF08",
INIT_24 => X"000000155FFD1400AA5D7FC01EFA2FFE8BEFFFFFEAB55002ABFE10080028BFFF",
INIT_25 => X"D1C71F8F7D147BEFBEFEBD152400000000000000000000000000000000000000",
INIT_26 => X"101C0005000E3D1401D71C7FC21EF5D75FFE10142EBAF7DE3D16DA0041209056",
INIT_27 => X"0BAAAD5420821C2EAAA10E3FFC0145F7A0801FFEBFBF8F6D417BC716DEBD1524",
INIT_28 => X"DE28F7F5D0545B6AAB8E38B68A3AFFF5551471FF1C2EB8F45555550545E3F5C2",
INIT_29 => X"021455D5B470925D51554AAE384001FF142E800AAFF802AA28AAAEAFABAE3D17",
INIT_2A => X"A9056D4924ADBD70820975FFA2A4BFFFF082E974BA4155401C7552097428550E",
INIT_2B => X"20BAE0008002ABFFF7DB505FFAAFBD7555417FEFA00495B52438F7FFEABFF412",
INIT_2C => X"00000000000000000000000145F7D147092557BC21D7BEF5EDBC7FFF1EFB6D14",
INIT_2D => X"AAD17DE100804001EF55516ABFF557BFDFEFA2D5400000000000000000000000",
INIT_2E => X"F007FD55FFA2D5400105D0417410AAD540155557FC01EF5D557DE105D2AA8BEF",
INIT_2F => X"455D5142155AAD1400AAA2D1420005D2EA9A00A2FBC0145FF84001EFA2FFEABF",
INIT_30 => X"ABAA2AEBDEAAAAD17DEBAFFD142155FFAAAAABAFFAAAABFF5551555FF552EAAB",
INIT_31 => X"01555D00154AA552E801455D7BD54105D55574BAA280021EF5D2E820BAF7842A",
INIT_32 => X"C00AAF7FBEABEF002E801EF00003FF550800155FFA2803CFFF002E954BA00514",
INIT_33 => X"57FF55F7D57FFEF550028A10000428BEFF7FFC01FFA2FFD5545007BFDE10087F",
INIT_34 => X"0000000000000000000000000000000000000000145FFD157410557FC0155F7D",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"1000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(9),        -- Port A data input
DOA(0)   => data_read_a_lo_256(9),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(9),        -- Port B data input
DOB(0)   => data_read_b_lo_256(9),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_10_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000B0001800002840002C0000281800020030000000033122000400992006",
INIT_01 => X"A140098018300848180060000C00424040000000080000080200000000110200",
INIT_02 => X"0801080200100000046558000080000041000000002402400800000009008010",
INIT_03 => X"0001000084000040842242000210810803006400088000003080054288C10000",
INIT_04 => X"0000100022008000000C08000800000400A83A2044200C840000000400001820",
INIT_05 => X"0400000080000000248080210044000402000025000800000004203010100800",
INIT_06 => X"00078000600000040410D4102850008024240001981024A82000010461052000",
INIT_07 => X"0800002430204084281000128100000300002040003124040D80204040000888",
INIT_08 => X"0005000108020220240030008000000000043E0408104C800000010000881100",
INIT_09 => X"0004010511100020200000400021004008808060400111080000200002008400",
INIT_0A => X"0000000000010000060210200008B20223048808000200000010024000000000",
INIT_0B => X"03C0411009808245010002000028000080002105010000000020A34249020801",
INIT_0C => X"8004480044800048000480044800448000440002400221008840009012104400",
INIT_0D => X"0000540100000020088000000100100013000400000800040062400200440004",
INIT_0E => X"4100820020000400020000400200204900800000000000000000000100120800",
INIT_0F => X"0000000000101400020401000000002804010401000000002804000000048010",
INIT_10 => X"0000000000000068010400200000002804010400200000002804005000000000",
INIT_11 => X"0050000000000000000000102800024000400000000000000011820010800100",
INIT_12 => X"4000010000000000D00000080004080000002000000000000000000009020000",
INIT_13 => X"00001A000000200000000681000000000000000008004A000400040000000003",
INIT_14 => X"A800040000080000000000000852000020000400000000000010024000002000",
INIT_15 => X"0000000200000000002000000000000000021802000020000000000000000020",
INIT_16 => X"00000040002800100004200009048005C0000080000400000000000000200654",
INIT_17 => X"0802008020080200802008020080200802008020080200800000000000000000",
INIT_18 => X"0000000000000000000080200802008020080200802008020080200802008020",
INIT_19 => X"2054282101000000000000000000000000000000000000000000000000000000",
INIT_1A => X"A28A28A28A28A28A355950666151451453D51A242A503F834E5C49851D243555",
INIT_1B => X"994CA6532994CA6532994CA65328A28A28A28A28A28A28A28A28A28A28A28A28",
INIT_1C => X"FFFFFFFE8E31DCAE532994CA6532995CAE572B94CA6532994CA6572B95CAE532",
INIT_1D => X"AAFFFBC2000000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"555007BFFF55087BE8BFFFFD557400FF842ABEFA2AAA8B5500003DF55F7D568A",
INIT_1F => X"FE0008556ABFFA2D16AB550000021FFF7D17FFEF08042AB55F7D168A00552E95",
INIT_20 => X"3FF55A2D557400557BC2010000000010F7D5421EF007BC01FF5D7FFFE10002AB",
INIT_21 => X"BC0145F7AE801EFF7FBFFF455D7BC0155F7D557545FFAE820AA007BFDFEF5500",
INIT_22 => X"D5400BA082AAAA00FFAE820AAAAAABDFEFF78028BEF005140145A2842AA10F7F",
INIT_23 => X"AD56AB55A2D157400552EBFFEF5D7BD75EF002ABDF555D5157555F7FBC00AAAA",
INIT_24 => X"0000000AAF7D17DE00FFFBD5555A2AABDE00AA803FFEF5D55420BA08557FEBAA",
INIT_25 => X"51C0E3AF55F7DF68ABAE3F1C0000000000000000000000000000000000000000",
INIT_26 => X"7DE3D16DA0041209056D1C71F8F7D147BEFBEFEBD152400F7842FBD7B6AAAAB5",
INIT_27 => X"1EF5D75FFE10142EBAE0008556FBD7B6DB6AB7D1C0A001D7FFD178FC71C0E28B",
INIT_28 => X"2092147BFAFEF49043AF45A2DF504285D71C00101C0005000E3D1401D71C7FC2",
INIT_29 => X"4017DA28428A10E3FFC0145F7A0801FFEBFBF8F6D417BC716DEBD15256DF7AA8",
INIT_2A => X"550545E3F5C20BAAAD5420821C2EAAA00E3AA82092A2AABAFD7EB8A2ABC70855",
INIT_2B => X"51470821C557AE92A2DF6AB7DA2DF50410412ABDFC75D7BD55FF1C2EB8F45555",
INIT_2C => X"000000000000000000000000BAE3D17DE28F7F5D0545B6AAB8E38B68A3AFFF55",
INIT_2D => X"FF803DF45FFAEA8B555D2EAAB45F7FBE8ABAAAD5400000000000000000000000",
INIT_2E => X"5FFD168B55552AA8BEFAAD17DE100804001EF55516ABFF557BFDFEFA2D540010",
INIT_2F => X"10AAD540155557FC01EF5D557DE105D2AA8A0008557FF45FFFFE8BEF5D2E8015",
INIT_30 => X"5FFA2D5401FFF7AA800105D7FE8BEF08002AB45AAFFC00AA5D51400105D04174",
INIT_31 => X"AB55AAAEAAB450055421FFAA8428A00A2FBC0145FF84001EFA2FFEABFF007FD5",
INIT_32 => X"D55FF552EAAB455D5142155AAD1400AAA2D1420005D2EA9A10A2AA82010AAAEA",
INIT_33 => X"AAAABAFFAAAABFF555155400555568A10AAFBEABEFA2FFC0010082ABFF55557B",
INIT_34 => X"00000000000000000000000000000000000000000AAAAD17DEBAFFD142155FFA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"11FFFFFFFFE00000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(10),        -- Port A data input
DOA(0)   => data_read_a_lo_256(10),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(10),        -- Port B data input
DOB(0)   => data_read_b_lo_256(10),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_11_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10180B05A0010402840602C2D001019000000300000000330A20080EC180002",
INIT_01 => X"AB400984B83008481800E0000C26426040000000080000088200000802112220",
INIT_02 => X"8801081438106400A4F55800008000004100000040CCE24208005000C9060032",
INIT_03 => X"000406A492E6E440842254D002108153422004800880000030C0315688C00006",
INIT_04 => X"00001201200090001205400000000094108C322644240C840008030440111800",
INIT_05 => X"444000888008010028404002A002009402400025080880000C04223000170900",
INIT_06 => X"40871408620B00801410D94CAAD0018024242008A8102CA88A44010401042200",
INIT_07 => X"08320054B624408428100094ADD080011721A04000316C140CA1A8A1F9001889",
INIT_08 => X"140500090B02C2E0EC04D1C08000000000647E858A104C920C81A5011088A61C",
INIT_09 => X"002481041F165820000101024061004004800567603592A801014C4642601100",
INIT_0A => X"01002020000101B0070310200008B60A23A51B28020CE24E4010026004000440",
INIT_0B => X"03404110230CBA457670820140212100C0692644010001420038935269093161",
INIT_0C => X"2A0872A0C72A0872A0C72A0C72A0872A0C595043950421400800009010104280",
INIT_0D => X"8852141110244066C0820221480010AA73000420808CAC040464D280144050C7",
INIT_0E => X"410082022C000C0002020094030220C960A0409020481024482501A004014100",
INIT_0F => X"6DA02836090540355D86C046619A54052A5B86A0466196940631682800048010",
INIT_10 => X"8B68AA2C60289802AB86A046619A54052A5B86C04661969406316AC018B0E293",
INIT_11 => X"1FC09CB0E1076D4A200B2AC611A3D0405886C6EB211550815A8A2686EC81E2A4",
INIT_12 => X"9C0418CE0C5E8F650E48000892B37885620C1E1A06D7016A90A4626D82B10F1B",
INIT_13 => X"F1E164E02144D335546F28724001B030A56140A184483000C410A2699A2E32AC",
INIT_14 => X"415AAE8018A0A01B2990242E278056AAA203920E0BAE2012C08281808319C186",
INIT_15 => X"9B80D44F9051C049B18A12CB481042AD140C227002A0A02066954E7540CCDB58",
INIT_16 => X"4090240902468118104408000904C0C0964200800200108010003A02272400C1",
INIT_17 => X"0902409024090240902409024090240902409024090240902409024090240902",
INIT_18 => X"1004010040100401004090240902409024090240902409024090240902409024",
INIT_19 => X"2014002840000000000000000004010040100401004010040100401004010040",
INIT_1A => X"0020820820820820A069105251C00000015418982201060302C4281390042104",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFE0FC1C000000000000040200000000000000000001008000000000000",
INIT_1D => X"55000015400000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"B5500003DF55F7D568AAAFFFBC2010557BEAA10AAFBE8A00557BFFFEF007BC21",
INIT_1F => X"75455D7FE8BFF5D7FD540055003FFEFFFD142145000000000FF842ABEFA2AAA8",
INIT_20 => X"C0145557FC2010557FFDF55F7D168A00552E95555007BFFF55087BE8BFFFFD55",
INIT_21 => X"56ABFFA2D16AB550000021FFF7D17FFEF08042AB55A2AAAAB4508517FE00557B",
INIT_22 => X"7FFFE10002ABFE00AAFFE8AAAFF8402000550002145085555400F7FFE8A00085",
INIT_23 => X"8043FEBA002A975EFF7D17DFFFAA8000010000000010F7D5421EF007BC01FF5D",
INIT_24 => X"000000145FFAE820AA007BFDFEF55003FF55A2D557400557BC2145A2D1421450",
INIT_25 => X"8557BF8FEF1C7FC516D080E15400000000000000000000000000000000000000",
INIT_26 => X"00F7842FBD7B6AAAAB551C0E3AF55F7DF68ABAE3F1C00005D7BEDA00B6F1EFA2",
INIT_27 => X"F7D147BEFBEFEBD15257D5D7FEFBD7417BD5438550038FC7FFDF4216D080E070",
INIT_28 => X"DB4514517FE105575C216D5571C50104171FDF7DE3D16DA0041209056D1C71F8",
INIT_29 => X"52400FFF1EFA0008556FBD7B6DB6AB7D1C0A001D7FFD178FC71C0E28B6DA2AEA",
INIT_2A => X"1401D71C7FC21EF5D75FFE10142EBAE10A2FBEFA92F78A05028550E001451455",
INIT_2B => X"71C016DB6D54514500003FEBA1420905FFFFDF78FC7BE84050101C0005000E3D",
INIT_2C => X"0000000000000000000000016DF7AA82092147BFAFEF49043AF45A2DF504285D",
INIT_2D => X"5D7FFDE00F7D17FEBA557BEABEF557BD55EF082A974000000000000000000000",
INIT_2E => X"5F7FBC01FF082A97410FF803DF45FFAEA8B555D2EAAB45F7FBE8ABAAAD540010",
INIT_2F => X"100804001EF55516ABFF557BFDFEFA2D5401FF5D7FFDF55007BD74BA5D042AB4",
INIT_30 => X"B55552AA8BEFAAAABFF5555517FE005555401FF55515541000517FFEFAAD17DE",
INIT_31 => X"74BA5D2A801455D5140000FFD57FE0008557FF45FFFFE8BEF5D2E80155FFD168",
INIT_32 => X"174105D0417410AAD540155557FC01EF5D557DE105D2AA8A10AAFBFFE00F7AA9",
INIT_33 => X"02AB45AAFFC00AA5D51401FFFFD15555500003FEBA5D04001EFFFFFE8B55FF84",
INIT_34 => X"00000000000000000000000000000000000000001FFF7AA800105D7FE8BEF080",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"1000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(11),        -- Port A data input
DOA(0)   => data_read_a_lo_256(11),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(11),        -- Port B data input
DOB(0)   => data_read_b_lo_256(11),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_12_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50080B01BC002006940202C0DE041196A83183000000023322287E0FC000006",
INIT_01 => X"0E000C068000E04D40238000001702684000000008000008820009280A553231",
INIT_02 => X"2809AD0E7D180040945008040090000061800000C0E2F66009DA3D11CB148015",
INIT_03 => X"210D050012F6F8D2108216E24842005B8A20640008800000B8E0141C28851006",
INIT_04 => X"0080100022408000060DE0C00466630C70241837041000040800820480001AA4",
INIT_05 => X"04800018800000003C808003E0C8001401000000040900020904004000070800",
INIT_06 => X"00074000601300119E12D348438000803030800020100800AF08000261042400",
INIT_07 => X"8C53200CA4850224301807D1CB45900147E03040083124FC0CD0C8A1FF00198C",
INIT_08 => X"46050013081206A4A503A9E8C0812000001C7E11A24058B84D40E33992D98F7E",
INIT_09 => X"1004810491175C200000820018A5104010C01086003C13E000004EDF02040004",
INIT_0A => X"0000000000010000180018200408B27E234913E9004CFA09A818024800902109",
INIT_0B => X"014100580004304D267C06CCD0056600007827C00000008C00000000000219C0",
INIT_0C => X"2F0C32F0832F0832F0C32F0832F0832F0C197861978400040000208010120ACA",
INIT_0D => X"E0BF40403CFE7E03E8080382FD0018FE670004000006AE01180493C5BC1AF083",
INIT_0E => X"2000401EA0000440000800A0040028108000000000000000000000A74812DF00",
INIT_0F => X"C48DF8362F658A7E5F82CD23B6B0E403DBBE82C563B6A4E403DBB88C0E048200",
INIT_10 => X"454CFBE5403AB992F282C563B6B0E403DBBE82CD23B6A4E403DBBB1084E4B25A",
INIT_11 => X"851000E4B1D32BAB504BB74AD3F3FE04A8E0D0C319A7988B6F0C75CFD801A962",
INIT_12 => X"BEC4118D994B866E2E8C3808B6B63040328E7A33AF99B0AC20DE634D06C437BF",
INIT_13 => X"70CDC5F6214CA5991C6A7177402C49CA354D808D358A927EAD10A652CC8E3538",
INIT_14 => X"49F36E80083C3EAEB2003695430A7CDAA289553922990C11A4E494988231B325",
INIT_15 => X"3BC0FD5B304AD05A946D81616970A225658940BA7CDAA0A312666BD600E5550B",
INIT_16 => X"00000000001000000104200A89A4D0040000008003B81000000021CFEE02E280",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"8020080200802008020000000000000000000000000000000000000000000000",
INIT_19 => X"0544202101000000000000000000080200802008020080200802008020080200",
INIT_1A => X"4124924924924924481C040000B51451440146E518222204D82A5446021090CB",
INIT_1B => X"2C964B2190C86432190C86432190410410410410410410410410410410410410",
INIT_1C => X"FFFFFFFEF001D64B2592C964B2592C964B2592C964B2592C964B2592C964B259",
INIT_1D => X"00AAFBC2000000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"A00557BFFFEF007BC2155000015555087FC0010AAFBFFE100004020BAAAFFD54",
INIT_1F => X"2155AA8400000A2AABFF45550400000AAFBFFFEF550000010557BEAA10AAFBE8",
INIT_20 => X"C0010555155555FF8017400FF842ABEFA2AAA8B5500003DF55F7D568AAAFFFBC",
INIT_21 => X"FE8BFF5D7FD540055003FFEFFFD142145000000145A2AA821EFFFFFD7410007F",
INIT_22 => X"7BE8BFFFFD5574000051420BA557FC2145557FC20AAA2D57DEBAA2FBD55455D7",
INIT_23 => X"82EAAA00550415410AAFBFFFEF55042AB55F7D168A00552E95555007BFFF5508",
INIT_24 => X"000000155A2AAAAB4508517FE00557BC0145557FC2010557FFDE10AA84000000",
INIT_25 => X"0000A02092B6F5D2438A2FBC2000000000000000000000000000000000000000",
INIT_26 => X"005D7BEDA00B6F1EFA28557BF8FEF1C7FC516D080E1557D0075C7028B6F1FAE0",
INIT_27 => X"F55F7DF68ABAE3F1C017DAA8E07028B6A0BFF6D490E00000BEF5FAFEF4904070",
INIT_28 => X"51FFE3FBD0438007FC00385D555556DEB8410400F7842FBD7B6AAAAB551C0E3A",
INIT_29 => X"7DEBAA2FBD557D5D7FEFBD7417BD5438550038FC7FFDF4216D080E0716DAAA08",
INIT_2A => X"09056D1C71F8F7D147BEFBEFEBD152400005F450BA417BC51454971C20AAB6D1",
INIT_2B => X"71FDE10BE8E070280020AAA28410410400BEFBFAFEF49042AB7DE3D16DA00412",
INIT_2C => X"0000000000000000000000016DA2AEADB4514517FE105575C216D5571C501041",
INIT_2D => X"0055574BAFFD568A10002A82000FFD5400AAA2FBC00000000000000000000000",
INIT_2E => X"0FFD568BEF0004174105D7FFDE00F7D17FEBA557BEABEF557BD55EF082A975EF",
INIT_2F => X"45FFAEA8B555D2EAAB45F7FBE8ABAAAD5401EFA2AA974BAF7803FFFF002A8200",
INIT_30 => X"1FF082A975EFA280175FFAAFFC00BA087FC20AA5D55555FFA28000010FF803DF",
INIT_31 => X"75450851420BAFFD57DEAAAAFBD75FF5D7FFDF55007BD74BA5D042AB45F7FBC0",
INIT_32 => X"28BEFAAD17DE100804001EF55516ABFF557BFDFEFA2D540010007FD74AA007BD",
INIT_33 => X"5401FF55515541000517FE10F7AA954AA080428AAA000002010FFFFE8BEF0804",
INIT_34 => X"00000000000000000000000000000000000000001EFAAAABFF5555517FE00555",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"01FFFFFFFFE00000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(12),        -- Port A data input
DOA(0)   => data_read_a_lo_256(12),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(12),        -- Port B data input
DOB(0)   => data_read_b_lo_256(12),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_13_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10110A0441812402840402822007818000E00700000000330A3000000008042",
INIT_01 => X"A1400984B830C848180260000C0042404001000008220008A200100802110200",
INIT_02 => X"88010C02801040002475580400800000410000000064024608134C0CC9018034",
INIT_03 => X"00010100926220D084234212421085084300648A0880000630C0654288C10000",
INIT_04 => X"0004122122029100100C00001200009C40A83A2044360C84190BAC04E0101820",
INIT_05 => X"04E000008009050064C8C00104C10184034010250089C00EB004327064B60900",
INIT_06 => X"CA875CA8600000880410DA8C285001802424B008881024A8204E010461042700",
INIT_07 => X"08320014B02848A4A8100015C55500057801A04000712C040CB1F8806000088D",
INIT_08 => X"5005000908020220E40170008042000000557E048A144C800590010000882D00",
INIT_09 => X"00250104B5310020000100020821004016CC1C616401910801010100CA204000",
INIT_0A => X"0000000000010192072310200028B602234608080280074AC010025900100401",
INIT_0B => X"014100101118BA451000824150052110480121000140014200101352690BAC20",
INIT_0C => X"0000000040000000000000040000000000000020000000000000008010102A82",
INIT_0D => X"094040100000006C0802042501001C8017000C21908200028448400000000040",
INIT_0E => X"000000010C000C00081A08BC832A209AB0A85094284A14254A25510105130801",
INIT_0F => X"30BA901293C0F5012906A96DCD13042CE0C206E92DCD07042CE0C40D02048000",
INIT_10 => X"4CA4271CA2168ACB0E06E92DCD13042CE0C206A96DCD07042CE0C4408632C395",
INIT_11 => X"58408632C30D522CE80239CC2806AC44E954939AB299E000738F88296CA13B44",
INIT_12 => X"5145CD5306028F01990C080808494A64708B265CC4052B0F30302E060965EA00",
INIT_13 => X"51E0328A2CA9722094650CCAC0629112BA89C04A228568547B1654B9104A3286",
INIT_14 => X"A158BB80D4D8D48CB54012290470562EC29E44050B1DC60132282B68B9AA60C0",
INIT_15 => X"280000A5C11B9008FE2FA38F87804251CB0FAD40562EC0B426149D17E0044B10",
INIT_16 => X"509425094246A10A10441010090480C0964201800044109012001A000726E454",
INIT_17 => X"0942509425094250942509425094250942509425094250942509425094250942",
INIT_18 => X"9425094250942509425094250942509425094250942509425094250942509425",
INIT_19 => X"7E24502A80000000000000000005094250942509425094250942509425094250",
INIT_1A => X"AEBAEBAEBAEBAEBAFFD7F7F7F775555557DFBEEFBBFCFDF7DFFCF9F80089F7DF",
INIT_1B => X"BF5FAFD7EBF5FAFD7EBF5FAFD7EBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEB",
INIT_1C => X"FFFFFFFE0001DFAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7E",
INIT_1D => X"4500557DE00000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"E100004020BAAAFFD5400AAFBC2155AAAA97410FFFFEAAAAF7AA955EFF7803FF",
INIT_1F => X"5410F7AEBDE10FFFFFDEAAF7D568AAA5D002AB55005568B55087FC0010AAFBFF",
INIT_20 => X"555FF5D04154BAAAAEAAA10557BEAA10AAFBE8A00557BFFFEF007BC215500001",
INIT_21 => X"400000A2AABFF45550400000AAFBFFFEF550000155A28415410F7AEAABFFA2D1",
INIT_22 => X"D568AAAFFFBC21555D517FF45F7AEA8BFFA2AEAAA10A280021EF5D557FF55AA8",
INIT_23 => X"AAE974AAF7D142145082A975FF555568A00FF842ABEFA2AAA8B5500003DF55F7",
INIT_24 => X"000000145A2AA821EFFFFFD7410007FC0010555155555FF80174000055555EFA",
INIT_25 => X"2E3A0925C7E38E38F7D14557AE00000000000000000000000000000000000000",
INIT_26 => X"7D0075C7028B6F1FAE00000A02092B6F5D2438A2FBC2145B6A090428FFF5EAA9",
INIT_27 => X"FEF1C7FC516D080E15438E3A4BAE00FFF5FAE92F7D16AAAA41042FB7D145568B",
INIT_28 => X"2428FFA4AFBFFAAD1505FF490E174AABEA0ADA005D7BEDA00B6F1EFA28557BF8",
INIT_29 => X"001FF555F7FF7DAA8E07028B6A0BFF6D490E00000BEF5FAFEF490407155BE8E1",
INIT_2A => X"AAAB551C0E3AF55F7DF68ABAE3F1C0145415B78F45FFA4AFBC7BEA4AAA10A284",
INIT_2B => X"84104380055525FFBEAE90482E3D54216D0024975FF555F68A00F7842FBD7B6A",
INIT_2C => X"0000000000000000000000016DAAA0851FFE3FBD0438007FC00385D555556DEB",
INIT_2D => X"FF80020BAF7D16AA10A28402155A2AEA8BEF5D516AA000000000000000000000",
INIT_2E => X"A08003DFEF55516ABEF0055574BAFFD568A10002A82000FFD5400AAA2FBC0145",
INIT_2F => X"00F7D17FEBA557BEABEF557BD55EF082A974BAA28028A00F7D16AA10F7D56AAB",
INIT_30 => X"BEF000417545FFAA820BAFF843DFFFA2D5421FF002E954AAFF843DE105D7FFDE",
INIT_31 => X"DF55F7802AA10AA80001FF5D7FFDFEFA2AA974BAF7803FFFF002A82000FFD568",
INIT_32 => X"EAA10FF803DF45FFAEA8B555D2EAAB45F7FBE8ABAAAD540145007FE8B55FF843",
INIT_33 => X"FC20AA5D55555FFA280000BA0855401EFF7AA82010AAD1421FF0004155FF557F",
INIT_34 => X"00000000000000000000000000000000000000001EFA280175FFAAFFC00BA087",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"19FFFFFFFFE00000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(13),        -- Port A data input
DOA(0)   => data_read_a_lo_256(13),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(13),        -- Port B data input
DOB(0)   => data_read_b_lo_256(13),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_14_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10020A000180000284008280000281800000030000000033022000000580002",
INIT_01 => X"A140098018300848184860000C20C24040000000084000084200000000110200",
INIT_02 => X"88010C5A8010A600A4F558040080000041000000022C024008003CCCC9028030",
INIT_03 => X"000103A7A00904D0842242024210810803006480088000003081054288C10000",
INIT_04 => X"0000120122009000100C00000000000400A83A2044200C840000800400101820",
INIT_05 => X"040000008008010024C0C0010040000402000025000800020004207000100800",
INIT_06 => X"40870408600800800410D006A850018024240008881024A82040010461042000",
INIT_07 => X"08120054B42850B42A100010ED1500010001A040003164040CF5E20140000888",
INIT_08 => X"400500090A020220A40A7000800000000014FE8508144C924080C10000880140",
INIT_09 => X"0004010411110020000100020021004000800461600191080101000042200000",
INIT_0A => X"0000000000010190070310200008B202236D080802000002C010024000000000",
INIT_0B => X"0141001001088A45000082400000010040012100010000020000135249020820",
INIT_0C => X"0004000000000000004000000000000004000000000000000000008010100000",
INIT_0D => X"0840401000000044080200210100100017000420808200000440400000000040",
INIT_0E => X"0000000000000C00000000040302200800A04090204810244825010104130800",
INIT_0F => X"397468090008142014840100002C382800008401000038382800006402048000",
INIT_10 => X"83514072C000444C00840020002C38280000840020003838280002C09D010868",
INIT_11 => X"03C09D0104B01C57100440202900184414430534605E38048021800224804191",
INIT_12 => X"40049594C194000090450808802008830024F0E248C902AEF0024170CF180010",
INIT_13 => X"8000120020E5A08E6000048200196264BCF1C030C0604800001076C047300002",
INIT_14 => X"A00002003DEDE82C78900902A0D0000080019FAAA32D9602490302409292B832",
INIT_15 => X"2800D049100021171F6C34080240108AB292CA000000800AD1A19F6F000AA0C0",
INIT_16 => X"409024090246810810440000090480C096420080000010801001600001200454",
INIT_17 => X"0902409024090240902409024090240902409024090240902409024090240902",
INIT_18 => X"9024090240902409024090240902409024090240902409024090240902409024",
INIT_19 => X"6504002800000000000000000004090240902409024090240902409024090240",
INIT_1A => X"E79E79E79E79E79E7FDDF77777F3CF3CF7D55E6D39723FC3DEFA75D77B75F7DF",
INIT_1B => X"9FCFE7F3F9FCFE7F3F9FCFE7F3F9E79E79E79E79E79E79E79E79E79E79E79E79",
INIT_1C => X"FFFFFFFEFFFE0FE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F",
INIT_1D => X"55A28417400000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"AAAF7AA955EFF7803FF4500557DF45F7D16AB455D00001EFAAAAAAABA5555575",
INIT_1F => X"214555003FF450804001555D2AA8AAA002ABDE10082ABDF55AAAA97410FFFFEA",
INIT_20 => X"175EF5D5168A10082E80155087FC0010AAFBFFE100004020BAAAFFD5400AAFBC",
INIT_21 => X"EBDE10FFFFFDEAAF7D568AAA5D002AB55005568A00A2D5401455D00175FFFF84",
INIT_22 => X"7BC2155000015400AAD157545080402145087FD75FFF7AE82145A2D17FE10F7A",
INIT_23 => X"000000BAFFFBE8AAAA2FBFDE00087FD5410557BEAA10AAFBE8A00557BFFFEF00",
INIT_24 => X"000000155A28415410F7AEAABFFA2D1555FF5D04154BAAAAEAAA005D002AB450",
INIT_25 => X"7B6A0AAA82555157555B68012400000000000000000000000000000000000000",
INIT_26 => X"45B6A090428FFF5EAA92E3A0925C7E38E38F7D14557AF45FFDB6AB6D4100071C",
INIT_27 => X"092B6F5D2438A2FBC21455D0A3FF6D080407155552AAAA920020BFE10002EBAF",
INIT_28 => X"01454100175C7E380125D7555B6DA1014248217D0075C7028B6F1FAE00000A02",
INIT_29 => X"82145AAD178E38E3A4BAE00FFF5FAE92F7D16AAAA41042FB7D145568A38AADF4",
INIT_2A => X"1EFA28557BF8FEF1C7FC516D080E15400A2DB5754508040716D007BD05EFEBAA",
INIT_2B => X"A0ADA0055002AB6D0000020BAFFF1E8ABABEF1FAE001C7FD54005D7BEDA00B6F",
INIT_2C => X"00000000000000000000000155BE8E12428FFA4AFBFFAAD1505FF490E174AABE",
INIT_2D => X"F7FFEABFF080015555F78028A00555155555FF84000000000000000000000000",
INIT_2E => X"000003DE10082EAAB45FF80020BAF7D16AA10A28402155A2AEA8BEF5D516AB45",
INIT_2F => X"BAFFD568A10002A82000FFD5400AAA2FBC0145552ABFFFF000417555552EA8A1",
INIT_30 => X"FEF55516AABAAAFFC0145000417555A280001455D7FFDE105504021EF0055574",
INIT_31 => X"55FF007BC01FFAAAE80155AAD568ABAA28028A00F7D16AA10F7D56AABA08003D",
INIT_32 => X"D74105D7FFDE00F7D17FEBA557BEABEF557BD55EF082A97410AAFFD554508001",
INIT_33 => X"5421FF002E954AAFF843DE10550028BEF0004020BAF7D568AAAF7D168A105D7F",
INIT_34 => X"0000000000000000000000000000000000000000145FFAA820BAFF843DFFFA2D",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"01FFFFFFFFE00000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(14),        -- Port A data input
DOA(0)   => data_read_a_lo_256(14),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(14),        -- Port B data input
DOB(0)   => data_read_b_lo_256(14),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_15_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000A000000000284000280000001800020030000000033022000000180002",
INIT_01 => X"A140098018300848180060000C00424040000000080000080200000000110200",
INIT_02 => X"080108000010E60004E55800008000004100000000040240080000C009170016",
INIT_03 => X"0000000080000040842240000210810002000400888000003080014288C00000",
INIT_04 => X"0001100024A0800000440000000000040088322044200C840000011400151800",
INIT_05 => X"440002988000000020000000000B8094020000254C8800000514203000108800",
INIT_06 => X"00070000620040880410D00C285000802424000AA81024A80040010C01062001",
INIT_07 => X"086100043224489428100010811100010001A040003124040CAC600040000888",
INIT_08 => X"160500090A0282A06400100080C300000005BE0488104C800000010000880000",
INIT_09 => X"000581041110022000000002002100400080046140011008010100008A040000",
INIT_0A => X"0000000000010180060210200008B2022304080800000007C010024000000000",
INIT_0B => X"4140001001088A45000082000000010000002000010000020000034249000020",
INIT_0C => X"0004000040000400000000000000000004000020000200000000008010100000",
INIT_0D => X"094000100000004C000200250000188016000400000000000440400000000040",
INIT_0E => X"0000000108000C00000000000200200800800000000000004020000000000000",
INIT_0F => X"0000000000000000000404200000000000000404200000000000008C00048000",
INIT_10 => X"4000000000000000000405000000000000000405000000000000004000001000",
INIT_11 => X"0040000010000000000000000000004000201000000000000000000000800002",
INIT_12 => X"0004000110000000000C00080010180000000001A10240500000000000000000",
INIT_13 => X"0000000020080400000000020000008040020000000000000010001200000000",
INIT_14 => X"0000020000000611002800000000000080000011044220000000000080200200",
INIT_15 => X"8800000100000000009080E2E0A0000000000000000080000040000000000000",
INIT_16 => X"0000000000460000004400000904808094020080000010000000000000000041",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0004002800000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000004000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFE00000000000000000000000000000000000000000000000000000000",
INIT_1D => X"EF08517DE00000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"1EFAAAAAAABA555557555A284175FF000002010552A97400007BFDE10A2AA801",
INIT_1F => X"DFEF5D2AAAB45F7D17DF45087BC0155002A801FF08003DF45F7D16AB455D0000",
INIT_20 => X"C2145F7D568BEFAAD557555AAAA97410FFFFEAAAAF7AA955EFF7803FF4500557",
INIT_21 => X"03FF450804001555D2AA8AAA002ABDE10082ABDFFFF7D17FE10002E954AAF7FB",
INIT_22 => X"FFD5400AAFBC21EFA2AE95545A2D56ABFFAAD17DE10FFD1420AA007FC0145550",
INIT_23 => X"02A801550055401555D00174BA002AA8B55087FC0010AAFBFFE100004020BAAA",
INIT_24 => X"000000000A2D5401455D00175FFFF84175EF5D5168A10082E801FFFF8428A100",
INIT_25 => X"80871FAE00A2A0871EF145B7FE00000000000000000000000000000000000000",
INIT_26 => X"45FFDB6AB6D4100071C7B6A0AAA82555157555B680125C71C0E0500049209543",
INIT_27 => X"5C7E38E38F7D14557AFC75524AFB45FFD178F7D1C71C2145002E801C7140A3FF",
INIT_28 => X"AE000024954AAFFFBC2145F7DB6DBEFA2D557545B6A090428FFF5EAA92E3A092",
INIT_29 => X"470820071C71455D0A3FF6D080407155552AAAA920020BFE10002EBAFC7FFDF7",
INIT_2A => X"1FAE00000A02092B6F5D2438A2FBC21FFBEA090545B6D568BFFAADB7AE10F7D5",
INIT_2B => X"24821FFE3802FA2808208017D1C5142155410A104AA1420AFB7D0075C7028B6F",
INIT_2C => X"00000000000000000000000038AADF401454100175C7E380125D7555B6DA1014",
INIT_2D => X"552E954100004174AA00516AA10AA80155EF5D7BFDE000000000000000000000",
INIT_2E => X"5082E801555D2EBDF45F7FFEABFF080015555F78028A00555155555FF8400155",
INIT_2F => X"BAF7D16AA10A28402155A2AEA8BEF5D516AB555D043DF55F7D56ABEF55514015",
INIT_30 => X"E10082EAAB55FFFBE8A100804154AAF7FFC2145FFFFFDFEFAAD157545FF80020",
INIT_31 => X"ABEFA2FBE8A00FFD155410005555545552ABFFFF000417555552EA8A1000003D",
INIT_32 => X"3DFEF0055574BAFFD568A10002A82000FFD5400AAA2FBC01FFF78400155F7D16",
INIT_33 => X"0001455D7FFDE105504021FFAA843DEBA0000021EF555142155002E800AA5500",
INIT_34 => X"00000000000000000000000000000000000000000BAAAFFC0145000417555A28",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"1800000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(15),        -- Port A data input
DOA(0)   => data_read_a_lo_256(15),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(15),        -- Port B data input
DOB(0)   => data_read_b_lo_256(15),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_16_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"DA22C618B1000482B688B186588884862A400438255FC38381441205BA803003",
INIT_01 => X"8645A80028404C211203A952A90341080B173340412000E1005D628000820484",
INIT_02 => X"A101A9006DC1084833011850AAC55001349B10881802821808B4110007005E11",
INIT_03 => X"010108A802BB00080080006020020001A61036202800000D2410104200404550",
INIT_04 => X"8BFA58800005C40A46240252145148B38248030356415A4E62B6FC660F287240",
INIT_05 => X"1E0BD423CAC0000D610000000710296E542B6E3A825C15FB30A643695BFC2D56",
INIT_06 => X"000D0000C8008820CAE16020619156A5815006028179808C00A0D2152B90707A",
INIT_07 => X"F500240510A00205F0A407D0021A155378900002A002433A0AA00EE6E7956108",
INIT_08 => X"015995440C8327241440096A2800002828123D542910380004E0310362404076",
INIT_09 => X"10222D90409A05B2CB2CA400200209E5601044A24000000462A6001888010000",
INIT_0A => X"0000000000259200140001A15000017F0051D0F837248C005514AC40C0820500",
INIT_0B => X"01200848002912300200092BA80325A2000000000001514B5500030241C000CC",
INIT_0C => X"0001100011000110001100011000110001080008800080005202280801080395",
INIT_0D => X"17680002815014B90000205DA00880100095A64800008003561180063DB4F611",
INIT_0E => X"0280080922554515512174000000490009000000000000004010042A204A0C58",
INIT_0F => X"2DA0063EAA9C238B2D4C800632B266E828EE4C800632AAAB6830D0FC6B06C041",
INIT_10 => X"0839AA149339E8FB964C800632B266E82B2E4C800632AAAB683310872800EDA5",
INIT_11 => X"C087A800EB090D4AAC91268FFCBE81397826C4A20D2B6C510E8624792A4A30A4",
INIT_12 => X"3638E8849D5C532408DD6E004C90C06AC019D88B9795012CA96902C799912BC3",
INIT_13 => X"78706531C74485BD42A30906057FADAA456218FD8E3ED83B60E3A242DC0F1898",
INIT_14 => X"51727A06FB555793057C444CF45C5C9E89543B8BC6E80193DC36F6C71D1093A4",
INIT_15 => X"10DCD45DC02B331650CA8ACB4007E00D1C6A6A58395C917F7E74D936F650D69B",
INIT_16 => X"000000000012000081500008A422150884081ACAAC0542054004FC5884640508",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"3604000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"45145145145145147A7797E1E1A79E79E15634455131A436993071A616D4F68A",
INIT_1B => X"3E9F4FA7D1E9F47A7D1E9F47A7D3453453453453453453453453453453453453",
INIT_1C => X"FFFFFFFE00001F4FA7D3E9F4FA3D1E8F47A3D1E8F47A3D1E9F4FA7D3E9F4FA7D",
INIT_1D => X"00FF8015400000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"400007BFDE10A2AA801EF08517DE10FFFFFDFEFA2D16AB55A2FFFFEAA5D7FC00",
INIT_1F => X"74BA5D2EBDFEFAAD17FFFF002EBDE000800174AA55043FFFF000002010552A97",
INIT_20 => X"E8AAAAA80000105D557FF45F7D16AB455D00001EFAAAAAAABA555557555A2841",
INIT_21 => X"AAAB45F7D17DF45087BC0155002A801FF08003DE000004154BA002A800BA087F",
INIT_22 => X"803FF4500557DEAAF7D57DEBA082A82010FFAE975555D7FFDEAAFF80155EF5D2",
INIT_23 => X"2D57FFFF557FD55FF08003FE0055043FF55AAAA97410FFFFEAAAAF7AA955EFF7",
INIT_24 => X"0000001FFF7D17FE10002E954AAF7FBC2145F7D568BEFAAD557410552EA8BEFA",
INIT_25 => X"DB6FFFDEAA5571C7010FF8412400000000000000000000000000000000000000",
INIT_26 => X"C71C0E050004920954380871FAE00A2A0871EF145B7FE10E3F1F8FC7AAD56DB7",
INIT_27 => X"A82555157555B680124924124BDFEFA2D57FFC71C2EBDE280000174825D0E3FF",
INIT_28 => X"74821424800AA007FEDAAAA284020385D5F7AF45FFDB6AB6D4100071C7B6A0AA",
INIT_29 => X"F8EAAFF80175C75524AFB45FFD178F7D1C71C2145002E801C7140A3FE10080A1",
INIT_2A => X"5EAA92E3A0925C7E38E38F7D14557AE92EBDB78EAA1C2482010FFAE9556D557F",
INIT_2B => X"D557410492EADBEFA2D178FEF5575D55EF000A38E10490A3AF45B6A090428FFF",
INIT_2C => X"000000000000000000000001C7FFDF7AE000024954AAFFFBC2145F7DB6DBEFA2",
INIT_2D => X"A2D56AB45A2D57DFFFF7FBFFEAA555555400F780000000000000000000000000",
INIT_2E => X"A080415400552ABDF55552E954100004174AA00516AA10AA80155EF5D7BFDE10",
INIT_2F => X"FF080015555F78028A00555155555FF840000000043DFEFAAD17FF45552ABFEB",
INIT_30 => X"1555D2EBDE10002E974005D04020BA007BFDEBAA284000BA557FE8B45F7FFEAB",
INIT_31 => X"0000F7AE955EF5D7BE8ABAF784175555D043DF55F7D56ABEF555140155082E80",
INIT_32 => X"AAB45FF80020BAF7D16AA10A28402155A2AEA8BEF5D516AA00AAFBE8AAA55040",
INIT_33 => X"FC2145FFFFFDFEFAAD157410082ABFFEFAAD16ABFF5555575FF082AA8A00002A",
INIT_34 => X"0000000000000000000000000000000000000000155FFFBE8A100804154AAF7F",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0800000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(16),        -- Port A data input
DOA(0)   => data_read_a_lo_256(16),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(16),        -- Port B data input
DOB(0)   => data_read_b_lo_256(16),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_17_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"5284CE4FB7BD2C8994A13392DBD02E14006B82AC7E800D44D3DD2FD5F9B961C0",
INIT_01 => X"F8ACD01F7E03FC6793F2199B39FC233C11D93AE6F3BB92B32091DBC339B24542",
INIT_02 => X"8F333007FD6808092A2AFA6667033DB50853379C10BFF70F1BD011110F205F18",
INIT_03 => X"294ADB4AFFCBF0DAD63ABF836B58EAFE060478202022234B2E0303FDC9E18339",
INIT_04 => X"DB7A40806FE4040840EBC563A0150A0926146FECB04196482236FC2005282AE1",
INIT_05 => X"0807B4070670083DC68206D7E6D0250834336D1E81500FDB306045255BFC2076",
INIT_06 => X"00000000141C5AF3EA6AB187F7F8CE039786062C6CE092F5FE005236781C402A",
INIT_07 => X"1684248A38B022475DCA9BD00116E33CC3821774BB55F53BB42329AA3C0CEF60",
INIT_08 => X"60700CE0641527241060AD844E1C0088001223022D189A2800542219204903F8",
INIT_09 => X"D94C1C1C51DFF881861CBE0305A12A0321810217C01D34EDC98FFA1C8E000016",
INIT_0A => X"7E7D8F8FBDE40E001E000B3A5DAADAFDDA5DA79350DF70027CE86F047BEF19B6",
INIT_0B => X"814102F800633F1D0A7CC9AE74117FE0003A6AD055819D1F9984014B37BA5FFC",
INIT_0C => X"CF4FBCF4FBCF4FBCF4FBCF4FBCF4FBCF4FBE7A7DE7A7800617112E46F05D02DD",
INIT_0D => X"D7FE4A5A99FD6D3FEF4BEB5FF994F0FEFFCCF8430006CE8A3F06ABD73DBCF4FB",
INIT_0E => X"B29760593F33FA0CF170F40006001B1A05C0000000000000008004BA78428C7A",
INIT_0F => X"EDA57E46444357B3950A9BFBAC94CFA8581E0A9BFBAC8CCFA8580C7CAF51EF68",
INIT_10 => X"7DF76B5DB54A09003E0A9BFBAC94CFA8581E0A9BFBAC8CCFA8580E46FBFCB0CB",
INIT_11 => X"E7467BFCB1D5CFEB56A1A100D5345C1BFFE8FBDB892DB463034198E2881F3F78",
INIT_12 => X"4E0ADD39387F92B2935DFEAADDF38EBCFB9E3D636DCDF9B90F966BF92966D5D9",
INIT_13 => X"F256527055EB6D555CB294981B7FB5B2954CD3013013FDF5E82AF5B6AAAE594A",
INIT_14 => X"F7D7E835C67E655BAA868610117575EA1C34BD6975D48B44A0405FC15BA7270F",
INIT_15 => X"BD07F6CD2A47D0CBA96252756D7217E5E1C61DBDF5FA167F7AE5D3D21A414007",
INIT_16 => X"00000000005F08000179C16DECF67F08BC02F9067ED55805600545DFE45A80E7",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"F981800C00000000000000000000000000000000000000000000000000000000",
INIT_1A => X"A69A69A69A69A69A919261A1A6075D75D10DC800C027B731014BA4B864617114",
INIT_1B => X"8341A0D068351A8D068351A8D069A6BAE9A69A6BAE9A6BAE9A69A6BAE9A6BAE9",
INIT_1C => X"FFFFFFFE000011A8D46A351A8D46A351A8D46A351A8D46A341A0D068341A0D06",
INIT_1D => X"55AAFFD5400000000000000000000000000000000000000000000001FFFFFFFF",
INIT_1E => X"B55A2FFFFEAA5D7FC0000FF8015410FFFFFFFFFFFFFFDFEFF7D568A1008003DF",
INIT_1F => X"DF55A2D1400000804154BAF7D168A00A2803DE10FFAE95410FFFFFDFEFA2D16A",
INIT_20 => X"2AABAFFD56ABFF002EBDFFF000002010552A97400007BFDE10A2AA801EF08517",
INIT_21 => X"EBDFEFAAD17FFFF002EBDE000800174AA55043FEBA0004174AA5504000AA5504",
INIT_22 => X"5557555A284175FFFFFBE8B55A2FFFFF55F7803DEBA002AAAAAAF7FBD74BA5D2",
INIT_23 => X"D0417400FFD57DE00AAAAAAB45A2AA97545F7D16AB455D00001EFAAAAAAABA55",
INIT_24 => X"0000000000004154BA002A800BA087FE8AAAAA80000105D557FE00A2D5420AA5",
INIT_25 => X"7EBD16AA00000E3DF6DBEF5D2400000000000000000000000000000000000000",
INIT_26 => X"10E3F1F8FC7AAD56DB7DB6FFFDEAA5571C7010FF8412428FFFFFFFFFF7FBF8FD",
INIT_27 => X"E00A2A0871EF145B7FF7DA2D547038140E10492FFDF6DA28A28E3DE00F7A0924",
INIT_28 => X"2492550A020BA55002AA82F7DF6DBD71C2EBFFC71C0E050004920954380871FA",
INIT_29 => X"ADABAF7F5D74924124BDFEFA2D57FFC71C2EBDE280000174825D0E3FEAA14001",
INIT_2A => X"0071C7B6A0AAA82555157555B680125FFEBFFEDB55BEFFFAF6DE38E3DEAA002E",
INIT_2B => X"5F7AE28B6D545092490E10400FFDB7AE00A2AAADB45BEA092545FFDB6AB6D410",
INIT_2C => X"00000000000000000000000010080A174821424800AA007FEDAAAA284020385D",
INIT_2D => X"FFFBFDFEFF7FFEAB45A2D56AA00002EBDFFFF7D5400000000000000000000000",
INIT_2E => X"AA2AABDE10FF8400010A2D56AB45A2D57DFFFF7FBFFEAA555555400F780000AA",
INIT_2F => X"100004174AA00516AA10AA80155EF5D7BFDFEFAAD1554BA552E82000F7FFFFEA",
INIT_30 => X"400552ABDEBA5D0002000552A800BA55042AA10FFFFFDF55552EBDF55552E954",
INIT_31 => X"ABFFA2AEBFEAA082EBDEBAFFD55540000043DFEFAAD17FF45552ABFEBA080415",
INIT_32 => X"00145F7FFEABFF080015555F78028A00555155555FF84001FFAAFBFFF55FFFBE",
INIT_33 => X"BFDEBAA284000BA557FE8AAAFFD155400082A82000F7FFE8A00A2AABDF45F780",
INIT_34 => X"0000000000000000000000000000000000000000010002E974005D04020BA007",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"19FFFFFFFFE00000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(17),        -- Port A data input
DOA(0)   => data_read_a_lo_256(17),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(17),        -- Port B data input
DOB(0)   => data_read_b_lo_256(17),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_18_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"69844019080000A21A611406840014122A641074155FC28A2024001001801003",
INIT_01 => X"A643D920034004180005E9E3C90360C0041C0181002001602025800008440084",
INIT_02 => X"B7333980808408103F2000F81FC0FEDEAC2161B0B84D0002188011110C018041",
INIT_03 => X"0405D434003F2C020081587008020561E55116B0290000042B71240C800440F8",
INIT_04 => X"50805AC31007D6125724029216554A9847669903D640EC8E2001002604503004",
INIT_05 => X"0E010001C1CA11803850C800010022660C1C0065003C0404002646DC20A02D40",
INIT_06 => X"50AD050AC00000002A4F612449903FE080000000005889AC41E04508A9907020",
INIT_07 => X"5584280B10014003A8067400920810FF3C72024300A0030048221ACEE383E518",
INIT_08 => X"00C983E6041505253500F66E620428000B1804000152E52801A2020084090040",
INIT_09 => X"20500B90419005B0C309402030060860E01004A828408800440405E350294010",
INIT_0A => X"008010100007865421432121804021C20452880C2D200000045C18C0E0000A08",
INIT_0B => X"09700C04C44C92A88DC42215C882E82250811000000C1AE061861710A401A4E8",
INIT_0C => X"308003080030800308003080030800308001840018400400602A018809800371",
INIT_0D => X"0801010202021000780004200408C1002003F66CA1B13111C0D95C20C2030A00",
INIT_0E => X"02900806400FC503F08180050942E4200020C1B060D8306C182701404C197301",
INIT_0F => X"22AABABAF377DF1CA160820520EB3057E70E60820520F33057E72E9154159000",
INIT_10 => X"8A2AD5D48F37FAFEFE60820520EB3057E7CE60820520F33057E7EC658BF2DA78",
INIT_11 => X"32658BF2D4B2A80BF8FE39FD78EB0D882014A62C568FFAFC73FFDD9C2B30E046",
INIT_12 => X"C728C800DFC06F59F710107533C0C4E37619440FBFBAB2400AFC1600361D798F",
INIT_13 => X"0DEBBEB9454005BAA36DEFF894823A3D1A88A2FE29D5FC6DCAA2A002DD51B6E7",
INIT_14 => X"F3B7092A78606A28A5427AAB9FF4EDD251C7123E291660733EBF6FE519001BF4",
INIT_15 => X"82202AB58AFBFD5DE200A8EBE3A3EC110339E1DCEDC2590495BB2112E2BE4BF5",
INIT_16 => X"C1B06C1B06808348340000020301805002D008C1F92000A5F421B8000DB49103",
INIT_17 => X"1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06",
INIT_18 => X"B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C",
INIT_19 => X"16000000000000000000000000041B06C1B06C1B06C1B06C1B06C1B06C1B06C1",
INIT_1A => X"A28A28A28A28A28A244C16454170410412CA2EFB3AE03B85CF08C03F1A30F7DF",
INIT_1B => X"8944A25128954AA552A944A2512AAA8A28A28A2AAAAAA8A28A28A2AAAAAA8A28",
INIT_1C => X"FFFFFFFE000004A25128944A25128944A25128944A25128944A25128944A2512",
INIT_1D => X"105D2A80000000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"FEFF7D568A1008003DF55AAFFD5410FFFFFFFFFFFFFFFFFFFFFBFDEBA552E974",
INIT_1F => X"5410FFFFFFFFFF7FBE8B55AAD16AA1000516AA005D0400010FFFFFFFFFFFFFFD",
INIT_20 => X"FFE00087BC2155087BC0010FFFFFDFEFA2D16AB55A2FFFFEAA5D7FC0000FF801",
INIT_21 => X"1400000804154BAF7D168A00A2803DE10FFAE95555FFFBE8B45A2D56ABEFFFFF",
INIT_22 => X"AA801EF08517DF55000000010082A974AA08557DEBAFFAEBFF55AA8028B55A2D",
INIT_23 => X"52E800105D2AAAA10A2D1420AAFFAEA8BFF000002010552A97400007BFDE10A2",
INIT_24 => X"0000000BA0004174AA5504000AA55042AABAFFD56ABFF002EBDEBA0004020BA5",
INIT_25 => X"FF7FBFFEBA552A95410552485000000000000000000000000000000000000000",
INIT_26 => X"28FFFFFFFFFF7FBF8FD7EBD16AA00000E3DF6DBEF5D2438FFFFFFFFFFFFFFFFE",
INIT_27 => X"EAA5571C7010FF8412410FFFBF8FC7E3F5EAB45BEDB6FA3800556FA005504050",
INIT_28 => X"AB55BEDB6FBC7EBF5F8E10007BC516D1C71C5010E3F1F8FC7AAD56DB7DB6FFFD",
INIT_29 => X"BFF55BE8A2DB7DA2D547038140E10492FFDF6DA28A28E3DE00F7A09256DE3F1E",
INIT_2A => X"0954380871FAE00A2A0871EF145B7FF45080E070280820924AA145578E92F7A4",
INIT_2B => X"2EBFEBA1C0A00092412E850005D2AAFA38A2DF45082F7AAA8BC71C0E05000492",
INIT_2C => X"000000000000000000000000AA140012492550A020BA55002AA82F7DF6DBD71C",
INIT_2D => X"FFFFFFFFFFFFBFDFEFF7FFFDEAA5D2E954105504154000000000000000000000",
INIT_2E => X"A08557DE005500154AAFFFBFDFEFF7FFEAB45A2D56AA00002EBDFFFF7D5400AA",
INIT_2F => X"45A2D57DFFFF7FBFFEAA555555400F78000010F7FBE8B55AAD16AB55F7FBFDEA",
INIT_30 => X"E10FF84001FFAAD568B45FFFBFFF55A2D568A00087BD55FF5D5555410A2D56AB",
INIT_31 => X"00AA555168A10FF803DF45FFAABDFEFAAD1554BA552E82000F7FFFFEAAA2AABD",
INIT_32 => X"A8B55552E954100004174AA00516AA10AA80155EF5D7BFDF45002A974AA08000",
INIT_33 => X"42AA10FFFFFDF55552EBDEBA5D2E80010082A97410552EBDEBAA2FBD5400F7AA",
INIT_34 => X"00000000000000000000000000000000000000000BA5D0002000552A800BA550",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0800000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(18),        -- Port A data input
DOA(0)   => data_read_a_lo_256(18),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(18),        -- Port B data input
DOB(0)   => data_read_b_lo_256(18),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_19_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"042200000000000041088001001AA00000000000000000000000500802000003",
INIT_01 => X"200048000024000000000404000000000A22000800000800004A200000000001",
INIT_02 => X"032210008DEF00400060000001C008002489E0F0004037B00010101010000000",
INIT_03 => X"0000008128000000000000000000000024001620280000000000354200004008",
INIT_04 => X"000058800004C4024024001210001054B1C822009640000E2000002604003000",
INIT_05 => X"0E010001C0400000000000000000200604000000001C04000026400000002C40",
INIT_06 => X"000000000000000001800166A84004A080000000005884020020400009907020",
INIT_07 => X"E200201C00A14080082B26208008A00900120101402240440280040840802000",
INIT_08 => X"004180261C81210031000004340000200008105428020568040213003499C006",
INIT_09 => X"00000990000000B0C30800000000086020016000000000003838000000000000",
INIT_0A => X"000000000005860000000080A000206020408000000000000454080000000000",
INIT_0B => X"00000000000040002000044000000000000000000005E0003E00004049640004",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"00000000210001D8000000000000000020009640000000000000000000000000",
INIT_0E => X"040000000000C500300080000000000000000000000000000000000000000000",
INIT_0F => X"50500101088A37034E156600D740022800EC156600D740022800D01E0412D069",
INIT_10 => X"E61700224081044914156600D7400228002C156600D7400228001098F00D0FB7",
INIT_11 => X"CC98F00D0F2DD014010046037814EA63DBB31CE7605001008C41A061F0E7D693",
INIT_12 => X"361526D600000004089E12350C0E01FF23315422BABB46FEF5019146C0800380",
INIT_13 => X"00000130AA3592000000000629C03F3E60330C00C628908214551AC900000010",
INIT_14 => X"4208D65C006070845039014460088235ACC3123E2A29148841008482A4DAC000",
INIT_15 => X"6CD4953A66BE7A5040018D8A8AD9090A1EC20A188235AC509FB50C2D0500B409",
INIT_16 => X"00000000000000000000000000000000000008C0180027000006110008404608",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"9200000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"61861861861861861A2882313054D34D301C822EE8FC31C043198028002C7441",
INIT_1B => X"84C261349A4C26130984C261309861861861A69861861861861A698618618618",
INIT_1C => X"FFFFFFFE0000026130984C26130984C26130984C26130984C26130984C261309",
INIT_1D => X"00082E97400000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"FFFFFFBFDEBA552E974105D2A801EFFFFFFFFFFFFFFFFFFFFFFFFFEAA552E954",
INIT_1F => X"55EFFFFFFFFFFFFFFFFFEFF7FBFFEAA5D2E97545FFFFC2010FFFFFFFFFFFFFFF",
INIT_20 => X"6AA0008003DF555D5157410FFFFFFFFFFFFFFDFEFF7D568A1008003DF55AAFFD",
INIT_21 => X"FFFFFFF7FBE8B55AAD16AA1000516AA005D04001EFFFFFFFFFFFFFBFDF45AAD1",
INIT_22 => X"7FC0000FF80155EFFFFFFFFEFF7D16AB55A2D57DEBA557FEAA10080402010FFF",
INIT_23 => X"2D56AB45FFFBFDEBA5D7FC0155FFFFD7410FFFFFDFEFA2D16AB55A2FFFFEAA5D",
INIT_24 => X"000000155FFFBE8B45A2D56ABEFFFFFFFE00087BC2155087BC00AAFFFBFDF45A",
INIT_25 => X"FFFFFFDEAA552E95400002095400000000000000000000000000000000000000",
INIT_26 => X"38FFFFFFFFFFFFFFFFEFF7FBFFEBA552A954105524851C7FFFFFFFFFFFFFFFFF",
INIT_27 => X"A00000E3DF6DBEF5D25D7FFFFFFFFFFFFBFDFEFEBF5F8E92552E9556DEBF1C20",
INIT_28 => X"DFEFE3F1FAF55A2D568A0000003FF7D495155428FFFFFFFFFF7FBF8FD7EBD16A",
INIT_29 => X"EFA00000002010FFFBF8FC7E3F5EAB45BEDB6FA3800556FA005504051FFFFFFF",
INIT_2A => X"56DB7DB6FFFDEAA5571C7010FF84125EFF7F1F8FC7EBD568B6DBEDF7DEBA5571",
INIT_2B => X"71C5092E3F1F8F55AADB6DB7DEBF1FAE82557FC516DEBF1D0410E3F1F8FC7AAD",
INIT_2C => X"0000000000000000000000016DE3F1EAB55BEDB6FBC7EBF5F8E10007BC516D1C",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFBFDEAA5D2A954000800154000000000000000000000",
INIT_2E => X"0552A955EFAAD1400AAFFFFFFFFFFFFBFDFEFF7FFFDEAA5D2E95410550415545",
INIT_2F => X"EFF7FFEAB45A2D56AA00002EBDFFFF7D540145FFFFFFFEFF7FBFFFFFAAD16AA0",
INIT_30 => X"E005500155EFF7FBFDFEFAAD568B55AAD568A0008003DFFF0855554AAFFFBFDF",
INIT_31 => X"ABEFFFFFFFEAA55517DE10080400010F7FBE8B55AAD16AB55F7FBFDEAA08557D",
INIT_32 => X"40010A2D56AB45A2D57DFFFF7FBFFEAA555555400F780001FFF7D16AB55A2D16",
INIT_33 => X"568A00087BD55FF5D5555410AAD56AB45AAFFFFFEFAAD168A00557BD55FFA2D5",
INIT_34 => X"00000000000000000000000000000000000000001FFAAD568B45FFFBFFF55A2D",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"1000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(19),        -- Port A data input
DOA(0)   => data_read_a_lo_256(19),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(19),        -- Port B data input
DOB(0)   => data_read_b_lo_256(19),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_20_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000003",
INIT_01 => X"A75FF80000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"14088080800008400F655001FFCFF80018FA8044000000000000011000000007",
INIT_03 => X"0000000000000000000000000000000024001660380000000000000000004FF8",
INIT_04 => X"000079800014CC02C034001600000000000000101EC0012EE0C0026E1E80F000",
INIT_05 => X"3E1FE867DFC044003902100002203F2EFC040388137C3E20C8EEC00284033CC0",
INIT_06 => X"001F0001E0020002E80020000005FEAF91D10802ABFB80000021C8010FB0F0F4",
INIT_07 => X"00040007700000000000000001080FF900160000000200C00080001840BFE538",
INIT_08 => X"09FFBFE5181606000410A4000004202AA8043E0000000000000001209244C040",
INIT_09 => X"01227FB0000000F7DF78020004011FEFE0000000002003150200008388020000",
INIT_0A => X"000000000015BE0000004000000100000100506002008C2007D5FC8000002400",
INIT_0B => X"0000000000000000000000000000000400400520000000000000000400000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000020002",
INIT_0D => X"00010000000200000020000004000100203FF6C0000000000000000000000000",
INIT_0E => X"0000000600FFC53FF001800000002004080000000000000040900005C8485380",
INIT_0F => X"8000000009A9C300020080000800000003CC0080000800000003CC0200078000",
INIT_10 => X"00800000000012963C0080000800000003CC0080000800000003CC1008000000",
INIT_11 => X"00100800004000000000066C5000020020000000800000000C2E180010002000",
INIT_12 => X"96004000000000052B0200000014200040C2829000400000000000860F987980",
INIT_13 => X"0000A4B00400000000002958000240400000000007E1B0000402000000000014",
INIT_14 => X"400004004181800000000005C5A00000200C40808000000000AF0D8008000000",
INIT_15 => X"000800020141812737DC3020100400001C19C1D80000200400000000000015D1",
INIT_16 => X"0000004010080800801810100000000000093EDFF80200000000000010010010",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"4D20400200000000000000000000000000000000000000000000000000000000",
INIT_1A => X"CB0C30C30C30C30C8192608486879E79E681C000C00E08000402241560412010",
INIT_1B => X"2190C86432190C86432190C86432CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2",
INIT_1C => X"FFFFFFFE000010C86432190C86432190C86432190C86432190C86432190C8643",
INIT_1D => X"10080402000000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"FFFFFFFFFEAA552E95400082E975FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2A954",
INIT_1F => X"0000FFFFFFFFFFFFFFFFFFFFFFFDEAA5D2A954000800001EFFFFFFFFFFFFFFFF",
INIT_20 => X"FFEBA5D2A97400FF8017410FFFFFFFFFFFFFFFFFFFFFBFDEBA552E974105D2A8",
INIT_21 => X"FFFFFFFFFFFFFEFF7FBFFEAA5D2E97545FFFFC21FFFFFFFFFFFFFFFFFFFFF7FB",
INIT_22 => X"003DF55AAFFD5400FFFFFFFFFFFFFFDFEFF7FFEAA10000417555AAD5555EFFFF",
INIT_23 => X"FFBFDFEFAAD568A0000043DF45AAFBC2010FFFFFFFFFFFFFFDFEFF7D568A1008",
INIT_24 => X"0000001EFFFFFFFFFFFFFBFDF45AAD16AA0008003DF555D51574BAFFFFFFFFFF",
INIT_25 => X"FFFFFFFEBA5D2A95410000A00000000000000000000000000000000000000000",
INIT_26 => X"C7FFFFFFFFFFFFFFFFFFFFFFFDEAA552E954000020955FFFFFFFFFFFFFFFFFFF",
INIT_27 => X"EBA552A95410552485010FFFFFFFFFFFFFFFFFFF7FBFDEBA5D2E95400140E001",
INIT_28 => X"FFFFFFFFFDFEFF7FFFFEAA5D2E95400E38A17438FFFFFFFFFFFFFFFFEFF7FBFF",
INIT_29 => X"1557DBEDF575D7FFFFFFFFFFFFBFDFEFEBF5F8E92552E9556DEBF1C21C7FFFFF",
INIT_2A => X"BF8FD7EBD16AA00000E3DF6DBEF5D2438FFFFFFFFFF7FBFDFC7EBF1E8A00080A",
INIT_2B => X"5155492FFFFFFFEFF7F1F8FD7A2D168A1008043FF6DAAFBC5028FFFFFFFFFF7F",
INIT_2C => X"000000000000000000000001FFFFFFFDFEFE3F1FAF55A2D568A0000003FF7D49",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFEBA552A95410002E820000000000000000000000",
INIT_2E => X"A552E954005D2A82145FFFFFFFFFFFFFFFFFFFFFBFDEAA5D2A954000800155FF",
INIT_2F => X"FFFFFBFDFEFF7FFFDEAA5D2E95410550415410FFFFFFFFFFFFFFDFEFF7FBFFEB",
INIT_30 => X"5EFAAD140155FFFFFFFFFF7FBFDFFFFFFBFDEBA5D2A95400A2AA974AAFFFFFFF",
INIT_31 => X"FF55A2D568A10082E955FFFFFFD7545FFFFFFFEFF7FBFFFFFAAD16AA00552A95",
INIT_32 => X"D74AAFFFBFDFEFF7FFEAB45A2D56AA00002EBDFFFF7D5400BAFFFFFDFEFF7FBF",
INIT_33 => X"568A0008003DFFF085555410F7FBFDFEFFFD568B45AAD16AA1008003DFEFAAFB",
INIT_34 => X"00000000000000000000000000000000000000001EFF7FBFDFEFAAD568B55AAD",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"01FFFFFFFFE00000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(20),        -- Port A data input
DOA(0)   => data_read_a_lo_256(20),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(20),        -- Port B data input
DOB(0)   => data_read_b_lo_256(20),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_21_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"4A302428B824900A128C090A5C1800261500213C005FE812D10420054085A202",
INIT_01 => X"081FFE3440B609703B0427F801A40B8115BC4F655300340288A40D30040E4DD8",
INIT_02 => X"0109095C30C98809800000F9FFFFFFFF149FF1FCA4C0421B182E3490DF145FE4",
INIT_03 => X"084A76341244919000099486400026523C041660BA000100CC12701015007FF8",
INIT_04 => X"000079800014CC03C075161E001118653D2408041FC004AEF000816E1C11F541",
INIT_05 => X"7E1F00F7FFC000240100004683103E7FFE02482553FC3C0204EFC25010143CC0",
INIT_06 => X"801008011010421960E339A20205FEBF8140000203FFC806C8A1C1048FF0F0E0",
INIT_07 => X"750504800680102542AD800504530FF9061E8026998E9A00402CC25BD0FFF800",
INIT_08 => X"11FBFFE04691A5A00101818A6800088228000001A044C8168480D010F200AA08",
INIT_09 => X"E85A7FF080AC70FFDF78220010841EFFE7116E144071268DFD3E4C2404010000",
INIT_0A => X"54518A8A31B7FE00040009814C089202225412115428C03BC7D7FC15025B1AB6",
INIT_0B => X"88300E20806520398C682157A493896600E24E10100DFF22FF86002020ED110C",
INIT_0C => X"28D9228D9228D9228D9228D9228D9228D99146C9146C84006309044081A001B1",
INIT_0D => X"890000403000A01282088624001201A8C43FF7C0011529904595123203040D92",
INIT_0E => X"06102C4053FFD5BFF00A04A00200602CA5200110008800444021048034004001",
INIT_0F => X"2A00263009140094D81A5040605800B506901A30406054013605620272181965",
INIT_10 => X"890A202811209062801A3040605800B506901A50406054013605604350B81282",
INIT_11 => X"3F4350B811068C00049A0A5820A3C1725A8006C0A40404D058320496C2C9C600",
INIT_12 => X"98361AC808127C454402483153A3A895BB3C1E2E820704020381702C1AAA2C4B",
INIT_13 => X"4D910CC1B154510413CC2A200501B400A40018A00C80400040D8AA288209AA21",
INIT_14 => X"0048A0141AA00418080460678A4012288463B2050302019200B00206C3590102",
INIT_15 => X"233142440470C8A9310280C0180302A01427D060022011606E800E00169C19A0",
INIT_16 => X"4010040100448008004000000E07008010003EFFFE0373056024B01118011988",
INIT_17 => X"0100401004010040100401004010040100401004010040100401004010040100",
INIT_18 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_19 => X"7E00000000000000000000000004010040100401004010040100401004010040",
INIT_1A => X"EFBEFBEFBEFBEFBEFFFFF7F7FFF3CF3CFFFFBE7FBBFDFFF7DFFCFBF08103DFDF",
INIT_1B => X"FFFFFFF7FBFDFEFF7FBFDFEFF7FBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFB",
INIT_1C => X"FFFFFFFE00003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"00080002000000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"FFFFFFFFFEBA5D2A954100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_1F => X"75FFFFFFFFFFFFFFFFFFFFFFFFFFEBA552A97400082A975FFFFFFFFFFFFFFFFF",
INIT_20 => X"FDEAA5D2E974100800155EFFFFFFFFFFFFFFFFFFFFFFFFFEAA552E95400082E9",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFDEAA5D2A95400080000000FFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"2E974105D2A80000FFFFFFFFFFFFFFFFFFFFFBFDEBA5D2E974005D2E80000FFF",
INIT_23 => X"FFFFFFFFF7FBFDEBA552A954005D2E97410FFFFFFFFFFFFFFFFFFFFFBFDEBA55",
INIT_24 => X"0000001FFFFFFFFFFFFFFFFFFFFF7FBFFEBA5D2A97400FF80174BAFFFFFFFFFF",
INIT_25 => X"FFFFFFFEBA5D2E97400000400000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2A95410000A001FFFFFFFFFFFFFFFFFFF",
INIT_27 => X"EAA552E954000020955EFFFFFFFFFFFFFFFFFFFFFFFFFEAA552E97400002E955",
INIT_28 => X"FFFFFFFFFFFFFFFFBFDEAA5D2A974101400155C7FFFFFFFFFFFFFFFFFFFFFFFD",
INIT_29 => X"97400552A80010FFFFFFFFFFFFFFFFFFF7FBFDEBA5D2E95400140E00000FFFFF",
INIT_2A => X"FFFFEFF7FBFFEBA552A95410552485038FFFFFFFFFFFFFFFFFFF7FBFDEBA552E",
INIT_2B => X"8A174AAFFFFFFFFFFFFFFFFEFF7FBFFEAA5D2E97400412497438FFFFFFFFFFFF",
INIT_2C => X"000000000000000000000001C7FFFFFFFFFFFFFFDFEFF7FFFFEAA5D2E95400E3",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974000004000000000000000000000000",
INIT_2E => X"A552E97400002E975FFFFFFFFFFFFFFFFFFFFFFFFFFEBA552A95410002E821FF",
INIT_2F => X"FFFFFFFFFFFFFFBFDEAA5D2A954000800155EFFFFFFFFFFFFFFFFFFFFFFFFDEA",
INIT_30 => X"4005D2A82010FFFFFFFFFFFFFFFFEFF7FBFDEBA552A974105D0015545FFFFFFF",
INIT_31 => X"DFEFF7FFFFEAA5D2A974005D2E82010FFFFFFFFFFFFFFDFEFF7FBFFEBA552E95",
INIT_32 => X"154AAFFFFFFFFFFFFBFDFEFF7FFFDEAA5D2E954105504154AAFFFFFFFFFFFFFF",
INIT_33 => X"BFDEBA5D2A95400A2AA974BAFFFFFFFFFF7FBFDFEFFFFFFDEBA552E974000004",
INIT_34 => X"0000000000000000000000000000000000000000155FFFFFFFFFF7FBFDFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(21),        -- Port A data input
DOA(0)   => data_read_a_lo_256(21),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(21),        -- Port B data input
DOB(0)   => data_read_b_lo_256(21),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_22_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"5290F4CDE914905A14A43D33F488243E17122300F55FEB189B343A1140548380",
INIT_01 => X"A94007B259F6A975386262000C344BA9573C6FF57B18A5FB0ABFCD3C2C5F4F0C",
INIT_02 => X"877FE30EB378008D202551040030071869D0040180AC4B685F6E26FAA0810006",
INIT_03 => X"431965109E4481D6B5AAD6875AD6AB5A1815600802888808DEA83552954D3000",
INIT_04 => X"492C0020220001010E4916C884DCD607E5EC2A344103E48003D0800023D0072C",
INIT_05 => X"0020F8882001102D620A06D683018001023D37E5088043620101179092540112",
INIT_06 => X"0803008022385AAA447A3306AA50001035B41C0A88046CAEE8C23C08E040011C",
INIT_07 => X"1EC04ED017AB5497EB923F08182E20020689B735011FBFE7BC06260294401CA8",
INIT_08 => X"4A00401D4425ADA9035BE19C8F9442A8801200F4C9D7AC8093A051727B2AC349",
INIT_09 => X"50020040E48D50080002B00A0C00801014541E9504703680017F6CB405070015",
INIT_0A => X"54538A8A738041C23020131A80CFDFF3FE509A907C6AC050402204090090319A",
INIT_0B => X"40050220103D2A512C6A8C4F0011550008E06E000140009A000000424DE61920",
INIT_0C => X"A81C2A81C2A81C2A81C2A81C2A81C2A81C9540E1540E001400006100003202D0",
INIT_0D => X"8B2940D0E153941A8B1A262CA542A9A8D6C0010A101628013456520CA09281C2",
INIT_0E => X"80410089180008800143D83888281A2034A85014280A14050A01509E05085449",
INIT_0F => X"000C26706B3C189CD84ACD20B03001E387D04AC560B02401E387E1028AC04500",
INIT_10 => X"458870201570B036C04AC560B03001E387D04ACD20B02401E387E24708E7E242",
INIT_11 => X"044708E7E1C20A0106EA167C84EBF052A8E010C0180606E86C3F459DC08DA902",
INIT_12 => X"98225189980254CDEC22A98032A22C50EAC462030A01800407C2700C2ACA2C0F",
INIT_13 => X"4A99BCC1154C258012D86F601A2E49003400138C0DA2443A208AA612C0096C37",
INIT_14 => X"90E16025483C1E0C0006B085CEC03858958D15310201015504B512044A313300",
INIT_15 => X"6B0469512C6FC01A1421006028038720640310643858162712020B001AA415F2",
INIT_16 => X"11044110445E22022365034A8EA754008004C0200323001182122548881649D1",
INIT_17 => X"1044110441104411044110441104411044110441104411044110441104411044",
INIT_18 => X"0401004010040100401004010040100401004010040100401004411044110441",
INIT_19 => X"7D05122890000000003FFFFFFFF9004010040100401004010040100401004010",
INIT_1A => X"E79E79E79E79E79EFFDFF7F5F777DF7DF7DF7EFF7BFA3FC7DF7AF5BF7EFDF7DF",
INIT_1B => X"9FCFE7F3F9FCFE7F3F9FCFE7F3F9E79E79E79E79E79E79E79E79E79E79E79E79",
INIT_1C => X"FFFFFFFE00000FE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F",
INIT_1D => X"10000000000000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"FFFFFFFFFEBA5D2E974000800021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_1F => X"21FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E954000004001FFFFFFFFFFFFFFFFF",
INIT_20 => X"FFEBA552A97400002A801FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2A9541008040",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFEBA552A97400082A975FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"2E95400082E975FFFFFFFFFFFFFFFFFFFFFFFFFFEAA552E95410002A955FFFFF",
INIT_23 => X"FFFFFFFFFFFFFFEAA552E95400002E975EFFFFFFFFFFFFFFFFFFFFFFFFFEAA55",
INIT_24 => X"000000000FFFFFFFFFFFFFFFFFFFFFFFDEAA5D2E97410080015545FFFFFFFFFF",
INIT_25 => X"FFFFFFFEBA5D2E97410080002000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974000004001FFFFFFFFFFFFFFFFFFF",
INIT_27 => X"EBA5D2A95410000A001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2A954000804021",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFEBA552A97400082E821FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"95410082A975EFFFFFFFFFFFFFFFFFFFFFFFFFEAA552E97400002E955FFFFFFF",
INIT_2A => X"FFFFFFFFFFFDEAA552E954000020955C7FFFFFFFFFFFFFFFFFFFFFFFFEAA552E",
INIT_2B => X"0015545FFFFFFFFFFFFFFFFFFFFFFFDEAA5D2A974001C24975C7FFFFFFFFFFFF",
INIT_2C => X"00000000000000000000000000FFFFFFFFFFFFFFFFFFFFFBFDEAA5D2A9741014",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800020000000000000000000000",
INIT_2E => X"A5D2A954000800021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974000004001FF",
INIT_2F => X"FFFFFFFFFFFFFFFFFEBA552A95410002E821FFFFFFFFFFFFFFFFFFFFFFFFFFEB",
INIT_30 => X"400002E975EFFFFFFFFFFFFFFFFFFFFFFFFFEAA552A97400082A801FFFFFFFFF",
INIT_31 => X"FFFFFFFBFDEAA5D2E95410082E955EFFFFFFFFFFFFFFFFFFFFFFFFDEAA552E97",
INIT_32 => X"17545FFFFFFFFFFFFFFFFFFFFFBFDEAA5D2A95400080015545FFFFFFFFFFFFFF",
INIT_33 => X"BFDEBA552A974105D0015555FFFFFFFFFFFFFFFFFFF7FBFDEBA5D2A974005504",
INIT_34 => X"0000000000000000000000000000000000000000010FFFFFFFFFFFFFFFFEFF7F",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"01FFFFFFFFE00000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(22),        -- Port A data input
DOA(0)   => data_read_a_lo_256(22),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(22),        -- Port B data input
DOB(0)   => data_read_b_lo_256(22),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_23_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"EF20906D902424807BC8241BC81801B97D38AD3C0800103362A6741C80A12A02",
INIT_01 => X"001FFF8409F089003B4422000D80C80106804A7951C5B9D1C828043EA28838F9",
INIT_02 => X"073B8858218C2C50801000F9FFEFF8E72CA7F5FC2E048026496834D84721DFE0",
INIT_03 => X"2C4360101A4001001005080400401420350016E0BB222341C312000014006FF8",
INIT_04 => X"00017B810015DC03D034201E14000036486008101FC0002EE006297E1C05F561",
INIT_05 => X"7E1F02FFFFC80100004044800080BEFFFC0248005FFC3C18A5FFC2444484BCC0",
INIT_06 => X"4082040800000811224DE0A00005FFBF8000000003FF810640A1C0008FF2F0E1",
INIT_07 => X"D1D72040048D00388387D03D0E591FFD201F862691DFBE077C2BC45B40FFE458",
INIT_08 => X"1FFBFFEC440501A5604B31062356282AA84200D12342113EDC40000004582800",
INIT_09 => X"A890FFF0002023FFDF79000000000EFFE309606020008005FC00000040200000",
INIT_0A => X"000000000037FF50010103134CAFDF03BA18000F39A0106F87D7FA84024B0225",
INIT_0B => X"88300C48907120AC81083315A493886640030010540DFF20FF8610302409000C",
INIT_0C => X"10C1010C1010C1010C1010C1010C1010C10086080860840063090442A18001B1",
INIT_0D => X"0000280600020040030090000012A500003FF7E08181119A41C1443243050C10",
INIT_0E => X"06542C7043FFD5FFF00A04BC010A7724B1000080004000200004150030010004",
INIT_0F => X"B2080290C2909080A872BC4FC8500054840072FC0FC8440054840200705F9861",
INIT_10 => X"0C8220180F1082E00072FC0FC8500054840072BC4FC84400548402214A380380",
INIT_11 => X"19214A380344920080B21810240AB182EB37C380B40800707011001B43253EE5",
INIT_12 => X"0019CE4000026C00C00042BD4149067465910640A0050C060A0028063672A000",
INIT_13 => X"4D801800CCB050001344060211629580B80022480A444111706658280009A203",
INIT_14 => X"944CB232D6D0100C040250200845132C10BE200403018061101A220339C80000",
INIT_15 => X"402102A5493B8E287E03808480060E40C83C1405132C90742E408D0082140820",
INIT_16 => X"0080200802000100100000000000004002403EFFF8002385F034901019465001",
INIT_17 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_18 => X"8020080200802008020080200802008020080200802008020080200802008020",
INIT_19 => X"0000000000000000000000000000080200802008020080200802008020080200",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000004000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFE00000000000000000000000000000000000000000000000000000000",
INIT_1D => X"10080400000000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"FFFFFFFFFEBA5D2E974100000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_1F => X"21FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100004021FFFFFFFFFFFFFFFFF",
INIT_20 => X"FFEBA5D2E954000800001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9740008000",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E954000004001FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"2A954100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2A954100000021FFFFF",
INIT_23 => X"FFFFFFFFFFFFFFEBA5D2A954100800021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_24 => X"0000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA552A97400002A801FFFFFFFFFFFF",
INIT_25 => X"FFFFFFFEBA5D2E97410080400000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800021FFFFFFFFFFFFFFFFFFF",
INIT_27 => X"EBA5D2E974000004001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100004021",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFEBA5D2E954000800001FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"954100004021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2A954000804021FFFFFFF",
INIT_2A => X"FFFFFFFFFFFFEBA5D2A95410000A001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2A",
INIT_2B => X"2E821FFFFFFFFFFFFFFFFFFFFFFFFFFEBA552A97410080E001FFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA552A9740008",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804000000000000000000000000",
INIT_2E => X"A5D2E974100000021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800021FF",
INIT_2F => X"FFFFFFFFFFFFFFFFFEBA5D2E974000004001FFFFFFFFFFFFFFFFFFFFFFFFFFEB",
INIT_30 => X"4000800021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E954000804021FFFFFFFFF",
INIT_31 => X"FFFFFFFFFFEBA552A954100004001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2A95",
INIT_32 => X"821FFFFFFFFFFFFFFFFFFFFFFFFFFEBA552A95410002E821FFFFFFFFFFFFFFFF",
INIT_33 => X"FFFEAA552A97400082A801EFFFFFFFFFFFFFFFFFFFFFFFFFEAA552A97410002A",
INIT_34 => X"00000000000000000000000000000000000000001EFFFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"01FFFFFFFFE00000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(23),        -- Port A data input
DOA(0)   => data_read_a_lo_256(23),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(23),        -- Port B data input
DOB(0)   => data_read_b_lo_256(23),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_24_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100600007FFF000080108004000800020000840041000080808",
INIT_02 => X"172A00D000EF8210000000F9FFEFF8E7240FF1FC224087B1000639401D005FC0",
INIT_03 => X"00003A2E200811000000000400000000340016603A0000004860400014006FFF",
INIT_04 => X"000079800014CC03C034001E04010850300000101FC0002EE000006E1C00F500",
INIT_05 => X"3E1F0067FFC000000000000000003E2FFC024800137C3C0000EFC00000003CC0",
INIT_06 => X"000000000000001123820AA00005FEBF8000000003FF80000021C0000FF0F0E0",
INIT_07 => X"E600084002040A10812A000500590FF9001F95406A8000037230C01840FFE000",
INIT_08 => X"01FBFFEC4695A501604A000C7585080002C200408102F16C0184800026C92C10",
INIT_09 => X"A8107FF0000000FFDF78000000000EFFE001600000000005FC00000000000000",
INIT_0A => X"000000000037FF4000000AA0354000019C4000012800002387D7F804024B0224",
INIT_0B => X"88300C0081408000800001002482886600020010100DFA20FF8600000000000C",
INIT_0C => X"00C1000C1000C1000C1000C1000C1000C1000608006084006301044081800121",
INIT_0D => X"00000000900160000000000000000000003FF7C0010101904181003003000C10",
INIT_0E => X"16100C4043FFD5BFF00004100000000411000000000000000000040030000000",
INIT_0F => X"3A0421080012302010049400086C022004200494000878022004120270599965",
INIT_10 => X"C19240300081406100049400086C022004200494000878022004124819081840",
INIT_11 => X"2348190814C09C01010400132100106836001504240E01040051200200D06410",
INIT_12 => X"202CD680C0100010408240BD80008983596CD86EA84104060503C0B000020250",
INIT_13 => X"0002090164F40086000082062C1B6600BC000C300818044000B27A0043000041",
INIT_14 => X"110002577FE4080C08010842180C40018545BBA00301808A0810C0059AD01802",
INIT_15 => X"4820C04100852B931F00800010081980B042D2044001850ED8808F00050A002C",
INIT_16 => X"0000000000000000000000000000000000003EFFF80037046031E0110001100A",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"9900000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"EFBE7BE7BE7BE7BEC99E61848655D75D7FCB42BBABDB9F3044CB35CF612B4441",
INIT_1B => X"83C1E0F0783C1E0F0783C1E0F07BEFBEFBEF9E79E79E79E79E7BEFBEFBEFBEFB",
INIT_1C => X"FFFFFFFE000001E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F07",
INIT_1D => X"10080402000000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"FFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_1F => X"01FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800021FFFFFFFFFFFFFFFFF",
INIT_20 => X"FFEBA5D2E974100000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741000000",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974100004021FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"2E974000800021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974000004001FFFFF",
INIT_23 => X"FFFFFFFFFFFFFFEBA5D2E974000800001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_24 => X"0000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E954000800001FFFFFFFFFFFF",
INIT_25 => X"FFFFFFFEBA5D2E97410080402000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFF",
INIT_27 => X"EBA5D2E974100800021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800021",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFEBA5D2E974100000001FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974000004001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100004021FFFFFFF",
INIT_2A => X"FFFFFFFFFFFFEBA5D2E974000004001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E",
INIT_2B => X"00001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E954000800021FFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9540008",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804020000000000000000000000",
INIT_2E => X"A5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FF",
INIT_2F => X"FFFFFFFFFFFFFFFFFEBA5D2E974100800021FFFFFFFFFFFFFFFFFFFFFFFFFFEB",
INIT_30 => X"4100000021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100000001FFFFFFFFF",
INIT_31 => X"FFFFFFFFFFEBA5D2E974000004021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E97",
INIT_32 => X"021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974000004001FFFFFFFFFFFFFFFF",
INIT_33 => X"FFFEBA5D2E954000804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E954000004",
INIT_34 => X"00000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(24),        -- Port A data input
DOA(0)   => data_read_a_lo_256(24),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(24),        -- Port B data input
DOB(0)   => data_read_b_lo_256(24),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_25_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100200002000000080100004000000020000800041000080808",
INIT_02 => X"1000218000000800000000F9FFEFF8E738FFF1FC20400400000004455A375FE0",
INIT_03 => X"00002000000001000000000400000000340016623A0000004000000014006FFF",
INIT_04 => X"924279824C94CC1BE0B4001F20000000020380401FE0082EF000106E1C00F500",
INIT_05 => X"3E1F0067FFE048002582800100523E2FFE024820137C3C0040EFE02000003CE4",
INIT_06 => X"821B0821B8019819200020200005FEBF81C1002203FF80000021C1140FF8F0E0",
INIT_07 => X"00040000000000000000000500590FF9001F0000000000033020C01840FFFC78",
INIT_08 => X"01FBFFFD0004000100502000011400000282004001020000000001009015C000",
INIT_09 => X"B8DA7FF8004000FFDF7C062031863EFFF75D78004001010DFC00002005010000",
INIT_0A => X"000000000037FFC00602000000000001980400002800032387D7FE94FBEF2B2C",
INIT_0B => X"88300C0080400000800001002486887600020110100DFA20FF8603000000000C",
INIT_0C => X"00C1000C1000C1000C1000C1000C1000C10006080060840077330C4889CC2925",
INIT_0D => X"00000000000000000000000000002500003FF7C0010101904189003003000C10",
INIT_0E => X"06140C6043FFD5BFF00A04B80608003CB120C110608830445821140134120800",
INIT_0F => X"02000000000200200000900000400200000000900000400200000200701E1861",
INIT_10 => X"0002000000010000000090000040020000000090000040020000000008080000",
INIT_11 => X"0000080800008000000000010100000022000000040000000040000000002400",
INIT_12 => X"0000420000000010000040318020000041000001000244000000008008000010",
INIT_13 => X"0002000004100000000080000002040040000000001000400002080000000040",
INIT_14 => X"0100000042000010002000001000400000042000040200000000400008400000",
INIT_15 => X"0030800000010800000000C0A000000000400000400000040800000000000004",
INIT_16 => X"41104451044C82082068C0200000008014023EFFFC0063046020801000001000",
INIT_17 => X"1104411044110441104411044110441104411044110441104411044110441104",
INIT_18 => X"1044110441104411044110441104411044110441104411044110441104411044",
INIT_19 => X"A080800002FFFFFFFFFFFFFFFFFC110441104411044110441104411044110441",
INIT_1A => X"41041249041249042824014C48569A69AFEE8A252865AA3168A4CBDF860EC15D",
INIT_1B => X"58AC56231188C46231188C462312492492492492492492492490410410410410",
INIT_1C => X"FFFFFFFE00002C562B158AC562B158AC562B158AC562B158AC562B158AC562B1",
INIT_1D => X"10080400000000000000000000000000000000000000000000000001FFFFFFFF",
INIT_1E => X"FFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_1F => X"01FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFF",
INIT_20 => X"FFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008040",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800021FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"2E974100000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800001FFFFF",
INIT_23 => X"FFFFFFFFFFFFFFEBA5D2E974100000021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_24 => X"0000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100000001FFFFFFFFFFFF",
INIT_25 => X"FFFFFFFEBA5D2E97410080400000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFF",
INIT_27 => X"EBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974100800001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800021FFFFFFF",
INIT_2A => X"FFFFFFFFFFFFEBA5D2E974100800021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E",
INIT_2B => X"00001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100000021FFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741000",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804000000000000000000000000",
INIT_2E => X"A5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FF",
INIT_2F => X"FFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEB",
INIT_30 => X"4100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFF",
INIT_31 => X"FFFFFFFFFFEBA5D2E974100800001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E97",
INIT_32 => X"021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800021FFFFFFFFFFFFFFFF",
INIT_33 => X"FFFEBA5D2E974100000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800",
INIT_34 => X"00000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"01FFFFFFFFE00000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(25),        -- Port A data input
DOA(0)   => data_read_a_lo_256(25),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(25),        -- Port B data input
DOB(0)   => data_read_b_lo_256(25),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_26_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"E9264EAB20190CA3BA4997AA9002AE9C001006B0778015CFA17E0811039879C7",
INIT_01 => X"F1FFF9BB1F773C7F9BB07DFFFDD863FC5FFF3FEFFBBF9FFB22FFFBC7B9F30686",
INIT_02 => X"1B33188302E708180F6FFBFFFFCFFFFF9C7FF7FC24350B99082400001D00DFD8",
INIT_03 => X"4A53D958C50000DCE7366303739CD98C27C57EF57980014F271807E3C9E9CFF8",
INIT_04 => X"DBFAFBD7FB1CDEBEF1BE17F7AC88042787FBFFF8FEE9FF7EE6F4C0EE1FFAF869",
INIT_05 => X"BE1FFD67DFFEFFBDA7F7FED508707E2EFEBF6FFEB37C3FF302EEEDFF9B487CF6",
INIT_06 => X"75F7275F7CAC98E261EDF0253C7FFFEF87C74E8CCFFBB6FF70E1FE61FFBDF0FE",
INIT_07 => X"73840C07783060C72DF7D828912E6FFB80162776F3BFB7077E82255E40BFEEBA",
INIT_08 => X"69FFBFE43C872321367036163F1C0820A3063F460D1AEFC000060042648C4181",
INIT_09 => X"FB967FBD13D981F7DF7D7E6171AF3FEFE8A3E679FAC1FD1FFFBEB000763A8447",
INIT_0A => X"6AED1D1DAD7FBE7D67D7F3BB79CFFB83BF14EC1E7D7300B017F5FFE6FBEF73BE",
INIT_0B => X"99F51EDDCDEBCFF589807B70AD9A99EE7583F931109FFE33FF8E3FDFDAF64A3C",
INIT_0C => X"C0D78C0D78C0D78C0D78C0D78C0D78C0D7A606BC606B8C56F7730ECCDBDF1521",
INIT_0D => X"1D406B9EC20181CC1F73F87501DED3409BFFFEFFEBF341B867D3683A03A40F78",
INIT_0E => X"86D70CE04FFFFF3FF1F5F5475BD7F72E4D75EBFAF5FD7AFEFDFFAF59B6FF28FE",
INIT_0F => X"020007C040101480807D17B0004001F804007D17B0004001F8040212F35FFC6D",
INIT_10 => X"700200001DC00068007D17B0004001F804007D17B0004001F804006F60081400",
INIT_11 => X"206F60081800800007B000102C0801FB02683800040007700011801003DE050A",
INIT_12 => X"403E232130207080D012CEFF41008D188D502100B02004000F01900039020040",
INIT_13 => X"0E101A01F21A2C40039006823F80048100003F0008004D8100F90D162001C803",
INIT_14 => X"B604027F020A07400007C040085581019D602451500001EC00100247C4642608",
INIT_15 => X"CC3F02010EA40EA00020C830100F0D000022180581019F40084800001F100020",
INIT_16 => X"EBFAFEFFBFEFDFDDFE7DD87FEFF7FF796FFFFFDFFC017FEFFD7E841001D8197D",
INIT_17 => X"BFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAF",
INIT_18 => X"FAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFE",
INIT_19 => X"EDB5C88646FFFFFFFFFFFFFFFFFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEB",
INIT_1A => X"61861A69A6986186EBCAF55357E1C71C751D6C56F3D247859B3214FA76953F86",
INIT_1B => X"84C26130984C26130984C2613098618618618618618618618618618618618618",
INIT_1C => X"FFFFFFFE0000026130984C26130984C26130984C26130984C26130984C261309",
INIT_1D => X"10080400000000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"FFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_1F => X"21FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFF",
INIT_20 => X"FFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008040",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFF",
INIT_23 => X"FFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_24 => X"0000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFF",
INIT_25 => X"FFFFFFFEBA5D2E97410080400000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFF",
INIT_27 => X"EBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFF",
INIT_2A => X"FFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E",
INIT_2B => X"04021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804000000000000000000000000",
INIT_2E => X"A5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FF",
INIT_2F => X"FFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEB",
INIT_30 => X"4100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFF",
INIT_31 => X"FFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E97",
INIT_32 => X"001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFF",
INIT_33 => X"FFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804",
INIT_34 => X"00000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(26),        -- Port A data input
DOA(0)   => data_read_a_lo_256(26),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(26),        -- Port B data input
DOB(0)   => data_read_b_lo_256(26),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_27_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"00080A40000A41248002029000050A088000008242A0004404480002000A1155",
INIT_01 => X"F1FFF1C11F781C129C107DFFFE0860941E81258CA2B71C2220EC1B86E1A00002",
INIT_02 => X"4000002100000014400FF6FFFF0FFFFF8007F1FC211100014200800000887FC0",
INIT_03 => X"0842D85841000098C63061026318C18404C459757000015F00088BE3C0618FF8",
INIT_04 => X"DBEAE5D6D91C2EBCE1B21EA72C00000007FBE7C8F8E9EF79E6D440E91FDAE061",
INIT_05 => X"B91FF9671FE6B68984B5BCE408347E28FEBF6FEEB3723F7102E8EDBF8A4872F6",
INIT_06 => X"3573A357308418E40000D4113C7FFE4F86064C8DDFE3B6FF50D1FC61DE39C8FC",
INIT_07 => X"00000A20083060C00C81882A008C6FF880060424B39FB6037F00051C003FE04A",
INIT_08 => X"61FA3FE4010440410844060001040A00002200460D1A06000005040000001080",
INIT_09 => X"EB027E390A4881C7BEFC5F6171CE2F8FE823E778DAC16C1FFBBC900031589547",
INIT_0A => X"03813030213C3E2D62D6E21259CFDB039E806C024531008017C1F826FFEF41FE",
INIT_0B => X"9AB55F0DEFABC705488069302DBA98EAB582D835109FFC31FFAEAFCFDAF4423D",
INIT_0C => X"40C3440C3440C3440C3440C3440C3440C3C2061A2061AD46FF730E5CCBCD5521",
INIT_0D => X"0C407D1F820101441DA3A8310198C34089BFF8DD6B7941BC63F1683803C00E34",
INIT_0E => X"5710AE4047FFD23FF315D54358D593474955AB6AD5B56ADAB5FAAE58B2F628EA",
INIT_0F => X"020007C0400004C080791290004001D80001791290004001D8000210F1587971",
INIT_10 => X"300200001DC0000801791290004001D80001791290004001D800012F60080400",
INIT_11 => X"202F60080800800007B000000E0801BB020828000400077000008210035E0408",
INIT_12 => X"40BA2220202070801010C6F1410085188D500100102004000F01900031000060",
INIT_13 => X"0E100205D2120840039000813F80040100003F0000000F8100E909042001C800",
INIT_14 => X"3E04007F020201400007C040001781011D602040500001EC0000005744440408",
INIT_15 => X"C43F02000EA40EA000004810100F0D000020080781011F40080800001F100000",
INIT_16 => X"AB6ADAB6BDE75ED5EC71385FC2512E3565BBBF1FFC00636EED7E841000D81924",
INIT_17 => X"B6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6AD",
INIT_18 => X"6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADA",
INIT_19 => X"A471688747FFFFFFFFFFFFFFFFFAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB",
INIT_1A => X"0020800000000000780401CBC840000005243885A04012072A1810DA84002104",
INIT_1B => X"5028140201008040201008040200000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFE000028140A05028140A05028140A05028140A05028140A05028140A0",
INIT_1D => X"10080400000000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"FFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_1F => X"01FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFF",
INIT_20 => X"FFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008040",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFF",
INIT_23 => X"FFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_24 => X"0000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFF",
INIT_25 => X"FFFFFFFEBA5D2E97410080400000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFF",
INIT_27 => X"EBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFF",
INIT_2A => X"FFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E",
INIT_2B => X"04021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804000000000000000000000000",
INIT_2E => X"A5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FF",
INIT_2F => X"FFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEB",
INIT_30 => X"4100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFF",
INIT_31 => X"FFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E97",
INIT_32 => X"021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFF",
INIT_33 => X"FFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804",
INIT_34 => X"00000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"01FFFFFFFFE00000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(27),        -- Port A data input
DOA(0)   => data_read_a_lo_256(27),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(27),        -- Port B data input
DOB(0)   => data_read_b_lo_256(27),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_28_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"02200AA400180030808802A900002A08001280A08A801044104A1000001818C3",
INIT_01 => X"50A00011460214428114180000882214413D0A71592A01D92213D28005210202",
INIT_02 => X"1444428102100884000AA30200000000C1000401041108404400022220800000",
INIT_03 => X"461080404900000C6314A900318C52A40051081000888806108802A141288001",
INIT_04 => X"00800040110102000902002000888400081045A8A00003C00000500000080008",
INIT_05 => X"0000000000024CA0A0101800032000400000000B800000014000000B08180000",
INIT_06 => X"10280102802C0240041000011428004022220024440013511000013510000000",
INIT_07 => X"0804420009122448451020100020400080002041000000008000010400000880",
INIT_08 => X"2800000140200808021006108010422AAA800022448902849220114009224081",
INIT_09 => X"01C800004080A0000002480B04008100011000088800081002C19020150B0013",
INIT_0A => X"56D29A9A52800004004070208000000040006408001100105000020000001800",
INIT_0B => X"00040024440245400082D0220800008010001020458000010000040D96104210",
INIT_0C => X"50160501605016050160501605016050160280B0280B00120008430660210014",
INIT_0D => X"054001884200810C1631181500CA60400B4008072020500002002C0040010360",
INIT_0E => X"104420A00C000200005000010040A0020CC000200010000800920040804020A6",
INIT_0F => X"0000000000001400000102900000002800000102900000002800001001802104",
INIT_10 => X"3000000000000048000102900000002800000102900000002800000020000400",
INIT_11 => X"0000200008000000000000002800000100082800000000000001800000020008",
INIT_12 => X"4000202020200000901005480000000800000100102000000000000009000000",
INIT_13 => X"0000120002020840000004800080000100000000000048800001010420000002",
INIT_14 => X"A200000800020140000000000050800008000040500000000000024004040408",
INIT_15 => X"840A000002000000000048100000000000020800800008000008000000000000",
INIT_16 => X"8020080210810840861CD33548542A10209D4100000010200400000000880035",
INIT_17 => X"0200802008020080200802008020080200802008020080200802008020080200",
INIT_18 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_19 => X"40A0C22E10000000000000000000020080200802008020080200802008020080",
INIT_1A => X"08208208208208200360D4141D630C30C7788440B044280091A5CB03D01BD89A",
INIT_1B => X"582C16030180C06030180C060302082082082082082082082082082082082082",
INIT_1C => X"FFFFFFFE00002C160B0582C160B0582C160B0582C160B0582C160B0582C160B0",
INIT_1D => X"10080400000000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"FFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_1F => X"01FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFF",
INIT_20 => X"FFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008040",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFF",
INIT_23 => X"FFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_24 => X"0000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFF",
INIT_25 => X"FFFFFFFEBA5D2E97410080400000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFF",
INIT_27 => X"EBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFF",
INIT_2A => X"FFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E",
INIT_2B => X"04001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804000000000000000000000000",
INIT_2E => X"A5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FF",
INIT_2F => X"FFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEB",
INIT_30 => X"4100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFF",
INIT_31 => X"FFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E97",
INIT_32 => X"001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFF",
INIT_33 => X"FFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804",
INIT_34 => X"00000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"01FFFFFFFFE00000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(28),        -- Port A data input
DOA(0)   => data_read_a_lo_256(28),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(28),        -- Port B data input
DOB(0)   => data_read_b_lo_256(28),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_29_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"79964E4BA01DACAB9E659792D00AAE160002829C7FDFEFCEE97C2815039D70C3",
INIT_01 => X"50BFF9AB0775343F9AB01DF80D5821FC0FFF3FEFD1AF9FF1207FFBC7B9720586",
INIT_02 => X"0B33180300E700080F6AAA7BFFC007189C7FF2FC003503980A0000001D00DFD8",
INIT_03 => X"0401D940CD0000C8421A2B03210868AC23403E903900010E271006A148A0C000",
INIT_04 => X"49B87A417315D20A313E17F1800000058013DDF8BE21F36E02F0D06E03E8F800",
INIT_05 => X"3E00FC67C03A4D9C87525E5101603E6E023D27DA937C03E340EE25CB9B483C12",
INIT_06 => X"50B5050B540C004261EDE025142DFFE003C30E0447F877F930203E213F8CF01E",
INIT_07 => X"73800407781020476467D008910A4FFB80100332D1AE93059282215E40800678",
INIT_08 => X"21FF80003C832320342036063F08000001063F42050AEB4000221000248C0180",
INIT_09 => X"51547F8C1111A0F041056A0100A11FE000916249A800B915FE82B02052290002",
INIT_0A => X"2AAD1515AD5780540541619968C76980E914E4163D53002017F405C409A42A9A",
INIT_0B => X"014002D445624DB481806A6288100184500171200085FE030000157FDF124A10",
INIT_0C => X"D0068D0068D0068D0068D0068D0068D006A68034680300021410028450530014",
INIT_0D => X"15402B0E8201018C1561E855008C50401B7FFE27A0B2500806522C0A40A50268",
INIT_0E => X"928324400DFFFF0001F1F0050342D42A086040B02058102C48970541944B20FA",
INIT_0F => X"0000000000101480000507B00000002804000507B000000028040212034FAD28",
INIT_10 => X"7000000000000068000507B00000002804000507B00000002804004020001400",
INIT_11 => X"0040200018000000000000102C0000410068380000000000001180000082010A",
INIT_12 => X"4004212130200000D0120ED64000080800002100B02000000000000009020040",
INIT_13 => X"00001A00220A2C4000000682008000810000000008004D800011051620000003",
INIT_14 => X"B6000208000A0740000000000855800088000451500000000010024084242608",
INIT_15 => X"8C0F0001020000000020C8300000000000021805800088000048000000000020",
INIT_16 => X"C0B02C4B12C989489418D13FE7F3FFD8BADB7FC004012CA5141600000198087D",
INIT_17 => X"0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02",
INIT_18 => X"B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C",
INIT_19 => X"FEA0C00602FFFFFFFFFFFFFFFFFC0B02C0B02C0B02C0B02C0B02C0B02C0B02C0",
INIT_1A => X"FBAEBAEBAEBAEBAEFFFFF7E7EFBFFFFFFAEF3E7E5BB9FFF7DFF9E3F08843FFDF",
INIT_1B => X"FDFEFF7FBFDFEFF7FBFDFEFF7FBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBE",
INIT_1C => X"FFFFFFFE00003EFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FB",
INIT_1D => X"10080400000000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"FFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_1F => X"01FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFF",
INIT_20 => X"FFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008040",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFF",
INIT_23 => X"FFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_24 => X"0000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFF",
INIT_25 => X"FFFFFFFEBA5D2E97410080400000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFF",
INIT_27 => X"EBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFF",
INIT_2A => X"FFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E",
INIT_2B => X"04001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804000000000000000000000000",
INIT_2E => X"A5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FF",
INIT_2F => X"FFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEB",
INIT_30 => X"4100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFF",
INIT_31 => X"FFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E97",
INIT_32 => X"001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFF",
INIT_33 => X"FFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804",
INIT_34 => X"00000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(29),        -- Port A data input
DOA(0)   => data_read_a_lo_256(29),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(29),        -- Port B data input
DOB(0)   => data_read_b_lo_256(29),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_30_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"FD00000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"E79E79E79E79E79EEBFEF5D7D7F7DF7DFFDFFEFFFBFE7F87DFFEFFBF77BFFFDF",
INIT_1B => X"9FCFE7F3F9FCFE7F3F9FCFE7F3F9E79E79E79E79E79E79E79E79E79E79E79E79",
INIT_1C => X"FFFFFFFE00000FE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F",
INIT_1D => X"10080400000000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"FFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_1F => X"01FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFF",
INIT_20 => X"FFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008040",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFF",
INIT_23 => X"FFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_24 => X"0000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFF",
INIT_25 => X"FFFFFFFEBA5D2E97410080400000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFF",
INIT_27 => X"EBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFF",
INIT_2A => X"FFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E",
INIT_2B => X"04001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804000000000000000000000000",
INIT_2E => X"A5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FF",
INIT_2F => X"FFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEB",
INIT_30 => X"4100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFF",
INIT_31 => X"FFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E97",
INIT_32 => X"001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFF",
INIT_33 => X"FFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804",
INIT_34 => X"00000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(30),        -- Port A data input
DOA(0)   => data_read_a_lo_256(30),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(30),        -- Port B data input
DOB(0)   => data_read_b_lo_256(30),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_31_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"129000008004A00804A40000400800020000000C005FEA005800200400050100",
INIT_01 => X"A15FF18019700810180065FFFC0040801E80258CA2951C2200EC0906A0804140",
INIT_02 => X"0000000000000011000550FDFF0FFFFF0007F1FC200000011000000000205FC0",
INIT_03 => X"08425818000000908428C0024210A30004045060302223490002014280410FF8",
INIT_04 => X"DB6A618248140C18E0B016872400000007EBA24058E1ECA8E2D400681FD0E061",
INIT_05 => X"381FF8671FE01009048084C400103E28FE3F6FE513703F7000E8E5B4825030F6",
INIT_06 => X"00130001300018A00000D0002855FE0F84040C088BE3E4AE40C1FD04CE38C0FC",
INIT_07 => X"000008800020408008818838000C2FF800060424B39FB6037E000418003FE008",
INIT_08 => X"41FA3FE400040001004000000104088000020044091204000004000000000000",
INIT_09 => X"E8027E38004801C79E7C162231862E8FE00166704041240DF93D000000000004",
INIT_0A => X"0000000000343E002202021259CFDB039E0008024520000047C1F804FBEF01BE",
INIT_0B => X"88310E08812982050800A9102492986200824810110DFC30FF86036249E4002C",
INIT_0C => X"00C1000C1000C1000C1000C1000C1000C18006080060840477330C4889CC0121",
INIT_0D => X"08006816800100400902A0200110810080BFF0C80111019861D1403803800C10",
INIT_0E => X"06100C4043FFD03FF101D4000800130401808100408020401020041830120848",
INIT_0F => X"020007C04000008080781000004001D00000781000004001D0000200F0185861",
INIT_10 => X"000200001DC0000000781000004001D00000781000004001D000002F40080000",
INIT_11 => X"202F40080000800007B00000040801BA020000000400077000000010035C0400",
INIT_12 => X"003A0200000070800000C231410085108D500000000004000F01900030000040",
INIT_13 => X"0E100001D0100000039000003F00040000003F000000050100E808000001C800",
INIT_14 => X"14040077020000000007C0400005010115602000000001EC0000000740400000",
INIT_15 => X"403502000CA40EA000000000100F0D000020000501011740080000001F100000",
INIT_16 => X"01004010044602002061004A820104809402BE1FFC006304E036841000501900",
INIT_17 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_18 => X"0040100401004010040100401004010040100401004010040100401004010040",
INIT_19 => X"0001000802FFFFFFFFFFFFFFFFF8100401004010040100401004010040100401",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFE00000000000000000000000000000000000000000000000000000000",
INIT_1D => X"10080400000000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"FFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_1F => X"01FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFF",
INIT_20 => X"FFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008040",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFF",
INIT_23 => X"FFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_24 => X"0000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFF",
INIT_25 => X"FFFFFFFEBA5D2E97410080400000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFF",
INIT_27 => X"EBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFF",
INIT_2A => X"FFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E",
INIT_2B => X"04001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804000000000000000000000000",
INIT_2E => X"A5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FF",
INIT_2F => X"FFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEB",
INIT_30 => X"4100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFF",
INIT_31 => X"FFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E97",
INIT_32 => X"001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFF",
INIT_33 => X"FFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804",
INIT_34 => X"00000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(31),        -- Port A data input
DOA(0)   => data_read_a_lo_256(31),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(31),        -- Port B data input
DOB(0)   => data_read_b_lo_256(31),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_0_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"ED39BA795990D275FB4A6E96ACC4731DEA4598B0AFB54867F6EE4618C3749807",
INIT_01 => X"58A0047D8607944AC7DA180001ECA2544042106208408208C20022E9173734B3",
INIT_02 => X"9F775E7CB273E6CCA7DAAF00001000000478020113C9C38E09FB7CCCDD9F203E",
INIT_03 => X"441406267B4CB04443163C91110C58F24A31000B8028A810A3D0F8B169A01006",
INIT_04 => X"0005802424830120024121209088809DF81454ACA01E03501D0A3B91E00F0A00",
INIT_05 => X"C1E0039800112014C20B0232838F80D001C0100AEC83C008EF101A034C8CC300",
INIT_06 => X"8B0478B04A83405954592F9B9628000002C3F08754001B51881E007900060F01",
INIT_07 => X"39F36677EE1C387777622717EF711004A6818111086008E080FDC30594001017",
INIT_08 => X"160400195E83A3A0F61BC3929ECB622AABF5FF83860CEB164833F179B48CEE59",
INIT_09 => X"036D8004FDB47600000229410C61010016DC998C84B0128202C0DCB48F05D513",
INIT_0A => X"204122A033000182502440888420247041E876810099D35F900002DB00105C01",
INIT_0B => X"41C000947E16656074EA560F080544900960260144D201890018080D36191110",
INIT_0C => X"781EA781E2781EA781E2781EA781E2781C33C0613C0E00120800239450112ED4",
INIT_0D => X"872917095352BD2A90515A1CA44E7EA84B00001010043803120C3E04E03383E2",
INIT_0E => X"70C7E0B92800224008AE09B8942C48D1FC491204890244812250588601285432",
INIT_0F => X"B80C2038ABACB83C7E03EA5FF83C002783F103EA5FF83C002783F0120847A704",
INIT_10 => X"BD9870380230F2D7C103EACFF83C002783F103EACFF83C002783F310BBF7EFC2",
INIT_11 => X"1F10BBF7EFC61E01804E1E6EA1E3FA01FD97EFC4B80E008C7C2F678FF023FAF5",
INIT_12 => X"B801FCC8E8320C4DAC9220C6B2FF22EF72ADDE6F1A67C80600C2683E0EF8AE1F",
INIT_13 => X"4189B5C00FE651C6104C6D6400FFFB01FC0000FC07EE42FA7C07F22CE3082636",
INIT_14 => X"8BE9FC08FDF4195C0C2038A7C6CAFA7E289F9BA4570380131CAFB2003F9D190A",
INIT_15 => X"270AE9FE635BE11B7F0308D4A80092E0FC1FC662FA7E283FF68A8F0080AE1DDA",
INIT_16 => X"1204812058112C12411402056954AB0C280D000003350013024179498C2EC6B9",
INIT_17 => X"2048120481204812048120481204812048120481204812048120481204812048",
INIT_18 => X"0481204812048120481204812048120481204812048120481204812048120481",
INIT_19 => X"13043A85D4000000000000000001204812048120481204812048120481204812",
INIT_1A => X"82082082082082082218821390771C71C557CE263826D5B1D36AC59E0765D1CF",
INIT_1B => X"1F0F87C3E1F0F87C3E1F0F87C3E0820820820820820820820820820820820820",
INIT_1C => X"FFFFFFFE00000F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E",
INIT_1D => X"EF5D7BD7400000000000000000000000000000000000000000000061F007FFFF",
INIT_1E => X"A10A2D1574005D0428A10A2AAA8BEF552EBDFFF557BC01FF5D7BFFEBA5D55555",
INIT_1F => X"DEBAFFFFC2000AA8428AAAFFAAA8BFF00002AA10FF802ABEFA2D16AA00F7FBE8",
INIT_20 => X"975EFFF8002010002EAAAAAAAD1555FFFFAEA8B550051401450055575FF00517",
INIT_21 => X"4155FF0855575455D2AA8BFFA2D1575EF5D5555545FFFBE8A00087FC20BA5D2A",
INIT_22 => X"8028A00FFAE800AA082A820005D2E974BAA2D140145A2842AA00A284021FF5D0",
INIT_23 => X"2D17FFEF000017400FFD1555FF007FFFEBA55042AA00000017400FFAABFEBAFF",
INIT_24 => X"000000155F7D540000F7FBFFE105D7BE8ABAA284000105D0428BFFA2FBFDFFFA",
INIT_25 => X"75D7BFAEBA5551501D51C5FC7E00000000000000000000000000000000000000",
INIT_26 => X"28B6D16AA28EBF5EDA38AADE1543849557D492BF8E2DE00552EBFFC7552BC01D",
INIT_27 => X"000A85400E00E38A175FDE3F5C002DAAD42DAAAF784AFA82BC042DF47E3D1F80",
INIT_28 => X"AA150021C0092490E904BAFFD550A90FFA495FC7A05B555C257AAA8B45007540",
INIT_29 => X"2DA02402ABD4AD1D0E175D7140B455D516A1EAB45E2A000B4748717A095F571E",
INIT_2A => X"4004A8BC0ABFF7D03A17D1D5147540B454AA080038E9748542AE3D0051C7B6F0",
INIT_2B => X"FB6D4B8FC7BFFFD2168B68F57492F505FF5FA550490BFA482B420B8428A3DA85",
INIT_2C => X"0000000000000000000000016ABD554201543A1EDE9016D4AAB454AF400547AB",
INIT_2D => X"5D2EBDF55556BC35E7557FE8AB25D11415FD0151614000000000000000000000",
INIT_2E => X"9596CBEA41D7D3DECFAF7D43FABAAAD57DEBAAAFFD74AA04547EE18D680BE9A5",
INIT_2F => X"47D78228E5000EA422E10439C1FBCD282351BDAAF9C20AAAABCBEB1DFF803FC5",
INIT_30 => X"1E6284683ABBDD7DEAA100069C14B25495A00F38EBAC0E198B97605018053575",
INIT_31 => X"4408FE6A755ED8EFEFE41B2D17EAF02552BC0545556BD61E501001DF5DD3EBA3",
INIT_32 => X"556F922ACA8AB8283C8310FAB1588916D3861C0422C44082B52A81550A828141",
INIT_33 => X"A5FDBCD7D262E5AFAC4B6AADDD562AF57D7C369AF25495A23068A8301BA7FB95",
INIT_34 => X"003FE0000003FE0000003FE0000003FE0000003FE03D5789700282E9FEFB501E",
INIT_35 => X"0003FE0000003FE0000003FE0000003FE0000003FE0000003FE0000003FE0000",
INIT_36 => X"00000000000000000000000000000000000000000000000000000000003FE000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(0),        -- Port A data input
DOA(0)   => data_read_a_hi_256(0),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(0),        -- Port B data input
DOB(0)   => data_read_b_hi_256(0),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_1_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"212C001411984004084D000508C53810A03D1450E839B003342114428A000807",
INIT_01 => X"08000010400A0008010600000084004000400002000000000000000000140000",
INIT_02 => X"484DEBA0111800C004400D000000000028800001CC404E6008B4933336880010",
INIT_03 => X"650C00000848A0423183089008C604224200000100A200002C280810098C0001",
INIT_04 => X"00000004208B00200E010800006667BE7000102C00080000040012010000080C",
INIT_05 => X"0100000000002000600100208D04414000800000000200004800080000800200",
INIT_06 => X"010420104032C204071200000200000010104020000001000910000000040800",
INIT_07 => X"8C0060242183060CF118011281B00000220010400020002081A0008210000802",
INIT_08 => X"000400014812466427040098C000622AAAA43E3060C158AC97F0356BDBFBD008",
INIT_09 => X"026C000559102400200281400469000008B0800000901080004004308B434040",
INIT_0A => X"50502A2800800000400408200000201041000208000040020820034200005C00",
INIT_0B => X"13C051112A800008402002021128000081202205001000000028880004010500",
INIT_0C => X"191AC191A4191A4191AC191AC191A4191A00C8560C8D2940804060901210441E",
INIT_0D => X"C1C114417882F82C00181707044212080300001002081224002006406401918C",
INIT_0E => X"60C0C0B92C000000000400001004200044010200810040802040080200284401",
INIT_0F => X"380C200000043C2016000000F03C00280030000000F03C00280030000004860C",
INIT_10 => X"8D18703800000049C0000000F03C00280030000000F03C002800321080000BC2",
INIT_11 => X"0110800007861E0180000002A9001A00000007C4380E00000001E00230000000",
INIT_12 => X"688004C0C81200009480010280340000008082430A07C80600C0000009008610",
INIT_13 => X"4000134400241186100004A500007B00FC000000000E4A402C001208C3080002",
INIT_14 => X"A9002C0001E0181C0C200000025A400A200812A4070380000000B25000981902",
INIT_15 => X"0000804A0002410A170300C4A800800000020E22400A200096828F008000000A",
INIT_16 => X"020080200820040041002000010080000000000002340002004118010C228614",
INIT_17 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_18 => X"0080200802008020080200802008020080200802008020080200802008020080",
INIT_19 => X"2B5000A000000000000000000000200802008020080200802008020080200802",
INIT_1A => X"AA8A28A28A28A28AB2048634B03249249604CA291AEAFBF1528205C00020C745",
INIT_1B => X"974BA5D6EB75BADD6EB75BADD6EAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA",
INIT_1C => X"FFFFFFFF00000BA5D2E974BA5D2E974BA5D2E974BA5D2E974BA5D2E974BA5D2E",
INIT_1D => X"55AAAAAAA00000000000000000000000000000000000000000000181FFFFFFFF",
INIT_1E => X"BEF5D7BE8ABA5D557DFEFFFD17FEBA00042AAAAFFFFFFE00FF843DF45FFAE955",
INIT_1F => X"DFEF552A800AA5555575FFA2AE820BAFFAEBFF555500155EF552E975FFF7D168",
INIT_20 => X"6AA00A2FBEAABA5D55420AA00002AA00AAFBE8B55A280175455D002AA00A2AAB",
INIT_21 => X"BD75FFAA802AAAAFFAA801EF00517FFFFF7D56ABEF0004155550004154105D55",
INIT_22 => X"55575FF08557DEBAA2FBEAAAA552E955EF5D0415410A2AE97545A2AE954BAF7F",
INIT_23 => X"7D17DF55A2AEBDEAAFFFFC20AAFFFFFFFFFAAD5555FFFFAEAAB55A2D168B555D",
INIT_24 => X"0000000BAFFFBE8A00087FC20BA5D2A975EF5D0002010552E820AAFFD57FF55F",
INIT_25 => X"8FF8A38F45F7AA9217FA380AD400000000000000000000000000000000000000",
INIT_26 => X"D7552E975EFFFDF68BFF557BEAA925551785D7BFD5EFE3F08002FA92EBA5FDE2",
INIT_27 => X"43841017DE92BF8E3AA824924870BF5551555C7A28A821EFE3AABAE38005B575",
INIT_28 => X"0568005A1041055716DB7DB6FBEFEA81C55D0A0516802AA28BEF5EDB7DAA8A15",
INIT_29 => X"C7FEF1C043FE28E3FBD55FFAADE2DAAAE3A5C51C71C042DF45A3D1D00281E8A1",
INIT_2A => X"AA8B45B47F6FB55A95555E90F78E17F52FEF5EDA82FD249057F080417492AAAF",
INIT_2B => X"5FF8AAAA95B7AF45FF8F7DFEDFFAFF8E005FAE92A3AE3DBFF57FA2DF555D257A",
INIT_2C => X"000000000000000000000000A8F571EAA150021C0092490E905FFFD0550BD75C",
INIT_2D => X"00043DE00A2C57DE08FFAAA8B55F7EE801F7F2849EE000000000000000000000",
INIT_2E => X"6AAAE29F067155543A15D2E955EFFFFBEABEF557FEAA10595169BED83D1EBCA8",
INIT_2F => X"BAFFD57DEEAAA15976EB0444BFEB086808A8E3082C954BA5D7DD6145AAAA821A",
INIT_30 => X"B47FFD55D6107782001FF0812000A255D57FFBEF3B97EEAB2C40217B9778428A",
INIT_31 => X"35FF003F17418AEE817B540D11CA80BAAFA825EFAABEBCA18FE803755D08079E",
INIT_32 => X"8BDEBA2D757547D7862AF57ABFFCABE5553FD5FBEFE86353EFFFD03FE0275000",
INIT_33 => X"5A01F70C6AA04537957D6FB4807FFFB45F7EFFDA58FF2AA88A0F3C5014018AC2",
INIT_34 => X"00000000000000000000000000000000000000000B2DD7DEAA100069C14B2549",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(1),        -- Port A data input
DOA(0)   => data_read_a_hi_256(1),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(1),        -- Port B data input
DOB(0)   => data_read_b_hi_256(1),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_2_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10E006600180111284380310006289800480032283E000A34301002001A0816",
INIT_01 => X"0005A00810790848048044A54E404340404000720885800802000806EC910200",
INIT_02 => X"5C010802020408040C400850AA055254090541A111200A104A0000000908B510",
INIT_03 => X"0C1101100C00004401060A0010041028021560A0218808002440840008880550",
INIT_04 => X"8840C2802205140048281202180804040960986850688C99444090C10A124A69",
INIT_05 => X"910A21220A880010214000010340086856B141252252142242A068B090106372",
INIT_06 => X"4007A400E8A40086213090040001520500204088012121026050A54CE2154840",
INIT_07 => X"0204022420000004601120108108055200022025A83AA3008882004A001542CA",
INIT_08 => X"091C154429220A2824642010A010020282843E00000248000021100000884101",
INIT_09 => X"80442C1411D120828A2A116A24632885419244606001110AE11B202046439511",
INIT_0A => X"644022201204145003031012D40D718241108815384200904160AE42CE2818E2",
INIT_0B => X"1BF047118108829501009202A5A20068C003211551163A00E522B3000562082D",
INIT_0C => X"90D0490D2C90D0C90D2C90D0C90D2490D04486124868294032384890B8985534",
INIT_0D => X"184014960000008402028041005232001715A040820B11A401E2443243450D04",
INIT_0E => X"9306260000554015520481040100004504A08110000820440001009134000004",
INIT_0F => X"02000000001014000028052000400028040050052000400028040200501C8D38",
INIT_10 => X"4002000000000068005005200040002804002805200040002804000E00001000",
INIT_11 => X"0028400010008000000000102800009800601000040000000011820002140102",
INIT_12 => X"4022010110000000D00008310000801080102000A00004000000000009020000",
INIT_13 => X"00001A00C0082400000006802500008000000000080048000060041200000003",
INIT_14 => X"A000005400080600000000000850000014200411000000000010024440202200",
INIT_15 => X"0000000008840600002080200000000000021800000013000040000000000020",
INIT_16 => X"40902449022A800800002208090684819402120AA8001C800000000000100014",
INIT_17 => X"1902409024090240906419064190641902409024090240906419064190641902",
INIT_18 => X"9044190440900409004090041904419044190440900409004090641906419064",
INIT_19 => X"7D402A2953F81F81F83F03F03F04190441904419044090040900409004190441",
INIT_1A => X"4104104104104104609D21808205965965D65801004E35C300C2D50A22B1C50C",
INIT_1B => X"128944A25128944A25128944A250410410410410410410410410410410410410",
INIT_1C => X"FFFFFFFFE3F00944A25128944A25128944A25128944A25128944A25128944A25",
INIT_1D => X"100055400000000000000000000000000000000000000000000001E1F007FFFF",
INIT_1E => X"400FF843DF45FFAEBDF55082A82155082AAAA10F7FFEAB455500175FF5D2A800",
INIT_1F => X"ABEF082ABDF455D7BD5545F7D5574BAFFD16AAAAA28428ABA000428AAA5D7FD7",
INIT_20 => X"EAB455D7BEAABA5D2A97545552E975FFFFD168AAA5D7BE8BFF5D557FFEFFFD16",
INIT_21 => X"A955555555555FFA2AE820BAFFFFEAABA5555554BA5D0417545F7D56AAAAAAFB",
INIT_22 => X"002AA00AAAEBDFFF08042AABA087BD54BA08043DEAAFF843FF5508517FF55552",
INIT_23 => X"02A82010AAD1401FF002EBFF45A2FBFDFEF00042AA00AAFBEAB5500003FF5500",
INIT_24 => X"0000000BA0004155550004154105D556AA00A2FBEAABA085542145082A800BA0",
INIT_25 => X"D5500155FF552A87410007145400000000000000000000000000000000000000",
INIT_26 => X"9208002FABA4171D5400FF8A38F45F7AABA57D0000855FD1C2AAFA00EBA5E8B7",
INIT_27 => X"A92555178FD7BFD5FDFFA0020BFF78417BD5545F7F1554AAF7D16DABABFF57DE",
INIT_28 => X"756DFFDF6DAAAAAF1EFB6D417BEFA901C2E97F40552E975EFEBDF68ABA557BEA",
INIT_29 => X"2DB7DA3FBD21C7492E9256D555B555C7A2ABC20AAE3AABAE38005B574AA49041",
INIT_2A => X"5EDB7D1E803AF6D400028E02AB8A3A012540E2AABABC75D043A00003FE10E380",
INIT_2B => X"0EB8B7D0AAA800AA147085000FFDA001C7B47BFABC7BFFF7AB4714042AA38BEF",
INIT_2C => X"000000000000000000000000821E8A10568005A1041055716DA38B6FBEFFEF1C",
INIT_2D => X"5D2EBDE00AAC16ABEF5500155EF552A954000855544000000000000000000000",
INIT_2E => X"AF7D57DE0AFAD1EBEB400043DEAA085555400FFAAAAB55F7AEA8BF77004147EF",
INIT_2F => X"EFAAFBEABAF557FEA8515951E8B4D83D1EBDFF082CBDFEF005756145FFD5574A",
INIT_30 => X"E005951550100004155EFF7FFFDE08AA557FFFF083FFCEB95104210405D2E955",
INIT_31 => X"00AA002A3FE18AE803CBE7A3C014351082E951FF5D7FD6145AAAA820A2AAAD29",
INIT_32 => X"EAD45550028ABAFFD17FFED01001FFEF5542ABEB2AA848AAA2552EA8ABA75514",
INIT_33 => X"57FEBAF3F95EEE95C00B7CF12AAA800BA551417105FFFFC21555556EAB4CD6D5",
INIT_34 => X"00000000000000000000000000000000000000000187782001FF0812000A255D",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0400000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(2),        -- Port A data input
DOA(0)   => data_read_a_hi_256(2),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(2),        -- Port B data input
DOB(0)   => data_read_b_hi_256(2),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_3_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"210C00A20020000108430020001600B8156021104940741B3530400E02B92202",
INIT_01 => X"A00C9BC058B00968240402C992000B61404040028804A0080A000D16A8990A08",
INIT_02 => X"4809A902031800444445089866E331352180D468B8200E600C0081110B80ACD0",
INIT_03 => X"6D0A601008000142B1A30A040AC68428320006010A80881068A80D401C846330",
INIT_04 => X"482218076809C03B24841CD92CDD5A4402091278072948042640102107102D04",
INIT_05 => X"0B063006A6402109000104E40B04644B32A86D20014A0D204063296082000E34",
INIT_06 => X"01072010703402800606D0102800CAB31434442810B4858060D0500008C52828",
INIT_07 => X"8C00222420A14204E01C581091020CC8000E3226413990008D80001A00CCC4AA",
INIT_08 => X"0874732009120665255420184000220002843E14294258E805E0116002D95101",
INIT_09 => X"BA546AC411102029A61C974014EDBA1320B1046100C0B4034928002002211145",
INIT_0A => X"1052088250A1CC2041051913208CE802438000082040008000F399406BC07998",
INIT_0B => X"19E416590908884D00020242A500090801806801041358222302084204460020",
INIT_0C => X"1019010190101B0101B01019010198101B20805C080C880080506990125E0514",
INIT_0D => X"03400040A101C05C0088242D0000320013339310018011A044414400400101B0",
INIT_0E => X"6514CA601CCCC8B33204C0401104244000018380818040A07060090000280009",
INIT_0F => X"0000000000020000006000000000020000011000000000020000010072CC9251",
INIT_10 => X"0000000000010000014000000000020000013800000000020000010700000000",
INIT_11 => X"002C000000000000000000010000001A00000000000000000040000002440000",
INIT_12 => X"00B2000000000010002049910000011000500000000000000000008000000000",
INIT_13 => X"00020005500000000000800133000000000000000010000000C0000000000040",
INIT_14 => X"0000005300000000000000001000000110600000000000000000401540000000",
INIT_15 => X"8000000008200620000000000000000000400000000107000000000000000004",
INIT_16 => X"0280C0280C0205104100000A8D06C404440230B9980210020040000010010003",
INIT_17 => X"280C0280C0280C0280803808038080380803808038080380C0280C0280C0280C",
INIT_18 => X"80E0200C0280E0200C0280E030080380A030080380A030080380C0280C0280C0",
INIT_19 => X"291008A004D54AAB556AA9556AA830080380A030080380A030080380A0200C02",
INIT_1A => X"4904104104104104A20E85800004924924054C0F031E31C190A285040164C586",
INIT_1B => X"1A8D46A753A9D4EA753A9D4EA752492492492492492492492492492492492492",
INIT_1C => X"FFFFFFFEB6FECD46A351A8D46A351A8D46A351A8D46A351A8D46A351A8D46A35",
INIT_1D => X"00AA8400000000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"B455500175FF5D2AA8A10005540155087BEABFF552ABDF45A2D16AAAAF7D5400",
INIT_1F => X"201000556AB55552ABDE00AAD140010F7D17FF45A2AA82155082AAAA10F7FFEA",
INIT_20 => X"42155557FEAA10007FEAABA000428AAA557FD7400FF843DE00FFAEBFF55082A8",
INIT_21 => X"AA8A105D7BD5545F7D5574BAFF802AA00A2D168ABA085568BEFFFAE820000855",
INIT_22 => X"557FFEFF7D56ABEF557BD74BAFF8402145A2AEBFFEF552EAAABA5D0028BEF082",
INIT_23 => X"5043DEAAAAAA95410F7803FFFF55556AAAA552A975FFFFD16AAAA5D7BC01EF5D",
INIT_24 => X"0000000105D0417545F7D56AAAAAAFBEAB455D7BEAABA5D2A974005D55574005",
INIT_25 => X"5B6DF6FABAFFD547010AA8407400000000000000000000000000000000000000",
INIT_26 => X"6D1C2AAFA28EBF5E8B7D5500155FF552AAF0100071455451C75EABC74174BAF5",
INIT_27 => X"F45F7AABAF7D00009543D1C556AB6D4124BAE10BED542010FFD57AF55AAF5D75",
INIT_28 => X"ABFFEBA0870281C5F4716D5D7FEDA3A0955FF48208002FABA4171D5400FF8A38",
INIT_29 => X"B8EBA15203FFFF002AAFA384171D5545F7D0154AAF7D16DABABFF57DE92005F6",
INIT_2A => X"F68ABA417BC01D7555178FD7BFD5FDF571575D24BA438E021D5B6A4BAFFF5D2E",
INIT_2B => X"24BFE005D5B52428410E3AE92E3A490410EB843ABD71551FFE02552A975FFEBD",
INIT_2C => X"0000000000000000000000003849041756DFFDF6DAAAAAF1EFB6D417BEFBD71C",
INIT_2D => X"5D556AB45081028B55FFFFFFEBAFFD557400A280144000000000000000000000",
INIT_2E => X"0FFD56ABF5AAD15455F5D2EBDEAAA2D16ABEF5500175EF552ABDE00085554545",
INIT_2F => X"AA085555400FFAAAAB14F7AE28BF77004146BA557DEABEF00002BE10FFD54000",
INIT_30 => X"E0AF2D1EAEBA007FEABEFAA84174BA557FD55EF5D3BFEEB35055DEE1000043DE",
INIT_31 => X"0155FFAA28BF7592EABE0A0804ABFFB082EBDEAA005556145FFD5574AAF7D47D",
INIT_32 => X"EB8105D2E955EFAAFBE8AAA547FE21550853E8B4FABD5EBFF75D55420AA82AA8",
INIT_33 => X"57FFFF087FFCEF90104B780A557FC20AA082AAAE10AA8000000A2AC2ABFD2151",
INIT_34 => X"00000000000000000000000000000000000000000AA0004155EFF7FFFDE08AA5",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(3),        -- Port A data input
DOA(0)   => data_read_a_hi_256(3),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(3),        -- Port B data input
DOB(0)   => data_read_b_hi_256(3),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_4_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10804002061080A284201081034809800A002303500078B3432C82904204002",
INIT_01 => X"810398000008004C0420050E12100368403008418984014902030806A0910204",
INIT_02 => X"480108A000000000446448E01E80F00A41043118680402000800000009882390",
INIT_03 => X"065040108C0000408406080002101020260012E03000000030808902088000F0",
INIT_04 => X"9100EB8368155C1AE0B01CD60433B944028A90385AC0D438E02010E81C32E801",
INIT_05 => X"B81E4166DE080029204044C401041C4CF01C489433483C8042EAC190100074C4",
INIT_06 => X"400F0400688002A22010D4342045C50F0004028993B3A5260041E4500EB4C0E2",
INIT_07 => X"000000243020008461000812810003C300060064012E00048C82005800BC2888",
INIT_08 => X"08CC8F0109064220240410008000002202043E44001048000020114000881000",
INIT_09 => X"F0DC1EB5131020C7BE7D172251E53E80E891E5016041B4083945202002419104",
INIT_0A => X"7D6025AC2A0982500302003200872003FB108808280200204400786612CE2B08",
INIT_0B => X"11D0025980480A458100930201820964408268101000F022D8083B4044A0002C",
INIT_0C => X"90C3490C1490C3490C1490C1490C3490C104869A48618800B66305989ABA0434",
INIT_0D => X"220000000500021002100088004010001370F030808110204581043243050C54",
INIT_0E => X"06100C40903C1C30F20025440102200541204090600830045825050034010000",
INIT_0F => X"000000000012000000BC04000000020004018C040000000200040000721CD861",
INIT_10 => X"000000000001002001A40400000002000401DC04000000020004014D44001000",
INIT_11 => X"0065040010000000000000110000007600200000000000000050000005D40002",
INIT_12 => X"00DE00001000001040004A3B0000180088500000200000000000008000020000",
INIT_13 => X"0002080760000400000082024300008000000000081006000170000200000041",
INIT_14 => X"180002B200000200000000001806000192000010000000000010401F80000200",
INIT_15 => X"0814000114A00200000000200000000000401006000085C00040000000000024",
INIT_16 => X"40102459044481081044880A0986D4C1560636C7840A61803000820012113042",
INIT_17 => X"1900411064090041102409044110240900401064190040106409004110640904",
INIT_18 => X"9064090240100411044090241902401044110041902409064110241904401024",
INIT_19 => X"04048028064B261934D964C3269C090641100401044090641902401044010041",
INIT_1A => X"AA8A28A28A28A28A74C132343334514513028A2818E01F81400050E130106345",
INIT_1B => X"8341A0D46A351A8D46A351A8D46AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA",
INIT_1C => X"FFFFFFFE58C001A0D068341A0D068341A0D068341A0D068341A0D068341A0D06",
INIT_1D => X"10550015400000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"F45A2D16AAAAF7D568A00AA8400000AAFFC21FFF7D542000FFAE821FF552EAAA",
INIT_1F => X"0000AAAE820BA550015400087FD74BAFFD540000F7D155555087BEABFF552ABD",
INIT_20 => X"A8AAAF78015545FFD555555082AAAA10F7FFEAB455500175FF5D2AAAA1000554",
INIT_21 => X"56AB45552ABDE00AAD140010F7D17FF45A2FBC2000A2FFC21555551554005D2E",
INIT_22 => X"AEBFF55082E82145A280001EFF78402145A2AE801555D2E95555552E97410005",
INIT_23 => X"D517DF45557BD5410F7D555545F7AA97410000428AAA557FD5400FF843DE00FF",
INIT_24 => X"0000000AA085568BEFFFAE82000085542155557FEAA10007FEABEFAAD1400AA5",
INIT_25 => X"8EBAA801EF4920AFA10490A17000000000000000000000000000000000000000",
INIT_26 => X"451C75EABEF4124BAF55B6DF6FABAFFD56F010AA8407428A2F1C01FFF7D14202",
INIT_27 => X"5FF552AAFA10007155428A2AE850925D0010400087FD24AAE3DF47010E38E051",
INIT_28 => X"01555D51524004920ADA82EB8A12555EBFB4717D1C2AAFA28EBF5E8B7D550015",
INIT_29 => X"92555492A850381C5F6AB6D4124BAE10BED542010FFD57AF55AAF5D7410A2FBC",
INIT_2A => X"1D5400FF8A38E00F7AABAF7D0000955FDB684051D7F7840517DA2A4871554124",
INIT_2B => X"55D75EFBED5400825D557FF55007BD7410EBDB5017DE38E8708008002FAAA417",
INIT_2C => X"00000000000000000000000082005F6ABFFEBA0870281C5F4716D5D7FEDB7D09",
INIT_2D => X"AAD1401FFFFD5420BAA2AA821FF08043DE10002A964000000000000000000000",
INIT_2E => X"AA2FBD7410A2AE965555D556ABEF080028B55FFFFFDEBAFFD57FE00A280144BA",
INIT_2F => X"AAA2D16ABEF5500175EF552ABDE000855544AAAA82174105D0402000087FC00B",
INIT_30 => X"BF5AAD154400AAFBC015555554001008003FE00AAEA81154AAFFD65FF5D2EBDE",
INIT_31 => X"75EFA2AA155550004021E5582A964BE557FEABEF00002BE10FFD540000FFD56A",
INIT_32 => X"9661000043DEAA085555400FFAAAAA10F7AC28BF558001454DF78017555F7801",
INIT_33 => X"FD55EF5D7BFEEF35055487EFF7D1400105D517FF55087FD7410A2FBC01E7F2AE",
INIT_34 => X"0000000000000000000000000000000000000000010007FEABEFAA84174BA557",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0400000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(4),        -- Port A data input
DOA(0)   => data_read_a_hi_256(4),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(4),        -- Port B data input
DOB(0)   => data_read_b_hi_256(4),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_5_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50DF0A0791B3FC1694378283C81FD996A091A32152007AB36B20E03C040C006",
INIT_01 => X"081FBDC49830884C5C6A60000C34C24841280A00084000C8C212892EEA953231",
INIT_02 => X"C809AD5CB118E640A4F008F8011FF0002080000082CCC66609DB7DDDCB1F2036",
INIT_03 => X"25080626BE4C904210831C80084204720B20048A88800000B8E0F8102885500E",
INIT_04 => X"4005122024899100064520C01444429C7804103C0416C007198A3916E0551A04",
INIT_05 => X"46E1829941C9000944C8C022898FE2F20D7D7A104CB5C208E51417C054848912",
INIT_06 => X"CA075CA0E63342991612DF9A8205C0A0B030B20B10480900886E220801073711",
INIT_07 => X"8C732074B68D1A34E3180717FFD13FC72691924098712CE481FDC241D43C1ACD",
INIT_08 => X"16053F180A1286A4E51BD18840C320000075FE91A24458BA4DE0D57992D9BE58",
INIT_09 => X"0A4D8105BF3472304100930258E510601EDE1D8524309285FD416CB402259504",
INIT_0A => X"3110AC0D11C901B2112109204C28B67061E8928920CAD3CFC0140079065A4A65",
INIT_0B => X"C3404959321C284D356A964F8125CD7AC8632614005DFBAACFBC800024091128",
INIT_0C => X"380D6380B6380F638096380F6380B6380D51C04B1C07AD10C14020D233127AD5",
INIT_0D => X"992940513052F4CA8A0A0664A5023CA8470FF000908C383755AF1604E0538096",
INIT_0E => X"200040194FFC044FFA4B08BC85282C91F028D094284A34054A25508605135C01",
INIT_0F => X"BA0C2038ABACBC7C7806F94FF87C002F83F106F94FF87C002F83F2000A04C200",
INIT_10 => X"8D9A70380230F2DFC106F86FF87C002F83F106F86FF87C002F83F3601BFFEBC2",
INIT_11 => X"1F401BFFE7C69E01804E1E6EABE3F040FFD7C7C4BC0E008C7C2FE58FC0A9FFF5",
INIT_12 => X"F8BFDFC8C8120C4DBC802208B2EB2AE777ADFE6F0A47CC0600C2683E0FF8AE3F",
INIT_13 => X"4189B7C56DF47186104C6DE7037FFF00FC0000FC07EE4E7A7076FE28C3082636",
INIT_14 => X"B9E9F272FFFC181C0C2038A7C6DE7A7D909FBFA4070380131CAFB257FBD93902",
INIT_15 => X"2B34E9F56DFBEB1B7F2300C4A80092E0FC1FCE667A7C877FFE828F0080AE1DDA",
INIT_16 => X"51142511405EA00A1344612A898494801602081F87204A9452217159891640D4",
INIT_17 => X"0942511425014450940519425114650140519405194650146511405194050946",
INIT_18 => X"1465114250146501465194051944509445094051146501465014251140509445",
INIT_19 => X"7ED430A983124B2DA6924965B4D5014650142511425094450940519405094450",
INIT_1A => X"EFBEFBEFBEFBEFBE5FDFF3F7F773CF3CF7D796ED39FDEE76DFFCE9F84801B6DB",
INIT_1B => X"BDDEEF77BBDDEEF77BBDDEEF77BBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFB",
INIT_1C => X"FFFFFFFE433B5EEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77B",
INIT_1D => X"AAFFFBFFE00000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"000FFAE821FF552E820105500155555D2AA8A00AA843FFFFF78002155AAAE974",
INIT_1F => X"0000FFAE80000AAAE974BAFFAEAAB45AAAEBDEAAA2FFEAA00AAFFC21FFF7D542",
INIT_20 => X"7FE000055574BA557FFFF55087BEABFF552ABDF45A2D16AAAAF7D56AA00AA840",
INIT_21 => X"E820BA550015400087FD74BAFFD540000F780155555D7BE8B45085168BFFA2D1",
INIT_22 => X"2AAAA10005140145FFFBC01EFAAFFD75FF002E97555A2AABDEAAAAAAAAA00AAA",
INIT_23 => X"A84174BA5D043FF45AAAA974AAF7AEBFF55082AAAA10F7FFEAB455500175FF5D",
INIT_24 => X"000000000A2FFC21555551554005D2EA8AAAF78015545FFD555410552EA8BEFA",
INIT_25 => X"FFF8E0217DBEA4954AAE3FBFDE00000000000000000000000000000000000000",
INIT_26 => X"28A2F1C01D7F7D142028EBAA801EF492087A10490A171455D2EADA28B6803FFF",
INIT_27 => X"ABAFFD56FA10AA8417428E3AE87010A2A4974AAE3AEAFB6DAAA4BDEAAA2F1EDA",
INIT_28 => X"8B6D14516DBD7BEDB7DE381451554AA497FFFF451C75EABEF4124BAF55B6DF6F",
INIT_29 => X"BDEAAAAA0AFA28A2A4850925D0010400087FD24AAE3DF47010E38E0516D5D7BE",
INIT_2A => X"5E8B7D5500155FF552AAFA10007155545F7F1C21D7AAF1D55FF082A9057DA2AA",
INIT_2B => X"FB470384124ADBFFBE84174AA55043FF6DBEAE950AAEB8ABDF7D1C2AAFA28EBF",
INIT_2C => X"00000000000000000000000010A2FBC01555D51524004920ADA82EB8A12410EB",
INIT_2D => X"552EBFEBAF7843DFEFF7AE801EFF780174AAAAFBFEE000000000000000000000",
INIT_2E => X"FA2803FEBAAAD17CEAAAAD140155FFD5420BAA2AA821FF080415410002A96555",
INIT_2F => X"EF080028B55FFFFFDEBAFFD57FE00A280144AAA2AA97400A280174AAA2AEBDFE",
INIT_30 => X"410A2AE965FF557FE8BFF55557FF55FFFBFFEAA5D51554AA087BFEF555D556AB",
INIT_31 => X"55FF0004821FFAAAEBDEAAAA843CEAAAA80174105D0402000087FC00BAA2FBD7",
INIT_32 => X"BEFFF5D2EBDEAAA2D16ABEF5500175EF552ABDE00005554545F7D140145A2D55",
INIT_33 => X"03FE00AAAA81114AAFFD64BA00043FFFFFF80174AA55043DFFFFFAE974BAA2AE",
INIT_34 => X"0000000000000000000000000000000000000000000AAFBC0155555540010080",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"1800000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(5),        -- Port A data input
DOA(0)   => data_read_a_hi_256(5),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(5),        -- Port B data input
DOB(0)   => data_read_b_hi_256(5),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_6_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10844B0061A258A2840112C03002C18000402322520070B303301C0381A0086",
INIT_01 => X"0600404820094048008100000042026041000000090800090210080008510204",
INIT_02 => X"080108220C1000004440080000C008010000000001203240080080000988A050",
INIT_03 => X"040000000823404000020A600000002983800584488000103080040C08C00000",
INIT_04 => X"00101610A029B08400044800000000040000102A040810040400100500101800",
INIT_05 => X"05000000800C8300306420002900404400820000000A00804004084001200A00",
INIT_06 => X"64472644640C00808C10D00401823F0020204209101001002650020001052800",
INIT_07 => X"080000242000000461100050818080380900224000200008818028804883E10A",
INIT_08 => X"01FE80E0090242602C0020608000000000043E00000048800021140000881106",
INIT_09 => X"12447E041B102020208000424029006FE0B085013204D0200101006862119140",
INIT_0A => X"4D540B0D916BBE39059191200000200441040108000020006FC5FA6000816908",
INIT_0B => X"8BF05D11A20808454010834225A28962E40AA05510180022FFA6A8800402A06D",
INIT_0C => X"16C1416C5416C5416C3416C3416C7416C500B60A0B60AD04EB4104C093904535",
INIT_0D => X"59802817888180E80112A1660050900003400430CB4911B445A105B05B016C14",
INIT_0E => X"000000062003C90000442006439324280034E85A742D1A16CD2DA30046848048",
INIT_0F => X"00000000000157000600000000000028000C00000000000028000CE800048000",
INIT_10 => X"00000000000000483C00000000000028000C00000000000028000D1080000000",
INIT_11 => X"00108000000000000000000078000A00000000000000000000019A0030000000",
INIT_12 => X"4604000000000000934909080014000000000000000000000000000009005180",
INIT_13 => X"00001230B00000000000049B3C000000000000000001FA000C98000000000002",
INIT_14 => X"E8000E05000000000000000001720002A56000000000000000000FC080000000",
INIT_15 => X"0840000B000404A000000000000000000002099A0003B0000000000000000001",
INIT_16 => X"69DA5685A146D19D084488080904C0A1172240C0781400C81908000205208614",
INIT_17 => X"85A1695A769DA3685A169DA768DA1685A169DA7685A1685A769DA7685A168DA7",
INIT_18 => X"5A368DA1685A769DA168DA3695A569DA3685A169DA5695A368DA1695A569DA36",
INIT_19 => X"7F10800846638C31C71C718638E685A769DA5685A3685A569DA7685A168DA769",
INIT_1A => X"E38E38E38E38E38E76DDB3B7B377DF7DF7D7DE2F39FE3FC3D3EA55FF37F5F7CF",
INIT_1B => X"9FCFE7F3F9FCFE7F3F9FCFE7F3F8E38E38E38E38E38E38E38E38E38E38E38E38",
INIT_1C => X"FFFFFFFF61AC8FE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F",
INIT_1D => X"EFAAAABFE00000000000000000000000000000000000000000000181F007FFFF",
INIT_1E => X"FFFF78002155AAAE974AAFFFBFFE10F7FBE8BEF552E95555552EAABEF082E975",
INIT_1F => X"5410A2AAAAA10087FC01EF552EAAB45F7AE821550851555555D2AA8A00AA843F",
INIT_20 => X"2ABEFA2AEBDFFF552AAAA00AAFFC21FFF7D542000FFAE821FF552E8001055001",
INIT_21 => X"E80000AAAE974BAFFAEAAB45AAAEBDEAAA2FFEAB45552E800AA555568A105D00",
INIT_22 => X"D56AA00AA8400000007BC21FFAA803FFEF5551420105D5568B45FF8400000FFA",
INIT_23 => X"7FBC2155007FC20BAA2D5575FF087FFFF55087BEABFF552ABDF45A2D16AAAAF7",
INIT_24 => X"0000001555D7BE8B45085168BFFA2D17FE000055574BA557FFFE10F7AAA8A00F",
INIT_25 => X"D4924ADBD70820975FFA2A4BFE00000000000000000000000000000000000000",
INIT_26 => X"455D2EADA28B6803FFFFFF8E0217DBEA4954AAE3FBFDE38F7FFEABFF412A9056",
INIT_27 => X"1EF492087010490A07038B6A0AFA38007BC51EF4920AFB55EBA4851450855555",
INIT_28 => X"5082555F68A3855002FBC7BEA4BFFFF492EADA28A2F1C01D7F7D142028EBAA80",
INIT_29 => X"6DB45E38A07028E3AE87010A2A4974AAE3AEAFB6DAAA4BDEAAA2F1EDB55492A8",
INIT_2A => X"4BAF55B6DF6FABAFFD56FA10AA84174381C7FC01C7B68E3DFC75555400105D51",
INIT_2B => X"7FFFE38F7A0AFA38E3FFC21450071C2092A2D5571FF0851FDF451C75EABEF412",
INIT_2C => X"0000000000000000000000016D5D7BE8B6D14516DBD7BEDB7DE381451554AA49",
INIT_2D => X"F7FBEABEF002E801EF00003FF550800155FFA2803CE000000000000000000000",
INIT_2E => X"5A28417555085154555552EBFEBAF7843DFEFF7AE801EFF780174AAAAFBFEEAA",
INIT_2F => X"55FFD5420BAA2AA821FF080415410002A964AAFF803DEAA087FD55FF00043DF4",
INIT_30 => X"EBAAAD17CF55002E95410557BEAABA55043DF55F7803FFEF002ABEEAAAAD1401",
INIT_31 => X"DF455D51420105D517DF55AAAA964AAA2AA97400A280174AAA2AEBDFEFA2803F",
INIT_32 => X"7CF555D556ABEF080028B55FFFFFDEBAFFD57FE00A280144BA5D7FC2155FFAAB",
INIT_33 => X"BFFEAA5D51554AA087BFEEAAF7803DEAAAAFBC0155085540000A2D5575FF0851",
INIT_34 => X"00000000000000000000000000000000000000001FF557FE8BFF55557FF55FFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"1200000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(6),        -- Port A data input
DOA(0)   => data_read_a_hi_256(6),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(6),        -- Port B data input
DOB(0)   => data_read_b_hi_256(6),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_7_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10844B00482258A2842112C02450418800002300500030B303300C018180002",
INIT_01 => X"0200084020084048040080000201026040000000080000080200090000510204",
INIT_02 => X"4801082048100000444008040080000041000000000222400800000009000010",
INIT_03 => X"0401018108A144D0000208424000002103006480088000003080000408C10000",
INIT_04 => X"0000120022419000000C80000000000400201829040000050001940400301820",
INIT_05 => X"04000000800840092CC080214144004400000000000800065004004020220800",
INIT_06 => X"40870408600000808C10D4500080008020200008001001000240000061052002",
INIT_07 => X"08000024200000046010005281848001494020400031240C8C8238A06A000988",
INIT_08 => X"40050001090242602C0408408000000000243E00000048800020154000881024",
INIT_09 => X"024401041B132820000011424069004000B20403200891420101026A42210440",
INIT_0A => X"013800A0281400300C0010200008B20663970148004424006818026200004800",
INIT_0B => X"01C1103022881845421082C2C0082300401121810012004600001010040028A0",
INIT_0C => X"1200112001120011204112041120411206089010890100408040008012101414",
INIT_0D => X"09146817802988694902A02451109006230006E0808294008C02848148092001",
INIT_0E => X"000000042C00040002000004020020490020401020081004482501010C120948",
INIT_0F => X"0130C807144102420700052000003C00780B00052000003C007808450484C000",
INIT_10 => X"400002C0E00E0D003300052000003C00780B00052000003C0078099080001000",
INIT_11 => X"80908000100000661801E18042100E000060100000B038038380124038000102",
INIT_12 => X"053A010111848322020512000414400000002000A1001058300C0741C0054120",
INIT_13 => X"90644029D008240864231011BF00008000C3C003F00186040EE8041204321188",
INIT_14 => X"18100D770008060130C807182106040375600411004C2600E3400C2740202230",
INIT_15 => X"9094100A8CA406A0002C812240B0201F0380211604037740004010472041E201",
INIT_16 => X"40100401006E8118104428088904C4C414420080049450801000088444300601",
INIT_17 => X"0906409004010040104409024090240906401004010040102409024090240100",
INIT_18 => X"1024090241900401004090240902401004010040902409004010440100409024",
INIT_19 => X"004420A945841040002082080004110240902409004110040902409024110040",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFEDD9EC000000000000000000000000000000000000000000000000000",
INIT_1D => X"BA082AAAA00000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"555552EAABEF082E975EFAAAABFFEF002ABDF555D5157555F7FBC00AAAAD5400",
INIT_1F => X"FEAAAAAABDF55FFFBFDF55555568ABAAAD5401FF5D2AAAA10F7FBE8BEF552E95",
INIT_20 => X"400005D55554105D51401555D2AA8A00AA843FFFFF78002155AAAE974AAFFFBF",
INIT_21 => X"AAAA10087FC01EF552EAAB45F7AE821550851554AAF7FBFFEAA007BFFFEFF7D5",
INIT_22 => X"2E800105500155EF5D2EBFF450000020AA5D7BC0000F7D555545A28000010A2A",
INIT_23 => X"FAAA8A10FFD568ABAA2D56AAAAF7AABFE00AAFFC21FFF7D542000FFAE821FF55",
INIT_24 => X"000000145552E800AA555568A105D002ABEFA2AEBDFFF552AAAABAA2AE95555F",
INIT_25 => X"5E3F5C20BAAAD5420821C2EAAA00000000000000000000000000000000000000",
INIT_26 => X"38F7FFEABFF412A9056D4924ADBD70820975FFA2A4BFFFF1C2EB8F4555555054",
INIT_27 => X"17DBEA4954AAE3FBFDE82B6AEBAF55E3FFFAF55555F6FA92BED5421C75D20AAA",
INIT_28 => X"FE920075FDFD7F7D5400385D51504385D55401455D2EADA28B6803FFFFFF8E02",
INIT_29 => X"5057DB68E02038B6A0AFA38007BC51EF4920AFB55EBA485145085555492F7F5F",
INIT_2A => X"142028EBAA801EF492087010490A071EF4920B8F45140E07082417BC2000EBD5",
INIT_2B => X"2EADA92A2A09257DE3A4AAA10F7D16FAAABED56AE82F780BAE28A2F1C01D7F7D",
INIT_2C => X"00000000000000000000000155492A85082555F68A3855002FBC7BEA4BFFFF49",
INIT_2D => X"552EAAB455D5142155AAD1400AAA2D1420005D2EA9A000000000000000000000",
INIT_2E => X"0F7D1421555D042BAAAF7FBEABEF002E801EF00003FF550800155FFA2803CFFF",
INIT_2F => X"BAF7843DFEFF7AE801EFF780174AAAAFBFEE00F7AAAAB55AAFBEAB555D7BFDE0",
INIT_30 => X"555085154400FFD17FE1000517FF55FFD5420BA5D55400BA555543155552EBFE",
INIT_31 => X"5400087BC0000A2D5421EFF7AE810AAFF803DEAA087FD55FF00043DF45A28417",
INIT_32 => X"2BAAAAAD140155FFD5420BAA2AA821FF080415410002A965FF080428B45552A9",
INIT_33 => X"43DF55F7803FFEF002ABEE00A280001FFA28028A00FFD17DEAAF7D56AA10FF84",
INIT_34 => X"0000000000000000000000000000000000000000155002E95410557BEAABA550",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"01FFFFFFFFE00000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(7),        -- Port A data input
DOA(0)   => data_read_a_hi_256(7),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(7),        -- Port B data input
DOB(0)   => data_read_b_hi_256(7),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_8_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00000648E2840112C00000418000002700500030B3032000000000082",
INIT_01 => X"000009C21838284D1C2160000E12424840000000180800080200000040110204",
INIT_02 => X"080108000090000004400C040080000051000000000002400800000009000010",
INIT_03 => X"00000100043008D0000200024000000003800504488000103080880008800000",
INIT_04 => X"00009410A028A084000440000000000400001022040800150400808500321800",
INIT_05 => X"8500010080048A09302420202804400400800010200A00020204084011014A00",
INIT_06 => X"2447A244608800840490D0040007FE0021204288001000000050024001042800",
INIT_07 => X"4800002420000004201000D281040003182020400031241C0D80004041BFE88A",
INIT_08 => X"4005000108020220240000048000000000043E00000048800000010000881000",
INIT_09 => X"0204010519110020008111020069004008A28501120450220101214122509140",
INIT_0A => X"0528A52291490029019190200008B20E23008028000208804010024000004000",
INIT_0B => X"13C151312A8808454104824001280108A409A044001200020020989000000061",
INIT_0C => X"0000000000000000000000000000000000400020000229508040008012105400",
INIT_0D => X"48022817880508602102A1200810B2020340043248CA00240420000000400040",
INIT_0E => X"4100820020000C0000442142419120000014684A34251A12CD2CA30042840248",
INIT_0F => X"45F3D80000000001020404000783FC0000010404000783FC000000880284C010",
INIT_10 => X"02658FC7E0000000010404000783FC0000010404000783FC000001500000103D",
INIT_11 => X"40500000103961FE78000000000402400020003B43F1F8000000022010800002",
INIT_12 => X"0080001617CD800000080B000804080000020090659833F9F03C000000000000",
INIT_13 => X"B000000400018639EC000000000000FE03FFC00000000600840000C31CF60000",
INIT_14 => X"180204000001E2A3F3D80000000600802000401AA8FC7E00000000100002C2F5",
INIT_15 => X"005404020000104480DC372B47F060000000000600802000017570FF60000000",
INIT_16 => X"28CA328CA34650850A4C000009A494A015624080044440481908000220308640",
INIT_17 => X"8CA328CA328CA328CA3284A1284A1284A1284A1284A1284A328CA328CA328CA3",
INIT_18 => X"CA1284A1284A1284A128CA328CA328CA328CA3284A1284A1284A1284A128CA32",
INIT_19 => X"64108088440000000000000000028CA1284A1284A1284A128CA328CA328CA328",
INIT_1A => X"E79E79E79E79E79EDFC8F33637D6CB6CB2900A282950FAF15E8428917C51E75D",
INIT_1B => X"87D3E1F0F87C3E1F0F87C3E1F0F9E79E79E79E79E79E79E79E79E79E79E79E79",
INIT_1C => X"FFFFFFFECB0593E1F4F87D3E1F4F87D3E1F4F87D3E1F4F87D3E1F4F87D3E1F4F",
INIT_1D => X"10002ABFE00000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"555F7FBC00AAAAD5400BA082AAAA10000000010F7D5421EF007BC01FF5D7FFFE",
INIT_1F => X"FEAA5551554AAFF80021EF002A820BAFF8428A00A2AAAABEF002ABDF555D5157",
INIT_20 => X"E8BEFFFFFEAB55002ABFE10F7FBE8BEF552E95555552EAABEF082E975EFAAAAB",
INIT_21 => X"ABDF55FFFBFDF55555568ABAAAD5401FF5D2AAAB55FFD1400AA5D7FC01EFA2FF",
INIT_22 => X"AE974AAFFFBFFEAA08001555555516ABEFA280020AA5D043DF55557BEAAAAAAA",
INIT_23 => X"8042AB55005140145AAFFE8AAAF7D1401555D2AA8A00AA843FFFFF78002155AA",
INIT_24 => X"0000000AAF7FBFFEAA007BFFFEFF7D5400005D55554105D51400005551421EF0",
INIT_25 => X"71C7FC21EF5D75FFE10142EBAE00000000000000000000000000000000000000",
INIT_26 => X"FF1C2EB8F45555550545E3F5C20BAAAD5420821C2EAAA101C0005000E3D1401D",
INIT_27 => X"BD70820975FFA2A4BFE925D51554AAE384001FF142E800AAFF802AA28AAAEAFB",
INIT_28 => X"7092557BC21D7BEF5EDBC7FFF1EFB6D1420BAE38F7FFEABFF412A9056D4924AD",
INIT_29 => X"3AF55417BEDA82B6AEBAF55E3FFFAF55555F6FA92BED5421C75D20AAB45F7D14",
INIT_2A => X"03FFFFFF8E0217DBEA4954AAE3FBFDEAA1C001056D415F6ABEFA284020824904",
INIT_2B => X"55400385D51401EF00002FB45085F4016DAAF1EDAAAFFFB401455D2EADA28B68",
INIT_2C => X"00000000000000000000000092F7F5FFE920075FDFD7F7D5400385D51504385D",
INIT_2D => X"5D0417410AAD540155557FC01EF5D557DE105D2AA8A000000000000000000000",
INIT_2E => X"AF7842AABAA2AEBDFFF552EAAB455D5142155AAD1400AAA2D1420005D2EA9A10",
INIT_2F => X"EF002E801EF00003FF550800155FFA2803CE105D55574BAA280021EF5D2E820B",
INIT_30 => X"1555D042BB45FFD157410557FC0155F7D57FF55F7D57FFEF550028AAAF7FBEAB",
INIT_31 => X"8BFFAA8000000080428B55087FFFE00F7AAAAB55AAFBEAB555D7BFDE00F7D142",
INIT_32 => X"C2155552EBFEBAF7843DFEFF7AE801EFF780174AAAAFBFEEBA5D04021EF087BE",
INIT_33 => X"5420BA5D55400BA5555430BA5555421EF00043FF45007BC21FFA2D57FEBAF7FB",
INIT_34 => X"0000000000000000000000000000000000000000000FFD17FE1000517FF55FFD",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0800000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(8),        -- Port A data input
DOA(0)   => data_read_a_hi_256(8),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(8),        -- Port B data input
DOB(0)   => data_read_b_hi_256(8),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_9_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00018248A2840112C00002C18000002300500030B3032000000000006",
INIT_01 => X"000008000000004C0020000000100268413C0A61590001D90213C00000110204",
INIT_02 => X"680108200010000054400C040080000041000000010002400800800009082011",
INIT_03 => X"00040100000020D0000200124000000043800504488000103081880008800000",
INIT_04 => X"00001410A00AA084000400000200000400001020040010050020820400101880",
INIT_05 => X"0400040080048A09202420000C00410400000000000800020804004000000800",
INIT_06 => X"24478244640800840410D4144002008020200009301000000140000201042000",
INIT_07 => X"0800002C20000004301000128104000100002040003164040D80000040000888",
INIT_08 => X"40050003080202202400000080000000000C3E00000048800010230000881000",
INIT_09 => X"0024010411110420008010020021004000A204011200500001010000AA10C000",
INIT_0A => X"7945282804010009009090200008B20223800008020000004010024204000440",
INIT_0B => X"114100112208084540008240110001002400A000001000020008288000000420",
INIT_0C => X"010400100001040010000104001000010400080000820800000000801010100A",
INIT_0D => X"08403C16800100640182A0210010921003400412484202200400004004001040",
INIT_0E => X"410082002C000C000240004240932041401468CA34651A32CD28A22002840048",
INIT_0F => X"000000000000144002000420000000280001000420000000280000000284C010",
INIT_10 => X"4000000000000048010005000000002800010005000000002800001000001000",
INIT_11 => X"0010000010000000000000002A00020000201000000000000001820010000002",
INIT_12 => X"40BA00011000000090000B000004000000000000A00000000000000009000020",
INIT_13 => X"00001205D0080400000004803F0000800000000000004C0004E8001200000002",
INIT_14 => X"B000047700000600000000000054000135600011000000000000025740200200",
INIT_15 => X"001400020CA406A0000080200000000000020804000137400040000000000000",
INIT_16 => X"28CA328CA36651951A4CA8000984D4E557220080040440481908000001300614",
INIT_17 => X"84A1284A1284A1284A1284A1284A1284A1284A1284A1284A328CA328CA328CA3",
INIT_18 => X"4A1284A1284A1284A128CA328CA328CA328CA328CA328CA328CA328CA3284A12",
INIT_19 => X"2540A809010000000000000000028CA328CA328CA328CA3284A1284A1284A128",
INIT_1A => X"4534D34D34D34D344A2D840100E4920824055CD13333D2379A2A24018615C38E",
INIT_1B => X"268341A0D068341A0D068341A0D1451451451451451451451451451451451451",
INIT_1C => X"FFFFFFFE6DA90341A4D268341A0D069349A0D069349A0D068341A4D268341A4D",
INIT_1D => X"FFFFD557400000000000000000000000000000000000000000000001FFFFFFFF",
INIT_1E => X"1EF007BC01FF5D7FFFE10002ABFF55F7D168A00552E95555007BFFF55087BE8B",
INIT_1F => X"AA10F7FBC0145F7AE801EFF7FBFFF455D7BC0155F7D557410000000010F7D542",
INIT_20 => X"BDE00AA803FFEF5D55421EF002ABDF555D5157555F7FBC00AAAAD5400BA082AA",
INIT_21 => X"1554AAFF80021EF002A820BAFF8428A00A2AAAAAAAF7D17DE00FFFBD5555A2AA",
INIT_22 => X"2E975EFAAAABFFEF002A954BA5551421EF552E954105D00021455555420AA555",
INIT_23 => X"7D5575EFA2FFD75455D7BE8A005D5557410F7FBE8BEF552E95555552EAABEF08",
INIT_24 => X"000000155FFD1400AA5D7FC01EFA2FFE8BEFFFFFEAB55002ABFE10080028BFFF",
INIT_25 => X"D1C71F8F7D147BEFBEFEBD152400000000000000000000000000000000000000",
INIT_26 => X"101C0005000E3D1401D71C7FC21EF5D75FFE10142EBAF7DE3D16DA0041209056",
INIT_27 => X"0BAAAD5420821C2EAAA10E3FFC0145F7A0801FFEBFBF8F6D417BC716DEBD1524",
INIT_28 => X"DE28F7F5D0545B6AAB8E38B68A3AFFF5551471FF1C2EB8F45555550545E3F5C2",
INIT_29 => X"021455D5B470925D51554AAE384001FF142E800AAFF802AA28AAAEAFABAE3D17",
INIT_2A => X"A9056D4924ADBD70820975FFA2A4BFFFF082E974BA4155401C7552097428550E",
INIT_2B => X"20BAE0008002ABFFF7DB505FFAAFBD7555417FEFA00495B52438F7FFEABFF412",
INIT_2C => X"00000000000000000000000145F7D147092557BC21D7BEF5EDBC7FFF1EFB6D14",
INIT_2D => X"AAD17DE100804001EF55516ABFF557BFDFEFA2D5400000000000000000000000",
INIT_2E => X"F007FD55FFA2D5400105D0417410AAD540155557FC01EF5D557DE105D2AA8BEF",
INIT_2F => X"455D5142155AAD1400AAA2D1420005D2EA9A00A2FBC0145FF84001EFA2FFEABF",
INIT_30 => X"ABAA2AEBDEAAAAD17DEBAFFD142155FFAAAAABAFFAAAABFF5551555FF552EAAB",
INIT_31 => X"01555D00154AA552E801455D7BD54105D55574BAA280021EF5D2E820BAF7842A",
INIT_32 => X"C00AAF7FBEABEF002E801EF00003FF550800155FFA2803CFFF002E954BA00514",
INIT_33 => X"57FF55F7D57FFEF550028A10000428BEFF7FFC01FFA2FFD5545007BFDE10087F",
INIT_34 => X"0000000000000000000000000000000000000000145FFD157410557FC0155F7D",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"1000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(9),        -- Port A data input
DOA(0)   => data_read_a_hi_256(9),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(9),        -- Port B data input
DOB(0)   => data_read_b_hi_256(9),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_10_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000B0001800002840002C0000281800020030000000033122000400992006",
INIT_01 => X"A140098018300848180060000C00424040000000080000080200000000110200",
INIT_02 => X"0801080200100000046558000080000041000000002402400800000009008010",
INIT_03 => X"0001000084000040842242000210810803006400088000003080054288C10000",
INIT_04 => X"0000100022008000000C08000800000400A83A2044200C840000000400001820",
INIT_05 => X"0400000080000000248080210044000402000025000800000004203010100800",
INIT_06 => X"00078000600000040410D4102850008024240001981024A82000010461052000",
INIT_07 => X"0800002430204084281000128100000300002040003124040D80204040000888",
INIT_08 => X"0005000108020220240030008000000000043E0408104C800000010000881100",
INIT_09 => X"0004010511100020200000400021004008808060400111080000200002008400",
INIT_0A => X"0000000000010000060210200008B20223048808000200000010024000000000",
INIT_0B => X"03C0411009808245010002000028000080002105010000000020A34249020801",
INIT_0C => X"8004480044800048000480044800448000440002400221008840009012104400",
INIT_0D => X"0000540100000020088000000100100013000400000800040062400200440004",
INIT_0E => X"4100820020000400020000400200204900800000000000000000000100120800",
INIT_0F => X"0000000000101400020401000000002804010401000000002804000000048010",
INIT_10 => X"0000000000000068010400200000002804010400200000002804005000000000",
INIT_11 => X"0050000000000000000000102800024000400000000000000011820010800100",
INIT_12 => X"4000010000000000D00000080004080000002000000000000000000009020000",
INIT_13 => X"00001A000000200000000681000000000000000008004A000400040000000003",
INIT_14 => X"A800040000080000000000000852000020000400000000000010024000002000",
INIT_15 => X"0000000200000000002000000000000000021802000020000000000000000020",
INIT_16 => X"00000040002800100004200009048005C0000080000400000000000000200654",
INIT_17 => X"0802008020080200802008020080200802008020080200800000000000000000",
INIT_18 => X"0000000000000000000080200802008020080200802008020080200802008020",
INIT_19 => X"2054282101000000000000000000000000000000000000000000000000000000",
INIT_1A => X"A28A28A28A28A28A355950666151451453D51A242A503F834E5C49851D243555",
INIT_1B => X"994CA6532994CA6532994CA65328A28A28A28A28A28A28A28A28A28A28A28A28",
INIT_1C => X"FFFFFFFE8E31DCAE532994CA6532995CAE572B94CA6532994CA6572B95CAE532",
INIT_1D => X"AAFFFBC2000000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"555007BFFF55087BE8BFFFFD557400FF842ABEFA2AAA8B5500003DF55F7D568A",
INIT_1F => X"FE0008556ABFFA2D16AB550000021FFF7D17FFEF08042AB55F7D168A00552E95",
INIT_20 => X"3FF55A2D557400557BC2010000000010F7D5421EF007BC01FF5D7FFFE10002AB",
INIT_21 => X"BC0145F7AE801EFF7FBFFF455D7BC0155F7D557545FFAE820AA007BFDFEF5500",
INIT_22 => X"D5400BA082AAAA00FFAE820AAAAAABDFEFF78028BEF005140145A2842AA10F7F",
INIT_23 => X"AD56AB55A2D157400552EBFFEF5D7BD75EF002ABDF555D5157555F7FBC00AAAA",
INIT_24 => X"0000000AAF7D17DE00FFFBD5555A2AABDE00AA803FFEF5D55420BA08557FEBAA",
INIT_25 => X"51C0E3AF55F7DF68ABAE3F1C0000000000000000000000000000000000000000",
INIT_26 => X"7DE3D16DA0041209056D1C71F8F7D147BEFBEFEBD152400F7842FBD7B6AAAAB5",
INIT_27 => X"1EF5D75FFE10142EBAE0008556FBD7B6DB6AB7D1C0A001D7FFD178FC71C0E28B",
INIT_28 => X"2092147BFAFEF49043AF45A2DF504285D71C00101C0005000E3D1401D71C7FC2",
INIT_29 => X"4017DA28428A10E3FFC0145F7A0801FFEBFBF8F6D417BC716DEBD15256DF7AA8",
INIT_2A => X"550545E3F5C20BAAAD5420821C2EAAA00E3AA82092A2AABAFD7EB8A2ABC70855",
INIT_2B => X"51470821C557AE92A2DF6AB7DA2DF50410412ABDFC75D7BD55FF1C2EB8F45555",
INIT_2C => X"000000000000000000000000BAE3D17DE28F7F5D0545B6AAB8E38B68A3AFFF55",
INIT_2D => X"FF803DF45FFAEA8B555D2EAAB45F7FBE8ABAAAD5400000000000000000000000",
INIT_2E => X"5FFD168B55552AA8BEFAAD17DE100804001EF55516ABFF557BFDFEFA2D540010",
INIT_2F => X"10AAD540155557FC01EF5D557DE105D2AA8A0008557FF45FFFFE8BEF5D2E8015",
INIT_30 => X"5FFA2D5401FFF7AA800105D7FE8BEF08002AB45AAFFC00AA5D51400105D04174",
INIT_31 => X"AB55AAAEAAB450055421FFAA8428A00A2FBC0145FF84001EFA2FFEABFF007FD5",
INIT_32 => X"D55FF552EAAB455D5142155AAD1400AAA2D1420005D2EA9A10A2AA82010AAAEA",
INIT_33 => X"AAAABAFFAAAABFF555155400555568A10AAFBEABEFA2FFC0010082ABFF55557B",
INIT_34 => X"00000000000000000000000000000000000000000AAAAD17DEBAFFD142155FFA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"11FFFFFFFFE00000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(10),        -- Port A data input
DOA(0)   => data_read_a_hi_256(10),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(10),        -- Port B data input
DOB(0)   => data_read_b_hi_256(10),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_11_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10180B05A0010402840602C2D001019000000300000000330A20080EC180002",
INIT_01 => X"AB400984B83008481800E0000C26426040000000080000088200000802112220",
INIT_02 => X"8801081438106400A4F55800008000004100000040CCE24208005000C9060032",
INIT_03 => X"000406A492E6E440842254D002108153422004800880000030C0315688C00006",
INIT_04 => X"00001201200090001205400000000094108C322644240C840008030440111800",
INIT_05 => X"444000888008010028404002A002009402400025080880000C04223000170900",
INIT_06 => X"40871408620B00801410D94CAAD0018024242008A8102CA88A44010401042200",
INIT_07 => X"08320054B624408428100094ADD080011721A04000316C140CA1A8A1F9001889",
INIT_08 => X"140500090B02C2E0EC04D1C08000000000647E858A104C920C81A5011088A61C",
INIT_09 => X"002481041F165820000101024061004004800567603592A801014C4642601100",
INIT_0A => X"01002020000101B0070310200008B60A23A51B28020CE24E4010026004000440",
INIT_0B => X"03404110230CBA457670820140212100C0692644010001420038935269093161",
INIT_0C => X"2A0872A0C72A0872A0C72A0C72A0872A0C595043950421400800009010104280",
INIT_0D => X"8852141110244066C0820221480010AA73000420808CAC040464D280144050C7",
INIT_0E => X"410082022C000C0002020094030220C960A0409020481024482501A004014100",
INIT_0F => X"6DA02836090540355D86C046619A54052A5B86A0466196940631682800048010",
INIT_10 => X"8B68AA2C60289802AB86A046619A54052A5B86C04661969406316AC018B0E293",
INIT_11 => X"1FC09CB0E1076D4A200B2AC611A3D0405886C6EB211550815A8A2686EC81E2A4",
INIT_12 => X"9C0418CE0C5E8F650E48000892B37885620C1E1A06D7016A90A4626D82B10F1B",
INIT_13 => X"F1E164E02144D335546F28724001B030A56140A184483000C410A2699A2E32AC",
INIT_14 => X"415AAE8018A0A01B2990242E278056AAA203920E0BAE2012C08281808319C186",
INIT_15 => X"9B80D44F9051C049B18A12CB481042AD140C227002A0A02066954E7540CCDB58",
INIT_16 => X"4090240902468118104408000904C0C0964200800200108010003A02272400C1",
INIT_17 => X"0902409024090240902409024090240902409024090240902409024090240902",
INIT_18 => X"1004010040100401004090240902409024090240902409024090240902409024",
INIT_19 => X"2014002840000000000000000004010040100401004010040100401004010040",
INIT_1A => X"0020820820820820A069105251C00000015418982201060302C4281390042104",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFE0FC1C000000000000040200000000000000000001008000000000000",
INIT_1D => X"55000015400000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"B5500003DF55F7D568AAAFFFBC2010557BEAA10AAFBE8A00557BFFFEF007BC21",
INIT_1F => X"75455D7FE8BFF5D7FD540055003FFEFFFD142145000000000FF842ABEFA2AAA8",
INIT_20 => X"C0145557FC2010557FFDF55F7D168A00552E95555007BFFF55087BE8BFFFFD55",
INIT_21 => X"56ABFFA2D16AB550000021FFF7D17FFEF08042AB55A2AAAAB4508517FE00557B",
INIT_22 => X"7FFFE10002ABFE00AAFFE8AAAFF8402000550002145085555400F7FFE8A00085",
INIT_23 => X"8043FEBA002A975EFF7D17DFFFAA8000010000000010F7D5421EF007BC01FF5D",
INIT_24 => X"000000145FFAE820AA007BFDFEF55003FF55A2D557400557BC2145A2D1421450",
INIT_25 => X"8557BF8FEF1C7FC516D080E15400000000000000000000000000000000000000",
INIT_26 => X"00F7842FBD7B6AAAAB551C0E3AF55F7DF68ABAE3F1C00005D7BEDA00B6F1EFA2",
INIT_27 => X"F7D147BEFBEFEBD15257D5D7FEFBD7417BD5438550038FC7FFDF4216D080E070",
INIT_28 => X"DB4514517FE105575C216D5571C50104171FDF7DE3D16DA0041209056D1C71F8",
INIT_29 => X"52400FFF1EFA0008556FBD7B6DB6AB7D1C0A001D7FFD178FC71C0E28B6DA2AEA",
INIT_2A => X"1401D71C7FC21EF5D75FFE10142EBAE10A2FBEFA92F78A05028550E001451455",
INIT_2B => X"71C016DB6D54514500003FEBA1420905FFFFDF78FC7BE84050101C0005000E3D",
INIT_2C => X"0000000000000000000000016DF7AA82092147BFAFEF49043AF45A2DF504285D",
INIT_2D => X"5D7FFDE00F7D17FEBA557BEABEF557BD55EF082A974000000000000000000000",
INIT_2E => X"5F7FBC01FF082A97410FF803DF45FFAEA8B555D2EAAB45F7FBE8ABAAAD540010",
INIT_2F => X"100804001EF55516ABFF557BFDFEFA2D5401FF5D7FFDF55007BD74BA5D042AB4",
INIT_30 => X"B55552AA8BEFAAAABFF5555517FE005555401FF55515541000517FFEFAAD17DE",
INIT_31 => X"74BA5D2A801455D5140000FFD57FE0008557FF45FFFFE8BEF5D2E80155FFD168",
INIT_32 => X"174105D0417410AAD540155557FC01EF5D557DE105D2AA8A10AAFBFFE00F7AA9",
INIT_33 => X"02AB45AAFFC00AA5D51401FFFFD15555500003FEBA5D04001EFFFFFE8B55FF84",
INIT_34 => X"00000000000000000000000000000000000000001FFF7AA800105D7FE8BEF080",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"1000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(11),        -- Port A data input
DOA(0)   => data_read_a_hi_256(11),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(11),        -- Port B data input
DOB(0)   => data_read_b_hi_256(11),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_12_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50080B01BC002006940202C0DE041196A83183000000023322287E0FC000006",
INIT_01 => X"0E000C068000E04D40238000001702684000000008000008820009280A553231",
INIT_02 => X"2809AD0E7D180040945008040090000061800000C0E2F66009DA3D11CB148015",
INIT_03 => X"210D050012F6F8D2108216E24842005B8A20640008800000B8E0141C28851006",
INIT_04 => X"0080100022408000060DE0C00466630C70241837041000040800820480001AA4",
INIT_05 => X"04800018800000003C808003E0C8001401000000040900020904004000070800",
INIT_06 => X"00074000601300119E12D348438000803030800020100800AF08000261042400",
INIT_07 => X"8C53200CA4850224301807D1CB45900147E03040083124FC0CD0C8A1FF00198C",
INIT_08 => X"46050013081206A4A503A9E8C0812000001C7E11A24058B84D40E33992D98F7E",
INIT_09 => X"1004810491175C200000820018A5104010C01086003C13E000004EDF02040004",
INIT_0A => X"0000000000010000180018200408B27E234913E9004CFA09A818024800902109",
INIT_0B => X"014100580004304D267C06CCD0056600007827C00000008C00000000000219C0",
INIT_0C => X"2F0C32F0832F0832F0C32F0832F0832F0C197861978400040000208010120ACA",
INIT_0D => X"E0BF40403CFE7E03E8080382FD0018FE670004000006AE01180493C5BC1AF083",
INIT_0E => X"2000401EA0000440000800A0040028108000000000000000000000A74812DF00",
INIT_0F => X"C48DF8362F658A7E5F82CD23B6B0E403DBBE82C563B6A4E403DBB88C0E048200",
INIT_10 => X"454CFBE5403AB992F282C563B6B0E403DBBE82CD23B6A4E403DBBB1084E4B25A",
INIT_11 => X"851000E4B1D32BAB504BB74AD3F3FE04A8E0D0C319A7988B6F0C75CFD801A962",
INIT_12 => X"BEC4118D994B866E2E8C3808B6B63040328E7A33AF99B0AC20DE634D06C437BF",
INIT_13 => X"70CDC5F6214CA5991C6A7177402C49CA354D808D358A927EAD10A652CC8E3538",
INIT_14 => X"49F36E80083C3EAEB2003695430A7CDAA289553922990C11A4E494988231B325",
INIT_15 => X"3BC0FD5B304AD05A946D81616970A225658940BA7CDAA0A312666BD600E5550B",
INIT_16 => X"00000000001000000104200A89A4D0040000008003B81000000021CFEE02E280",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"8020080200802008020000000000000000000000000000000000000000000000",
INIT_19 => X"0544202101000000000000000000080200802008020080200802008020080200",
INIT_1A => X"4124924924924924481C040000B51451440146E518222204D82A5446021090CB",
INIT_1B => X"2C964B2190C86432190C86432190410410410410410410410410410410410410",
INIT_1C => X"FFFFFFFEF001D64B2592C964B2592C964B2592C964B2592C964B2592C964B259",
INIT_1D => X"00AAFBC2000000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"A00557BFFFEF007BC2155000015555087FC0010AAFBFFE100004020BAAAFFD54",
INIT_1F => X"2155AA8400000A2AABFF45550400000AAFBFFFEF550000010557BEAA10AAFBE8",
INIT_20 => X"C0010555155555FF8017400FF842ABEFA2AAA8B5500003DF55F7D568AAAFFFBC",
INIT_21 => X"FE8BFF5D7FD540055003FFEFFFD142145000000145A2AA821EFFFFFD7410007F",
INIT_22 => X"7BE8BFFFFD5574000051420BA557FC2145557FC20AAA2D57DEBAA2FBD55455D7",
INIT_23 => X"82EAAA00550415410AAFBFFFEF55042AB55F7D168A00552E95555007BFFF5508",
INIT_24 => X"000000155A2AAAAB4508517FE00557BC0145557FC2010557FFDE10AA84000000",
INIT_25 => X"0000A02092B6F5D2438A2FBC2000000000000000000000000000000000000000",
INIT_26 => X"005D7BEDA00B6F1EFA28557BF8FEF1C7FC516D080E1557D0075C7028B6F1FAE0",
INIT_27 => X"F55F7DF68ABAE3F1C017DAA8E07028B6A0BFF6D490E00000BEF5FAFEF4904070",
INIT_28 => X"51FFE3FBD0438007FC00385D555556DEB8410400F7842FBD7B6AAAAB551C0E3A",
INIT_29 => X"7DEBAA2FBD557D5D7FEFBD7417BD5438550038FC7FFDF4216D080E0716DAAA08",
INIT_2A => X"09056D1C71F8F7D147BEFBEFEBD152400005F450BA417BC51454971C20AAB6D1",
INIT_2B => X"71FDE10BE8E070280020AAA28410410400BEFBFAFEF49042AB7DE3D16DA00412",
INIT_2C => X"0000000000000000000000016DA2AEADB4514517FE105575C216D5571C501041",
INIT_2D => X"0055574BAFFD568A10002A82000FFD5400AAA2FBC00000000000000000000000",
INIT_2E => X"0FFD568BEF0004174105D7FFDE00F7D17FEBA557BEABEF557BD55EF082A975EF",
INIT_2F => X"45FFAEA8B555D2EAAB45F7FBE8ABAAAD5401EFA2AA974BAF7803FFFF002A8200",
INIT_30 => X"1FF082A975EFA280175FFAAFFC00BA087FC20AA5D55555FFA28000010FF803DF",
INIT_31 => X"75450851420BAFFD57DEAAAAFBD75FF5D7FFDF55007BD74BA5D042AB45F7FBC0",
INIT_32 => X"28BEFAAD17DE100804001EF55516ABFF557BFDFEFA2D540010007FD74AA007BD",
INIT_33 => X"5401FF55515541000517FE10F7AA954AA080428AAA000002010FFFFE8BEF0804",
INIT_34 => X"00000000000000000000000000000000000000001EFAAAABFF5555517FE00555",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"01FFFFFFFFE00000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(12),        -- Port A data input
DOA(0)   => data_read_a_hi_256(12),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(12),        -- Port B data input
DOB(0)   => data_read_b_hi_256(12),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_13_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10110A0441812402840402822007818000E00700000000330A3000000008042",
INIT_01 => X"A1400984B830C848180260000C0042404001000008220008A200100802110200",
INIT_02 => X"88010C02801040002475580400800000410000000064024608134C0CC9018034",
INIT_03 => X"00010100926220D084234212421085084300648A0880000630C0654288C10000",
INIT_04 => X"0004122122029100100C00001200009C40A83A2044360C84190BAC04E0101820",
INIT_05 => X"04E000008009050064C8C00104C10184034010250089C00EB004327064B60900",
INIT_06 => X"CA875CA8600000880410DA8C285001802424B008881024A8204E010461042700",
INIT_07 => X"08320014B02848A4A8100015C55500057801A04000712C040CB1F8806000088D",
INIT_08 => X"5005000908020220E40170008042000000557E048A144C800590010000882D00",
INIT_09 => X"00250104B5310020000100020821004016CC1C616401910801010100CA204000",
INIT_0A => X"0000000000010192072310200028B602234608080280074AC010025900100401",
INIT_0B => X"014100101118BA451000824150052110480121000140014200101352690BAC20",
INIT_0C => X"0000000040000000000000040000000000000020000000000000008010102A82",
INIT_0D => X"094040100000006C0802042501001C8017000C21908200028448400000000040",
INIT_0E => X"000000010C000C00081A08BC832A209AB0A85094284A14254A25510105130801",
INIT_0F => X"30BA901293C0F5012906A96DCD13042CE0C206E92DCD07042CE0C40D02048000",
INIT_10 => X"4CA4271CA2168ACB0E06E92DCD13042CE0C206A96DCD07042CE0C4408632C395",
INIT_11 => X"58408632C30D522CE80239CC2806AC44E954939AB299E000738F88296CA13B44",
INIT_12 => X"5145CD5306028F01990C080808494A64708B265CC4052B0F30302E060965EA00",
INIT_13 => X"51E0328A2CA9722094650CCAC0629112BA89C04A228568547B1654B9104A3286",
INIT_14 => X"A158BB80D4D8D48CB54012290470562EC29E44050B1DC60132282B68B9AA60C0",
INIT_15 => X"280000A5C11B9008FE2FA38F87804251CB0FAD40562EC0B426149D17E0044B10",
INIT_16 => X"509425094246A10A10441010090480C0964201800044109012001A000726E454",
INIT_17 => X"0942509425094250942509425094250942509425094250942509425094250942",
INIT_18 => X"9425094250942509425094250942509425094250942509425094250942509425",
INIT_19 => X"7E24502A80000000000000000005094250942509425094250942509425094250",
INIT_1A => X"AEBAEBAEBAEBAEBAFFD7F7F7F775555557DFBEEFBBFCFDF7DFFCF9F80089F7DF",
INIT_1B => X"BF5FAFD7EBF5FAFD7EBF5FAFD7EBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEB",
INIT_1C => X"FFFFFFFE0001DFAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7E",
INIT_1D => X"4500557DE00000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"E100004020BAAAFFD5400AAFBC2155AAAA97410FFFFEAAAAF7AA955EFF7803FF",
INIT_1F => X"5410F7AEBDE10FFFFFDEAAF7D568AAA5D002AB55005568B55087FC0010AAFBFF",
INIT_20 => X"555FF5D04154BAAAAEAAA10557BEAA10AAFBE8A00557BFFFEF007BC215500001",
INIT_21 => X"400000A2AABFF45550400000AAFBFFFEF550000155A28415410F7AEAABFFA2D1",
INIT_22 => X"D568AAAFFFBC21555D517FF45F7AEA8BFFA2AEAAA10A280021EF5D557FF55AA8",
INIT_23 => X"AAE974AAF7D142145082A975FF555568A00FF842ABEFA2AAA8B5500003DF55F7",
INIT_24 => X"000000145A2AA821EFFFFFD7410007FC0010555155555FF80174000055555EFA",
INIT_25 => X"2E3A0925C7E38E38F7D14557AE00000000000000000000000000000000000000",
INIT_26 => X"7D0075C7028B6F1FAE00000A02092B6F5D2438A2FBC2145B6A090428FFF5EAA9",
INIT_27 => X"FEF1C7FC516D080E15438E3A4BAE00FFF5FAE92F7D16AAAA41042FB7D145568B",
INIT_28 => X"2428FFA4AFBFFAAD1505FF490E174AABEA0ADA005D7BEDA00B6F1EFA28557BF8",
INIT_29 => X"001FF555F7FF7DAA8E07028B6A0BFF6D490E00000BEF5FAFEF490407155BE8E1",
INIT_2A => X"AAAB551C0E3AF55F7DF68ABAE3F1C0145415B78F45FFA4AFBC7BEA4AAA10A284",
INIT_2B => X"84104380055525FFBEAE90482E3D54216D0024975FF555F68A00F7842FBD7B6A",
INIT_2C => X"0000000000000000000000016DAAA0851FFE3FBD0438007FC00385D555556DEB",
INIT_2D => X"FF80020BAF7D16AA10A28402155A2AEA8BEF5D516AA000000000000000000000",
INIT_2E => X"A08003DFEF55516ABEF0055574BAFFD568A10002A82000FFD5400AAA2FBC0145",
INIT_2F => X"00F7D17FEBA557BEABEF557BD55EF082A974BAA28028A00F7D16AA10F7D56AAB",
INIT_30 => X"BEF000417545FFAA820BAFF843DFFFA2D5421FF002E954AAFF843DE105D7FFDE",
INIT_31 => X"DF55F7802AA10AA80001FF5D7FFDFEFA2AA974BAF7803FFFF002A82000FFD568",
INIT_32 => X"EAA10FF803DF45FFAEA8B555D2EAAB45F7FBE8ABAAAD540145007FE8B55FF843",
INIT_33 => X"FC20AA5D55555FFA280000BA0855401EFF7AA82010AAD1421FF0004155FF557F",
INIT_34 => X"00000000000000000000000000000000000000001EFA280175FFAAFFC00BA087",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"19FFFFFFFFE00000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(13),        -- Port A data input
DOA(0)   => data_read_a_hi_256(13),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(13),        -- Port B data input
DOB(0)   => data_read_b_hi_256(13),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_14_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10020A000180000284008280000281800000030000000033022000000580002",
INIT_01 => X"A140098018300848184860000C20C24040000000084000084200000000110200",
INIT_02 => X"88010C5A8010A600A4F558040080000041000000022C024008003CCCC9028030",
INIT_03 => X"000103A7A00904D0842242024210810803006480088000003081054288C10000",
INIT_04 => X"0000120122009000100C00000000000400A83A2044200C840000800400101820",
INIT_05 => X"040000008008010024C0C0010040000402000025000800020004207000100800",
INIT_06 => X"40870408600800800410D006A850018024240008881024A82040010461042000",
INIT_07 => X"08120054B42850B42A100010ED1500010001A040003164040CF5E20140000888",
INIT_08 => X"400500090A020220A40A7000800000000014FE8508144C924080C10000880140",
INIT_09 => X"0004010411110020000100020021004000800461600191080101000042200000",
INIT_0A => X"0000000000010190070310200008B202236D080802000002C010024000000000",
INIT_0B => X"0141001001088A45000082400000010040012100010000020000135249020820",
INIT_0C => X"0004000000000000004000000000000004000000000000000000008010100000",
INIT_0D => X"0840401000000044080200210100100017000420808200000440400000000040",
INIT_0E => X"0000000000000C00000000040302200800A04090204810244825010104130800",
INIT_0F => X"397468090008142014840100002C382800008401000038382800006402048000",
INIT_10 => X"83514072C000444C00840020002C38280000840020003838280002C09D010868",
INIT_11 => X"03C09D0104B01C57100440202900184414430534605E38048021800224804191",
INIT_12 => X"40049594C194000090450808802008830024F0E248C902AEF0024170CF180010",
INIT_13 => X"8000120020E5A08E6000048200196264BCF1C030C0604800001076C047300002",
INIT_14 => X"A00002003DEDE82C78900902A0D0000080019FAAA32D9602490302409292B832",
INIT_15 => X"2800D049100021171F6C34080240108AB292CA000000800AD1A19F6F000AA0C0",
INIT_16 => X"409024090246810810440000090480C096420080000010801001600001200454",
INIT_17 => X"0902409024090240902409024090240902409024090240902409024090240902",
INIT_18 => X"9024090240902409024090240902409024090240902409024090240902409024",
INIT_19 => X"6504002800000000000000000004090240902409024090240902409024090240",
INIT_1A => X"E79E79E79E79E79E7FDDF77777F3CF3CF7D55E6D39723FC3DEFA75D77B75F7DF",
INIT_1B => X"9FCFE7F3F9FCFE7F3F9FCFE7F3F9E79E79E79E79E79E79E79E79E79E79E79E79",
INIT_1C => X"FFFFFFFEFFFE0FE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F",
INIT_1D => X"55A28417400000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"AAAF7AA955EFF7803FF4500557DF45F7D16AB455D00001EFAAAAAAABA5555575",
INIT_1F => X"214555003FF450804001555D2AA8AAA002ABDE10082ABDF55AAAA97410FFFFEA",
INIT_20 => X"175EF5D5168A10082E80155087FC0010AAFBFFE100004020BAAAFFD5400AAFBC",
INIT_21 => X"EBDE10FFFFFDEAAF7D568AAA5D002AB55005568A00A2D5401455D00175FFFF84",
INIT_22 => X"7BC2155000015400AAD157545080402145087FD75FFF7AE82145A2D17FE10F7A",
INIT_23 => X"000000BAFFFBE8AAAA2FBFDE00087FD5410557BEAA10AAFBE8A00557BFFFEF00",
INIT_24 => X"000000155A28415410F7AEAABFFA2D1555FF5D04154BAAAAEAAA005D002AB450",
INIT_25 => X"7B6A0AAA82555157555B68012400000000000000000000000000000000000000",
INIT_26 => X"45B6A090428FFF5EAA92E3A0925C7E38E38F7D14557AF45FFDB6AB6D4100071C",
INIT_27 => X"092B6F5D2438A2FBC21455D0A3FF6D080407155552AAAA920020BFE10002EBAF",
INIT_28 => X"01454100175C7E380125D7555B6DA1014248217D0075C7028B6F1FAE00000A02",
INIT_29 => X"82145AAD178E38E3A4BAE00FFF5FAE92F7D16AAAA41042FB7D145568A38AADF4",
INIT_2A => X"1EFA28557BF8FEF1C7FC516D080E15400A2DB5754508040716D007BD05EFEBAA",
INIT_2B => X"A0ADA0055002AB6D0000020BAFFF1E8ABABEF1FAE001C7FD54005D7BEDA00B6F",
INIT_2C => X"00000000000000000000000155BE8E12428FFA4AFBFFAAD1505FF490E174AABE",
INIT_2D => X"F7FFEABFF080015555F78028A00555155555FF84000000000000000000000000",
INIT_2E => X"000003DE10082EAAB45FF80020BAF7D16AA10A28402155A2AEA8BEF5D516AB45",
INIT_2F => X"BAFFD568A10002A82000FFD5400AAA2FBC0145552ABFFFF000417555552EA8A1",
INIT_30 => X"FEF55516AABAAAFFC0145000417555A280001455D7FFDE105504021EF0055574",
INIT_31 => X"55FF007BC01FFAAAE80155AAD568ABAA28028A00F7D16AA10F7D56AABA08003D",
INIT_32 => X"D74105D7FFDE00F7D17FEBA557BEABEF557BD55EF082A97410AAFFD554508001",
INIT_33 => X"5421FF002E954AAFF843DE10550028BEF0004020BAF7D568AAAF7D168A105D7F",
INIT_34 => X"0000000000000000000000000000000000000000145FFAA820BAFF843DFFFA2D",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"01FFFFFFFFE00000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(14),        -- Port A data input
DOA(0)   => data_read_a_hi_256(14),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(14),        -- Port B data input
DOB(0)   => data_read_b_hi_256(14),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_15_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000A000000000284000280000001800020030000000033022000000180002",
INIT_01 => X"A140098018300848180060000C00424040000000080000080200000000110200",
INIT_02 => X"080108000010E60004E55800008000004100000000040240080000C009170016",
INIT_03 => X"0000000080000040842240000210810002000400888000003080014288C00000",
INIT_04 => X"0001100024A0800000440000000000040088322044200C840000011400151800",
INIT_05 => X"440002988000000020000000000B8094020000254C8800000514203000108800",
INIT_06 => X"00070000620040880410D00C285000802424000AA81024A80040010C01062001",
INIT_07 => X"086100043224489428100010811100010001A040003124040CAC600040000888",
INIT_08 => X"160500090A0282A06400100080C300000005BE0488104C800000010000880000",
INIT_09 => X"000581041110022000000002002100400080046140011008010100008A040000",
INIT_0A => X"0000000000010180060210200008B2022304080800000007C010024000000000",
INIT_0B => X"4140001001088A45000082000000010000002000010000020000034249000020",
INIT_0C => X"0004000040000400000000000000000004000020000200000000008010100000",
INIT_0D => X"094000100000004C000200250000188016000400000000000440400000000040",
INIT_0E => X"0000000108000C00000000000200200800800000000000004020000000000000",
INIT_0F => X"0000000000000000000404200000000000000404200000000000008C00048000",
INIT_10 => X"4000000000000000000405000000000000000405000000000000004000001000",
INIT_11 => X"0040000010000000000000000000004000201000000000000000000000800002",
INIT_12 => X"0004000110000000000C00080010180000000001A10240500000000000000000",
INIT_13 => X"0000000020080400000000020000008040020000000000000010001200000000",
INIT_14 => X"0000020000000611002800000000000080000011044220000000000080200200",
INIT_15 => X"8800000100000000009080E2E0A0000000000000000080000040000000000000",
INIT_16 => X"0000000000460000004400000904808094020080000010000000000000000041",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0004002800000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000004000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFE00000000000000000000000000000000000000000000000000000000",
INIT_1D => X"EF08517DE00000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"1EFAAAAAAABA555557555A284175FF000002010552A97400007BFDE10A2AA801",
INIT_1F => X"DFEF5D2AAAB45F7D17DF45087BC0155002A801FF08003DF45F7D16AB455D0000",
INIT_20 => X"C2145F7D568BEFAAD557555AAAA97410FFFFEAAAAF7AA955EFF7803FF4500557",
INIT_21 => X"03FF450804001555D2AA8AAA002ABDE10082ABDFFFF7D17FE10002E954AAF7FB",
INIT_22 => X"FFD5400AAFBC21EFA2AE95545A2D56ABFFAAD17DE10FFD1420AA007FC0145550",
INIT_23 => X"02A801550055401555D00174BA002AA8B55087FC0010AAFBFFE100004020BAAA",
INIT_24 => X"000000000A2D5401455D00175FFFF84175EF5D5168A10082E801FFFF8428A100",
INIT_25 => X"80871FAE00A2A0871EF145B7FE00000000000000000000000000000000000000",
INIT_26 => X"45FFDB6AB6D4100071C7B6A0AAA82555157555B680125C71C0E0500049209543",
INIT_27 => X"5C7E38E38F7D14557AFC75524AFB45FFD178F7D1C71C2145002E801C7140A3FF",
INIT_28 => X"AE000024954AAFFFBC2145F7DB6DBEFA2D557545B6A090428FFF5EAA92E3A092",
INIT_29 => X"470820071C71455D0A3FF6D080407155552AAAA920020BFE10002EBAFC7FFDF7",
INIT_2A => X"1FAE00000A02092B6F5D2438A2FBC21FFBEA090545B6D568BFFAADB7AE10F7D5",
INIT_2B => X"24821FFE3802FA2808208017D1C5142155410A104AA1420AFB7D0075C7028B6F",
INIT_2C => X"00000000000000000000000038AADF401454100175C7E380125D7555B6DA1014",
INIT_2D => X"552E954100004174AA00516AA10AA80155EF5D7BFDE000000000000000000000",
INIT_2E => X"5082E801555D2EBDF45F7FFEABFF080015555F78028A00555155555FF8400155",
INIT_2F => X"BAF7D16AA10A28402155A2AEA8BEF5D516AB555D043DF55F7D56ABEF55514015",
INIT_30 => X"E10082EAAB55FFFBE8A100804154AAF7FFC2145FFFFFDFEFAAD157545FF80020",
INIT_31 => X"ABEFA2FBE8A00FFD155410005555545552ABFFFF000417555552EA8A1000003D",
INIT_32 => X"3DFEF0055574BAFFD568A10002A82000FFD5400AAA2FBC01FFF78400155F7D16",
INIT_33 => X"0001455D7FFDE105504021FFAA843DEBA0000021EF555142155002E800AA5500",
INIT_34 => X"00000000000000000000000000000000000000000BAAAFFC0145000417555A28",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"1800000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(15),        -- Port A data input
DOA(0)   => data_read_a_hi_256(15),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(15),        -- Port B data input
DOB(0)   => data_read_b_hi_256(15),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_16_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"DA22C618B1000482B688B186588884862A400438255FC38381441205BA803003",
INIT_01 => X"8645A80028404C211203A952A90341080B173340412000E1005D628000820484",
INIT_02 => X"A101A9006DC1084833011850AAC55001349B10881802821808B4110007005E11",
INIT_03 => X"010108A802BB00080080006020020001A61036202800000D2410104200404550",
INIT_04 => X"8BFA58800005C40A46240252145148B38248030356415A4E62B6FC660F287240",
INIT_05 => X"1E0BD423CAC0000D610000000710296E542B6E3A825C15FB30A643695BFC2D56",
INIT_06 => X"000D0000C8008820CAE16020619156A5815006028179808C00A0D2152B90707A",
INIT_07 => X"F500240510A00205F0A407D0021A155378900002A002433A0AA00EE6E7956108",
INIT_08 => X"015995440C8327241440096A2800002828123D542910380004E0310362404076",
INIT_09 => X"10222D90409A05B2CB2CA400200209E5601044A24000000462A6001888010000",
INIT_0A => X"0000000000259200140001A15000017F0051D0F837248C005514AC40C0820500",
INIT_0B => X"01200848002912300200092BA80325A2000000000001514B5500030241C000CC",
INIT_0C => X"0001100011000110001100011000110001080008800080005202280801080395",
INIT_0D => X"17680002815014B90000205DA00880100095A64800008003561180063DB4F611",
INIT_0E => X"0280080922554515512174000000490009000000000000004010042A204A0C58",
INIT_0F => X"2DA0063EAA9C238B2D4C800632B266E828EE4C800632AAAB6830D0FC6B06C041",
INIT_10 => X"0839AA149339E8FB964C800632B266E82B2E4C800632AAAB683310872800EDA5",
INIT_11 => X"C087A800EB090D4AAC91268FFCBE81397826C4A20D2B6C510E8624792A4A30A4",
INIT_12 => X"3638E8849D5C532408DD6E004C90C06AC019D88B9795012CA96902C799912BC3",
INIT_13 => X"78706531C74485BD42A30906057FADAA456218FD8E3ED83B60E3A242DC0F1898",
INIT_14 => X"51727A06FB555793057C444CF45C5C9E89543B8BC6E80193DC36F6C71D1093A4",
INIT_15 => X"10DCD45DC02B331650CA8ACB4007E00D1C6A6A58395C917F7E74D936F650D69B",
INIT_16 => X"000000000012000081500008A422150884081ACAAC0542054004FC5884640508",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"3604000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"45145145145145147A7797E1E1A79E79E15634455131A436993071A616D4F68A",
INIT_1B => X"3E9F4FA7D1E9F47A7D1E9F47A7D3453453453453453453453453453453453453",
INIT_1C => X"FFFFFFFE00001F4FA7D3E9F4FA3D1E8F47A3D1E8F47A3D1E9F4FA7D3E9F4FA7D",
INIT_1D => X"00FF8015400000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"400007BFDE10A2AA801EF08517DE10FFFFFDFEFA2D16AB55A2FFFFEAA5D7FC00",
INIT_1F => X"74BA5D2EBDFEFAAD17FFFF002EBDE000800174AA55043FFFF000002010552A97",
INIT_20 => X"E8AAAAA80000105D557FF45F7D16AB455D00001EFAAAAAAABA555557555A2841",
INIT_21 => X"AAAB45F7D17DF45087BC0155002A801FF08003DE000004154BA002A800BA087F",
INIT_22 => X"803FF4500557DEAAF7D57DEBA082A82010FFAE975555D7FFDEAAFF80155EF5D2",
INIT_23 => X"2D57FFFF557FD55FF08003FE0055043FF55AAAA97410FFFFEAAAAF7AA955EFF7",
INIT_24 => X"0000001FFF7D17FE10002E954AAF7FBC2145F7D568BEFAAD557410552EA8BEFA",
INIT_25 => X"DB6FFFDEAA5571C7010FF8412400000000000000000000000000000000000000",
INIT_26 => X"C71C0E050004920954380871FAE00A2A0871EF145B7FE10E3F1F8FC7AAD56DB7",
INIT_27 => X"A82555157555B680124924124BDFEFA2D57FFC71C2EBDE280000174825D0E3FF",
INIT_28 => X"74821424800AA007FEDAAAA284020385D5F7AF45FFDB6AB6D4100071C7B6A0AA",
INIT_29 => X"F8EAAFF80175C75524AFB45FFD178F7D1C71C2145002E801C7140A3FE10080A1",
INIT_2A => X"5EAA92E3A0925C7E38E38F7D14557AE92EBDB78EAA1C2482010FFAE9556D557F",
INIT_2B => X"D557410492EADBEFA2D178FEF5575D55EF000A38E10490A3AF45B6A090428FFF",
INIT_2C => X"000000000000000000000001C7FFDF7AE000024954AAFFFBC2145F7DB6DBEFA2",
INIT_2D => X"A2D56AB45A2D57DFFFF7FBFFEAA555555400F780000000000000000000000000",
INIT_2E => X"A080415400552ABDF55552E954100004174AA00516AA10AA80155EF5D7BFDE10",
INIT_2F => X"FF080015555F78028A00555155555FF840000000043DFEFAAD17FF45552ABFEB",
INIT_30 => X"1555D2EBDE10002E974005D04020BA007BFDEBAA284000BA557FE8B45F7FFEAB",
INIT_31 => X"0000F7AE955EF5D7BE8ABAF784175555D043DF55F7D56ABEF555140155082E80",
INIT_32 => X"AAB45FF80020BAF7D16AA10A28402155A2AEA8BEF5D516AA00AAFBE8AAA55040",
INIT_33 => X"FC2145FFFFFDFEFAAD157410082ABFFEFAAD16ABFF5555575FF082AA8A00002A",
INIT_34 => X"0000000000000000000000000000000000000000155FFFBE8A100804154AAF7F",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0800000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(16),        -- Port A data input
DOA(0)   => data_read_a_hi_256(16),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(16),        -- Port B data input
DOB(0)   => data_read_b_hi_256(16),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_17_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"5284CE4FB7BD2C8994A13392DBD02E14006B82AC7E800D44D3DD2FD5F9B961C0",
INIT_01 => X"F8ACD01F7E03FC6793F2199B39FC233C11D93AE6F3BB92B32091DBC339B24542",
INIT_02 => X"8F333007FD6808092A2AFA6667033DB50853379C10BFF70F1BD011110F205F18",
INIT_03 => X"294ADB4AFFCBF0DAD63ABF836B58EAFE060478202022234B2E0303FDC9E18339",
INIT_04 => X"DB7A40806FE4040840EBC563A0150A0926146FECB04196482236FC2005282AE1",
INIT_05 => X"0807B4070670083DC68206D7E6D0250834336D1E81500FDB306045255BFC2076",
INIT_06 => X"00000000141C5AF3EA6AB187F7F8CE039786062C6CE092F5FE005236781C402A",
INIT_07 => X"1684248A38B022475DCA9BD00116E33CC3821774BB55F53BB42329AA3C0CEF60",
INIT_08 => X"60700CE0641527241060AD844E1C0088001223022D189A2800542219204903F8",
INIT_09 => X"D94C1C1C51DFF881861CBE0305A12A0321810217C01D34EDC98FFA1C8E000016",
INIT_0A => X"7E7D8F8FBDE40E001E000B3A5DAADAFDDA5DA79350DF70027CE86F047BEF19B6",
INIT_0B => X"814102F800633F1D0A7CC9AE74117FE0003A6AD055819D1F9984014B37BA5FFC",
INIT_0C => X"CF4FBCF4FBCF4FBCF4FBCF4FBCF4FBCF4FBE7A7DE7A7800617112E46F05D02DD",
INIT_0D => X"D7FE4A5A99FD6D3FEF4BEB5FF994F0FEFFCCF8430006CE8A3F06ABD73DBCF4FB",
INIT_0E => X"B29760593F33FA0CF170F40006001B1A05C0000000000000008004BA78428C7A",
INIT_0F => X"EDA57E46444357B3950A9BFBAC94CFA8581E0A9BFBAC8CCFA8580C7CAF51EF68",
INIT_10 => X"7DF76B5DB54A09003E0A9BFBAC94CFA8581E0A9BFBAC8CCFA8580E46FBFCB0CB",
INIT_11 => X"E7467BFCB1D5CFEB56A1A100D5345C1BFFE8FBDB892DB463034198E2881F3F78",
INIT_12 => X"4E0ADD39387F92B2935DFEAADDF38EBCFB9E3D636DCDF9B90F966BF92966D5D9",
INIT_13 => X"F256527055EB6D555CB294981B7FB5B2954CD3013013FDF5E82AF5B6AAAE594A",
INIT_14 => X"F7D7E835C67E655BAA868610117575EA1C34BD6975D48B44A0405FC15BA7270F",
INIT_15 => X"BD07F6CD2A47D0CBA96252756D7217E5E1C61DBDF5FA167F7AE5D3D21A414007",
INIT_16 => X"00000000005F08000179C16DECF67F08BC02F9067ED55805600545DFE45A80E7",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"F981800C00000000000000000000000000000000000000000000000000000000",
INIT_1A => X"A69A69A69A69A69A919261A1A6075D75D10DC800C027B731014BA4B864617114",
INIT_1B => X"8341A0D068351A8D068351A8D069A6BAE9A69A6BAE9A6BAE9A69A6BAE9A6BAE9",
INIT_1C => X"FFFFFFFE000011A8D46A351A8D46A351A8D46A351A8D46A341A0D068341A0D06",
INIT_1D => X"55AAFFD5400000000000000000000000000000000000000000000001FFFFFFFF",
INIT_1E => X"B55A2FFFFEAA5D7FC0000FF8015410FFFFFFFFFFFFFFDFEFF7D568A1008003DF",
INIT_1F => X"DF55A2D1400000804154BAF7D168A00A2803DE10FFAE95410FFFFFDFEFA2D16A",
INIT_20 => X"2AABAFFD56ABFF002EBDFFF000002010552A97400007BFDE10A2AA801EF08517",
INIT_21 => X"EBDFEFAAD17FFFF002EBDE000800174AA55043FEBA0004174AA5504000AA5504",
INIT_22 => X"5557555A284175FFFFFBE8B55A2FFFFF55F7803DEBA002AAAAAAF7FBD74BA5D2",
INIT_23 => X"D0417400FFD57DE00AAAAAAB45A2AA97545F7D16AB455D00001EFAAAAAAABA55",
INIT_24 => X"0000000000004154BA002A800BA087FE8AAAAA80000105D557FE00A2D5420AA5",
INIT_25 => X"7EBD16AA00000E3DF6DBEF5D2400000000000000000000000000000000000000",
INIT_26 => X"10E3F1F8FC7AAD56DB7DB6FFFDEAA5571C7010FF8412428FFFFFFFFFF7FBF8FD",
INIT_27 => X"E00A2A0871EF145B7FF7DA2D547038140E10492FFDF6DA28A28E3DE00F7A0924",
INIT_28 => X"2492550A020BA55002AA82F7DF6DBD71C2EBFFC71C0E050004920954380871FA",
INIT_29 => X"ADABAF7F5D74924124BDFEFA2D57FFC71C2EBDE280000174825D0E3FEAA14001",
INIT_2A => X"0071C7B6A0AAA82555157555B680125FFEBFFEDB55BEFFFAF6DE38E3DEAA002E",
INIT_2B => X"5F7AE28B6D545092490E10400FFDB7AE00A2AAADB45BEA092545FFDB6AB6D410",
INIT_2C => X"00000000000000000000000010080A174821424800AA007FEDAAAA284020385D",
INIT_2D => X"FFFBFDFEFF7FFEAB45A2D56AA00002EBDFFFF7D5400000000000000000000000",
INIT_2E => X"AA2AABDE10FF8400010A2D56AB45A2D57DFFFF7FBFFEAA555555400F780000AA",
INIT_2F => X"100004174AA00516AA10AA80155EF5D7BFDFEFAAD1554BA552E82000F7FFFFEA",
INIT_30 => X"400552ABDEBA5D0002000552A800BA55042AA10FFFFFDF55552EBDF55552E954",
INIT_31 => X"ABFFA2AEBFEAA082EBDEBAFFD55540000043DFEFAAD17FF45552ABFEBA080415",
INIT_32 => X"00145F7FFEABFF080015555F78028A00555155555FF84001FFAAFBFFF55FFFBE",
INIT_33 => X"BFDEBAA284000BA557FE8AAAFFD155400082A82000F7FFE8A00A2AABDF45F780",
INIT_34 => X"0000000000000000000000000000000000000000010002E974005D04020BA007",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"19FFFFFFFFE00000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(17),        -- Port A data input
DOA(0)   => data_read_a_hi_256(17),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(17),        -- Port B data input
DOB(0)   => data_read_b_hi_256(17),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_18_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"69844019080000A21A611406840014122A641074155FC28A2024001001801003",
INIT_01 => X"A643D920034004180005E9E3C90360C0041C0181002001602025800008440084",
INIT_02 => X"B7333980808408103F2000F81FC0FEDEAC2161B0B84D0002188011110C018041",
INIT_03 => X"0405D434003F2C020081587008020561E55116B0290000042B71240C800440F8",
INIT_04 => X"50805AC31007D6125724029216554A9847669903D640EC8E2001002604503004",
INIT_05 => X"0E010001C1CA11803850C800010022660C1C0065003C0404002646DC20A02D40",
INIT_06 => X"50AD050AC00000002A4F612449903FE080000000005889AC41E04508A9907020",
INIT_07 => X"5584280B10014003A8067400920810FF3C72024300A0030048221ACEE383E518",
INIT_08 => X"00C983E6041505253500F66E620428000B1804000152E52801A2020084090040",
INIT_09 => X"20500B90419005B0C309402030060860E01004A828408800440405E350294010",
INIT_0A => X"008010100007865421432121804021C20452880C2D200000045C18C0E0000A08",
INIT_0B => X"09700C04C44C92A88DC42215C882E82250811000000C1AE061861710A401A4E8",
INIT_0C => X"308003080030800308003080030800308001840018400400602A018809800371",
INIT_0D => X"0801010202021000780004200408C1002003F66CA1B13111C0D95C20C2030A00",
INIT_0E => X"02900806400FC503F08180050942E4200020C1B060D8306C182701404C197301",
INIT_0F => X"22AABABAF377DF1CA160820520EB3057E70E60820520F33057E72E9154159000",
INIT_10 => X"8A2AD5D48F37FAFEFE60820520EB3057E7CE60820520F33057E7EC658BF2DA78",
INIT_11 => X"32658BF2D4B2A80BF8FE39FD78EB0D882014A62C568FFAFC73FFDD9C2B30E046",
INIT_12 => X"C728C800DFC06F59F710107533C0C4E37619440FBFBAB2400AFC1600361D798F",
INIT_13 => X"0DEBBEB9454005BAA36DEFF894823A3D1A88A2FE29D5FC6DCAA2A002DD51B6E7",
INIT_14 => X"F3B7092A78606A28A5427AAB9FF4EDD251C7123E291660733EBF6FE519001BF4",
INIT_15 => X"82202AB58AFBFD5DE200A8EBE3A3EC110339E1DCEDC2590495BB2112E2BE4BF5",
INIT_16 => X"C1B06C1B06808348340000020301805002D008C1F92000A5F421B8000DB49103",
INIT_17 => X"1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06",
INIT_18 => X"B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C",
INIT_19 => X"16000000000000000000000000041B06C1B06C1B06C1B06C1B06C1B06C1B06C1",
INIT_1A => X"A28A28A28A28A28A244C16454170410412CA2EFB3AE03B85CF08C03F1A30F7DF",
INIT_1B => X"8944A25128954AA552A944A2512AAA8A28A28A2AAAAAA8A28A28A2AAAAAA8A28",
INIT_1C => X"FFFFFFFE000004A25128944A25128944A25128944A25128944A25128944A2512",
INIT_1D => X"105D2A80000000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"FEFF7D568A1008003DF55AAFFD5410FFFFFFFFFFFFFFFFFFFFFBFDEBA552E974",
INIT_1F => X"5410FFFFFFFFFF7FBE8B55AAD16AA1000516AA005D0400010FFFFFFFFFFFFFFD",
INIT_20 => X"FFE00087BC2155087BC0010FFFFFDFEFA2D16AB55A2FFFFEAA5D7FC0000FF801",
INIT_21 => X"1400000804154BAF7D168A00A2803DE10FFAE95555FFFBE8B45A2D56ABEFFFFF",
INIT_22 => X"AA801EF08517DF55000000010082A974AA08557DEBAFFAEBFF55AA8028B55A2D",
INIT_23 => X"52E800105D2AAAA10A2D1420AAFFAEA8BFF000002010552A97400007BFDE10A2",
INIT_24 => X"0000000BA0004174AA5504000AA55042AABAFFD56ABFF002EBDEBA0004020BA5",
INIT_25 => X"FF7FBFFEBA552A95410552485000000000000000000000000000000000000000",
INIT_26 => X"28FFFFFFFFFF7FBF8FD7EBD16AA00000E3DF6DBEF5D2438FFFFFFFFFFFFFFFFE",
INIT_27 => X"EAA5571C7010FF8412410FFFBF8FC7E3F5EAB45BEDB6FA3800556FA005504050",
INIT_28 => X"AB55BEDB6FBC7EBF5F8E10007BC516D1C71C5010E3F1F8FC7AAD56DB7DB6FFFD",
INIT_29 => X"BFF55BE8A2DB7DA2D547038140E10492FFDF6DA28A28E3DE00F7A09256DE3F1E",
INIT_2A => X"0954380871FAE00A2A0871EF145B7FF45080E070280820924AA145578E92F7A4",
INIT_2B => X"2EBFEBA1C0A00092412E850005D2AAFA38A2DF45082F7AAA8BC71C0E05000492",
INIT_2C => X"000000000000000000000000AA140012492550A020BA55002AA82F7DF6DBD71C",
INIT_2D => X"FFFFFFFFFFFFBFDFEFF7FFFDEAA5D2E954105504154000000000000000000000",
INIT_2E => X"A08557DE005500154AAFFFBFDFEFF7FFEAB45A2D56AA00002EBDFFFF7D5400AA",
INIT_2F => X"45A2D57DFFFF7FBFFEAA555555400F78000010F7FBE8B55AAD16AB55F7FBFDEA",
INIT_30 => X"E10FF84001FFAAD568B45FFFBFFF55A2D568A00087BD55FF5D5555410A2D56AB",
INIT_31 => X"00AA555168A10FF803DF45FFAABDFEFAAD1554BA552E82000F7FFFFEAAA2AABD",
INIT_32 => X"A8B55552E954100004174AA00516AA10AA80155EF5D7BFDF45002A974AA08000",
INIT_33 => X"42AA10FFFFFDF55552EBDEBA5D2E80010082A97410552EBDEBAA2FBD5400F7AA",
INIT_34 => X"00000000000000000000000000000000000000000BA5D0002000552A800BA550",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0800000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(18),        -- Port A data input
DOA(0)   => data_read_a_hi_256(18),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(18),        -- Port B data input
DOB(0)   => data_read_b_hi_256(18),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_19_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"042200000000000041088001001AA00000000000000000000000500802000003",
INIT_01 => X"200048000024000000000404000000000A22000800000800004A200000000001",
INIT_02 => X"032210008DEF00400060000001C008002489E0F0004037B00010101010000000",
INIT_03 => X"0000008128000000000000000000000024001620280000000000354200004008",
INIT_04 => X"000058800004C4024024001210001054B1C822009640000E2000002604003000",
INIT_05 => X"0E010001C0400000000000000000200604000000001C04000026400000002C40",
INIT_06 => X"000000000000000001800166A84004A080000000005884020020400009907020",
INIT_07 => X"E200201C00A14080082B26208008A00900120101402240440280040840802000",
INIT_08 => X"004180261C81210031000004340000200008105428020568040213003499C006",
INIT_09 => X"00000990000000B0C30800000000086020016000000000003838000000000000",
INIT_0A => X"000000000005860000000080A000206020408000000000000454080000000000",
INIT_0B => X"00000000000040002000044000000000000000000005E0003E00004049640004",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"00000000210001D8000000000000000020009640000000000000000000000000",
INIT_0E => X"040000000000C500300080000000000000000000000000000000000000000000",
INIT_0F => X"50500101088A37034E156600D740022800EC156600D740022800D01E0412D069",
INIT_10 => X"E61700224081044914156600D7400228002C156600D7400228001098F00D0FB7",
INIT_11 => X"CC98F00D0F2DD014010046037814EA63DBB31CE7605001008C41A061F0E7D693",
INIT_12 => X"361526D600000004089E12350C0E01FF23315422BABB46FEF5019146C0800380",
INIT_13 => X"00000130AA3592000000000629C03F3E60330C00C628908214551AC900000010",
INIT_14 => X"4208D65C006070845039014460088235ACC3123E2A29148841008482A4DAC000",
INIT_15 => X"6CD4953A66BE7A5040018D8A8AD9090A1EC20A188235AC509FB50C2D0500B409",
INIT_16 => X"00000000000000000000000000000000000008C0180027000006110008404608",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"9200000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"61861861861861861A2882313054D34D301C822EE8FC31C043198028002C7441",
INIT_1B => X"84C261349A4C26130984C261309861861861A69861861861861A698618618618",
INIT_1C => X"FFFFFFFE0000026130984C26130984C26130984C26130984C26130984C261309",
INIT_1D => X"00082E97400000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"FFFFFFBFDEBA552E974105D2A801EFFFFFFFFFFFFFFFFFFFFFFFFFEAA552E954",
INIT_1F => X"55EFFFFFFFFFFFFFFFFFEFF7FBFFEAA5D2E97545FFFFC2010FFFFFFFFFFFFFFF",
INIT_20 => X"6AA0008003DF555D5157410FFFFFFFFFFFFFFDFEFF7D568A1008003DF55AAFFD",
INIT_21 => X"FFFFFFF7FBE8B55AAD16AA1000516AA005D04001EFFFFFFFFFFFFFBFDF45AAD1",
INIT_22 => X"7FC0000FF80155EFFFFFFFFEFF7D16AB55A2D57DEBA557FEAA10080402010FFF",
INIT_23 => X"2D56AB45FFFBFDEBA5D7FC0155FFFFD7410FFFFFDFEFA2D16AB55A2FFFFEAA5D",
INIT_24 => X"000000155FFFBE8B45A2D56ABEFFFFFFFE00087BC2155087BC00AAFFFBFDF45A",
INIT_25 => X"FFFFFFDEAA552E95400002095400000000000000000000000000000000000000",
INIT_26 => X"38FFFFFFFFFFFFFFFFEFF7FBFFEBA552A954105524851C7FFFFFFFFFFFFFFFFF",
INIT_27 => X"A00000E3DF6DBEF5D25D7FFFFFFFFFFFFBFDFEFEBF5F8E92552E9556DEBF1C20",
INIT_28 => X"DFEFE3F1FAF55A2D568A0000003FF7D495155428FFFFFFFFFF7FBF8FD7EBD16A",
INIT_29 => X"EFA00000002010FFFBF8FC7E3F5EAB45BEDB6FA3800556FA005504051FFFFFFF",
INIT_2A => X"56DB7DB6FFFDEAA5571C7010FF84125EFF7F1F8FC7EBD568B6DBEDF7DEBA5571",
INIT_2B => X"71C5092E3F1F8F55AADB6DB7DEBF1FAE82557FC516DEBF1D0410E3F1F8FC7AAD",
INIT_2C => X"0000000000000000000000016DE3F1EAB55BEDB6FBC7EBF5F8E10007BC516D1C",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFBFDEAA5D2A954000800154000000000000000000000",
INIT_2E => X"0552A955EFAAD1400AAFFFFFFFFFFFFBFDFEFF7FFFDEAA5D2E95410550415545",
INIT_2F => X"EFF7FFEAB45A2D56AA00002EBDFFFF7D540145FFFFFFFEFF7FBFFFFFAAD16AA0",
INIT_30 => X"E005500155EFF7FBFDFEFAAD568B55AAD568A0008003DFFF0855554AAFFFBFDF",
INIT_31 => X"ABEFFFFFFFEAA55517DE10080400010F7FBE8B55AAD16AB55F7FBFDEAA08557D",
INIT_32 => X"40010A2D56AB45A2D57DFFFF7FBFFEAA555555400F780001FFF7D16AB55A2D16",
INIT_33 => X"568A00087BD55FF5D5555410AAD56AB45AAFFFFFEFAAD168A00557BD55FFA2D5",
INIT_34 => X"00000000000000000000000000000000000000001FFAAD568B45FFFBFFF55A2D",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"1000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(19),        -- Port A data input
DOA(0)   => data_read_a_hi_256(19),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(19),        -- Port B data input
DOB(0)   => data_read_b_hi_256(19),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_20_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000003",
INIT_01 => X"A75FF80000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"14088080800008400F655001FFCFF80018FA8044000000000000011000000007",
INIT_03 => X"0000000000000000000000000000000024001660380000000000000000004FF8",
INIT_04 => X"000079800014CC02C034001600000000000000101EC0012EE0C0026E1E80F000",
INIT_05 => X"3E1FE867DFC044003902100002203F2EFC040388137C3E20C8EEC00284033CC0",
INIT_06 => X"001F0001E0020002E80020000005FEAF91D10802ABFB80000021C8010FB0F0F4",
INIT_07 => X"00040007700000000000000001080FF900160000000200C00080001840BFE538",
INIT_08 => X"09FFBFE5181606000410A4000004202AA8043E0000000000000001209244C040",
INIT_09 => X"01227FB0000000F7DF78020004011FEFE0000000002003150200008388020000",
INIT_0A => X"000000000015BE0000004000000100000100506002008C2007D5FC8000002400",
INIT_0B => X"0000000000000000000000000000000400400520000000000000000400000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000020002",
INIT_0D => X"00010000000200000020000004000100203FF6C0000000000000000000000000",
INIT_0E => X"0000000600FFC53FF001800000002004080000000000000040900005C8485380",
INIT_0F => X"8000000009A9C300020080000800000003CC0080000800000003CC0200078000",
INIT_10 => X"00800000000012963C0080000800000003CC0080000800000003CC1008000000",
INIT_11 => X"00100800004000000000066C5000020020000000800000000C2E180010002000",
INIT_12 => X"96004000000000052B0200000014200040C2829000400000000000860F987980",
INIT_13 => X"0000A4B00400000000002958000240400000000007E1B0000402000000000014",
INIT_14 => X"400004004181800000000005C5A00000200C40808000000000AF0D8008000000",
INIT_15 => X"000800020141812737DC3020100400001C19C1D80000200400000000000015D1",
INIT_16 => X"0000004010080800801810100000000000093EDFF80200000000000010010010",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"4D20400200000000000000000000000000000000000000000000000000000000",
INIT_1A => X"CB0C30C30C30C30C8192608486879E79E681C000C00E08000402241560412010",
INIT_1B => X"2190C86432190C86432190C86432CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2",
INIT_1C => X"FFFFFFFE000010C86432190C86432190C86432190C86432190C86432190C8643",
INIT_1D => X"10080402000000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"FFFFFFFFFEAA552E95400082E975FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2A954",
INIT_1F => X"0000FFFFFFFFFFFFFFFFFFFFFFFDEAA5D2A954000800001EFFFFFFFFFFFFFFFF",
INIT_20 => X"FFEBA5D2A97400FF8017410FFFFFFFFFFFFFFFFFFFFFBFDEBA552E974105D2A8",
INIT_21 => X"FFFFFFFFFFFFFEFF7FBFFEAA5D2E97545FFFFC21FFFFFFFFFFFFFFFFFFFFF7FB",
INIT_22 => X"003DF55AAFFD5400FFFFFFFFFFFFFFDFEFF7FFEAA10000417555AAD5555EFFFF",
INIT_23 => X"FFBFDFEFAAD568A0000043DF45AAFBC2010FFFFFFFFFFFFFFDFEFF7D568A1008",
INIT_24 => X"0000001EFFFFFFFFFFFFFBFDF45AAD16AA0008003DF555D51574BAFFFFFFFFFF",
INIT_25 => X"FFFFFFFEBA5D2A95410000A00000000000000000000000000000000000000000",
INIT_26 => X"C7FFFFFFFFFFFFFFFFFFFFFFFDEAA552E954000020955FFFFFFFFFFFFFFFFFFF",
INIT_27 => X"EBA552A95410552485010FFFFFFFFFFFFFFFFFFF7FBFDEBA5D2E95400140E001",
INIT_28 => X"FFFFFFFFFDFEFF7FFFFEAA5D2E95400E38A17438FFFFFFFFFFFFFFFFEFF7FBFF",
INIT_29 => X"1557DBEDF575D7FFFFFFFFFFFFBFDFEFEBF5F8E92552E9556DEBF1C21C7FFFFF",
INIT_2A => X"BF8FD7EBD16AA00000E3DF6DBEF5D2438FFFFFFFFFF7FBFDFC7EBF1E8A00080A",
INIT_2B => X"5155492FFFFFFFEFF7F1F8FD7A2D168A1008043FF6DAAFBC5028FFFFFFFFFF7F",
INIT_2C => X"000000000000000000000001FFFFFFFDFEFE3F1FAF55A2D568A0000003FF7D49",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFEBA552A95410002E820000000000000000000000",
INIT_2E => X"A552E954005D2A82145FFFFFFFFFFFFFFFFFFFFFBFDEAA5D2A954000800155FF",
INIT_2F => X"FFFFFBFDFEFF7FFFDEAA5D2E95410550415410FFFFFFFFFFFFFFDFEFF7FBFFEB",
INIT_30 => X"5EFAAD140155FFFFFFFFFF7FBFDFFFFFFBFDEBA5D2A95400A2AA974AAFFFFFFF",
INIT_31 => X"FF55A2D568A10082E955FFFFFFD7545FFFFFFFEFF7FBFFFFFAAD16AA00552A95",
INIT_32 => X"D74AAFFFBFDFEFF7FFEAB45A2D56AA00002EBDFFFF7D5400BAFFFFFDFEFF7FBF",
INIT_33 => X"568A0008003DFFF085555410F7FBFDFEFFFD568B45AAD16AA1008003DFEFAAFB",
INIT_34 => X"00000000000000000000000000000000000000001EFF7FBFDFEFAAD568B55AAD",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"01FFFFFFFFE00000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(20),        -- Port A data input
DOA(0)   => data_read_a_hi_256(20),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(20),        -- Port B data input
DOB(0)   => data_read_b_hi_256(20),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_21_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"4A302428B824900A128C090A5C1800261500213C005FE812D10420054085A202",
INIT_01 => X"081FFE3440B609703B0427F801A40B8115BC4F655300340288A40D30040E4DD8",
INIT_02 => X"0109095C30C98809800000F9FFFFFFFF149FF1FCA4C0421B182E3490DF145FE4",
INIT_03 => X"084A76341244919000099486400026523C041660BA000100CC12701015007FF8",
INIT_04 => X"000079800014CC03C075161E001118653D2408041FC004AEF000816E1C11F541",
INIT_05 => X"7E1F00F7FFC000240100004683103E7FFE02482553FC3C0204EFC25010143CC0",
INIT_06 => X"801008011010421960E339A20205FEBF8140000203FFC806C8A1C1048FF0F0E0",
INIT_07 => X"750504800680102542AD800504530FF9061E8026998E9A00402CC25BD0FFF800",
INIT_08 => X"11FBFFE04691A5A00101818A6800088228000001A044C8168480D010F200AA08",
INIT_09 => X"E85A7FF080AC70FFDF78220010841EFFE7116E144071268DFD3E4C2404010000",
INIT_0A => X"54518A8A31B7FE00040009814C089202225412115428C03BC7D7FC15025B1AB6",
INIT_0B => X"88300E20806520398C682157A493896600E24E10100DFF22FF86002020ED110C",
INIT_0C => X"28D9228D9228D9228D9228D9228D9228D99146C9146C84006309044081A001B1",
INIT_0D => X"890000403000A01282088624001201A8C43FF7C0011529904595123203040D92",
INIT_0E => X"06102C4053FFD5BFF00A04A00200602CA5200110008800444021048034004001",
INIT_0F => X"2A00263009140094D81A5040605800B506901A30406054013605620272181965",
INIT_10 => X"890A202811209062801A3040605800B506901A50406054013605604350B81282",
INIT_11 => X"3F4350B811068C00049A0A5820A3C1725A8006C0A40404D058320496C2C9C600",
INIT_12 => X"98361AC808127C454402483153A3A895BB3C1E2E820704020381702C1AAA2C4B",
INIT_13 => X"4D910CC1B154510413CC2A200501B400A40018A00C80400040D8AA288209AA21",
INIT_14 => X"0048A0141AA00418080460678A4012288463B2050302019200B00206C3590102",
INIT_15 => X"233142440470C8A9310280C0180302A01427D060022011606E800E00169C19A0",
INIT_16 => X"4010040100448008004000000E07008010003EFFFE0373056024B01118011988",
INIT_17 => X"0100401004010040100401004010040100401004010040100401004010040100",
INIT_18 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_19 => X"7E00000000000000000000000004010040100401004010040100401004010040",
INIT_1A => X"EFBEFBEFBEFBEFBEFFFFF7F7FFF3CF3CFFFFBE7FBBFDFFF7DFFCFBF08103DFDF",
INIT_1B => X"FFFFFFF7FBFDFEFF7FBFDFEFF7FBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFB",
INIT_1C => X"FFFFFFFE00003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"00080002000000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"FFFFFFFFFEBA5D2A954100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_1F => X"75FFFFFFFFFFFFFFFFFFFFFFFFFFEBA552A97400082A975FFFFFFFFFFFFFFFFF",
INIT_20 => X"FDEAA5D2E974100800155EFFFFFFFFFFFFFFFFFFFFFFFFFEAA552E95400082E9",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFDEAA5D2A95400080000000FFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"2E974105D2A80000FFFFFFFFFFFFFFFFFFFFFBFDEBA5D2E974005D2E80000FFF",
INIT_23 => X"FFFFFFFFF7FBFDEBA552A954005D2E97410FFFFFFFFFFFFFFFFFFFFFBFDEBA55",
INIT_24 => X"0000001FFFFFFFFFFFFFFFFFFFFF7FBFFEBA5D2A97400FF80174BAFFFFFFFFFF",
INIT_25 => X"FFFFFFFEBA5D2E97400000400000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2A95410000A001FFFFFFFFFFFFFFFFFFF",
INIT_27 => X"EAA552E954000020955EFFFFFFFFFFFFFFFFFFFFFFFFFEAA552E97400002E955",
INIT_28 => X"FFFFFFFFFFFFFFFFBFDEAA5D2A974101400155C7FFFFFFFFFFFFFFFFFFFFFFFD",
INIT_29 => X"97400552A80010FFFFFFFFFFFFFFFFFFF7FBFDEBA5D2E95400140E00000FFFFF",
INIT_2A => X"FFFFEFF7FBFFEBA552A95410552485038FFFFFFFFFFFFFFFFFFF7FBFDEBA552E",
INIT_2B => X"8A174AAFFFFFFFFFFFFFFFFEFF7FBFFEAA5D2E97400412497438FFFFFFFFFFFF",
INIT_2C => X"000000000000000000000001C7FFFFFFFFFFFFFFDFEFF7FFFFEAA5D2E95400E3",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974000004000000000000000000000000",
INIT_2E => X"A552E97400002E975FFFFFFFFFFFFFFFFFFFFFFFFFFEBA552A95410002E821FF",
INIT_2F => X"FFFFFFFFFFFFFFBFDEAA5D2A954000800155EFFFFFFFFFFFFFFFFFFFFFFFFDEA",
INIT_30 => X"4005D2A82010FFFFFFFFFFFFFFFFEFF7FBFDEBA552A974105D0015545FFFFFFF",
INIT_31 => X"DFEFF7FFFFEAA5D2A974005D2E82010FFFFFFFFFFFFFFDFEFF7FBFFEBA552E95",
INIT_32 => X"154AAFFFFFFFFFFFFBFDFEFF7FFFDEAA5D2E954105504154AAFFFFFFFFFFFFFF",
INIT_33 => X"BFDEBA5D2A95400A2AA974BAFFFFFFFFFF7FBFDFEFFFFFFDEBA552E974000004",
INIT_34 => X"0000000000000000000000000000000000000000155FFFFFFFFFF7FBFDFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(21),        -- Port A data input
DOA(0)   => data_read_a_hi_256(21),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(21),        -- Port B data input
DOB(0)   => data_read_b_hi_256(21),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_22_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"5290F4CDE914905A14A43D33F488243E17122300F55FEB189B343A1140548380",
INIT_01 => X"A94007B259F6A975386262000C344BA9573C6FF57B18A5FB0ABFCD3C2C5F4F0C",
INIT_02 => X"877FE30EB378008D202551040030071869D0040180AC4B685F6E26FAA0810006",
INIT_03 => X"431965109E4481D6B5AAD6875AD6AB5A1815600802888808DEA83552954D3000",
INIT_04 => X"492C0020220001010E4916C884DCD607E5EC2A344103E48003D0800023D0072C",
INIT_05 => X"0020F8882001102D620A06D683018001023D37E5088043620101179092540112",
INIT_06 => X"0803008022385AAA447A3306AA50001035B41C0A88046CAEE8C23C08E040011C",
INIT_07 => X"1EC04ED017AB5497EB923F08182E20020689B735011FBFE7BC06260294401CA8",
INIT_08 => X"4A00401D4425ADA9035BE19C8F9442A8801200F4C9D7AC8093A051727B2AC349",
INIT_09 => X"50020040E48D50080002B00A0C00801014541E9504703680017F6CB405070015",
INIT_0A => X"54538A8A738041C23020131A80CFDFF3FE509A907C6AC050402204090090319A",
INIT_0B => X"40050220103D2A512C6A8C4F0011550008E06E000140009A000000424DE61920",
INIT_0C => X"A81C2A81C2A81C2A81C2A81C2A81C2A81C9540E1540E001400006100003202D0",
INIT_0D => X"8B2940D0E153941A8B1A262CA542A9A8D6C0010A101628013456520CA09281C2",
INIT_0E => X"80410089180008800143D83888281A2034A85014280A14050A01509E05085449",
INIT_0F => X"000C26706B3C189CD84ACD20B03001E387D04AC560B02401E387E1028AC04500",
INIT_10 => X"458870201570B036C04AC560B03001E387D04ACD20B02401E387E24708E7E242",
INIT_11 => X"044708E7E1C20A0106EA167C84EBF052A8E010C0180606E86C3F459DC08DA902",
INIT_12 => X"98225189980254CDEC22A98032A22C50EAC462030A01800407C2700C2ACA2C0F",
INIT_13 => X"4A99BCC1154C258012D86F601A2E49003400138C0DA2443A208AA612C0096C37",
INIT_14 => X"90E16025483C1E0C0006B085CEC03858958D15310201015504B512044A313300",
INIT_15 => X"6B0469512C6FC01A1421006028038720640310643858162712020B001AA415F2",
INIT_16 => X"11044110445E22022365034A8EA754008004C0200323001182122548881649D1",
INIT_17 => X"1044110441104411044110441104411044110441104411044110441104411044",
INIT_18 => X"0401004010040100401004010040100401004010040100401004411044110441",
INIT_19 => X"7D05122890000000003FFFFFFFF9004010040100401004010040100401004010",
INIT_1A => X"E79E79E79E79E79EFFDFF7F5F777DF7DF7DF7EFF7BFA3FC7DF7AF5BF7EFDF7DF",
INIT_1B => X"9FCFE7F3F9FCFE7F3F9FCFE7F3F9E79E79E79E79E79E79E79E79E79E79E79E79",
INIT_1C => X"FFFFFFFE00000FE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F",
INIT_1D => X"10000000000000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"FFFFFFFFFEBA5D2E974000800021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_1F => X"21FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E954000004001FFFFFFFFFFFFFFFFF",
INIT_20 => X"FFEBA552A97400002A801FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2A9541008040",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFEBA552A97400082A975FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"2E95400082E975FFFFFFFFFFFFFFFFFFFFFFFFFFEAA552E95410002A955FFFFF",
INIT_23 => X"FFFFFFFFFFFFFFEAA552E95400002E975EFFFFFFFFFFFFFFFFFFFFFFFFFEAA55",
INIT_24 => X"000000000FFFFFFFFFFFFFFFFFFFFFFFDEAA5D2E97410080015545FFFFFFFFFF",
INIT_25 => X"FFFFFFFEBA5D2E97410080002000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974000004001FFFFFFFFFFFFFFFFFFF",
INIT_27 => X"EBA5D2A95410000A001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2A954000804021",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFEBA552A97400082E821FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"95410082A975EFFFFFFFFFFFFFFFFFFFFFFFFFEAA552E97400002E955FFFFFFF",
INIT_2A => X"FFFFFFFFFFFDEAA552E954000020955C7FFFFFFFFFFFFFFFFFFFFFFFFEAA552E",
INIT_2B => X"0015545FFFFFFFFFFFFFFFFFFFFFFFDEAA5D2A974001C24975C7FFFFFFFFFFFF",
INIT_2C => X"00000000000000000000000000FFFFFFFFFFFFFFFFFFFFFBFDEAA5D2A9741014",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800020000000000000000000000",
INIT_2E => X"A5D2A954000800021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974000004001FF",
INIT_2F => X"FFFFFFFFFFFFFFFFFEBA552A95410002E821FFFFFFFFFFFFFFFFFFFFFFFFFFEB",
INIT_30 => X"400002E975EFFFFFFFFFFFFFFFFFFFFFFFFFEAA552A97400082A801FFFFFFFFF",
INIT_31 => X"FFFFFFFBFDEAA5D2E95410082E955EFFFFFFFFFFFFFFFFFFFFFFFFDEAA552E97",
INIT_32 => X"17545FFFFFFFFFFFFFFFFFFFFFBFDEAA5D2A95400080015545FFFFFFFFFFFFFF",
INIT_33 => X"BFDEBA552A974105D0015555FFFFFFFFFFFFFFFFFFF7FBFDEBA5D2A974005504",
INIT_34 => X"0000000000000000000000000000000000000000010FFFFFFFFFFFFFFFFEFF7F",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"01FFFFFFFFE00000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(22),        -- Port A data input
DOA(0)   => data_read_a_hi_256(22),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(22),        -- Port B data input
DOB(0)   => data_read_b_hi_256(22),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_23_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"EF20906D902424807BC8241BC81801B97D38AD3C0800103362A6741C80A12A02",
INIT_01 => X"001FFF8409F089003B4422000D80C80106804A7951C5B9D1C828043EA28838F9",
INIT_02 => X"073B8858218C2C50801000F9FFEFF8E72CA7F5FC2E048026496834D84721DFE0",
INIT_03 => X"2C4360101A4001001005080400401420350016E0BB222341C312000014006FF8",
INIT_04 => X"00017B810015DC03D034201E14000036486008101FC0002EE006297E1C05F561",
INIT_05 => X"7E1F02FFFFC80100004044800080BEFFFC0248005FFC3C18A5FFC2444484BCC0",
INIT_06 => X"4082040800000811224DE0A00005FFBF8000000003FF810640A1C0008FF2F0E1",
INIT_07 => X"D1D72040048D00388387D03D0E591FFD201F862691DFBE077C2BC45B40FFE458",
INIT_08 => X"1FFBFFEC440501A5604B31062356282AA84200D12342113EDC40000004582800",
INIT_09 => X"A890FFF0002023FFDF79000000000EFFE309606020008005FC00000040200000",
INIT_0A => X"000000000037FF50010103134CAFDF03BA18000F39A0106F87D7FA84024B0225",
INIT_0B => X"88300C48907120AC81083315A493886640030010540DFF20FF8610302409000C",
INIT_0C => X"10C1010C1010C1010C1010C1010C1010C10086080860840063090442A18001B1",
INIT_0D => X"0000280600020040030090000012A500003FF7E08181119A41C1443243050C10",
INIT_0E => X"06542C7043FFD5FFF00A04BC010A7724B1000080004000200004150030010004",
INIT_0F => X"B2080290C2909080A872BC4FC8500054840072FC0FC8440054840200705F9861",
INIT_10 => X"0C8220180F1082E00072FC0FC8500054840072BC4FC84400548402214A380380",
INIT_11 => X"19214A380344920080B21810240AB182EB37C380B40800707011001B43253EE5",
INIT_12 => X"0019CE4000026C00C00042BD4149067465910640A0050C060A0028063672A000",
INIT_13 => X"4D801800CCB050001344060211629580B80022480A444111706658280009A203",
INIT_14 => X"944CB232D6D0100C040250200845132C10BE200403018061101A220339C80000",
INIT_15 => X"402102A5493B8E287E03808480060E40C83C1405132C90742E408D0082140820",
INIT_16 => X"0080200802000100100000000000004002403EFFF8002385F034901019465001",
INIT_17 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_18 => X"8020080200802008020080200802008020080200802008020080200802008020",
INIT_19 => X"0000000000000000000000000000080200802008020080200802008020080200",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000004000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFE00000000000000000000000000000000000000000000000000000000",
INIT_1D => X"10080400000000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"FFFFFFFFFEBA5D2E974100000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_1F => X"21FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100004021FFFFFFFFFFFFFFFFF",
INIT_20 => X"FFEBA5D2E954000800001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9740008000",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E954000004001FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"2A954100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2A954100000021FFFFF",
INIT_23 => X"FFFFFFFFFFFFFFEBA5D2A954100800021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_24 => X"0000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA552A97400002A801FFFFFFFFFFFF",
INIT_25 => X"FFFFFFFEBA5D2E97410080400000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800021FFFFFFFFFFFFFFFFFFF",
INIT_27 => X"EBA5D2E974000004001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100004021",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFEBA5D2E954000800001FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"954100004021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2A954000804021FFFFFFF",
INIT_2A => X"FFFFFFFFFFFFEBA5D2A95410000A001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2A",
INIT_2B => X"2E821FFFFFFFFFFFFFFFFFFFFFFFFFFEBA552A97410080E001FFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA552A9740008",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804000000000000000000000000",
INIT_2E => X"A5D2E974100000021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800021FF",
INIT_2F => X"FFFFFFFFFFFFFFFFFEBA5D2E974000004001FFFFFFFFFFFFFFFFFFFFFFFFFFEB",
INIT_30 => X"4000800021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E954000804021FFFFFFFFF",
INIT_31 => X"FFFFFFFFFFEBA552A954100004001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2A95",
INIT_32 => X"821FFFFFFFFFFFFFFFFFFFFFFFFFFEBA552A95410002E821FFFFFFFFFFFFFFFF",
INIT_33 => X"FFFEAA552A97400082A801EFFFFFFFFFFFFFFFFFFFFFFFFFEAA552A97410002A",
INIT_34 => X"00000000000000000000000000000000000000001EFFFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"01FFFFFFFFE00000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(23),        -- Port A data input
DOA(0)   => data_read_a_hi_256(23),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(23),        -- Port B data input
DOB(0)   => data_read_b_hi_256(23),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_24_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100600007FFF000080108004000800020000840041000080808",
INIT_02 => X"172A00D000EF8210000000F9FFEFF8E7240FF1FC224087B1000639401D005FC0",
INIT_03 => X"00003A2E200811000000000400000000340016603A0000004860400014006FFF",
INIT_04 => X"000079800014CC03C034001E04010850300000101FC0002EE000006E1C00F500",
INIT_05 => X"3E1F0067FFC000000000000000003E2FFC024800137C3C0000EFC00000003CC0",
INIT_06 => X"000000000000001123820AA00005FEBF8000000003FF80000021C0000FF0F0E0",
INIT_07 => X"E600084002040A10812A000500590FF9001F95406A8000037230C01840FFE000",
INIT_08 => X"01FBFFEC4695A501604A000C7585080002C200408102F16C0184800026C92C10",
INIT_09 => X"A8107FF0000000FFDF78000000000EFFE001600000000005FC00000000000000",
INIT_0A => X"000000000037FF4000000AA0354000019C4000012800002387D7F804024B0224",
INIT_0B => X"88300C0081408000800001002482886600020010100DFA20FF8600000000000C",
INIT_0C => X"00C1000C1000C1000C1000C1000C1000C1000608006084006301044081800121",
INIT_0D => X"00000000900160000000000000000000003FF7C0010101904181003003000C10",
INIT_0E => X"16100C4043FFD5BFF00004100000000411000000000000000000040030000000",
INIT_0F => X"3A0421080012302010049400086C022004200494000878022004120270599965",
INIT_10 => X"C19240300081406100049400086C022004200494000878022004124819081840",
INIT_11 => X"2348190814C09C01010400132100106836001504240E01040051200200D06410",
INIT_12 => X"202CD680C0100010408240BD80008983596CD86EA84104060503C0B000020250",
INIT_13 => X"0002090164F40086000082062C1B6600BC000C300818044000B27A0043000041",
INIT_14 => X"110002577FE4080C08010842180C40018545BBA00301808A0810C0059AD01802",
INIT_15 => X"4820C04100852B931F00800010081980B042D2044001850ED8808F00050A002C",
INIT_16 => X"0000000000000000000000000000000000003EFFF80037046031E0110001100A",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"9900000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"EFBE7BE7BE7BE7BEC99E61848655D75D7FCB42BBABDB9F3044CB35CF612B4441",
INIT_1B => X"83C1E0F0783C1E0F0783C1E0F07BEFBEFBEF9E79E79E79E79E7BEFBEFBEFBEFB",
INIT_1C => X"FFFFFFFE000001E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F07",
INIT_1D => X"10080402000000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"FFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_1F => X"01FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800021FFFFFFFFFFFFFFFFF",
INIT_20 => X"FFEBA5D2E974100000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741000000",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974100004021FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"2E974000800021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974000004001FFFFF",
INIT_23 => X"FFFFFFFFFFFFFFEBA5D2E974000800001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_24 => X"0000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E954000800001FFFFFFFFFFFF",
INIT_25 => X"FFFFFFFEBA5D2E97410080402000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFF",
INIT_27 => X"EBA5D2E974100800021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800021",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFEBA5D2E974100000001FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974000004001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100004021FFFFFFF",
INIT_2A => X"FFFFFFFFFFFFEBA5D2E974000004001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E",
INIT_2B => X"00001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E954000800021FFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9540008",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804020000000000000000000000",
INIT_2E => X"A5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FF",
INIT_2F => X"FFFFFFFFFFFFFFFFFEBA5D2E974100800021FFFFFFFFFFFFFFFFFFFFFFFFFFEB",
INIT_30 => X"4100000021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100000001FFFFFFFFF",
INIT_31 => X"FFFFFFFFFFEBA5D2E974000004021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E97",
INIT_32 => X"021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974000004001FFFFFFFFFFFFFFFF",
INIT_33 => X"FFFEBA5D2E954000804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E954000004",
INIT_34 => X"00000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(24),        -- Port A data input
DOA(0)   => data_read_a_hi_256(24),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(24),        -- Port B data input
DOB(0)   => data_read_b_hi_256(24),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_25_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100200002000000080100004000000020000800041000080808",
INIT_02 => X"1000218000000800000000F9FFEFF8E738FFF1FC20400400000004455A375FE0",
INIT_03 => X"00002000000001000000000400000000340016623A0000004000000014006FFF",
INIT_04 => X"924279824C94CC1BE0B4001F20000000020380401FE0082EF000106E1C00F500",
INIT_05 => X"3E1F0067FFE048002582800100523E2FFE024820137C3C0040EFE02000003CE4",
INIT_06 => X"821B0821B8019819200020200005FEBF81C1002203FF80000021C1140FF8F0E0",
INIT_07 => X"00040000000000000000000500590FF9001F0000000000033020C01840FFFC78",
INIT_08 => X"01FBFFFD0004000100502000011400000282004001020000000001009015C000",
INIT_09 => X"B8DA7FF8004000FFDF7C062031863EFFF75D78004001010DFC00002005010000",
INIT_0A => X"000000000037FFC00602000000000001980400002800032387D7FE94FBEF2B2C",
INIT_0B => X"88300C0080400000800001002486887600020110100DFA20FF8603000000000C",
INIT_0C => X"00C1000C1000C1000C1000C1000C1000C10006080060840077330C4889CC2925",
INIT_0D => X"00000000000000000000000000002500003FF7C0010101904189003003000C10",
INIT_0E => X"06140C6043FFD5BFF00A04B80608003CB120C110608830445821140134120800",
INIT_0F => X"02000000000200200000900000400200000000900000400200000200701E1861",
INIT_10 => X"0002000000010000000090000040020000000090000040020000000008080000",
INIT_11 => X"0000080800008000000000010100000022000000040000000040000000002400",
INIT_12 => X"0000420000000010000040318020000041000001000244000000008008000010",
INIT_13 => X"0002000004100000000080000002040040000000001000400002080000000040",
INIT_14 => X"0100000042000010002000001000400000042000040200000000400008400000",
INIT_15 => X"0030800000010800000000C0A000000000400000400000040800000000000004",
INIT_16 => X"41104451044C82082068C0200000008014023EFFFC0063046020801000001000",
INIT_17 => X"1104411044110441104411044110441104411044110441104411044110441104",
INIT_18 => X"1044110441104411044110441104411044110441104411044110441104411044",
INIT_19 => X"A080800002FFFFFFFFFFFFFFFFFC110441104411044110441104411044110441",
INIT_1A => X"41041249041249042824014C48569A69AFEE8A252865AA3168A4CBDF860EC15D",
INIT_1B => X"58AC56231188C46231188C462312492492492492492492492490410410410410",
INIT_1C => X"FFFFFFFE00002C562B158AC562B158AC562B158AC562B158AC562B158AC562B1",
INIT_1D => X"10080400000000000000000000000000000000000000000000000001FFFFFFFF",
INIT_1E => X"FFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_1F => X"01FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFF",
INIT_20 => X"FFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008040",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800021FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"2E974100000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800001FFFFF",
INIT_23 => X"FFFFFFFFFFFFFFEBA5D2E974100000021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_24 => X"0000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100000001FFFFFFFFFFFF",
INIT_25 => X"FFFFFFFEBA5D2E97410080400000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFF",
INIT_27 => X"EBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974100800001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800021FFFFFFF",
INIT_2A => X"FFFFFFFFFFFFEBA5D2E974100800021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E",
INIT_2B => X"00001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100000021FFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741000",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804000000000000000000000000",
INIT_2E => X"A5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FF",
INIT_2F => X"FFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEB",
INIT_30 => X"4100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFF",
INIT_31 => X"FFFFFFFFFFEBA5D2E974100800001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E97",
INIT_32 => X"021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800021FFFFFFFFFFFFFFFF",
INIT_33 => X"FFFEBA5D2E974100000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800",
INIT_34 => X"00000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"01FFFFFFFFE00000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(25),        -- Port A data input
DOA(0)   => data_read_a_hi_256(25),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(25),        -- Port B data input
DOB(0)   => data_read_b_hi_256(25),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_26_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"E9264EAB20190CA3BA4997AA9002AE9C001006B0778015CFA17E0811039879C7",
INIT_01 => X"F1FFF9BB1F773C7F9BB07DFFFDD863FC5FFF3FEFFBBF9FFB22FFFBC7B9F30686",
INIT_02 => X"1B33188302E708180F6FFBFFFFCFFFFF9C7FF7FC24350B99082400001D00DFD8",
INIT_03 => X"4A53D958C50000DCE7366303739CD98C27C57EF57980014F271807E3C9E9CFF8",
INIT_04 => X"DBFAFBD7FB1CDEBEF1BE17F7AC88042787FBFFF8FEE9FF7EE6F4C0EE1FFAF869",
INIT_05 => X"BE1FFD67DFFEFFBDA7F7FED508707E2EFEBF6FFEB37C3FF302EEEDFF9B487CF6",
INIT_06 => X"75F7275F7CAC98E261EDF0253C7FFFEF87C74E8CCFFBB6FF70E1FE61FFBDF0FE",
INIT_07 => X"73840C07783060C72DF7D828912E6FFB80162776F3BFB7077E82255E40BFEEBA",
INIT_08 => X"69FFBFE43C872321367036163F1C0820A3063F460D1AEFC000060042648C4181",
INIT_09 => X"FB967FBD13D981F7DF7D7E6171AF3FEFE8A3E679FAC1FD1FFFBEB000763A8447",
INIT_0A => X"6AED1D1DAD7FBE7D67D7F3BB79CFFB83BF14EC1E7D7300B017F5FFE6FBEF73BE",
INIT_0B => X"99F51EDDCDEBCFF589807B70AD9A99EE7583F931109FFE33FF8E3FDFDAF64A3C",
INIT_0C => X"C0D78C0D78C0D78C0D78C0D78C0D78C0D7A606BC606B8C56F7730ECCDBDF1521",
INIT_0D => X"1D406B9EC20181CC1F73F87501DED3409BFFFEFFEBF341B867D3683A03A40F78",
INIT_0E => X"86D70CE04FFFFF3FF1F5F5475BD7F72E4D75EBFAF5FD7AFEFDFFAF59B6FF28FE",
INIT_0F => X"020007C040101480807D17B0004001F804007D17B0004001F8040212F35FFC6D",
INIT_10 => X"700200001DC00068007D17B0004001F804007D17B0004001F804006F60081400",
INIT_11 => X"206F60081800800007B000102C0801FB02683800040007700011801003DE050A",
INIT_12 => X"403E232130207080D012CEFF41008D188D502100B02004000F01900039020040",
INIT_13 => X"0E101A01F21A2C40039006823F80048100003F0008004D8100F90D162001C803",
INIT_14 => X"B604027F020A07400007C040085581019D602451500001EC00100247C4642608",
INIT_15 => X"CC3F02010EA40EA00020C830100F0D000022180581019F40084800001F100020",
INIT_16 => X"EBFAFEFFBFEFDFDDFE7DD87FEFF7FF796FFFFFDFFC017FEFFD7E841001D8197D",
INIT_17 => X"BFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAF",
INIT_18 => X"FAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFE",
INIT_19 => X"EDB5C88646FFFFFFFFFFFFFFFFFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEB",
INIT_1A => X"61861A69A6986186EBCAF55357E1C71C751D6C56F3D247859B3214FA76953F86",
INIT_1B => X"84C26130984C26130984C2613098618618618618618618618618618618618618",
INIT_1C => X"FFFFFFFE0000026130984C26130984C26130984C26130984C26130984C261309",
INIT_1D => X"10080400000000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"FFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_1F => X"21FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFF",
INIT_20 => X"FFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008040",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFF",
INIT_23 => X"FFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_24 => X"0000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFF",
INIT_25 => X"FFFFFFFEBA5D2E97410080400000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFF",
INIT_27 => X"EBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFF",
INIT_2A => X"FFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E",
INIT_2B => X"04021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804000000000000000000000000",
INIT_2E => X"A5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FF",
INIT_2F => X"FFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEB",
INIT_30 => X"4100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFF",
INIT_31 => X"FFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E97",
INIT_32 => X"001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFF",
INIT_33 => X"FFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804",
INIT_34 => X"00000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(26),        -- Port A data input
DOA(0)   => data_read_a_hi_256(26),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(26),        -- Port B data input
DOB(0)   => data_read_b_hi_256(26),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_27_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"00080A40000A41248002029000050A088000008242A0004404480002000A1155",
INIT_01 => X"F1FFF1C11F781C129C107DFFFE0860941E81258CA2B71C2220EC1B86E1A00002",
INIT_02 => X"4000002100000014400FF6FFFF0FFFFF8007F1FC211100014200800000887FC0",
INIT_03 => X"0842D85841000098C63061026318C18404C459757000015F00088BE3C0618FF8",
INIT_04 => X"DBEAE5D6D91C2EBCE1B21EA72C00000007FBE7C8F8E9EF79E6D440E91FDAE061",
INIT_05 => X"B91FF9671FE6B68984B5BCE408347E28FEBF6FEEB3723F7102E8EDBF8A4872F6",
INIT_06 => X"3573A357308418E40000D4113C7FFE4F86064C8DDFE3B6FF50D1FC61DE39C8FC",
INIT_07 => X"00000A20083060C00C81882A008C6FF880060424B39FB6037F00051C003FE04A",
INIT_08 => X"61FA3FE4010440410844060001040A00002200460D1A06000005040000001080",
INIT_09 => X"EB027E390A4881C7BEFC5F6171CE2F8FE823E778DAC16C1FFBBC900031589547",
INIT_0A => X"03813030213C3E2D62D6E21259CFDB039E806C024531008017C1F826FFEF41FE",
INIT_0B => X"9AB55F0DEFABC705488069302DBA98EAB582D835109FFC31FFAEAFCFDAF4423D",
INIT_0C => X"40C3440C3440C3440C3440C3440C3440C3C2061A2061AD46FF730E5CCBCD5521",
INIT_0D => X"0C407D1F820101441DA3A8310198C34089BFF8DD6B7941BC63F1683803C00E34",
INIT_0E => X"5710AE4047FFD23FF315D54358D593474955AB6AD5B56ADAB5FAAE58B2F628EA",
INIT_0F => X"020007C0400004C080791290004001D80001791290004001D8000210F1587971",
INIT_10 => X"300200001DC0000801791290004001D80001791290004001D800012F60080400",
INIT_11 => X"202F60080800800007B000000E0801BB020828000400077000008210035E0408",
INIT_12 => X"40BA2220202070801010C6F1410085188D500100102004000F01900031000060",
INIT_13 => X"0E100205D2120840039000813F80040100003F0000000F8100E909042001C800",
INIT_14 => X"3E04007F020201400007C040001781011D602040500001EC0000005744440408",
INIT_15 => X"C43F02000EA40EA000004810100F0D000020080781011F40080800001F100000",
INIT_16 => X"AB6ADAB6BDE75ED5EC71385FC2512E3565BBBF1FFC00636EED7E841000D81924",
INIT_17 => X"B6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6AD",
INIT_18 => X"6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADA",
INIT_19 => X"A471688747FFFFFFFFFFFFFFFFFAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB",
INIT_1A => X"0020800000000000780401CBC840000005243885A04012072A1810DA84002104",
INIT_1B => X"5028140201008040201008040200000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFE000028140A05028140A05028140A05028140A05028140A05028140A0",
INIT_1D => X"10080400000000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"FFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_1F => X"01FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFF",
INIT_20 => X"FFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008040",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFF",
INIT_23 => X"FFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_24 => X"0000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFF",
INIT_25 => X"FFFFFFFEBA5D2E97410080400000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFF",
INIT_27 => X"EBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFF",
INIT_2A => X"FFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E",
INIT_2B => X"04021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804000000000000000000000000",
INIT_2E => X"A5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FF",
INIT_2F => X"FFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEB",
INIT_30 => X"4100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFF",
INIT_31 => X"FFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E97",
INIT_32 => X"021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFF",
INIT_33 => X"FFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804",
INIT_34 => X"00000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"01FFFFFFFFE00000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(27),        -- Port A data input
DOA(0)   => data_read_a_hi_256(27),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(27),        -- Port B data input
DOB(0)   => data_read_b_hi_256(27),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_28_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"02200AA400180030808802A900002A08001280A08A801044104A1000001818C3",
INIT_01 => X"50A00011460214428114180000882214413D0A71592A01D92213D28005210202",
INIT_02 => X"1444428102100884000AA30200000000C1000401041108404400022220800000",
INIT_03 => X"461080404900000C6314A900318C52A40051081000888806108802A141288001",
INIT_04 => X"00800040110102000902002000888400081045A8A00003C00000500000080008",
INIT_05 => X"0000000000024CA0A0101800032000400000000B800000014000000B08180000",
INIT_06 => X"10280102802C0240041000011428004022220024440013511000013510000000",
INIT_07 => X"0804420009122448451020100020400080002041000000008000010400000880",
INIT_08 => X"2800000140200808021006108010422AAA800022448902849220114009224081",
INIT_09 => X"01C800004080A0000002480B04008100011000088800081002C19020150B0013",
INIT_0A => X"56D29A9A52800004004070208000000040006408001100105000020000001800",
INIT_0B => X"00040024440245400082D0220800008010001020458000010000040D96104210",
INIT_0C => X"50160501605016050160501605016050160280B0280B00120008430660210014",
INIT_0D => X"054001884200810C1631181500CA60400B4008072020500002002C0040010360",
INIT_0E => X"104420A00C000200005000010040A0020CC000200010000800920040804020A6",
INIT_0F => X"0000000000001400000102900000002800000102900000002800001001802104",
INIT_10 => X"3000000000000048000102900000002800000102900000002800000020000400",
INIT_11 => X"0000200008000000000000002800000100082800000000000001800000020008",
INIT_12 => X"4000202020200000901005480000000800000100102000000000000009000000",
INIT_13 => X"0000120002020840000004800080000100000000000048800001010420000002",
INIT_14 => X"A200000800020140000000000050800008000040500000000000024004040408",
INIT_15 => X"840A000002000000000048100000000000020800800008000008000000000000",
INIT_16 => X"8020080210810840861CD33548542A10209D4100000010200400000000880035",
INIT_17 => X"0200802008020080200802008020080200802008020080200802008020080200",
INIT_18 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_19 => X"40A0C22E10000000000000000000020080200802008020080200802008020080",
INIT_1A => X"08208208208208200360D4141D630C30C7788440B044280091A5CB03D01BD89A",
INIT_1B => X"582C16030180C06030180C060302082082082082082082082082082082082082",
INIT_1C => X"FFFFFFFE00002C160B0582C160B0582C160B0582C160B0582C160B0582C160B0",
INIT_1D => X"10080400000000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"FFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_1F => X"01FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFF",
INIT_20 => X"FFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008040",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFF",
INIT_23 => X"FFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_24 => X"0000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFF",
INIT_25 => X"FFFFFFFEBA5D2E97410080400000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFF",
INIT_27 => X"EBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFF",
INIT_2A => X"FFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E",
INIT_2B => X"04001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804000000000000000000000000",
INIT_2E => X"A5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FF",
INIT_2F => X"FFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEB",
INIT_30 => X"4100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFF",
INIT_31 => X"FFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E97",
INIT_32 => X"001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFF",
INIT_33 => X"FFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804",
INIT_34 => X"00000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"01FFFFFFFFE00000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(28),        -- Port A data input
DOA(0)   => data_read_a_hi_256(28),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(28),        -- Port B data input
DOB(0)   => data_read_b_hi_256(28),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_29_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"79964E4BA01DACAB9E659792D00AAE160002829C7FDFEFCEE97C2815039D70C3",
INIT_01 => X"50BFF9AB0775343F9AB01DF80D5821FC0FFF3FEFD1AF9FF1207FFBC7B9720586",
INIT_02 => X"0B33180300E700080F6AAA7BFFC007189C7FF2FC003503980A0000001D00DFD8",
INIT_03 => X"0401D940CD0000C8421A2B03210868AC23403E903900010E271006A148A0C000",
INIT_04 => X"49B87A417315D20A313E17F1800000058013DDF8BE21F36E02F0D06E03E8F800",
INIT_05 => X"3E00FC67C03A4D9C87525E5101603E6E023D27DA937C03E340EE25CB9B483C12",
INIT_06 => X"50B5050B540C004261EDE025142DFFE003C30E0447F877F930203E213F8CF01E",
INIT_07 => X"73800407781020476467D008910A4FFB80100332D1AE93059282215E40800678",
INIT_08 => X"21FF80003C832320342036063F08000001063F42050AEB4000221000248C0180",
INIT_09 => X"51547F8C1111A0F041056A0100A11FE000916249A800B915FE82B02052290002",
INIT_0A => X"2AAD1515AD5780540541619968C76980E914E4163D53002017F405C409A42A9A",
INIT_0B => X"014002D445624DB481806A6288100184500171200085FE030000157FDF124A10",
INIT_0C => X"D0068D0068D0068D0068D0068D0068D006A68034680300021410028450530014",
INIT_0D => X"15402B0E8201018C1561E855008C50401B7FFE27A0B2500806522C0A40A50268",
INIT_0E => X"928324400DFFFF0001F1F0050342D42A086040B02058102C48970541944B20FA",
INIT_0F => X"0000000000101480000507B00000002804000507B000000028040212034FAD28",
INIT_10 => X"7000000000000068000507B00000002804000507B00000002804004020001400",
INIT_11 => X"0040200018000000000000102C0000410068380000000000001180000082010A",
INIT_12 => X"4004212130200000D0120ED64000080800002100B02000000000000009020040",
INIT_13 => X"00001A00220A2C4000000682008000810000000008004D800011051620000003",
INIT_14 => X"B6000208000A0740000000000855800088000451500000000010024084242608",
INIT_15 => X"8C0F0001020000000020C8300000000000021805800088000048000000000020",
INIT_16 => X"C0B02C4B12C989489418D13FE7F3FFD8BADB7FC004012CA5141600000198087D",
INIT_17 => X"0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02",
INIT_18 => X"B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C",
INIT_19 => X"FEA0C00602FFFFFFFFFFFFFFFFFC0B02C0B02C0B02C0B02C0B02C0B02C0B02C0",
INIT_1A => X"FBAEBAEBAEBAEBAEFFFFF7E7EFBFFFFFFAEF3E7E5BB9FFF7DFF9E3F08843FFDF",
INIT_1B => X"FDFEFF7FBFDFEFF7FBFDFEFF7FBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBE",
INIT_1C => X"FFFFFFFE00003EFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FB",
INIT_1D => X"10080400000000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"FFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_1F => X"01FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFF",
INIT_20 => X"FFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008040",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFF",
INIT_23 => X"FFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_24 => X"0000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFF",
INIT_25 => X"FFFFFFFEBA5D2E97410080400000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFF",
INIT_27 => X"EBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFF",
INIT_2A => X"FFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E",
INIT_2B => X"04001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804000000000000000000000000",
INIT_2E => X"A5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FF",
INIT_2F => X"FFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEB",
INIT_30 => X"4100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFF",
INIT_31 => X"FFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E97",
INIT_32 => X"001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFF",
INIT_33 => X"FFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804",
INIT_34 => X"00000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(29),        -- Port A data input
DOA(0)   => data_read_a_hi_256(29),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(29),        -- Port B data input
DOB(0)   => data_read_b_hi_256(29),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_30_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"FD00000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"E79E79E79E79E79EEBFEF5D7D7F7DF7DFFDFFEFFFBFE7F87DFFEFFBF77BFFFDF",
INIT_1B => X"9FCFE7F3F9FCFE7F3F9FCFE7F3F9E79E79E79E79E79E79E79E79E79E79E79E79",
INIT_1C => X"FFFFFFFE00000FE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F",
INIT_1D => X"10080400000000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"FFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_1F => X"01FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFF",
INIT_20 => X"FFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008040",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFF",
INIT_23 => X"FFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_24 => X"0000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFF",
INIT_25 => X"FFFFFFFEBA5D2E97410080400000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFF",
INIT_27 => X"EBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFF",
INIT_2A => X"FFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E",
INIT_2B => X"04001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804000000000000000000000000",
INIT_2E => X"A5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FF",
INIT_2F => X"FFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEB",
INIT_30 => X"4100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFF",
INIT_31 => X"FFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E97",
INIT_32 => X"001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFF",
INIT_33 => X"FFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804",
INIT_34 => X"00000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(30),        -- Port A data input
DOA(0)   => data_read_a_hi_256(30),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(30),        -- Port B data input
DOB(0)   => data_read_b_hi_256(30),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_31_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"129000008004A00804A40000400800020000000C005FEA005800200400050100",
INIT_01 => X"A15FF18019700810180065FFFC0040801E80258CA2951C2200EC0906A0804140",
INIT_02 => X"0000000000000011000550FDFF0FFFFF0007F1FC200000011000000000205FC0",
INIT_03 => X"08425818000000908428C0024210A30004045060302223490002014280410FF8",
INIT_04 => X"DB6A618248140C18E0B016872400000007EBA24058E1ECA8E2D400681FD0E061",
INIT_05 => X"381FF8671FE01009048084C400103E28FE3F6FE513703F7000E8E5B4825030F6",
INIT_06 => X"00130001300018A00000D0002855FE0F84040C088BE3E4AE40C1FD04CE38C0FC",
INIT_07 => X"000008800020408008818838000C2FF800060424B39FB6037E000418003FE008",
INIT_08 => X"41FA3FE400040001004000000104088000020044091204000004000000000000",
INIT_09 => X"E8027E38004801C79E7C162231862E8FE00166704041240DF93D000000000004",
INIT_0A => X"0000000000343E002202021259CFDB039E0008024520000047C1F804FBEF01BE",
INIT_0B => X"88310E08812982050800A9102492986200824810110DFC30FF86036249E4002C",
INIT_0C => X"00C1000C1000C1000C1000C1000C1000C18006080060840477330C4889CC0121",
INIT_0D => X"08006816800100400902A0200110810080BFF0C80111019861D1403803800C10",
INIT_0E => X"06100C4043FFD03FF101D4000800130401808100408020401020041830120848",
INIT_0F => X"020007C04000008080781000004001D00000781000004001D0000200F0185861",
INIT_10 => X"000200001DC0000000781000004001D00000781000004001D000002F40080000",
INIT_11 => X"202F40080000800007B00000040801BA020000000400077000000010035C0400",
INIT_12 => X"003A0200000070800000C231410085108D500000000004000F01900030000040",
INIT_13 => X"0E100001D0100000039000003F00040000003F000000050100E808000001C800",
INIT_14 => X"14040077020000000007C0400005010115602000000001EC0000000740400000",
INIT_15 => X"403502000CA40EA000000000100F0D000020000501011740080000001F100000",
INIT_16 => X"01004010044602002061004A820104809402BE1FFC006304E036841000501900",
INIT_17 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_18 => X"0040100401004010040100401004010040100401004010040100401004010040",
INIT_19 => X"0001000802FFFFFFFFFFFFFFFFF8100401004010040100401004010040100401",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFE00000000000000000000000000000000000000000000000000000000",
INIT_1D => X"10080400000000000000000000000000000000000000000000000001F007FFFF",
INIT_1E => X"FFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_1F => X"01FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFF",
INIT_20 => X"FFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008040",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFF",
INIT_23 => X"FFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_24 => X"0000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFF",
INIT_25 => X"FFFFFFFEBA5D2E97410080400000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFF",
INIT_27 => X"EBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFF",
INIT_2A => X"FFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E",
INIT_2B => X"04001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804000000000000000000000000",
INIT_2E => X"A5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FF",
INIT_2F => X"FFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEB",
INIT_30 => X"4100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFF",
INIT_31 => X"FFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E97",
INIT_32 => X"001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFF",
INIT_33 => X"FFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804",
INIT_34 => X"00000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(31),        -- Port A data input
DOA(0)   => data_read_a_hi_256(31),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(31),        -- Port B data input
DOB(0)   => data_read_b_hi_256(31),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


end;