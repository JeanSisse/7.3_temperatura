-------------------------------------------------------------------------------------
--	Partial Repository																
--		Contains the object codes of the tasks inserted on runtime						
-------------------------------------------------------------------------------------
--repository structure:																
--[/this structure is replicaded according the number of tasks]						
--number of tasks																	
--task id																			
--task code size																		
--processor (ffffffff means dynamic allocation)										
--task code start address															
--[/this structure is replicaded according the number of tasks]						
--tasks codes																		
-------------------------------------------------------------------------------------
library IEEE;																		
use IEEE.Std_Logic_1164.all;														  

package memory_pack is 															  

	constant NUMBER_OF_APPS			: integer := 50;
	type timearray is array(0 to NUMBER_OF_APPS) of time;
	constant appstime : timearray := (0 ms,0 ms,0 ms,0 ms,0 ms,0 ms,0 ms,0 ms,0 ms,0 ms,0 ms,0 ms,0 ms,0 ms,0 ms,0 ms,0 ms,0 ms,0 ms,0 ms,0 ms,0 ms,0 ms,0 ms,0 ms,0 ms,0 ms,0 ms,0 ms,0 ms,0 ms,0 ms,0 ms,0 ms,0 ms,0 ms,0 ms,0 ms,0 ms,0 ms,0 ms,0 ms,0 ms,0 ms,0 ms,0 ms,0 ms,0 ms,0 ms,0 ms,0 ms);
	constant REPOSITORY_SIZE	: integer := 3855;
	type ram is array (0 to REPOSITORY_SIZE) of std_logic_vector(31 downto 0);		  

	signal memory : ram := (		
														
		x"00000005",	 --application mpeg	#id 0
		x"00000004",	 --initial task id start.c
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"00000000",	 --idct.c
		x"00000532",	 --code size
		x"00000200",	 --data size
		x"00000093",	 --bss size
		x"00000234",	 --initial address
		x"00005536",	 --load
		x"00000001",
		x"00000500",
		x"00000003",
		x"00000500",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"00000001",	 --iquant.c
		x"000001d7",	 --code size
		x"00000010",	 --data size
		x"00000092",	 --bss size
		x"000016fc",	 --initial address
		x"00003815",	 --load
		x"00000002",
		x"00000500",
		x"00000000",
		x"00000500",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"00000002",	 --ivlc.c
		x"0000040b",	 --code size
		x"00000110",	 --data size
		x"00000094",	 --bss size
		x"00001e58",	 --initial address
		x"00039bc8",	 --load
		x"00000004",
		x"00000a00",
		x"00000001",
		x"00000500",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"00000003",	 --print.c
		x"00000153",	 --code size
		x"00000000",	 --data size
		x"00000092",	 --bss size
		x"00002e84",	 --initial address
		x"00000403",	 --load
		x"00000000",
		x"00000500",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"00000004",	 --start.c
		x"0000021b",	 --code size
		x"00000080",	 --data size
		x"00000092",	 --bss size
		x"000033d0",	 --initial address
		x"00000dd8",	 --load
		x"00000002",
		x"00000a00",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"241d3fff",	 --idct.c
		x"0c0002bc",
		x"00000000",
		x"00002021",
		x"0000000c",
		x"00000000",
		x"08000006",
		x"00000000",
		x"0000000c",
		x"00000000",
		x"03e00008",
		x"00000000",
		x"14800007",
		x"3c050000",
		x"24a31504",
		x"24020030",
		x"00602021",
		x"a0a21504",
		x"08000045",
		x"a0600001",
		x"3c02cccc",
		x"3442cccd",
		x"00820019",
		x"00404021",
		x"24a71504",
		x"24060001",
		x"2409000b",
		x"00001810",
		x"000318c2",
		x"000310c0",
		x"00031840",
		x"00621821",
		x"00831823",
		x"24630030",
		x"0800002f",
		x"a0a31504",
		x"00880019",
		x"24c60001",
		x"00001010",
		x"000210c2",
		x"000218c0",
		x"00021040",
		x"00431021",
		x"00821023",
		x"24420030",
		x"10c90006",
		x"a0e20000",
		x"00880019",
		x"00001010",
		x"000220c2",
		x"1480fff1",
		x"24e70001",
		x"3c020000",
		x"244214f8",
		x"24c4ffff",
		x"3c030000",
		x"00822821",
		x"24631504",
		x"00c21021",
		x"08000040",
		x"a0400000",
		x"9062ffff",
		x"2484ffff",
		x"a0a20001",
		x"24630001",
		x"0481fffb",
		x"24a5ffff",
		x"3c020000",
		x"244414f8",
		x"03e00008",
		x"00801021",
		x"3c020000",
		x"24050030",
		x"244314ec",
		x"a04514ec",
		x"24020078",
		x"a0620001",
		x"1480000a",
		x"a060000a",
		x"a0650009",
		x"a0650002",
		x"a0650003",
		x"a0650004",
		x"a0650005",
		x"a0650006",
		x"a0650007",
		x"08000068",
		x"a0650008",
		x"3c020000",
		x"244514f5",
		x"3c020000",
		x"244714ed",
		x"3082000f",
		x"24460030",
		x"24430057",
		x"2c42000a",
		x"10400003",
		x"00000000",
		x"08000065",
		x"a0a60000",
		x"a0a30000",
		x"24a5ffff",
		x"14a7fff5",
		x"00042102",
		x"3c020000",
		x"03e00008",
		x"244214ec",
		x"04810002",
		x"00801021",
		x"00041023",
		x"03e00008",
		x"00000000",
		x"30820001",
		x"00021023",
		x"3042b400",
		x"00042043",
		x"00822026",
		x"14c00002",
		x"0086001a",
		x"0007000d",
		x"00001010",
		x"03e00008",
		x"00451021",
		x"03e00008",
		x"00851021",
		x"03e00008",
		x"00851023",
		x"00801021",
		x"08000084",
		x"00801821",
		x"a0650000",
		x"24630001",
		x"1cc0fffd",
		x"24c6ffff",
		x"03e00008",
		x"00000000",
		x"0481003c",
		x"00801021",
		x"3c020000",
		x"244714dc",
		x"3c026666",
		x"00042823",
		x"344a6667",
		x"00003021",
		x"24090030",
		x"080000a3",
		x"2408000c",
		x"080000a0",
		x"a0e90000",
		x"00aa0018",
		x"00001010",
		x"00021083",
		x"00431023",
		x"00021840",
		x"000220c0",
		x"00641821",
		x"00a31823",
		x"24630030",
		x"00402821",
		x"a0e30000",
		x"24c60001",
		x"10c80006",
		x"24e70001",
		x"00051fc3",
		x"14a0fff0",
		x"28c20005",
		x"1440ffec",
		x"00000000",
		x"3c030000",
		x"246314cc",
		x"3c020000",
		x"24c40001",
		x"00604021",
		x"244714dc",
		x"00c31821",
		x"00002821",
		x"24090004",
		x"2406002e",
		x"080000be",
		x"a0600002",
		x"14a90003",
		x"00000000",
		x"a0460000",
		x"2484ffff",
		x"90e30000",
		x"00881021",
		x"24a50001",
		x"a0430000",
		x"2484ffff",
		x"24e70001",
		x"0481fff5",
		x"00881021",
		x"3c030000",
		x"2402002d",
		x"246514cc",
		x"08000104",
		x"a06214cc",
		x"10400005",
		x"3c040000",
		x"00402821",
		x"248714dc",
		x"080000e5",
		x"00003021",
		x"248314dc",
		x"24020030",
		x"00602821",
		x"a08214dc",
		x"08000104",
		x"a0600001",
		x"24020030",
		x"080000e1",
		x"a0e20000",
		x"3c026666",
		x"34426667",
		x"00a20018",
		x"00001010",
		x"00021083",
		x"00431023",
		x"00021840",
		x"000220c0",
		x"00641821",
		x"00a31823",
		x"24630030",
		x"00402821",
		x"a0e30000",
		x"24c60001",
		x"2402000c",
		x"10c20006",
		x"24e70001",
		x"00051fc3",
		x"14a0ffed",
		x"28c20005",
		x"1440ffe8",
		x"00000000",
		x"3c030000",
		x"246314cc",
		x"3c020000",
		x"00c02021",
		x"00604021",
		x"244714dc",
		x"00c31821",
		x"00002821",
		x"24090004",
		x"2406002e",
		x"08000100",
		x"a0600001",
		x"14a90003",
		x"00000000",
		x"a0460000",
		x"2484ffff",
		x"90e30000",
		x"00881021",
		x"24a50001",
		x"a0430000",
		x"2484ffff",
		x"24e70001",
		x"0481fff5",
		x"00881021",
		x"3c020000",
		x"244514cc",
		x"03e00008",
		x"00a01021",
		x"00801821",
		x"80a20000",
		x"24a50001",
		x"a0620000",
		x"1440fffc",
		x"24630001",
		x"03e00008",
		x"00801021",
		x"00801821",
		x"80620000",
		x"00000000",
		x"1440fffd",
		x"24630001",
		x"00641023",
		x"03e00008",
		x"2442ffff",
		x"27bdffc0",
		x"afbe0038",
		x"afb70034",
		x"afb40028",
		x"afb30024",
		x"afb1001c",
		x"afb60030",
		x"afb5002c",
		x"afb20020",
		x"afb00018",
		x"00809821",
		x"00a0a021",
		x"0005f080",
		x"00808821",
		x"0000b821",
		x"8e220010",
		x"8e390018",
		x"8e320008",
		x"8e300004",
		x"8e2e001c",
		x"0002aac0",
		x"8e380014",
		x"8e2f000c",
		x"02591025",
		x"004e1025",
		x"02b01825",
		x"00781825",
		x"004f1025",
		x"00621825",
		x"8e360000",
		x"1460000b",
		x"000e1180",
		x"001610c0",
		x"ae220000",
		x"ae22001c",
		x"ae220018",
		x"ae220014",
		x"ae220010",
		x"ae22000c",
		x"ae220008",
		x"080001ba",
		x"ae220004",
		x"000e28c0",
		x"030f5821",
		x"00a22821",
		x"020e3821",
		x"00ae2823",
		x"00101940",
		x"000b1100",
		x"00102080",
		x"000b3080",
		x"00c23021",
		x"00076100",
		x"000f4080",
		x"00832021",
		x"000749c0",
		x"00055080",
		x"001811c0",
		x"000f6a00",
		x"00181940",
		x"00621821",
		x"00902023",
		x"012c4823",
		x"01455023",
		x"01a86823",
		x"00066100",
		x"01274821",
		x"01866023",
		x"01af6823",
		x"00041180",
		x"00032880",
		x"000a50c0",
		x"00822021",
		x"014e5023",
		x"018b6021",
		x"00651821",
		x"00091080",
		x"000d6900",
		x"01224821",
		x"00902021",
		x"00781823",
		x"01af6821",
		x"000c60c0",
		x"000a5040",
		x"018d6823",
		x"012a5023",
		x"01836023",
		x"01244821",
		x"014d1023",
		x"012c7023",
		x"02597821",
		x"01c28023",
		x"000f2880",
		x"01c27021",
		x"000f21c0",
		x"00191080",
		x"00191980",
		x"00852023",
		x"00621823",
		x"000e2880",
		x"00101080",
		x"000e5900",
		x"00104100",
		x"01024023",
		x"01655823",
		x"008f2023",
		x"00121140",
		x"00791823",
		x"00123a00",
		x"00e23823",
		x"000b2900",
		x"000410c0",
		x"00083100",
		x"000318c0",
		x"00822021",
		x"00ab2823",
		x"00c83023",
		x"00791821",
		x"000740c0",
		x"001612c0",
		x"008f2021",
		x"01074023",
		x"24420080",
		x"000318c0",
		x"00ae2821",
		x"00d03021",
		x"00884021",
		x"00553823",
		x"00832023",
		x"00551021",
		x"24a50080",
		x"24c60080",
		x"00485823",
		x"00e41823",
		x"012c4821",
		x"014d5021",
		x"00481021",
		x"00e43821",
		x"00052a03",
		x"00063203",
		x"016a2023",
		x"00664023",
		x"00e56023",
		x"00496823",
		x"00e53821",
		x"00491021",
		x"00661821",
		x"016a5821",
		x"00021203",
		x"00073a03",
		x"00031a03",
		x"000b5a03",
		x"00042203",
		x"00084203",
		x"000c6203",
		x"000d6a03",
		x"ae220000",
		x"ae270004",
		x"ae230008",
		x"ae2b000c",
		x"ae240010",
		x"ae280014",
		x"ae2c0018",
		x"ae2d001c",
		x"26f70001",
		x"24020008",
		x"16e2ff68",
		x"023e8821",
		x"001438c0",
		x"00141840",
		x"00743021",
		x"00142080",
		x"00141100",
		x"00e31823",
		x"00f42823",
		x"00942021",
		x"02621021",
		x"00031880",
		x"027ef021",
		x"00052880",
		x"00042080",
		x"00063080",
		x"afa20008",
		x"02631821",
		x"3c020000",
		x"afbe0000",
		x"afa30004",
		x"0265f021",
		x"0264b821",
		x"0266b021",
		x"0260c821",
		x"24540cc8",
		x"0267a821",
		x"afa0000c",
		x"8fa30008",
		x"8fa80004",
		x"8c620000",
		x"8fa30000",
		x"8d180000",
		x"8eb20000",
		x"8c700000",
		x"8fce0000",
		x"00029a00",
		x"8ef10000",
		x"8ecf0000",
		x"02581025",
		x"004e1025",
		x"02701825",
		x"00711825",
		x"004f1025",
		x"8f280000",
		x"00621825",
		x"14600012",
		x"afa80010",
		x"25020020",
		x"00021183",
		x"00021040",
		x"00541021",
		x"84420400",
		x"8fa30004",
		x"afc20000",
		x"8fa80008",
		x"ac620000",
		x"8fa30000",
		x"aee20000",
		x"ad020000",
		x"aec20000",
		x"aea20000",
		x"ac620000",
		x"0800029d",
		x"af220000",
		x"022f5021",
		x"000e1180",
		x"000e20c0",
		x"020e3821",
		x"00822021",
		x"000a2880",
		x"000a1100",
		x"00a22821",
		x"008e2023",
		x"00073100",
		x"00101140",
		x"000749c0",
		x"00101880",
		x"000f4080",
		x"01264823",
		x"00621821",
		x"001131c0",
		x"00046080",
		x"00055900",
		x"00111140",
		x"000f6a00",
		x"01274821",
		x"00701823",
		x"00461021",
		x"01846023",
		x"01655823",
		x"01a86823",
		x"016a5821",
		x"01af6823",
		x"00092080",
		x"00032980",
		x"00023080",
		x"000c60c0",
		x"01244821",
		x"00651821",
		x"018e6023",
		x"00461021",
		x"000b58c0",
		x"000d6900",
		x"00701821",
		x"00511023",
		x"01af6821",
		x"25290004",
		x"256b0004",
		x"000c6040",
		x"012c6023",
		x"016d6823",
		x"01234821",
		x"01625823",
		x"000b58c3",
		x"000d68c3",
		x"000948c3",
		x"000c60c3",
		x"018d2823",
		x"02587821",
		x"012b7023",
		x"01c58023",
		x"000f1880",
		x"01c57021",
		x"000f11c0",
		x"00431023",
		x"000e3880",
		x"000e4100",
		x"01074023",
		x"00181880",
		x"004f1023",
		x"00123140",
		x"00182180",
		x"00125200",
		x"01465023",
		x"00832023",
		x"00102880",
		x"00083100",
		x"000288c0",
		x"00101900",
		x"00651823",
		x"00c83023",
		x"00982023",
		x"8fa80010",
		x"00511021",
		x"000a28c0",
		x"00033900",
		x"000420c0",
		x"004f1021",
		x"00aa2823",
		x"00e33823",
		x"24420004",
		x"00081a00",
		x"00982021",
		x"000420c0",
		x"00452821",
		x"24632000",
		x"000528c3",
		x"00441023",
		x"00732023",
		x"00731821",
		x"00655023",
		x"012b4821",
		x"00651821",
		x"00ce3021",
		x"000210c3",
		x"018d6021",
		x"24c60080",
		x"00696823",
		x"00691821",
		x"00824023",
		x"00063203",
		x"00822021",
		x"00f03821",
		x"00031b83",
		x"00865823",
		x"24e70080",
		x"00862021",
		x"00031840",
		x"00073a03",
		x"00042383",
		x"00741821",
		x"01072823",
		x"014c1023",
		x"01074021",
		x"84630400",
		x"014c5021",
		x"00042040",
		x"00084383",
		x"000a5383",
		x"00021383",
		x"00942021",
		x"af230000",
		x"00084040",
		x"8fa30000",
		x"000a5040",
		x"00021040",
		x"84840400",
		x"01144021",
		x"00052b83",
		x"000b5b83",
		x"000d6b83",
		x"01545021",
		x"00541021",
		x"ac640000",
		x"85060400",
		x"84420400",
		x"00052840",
		x"000b5840",
		x"000d6840",
		x"85470400",
		x"8fa30008",
		x"00b42821",
		x"01745821",
		x"01b46821",
		x"aea60000",
		x"84a50400",
		x"aec70000",
		x"85680400",
		x"ac620000",
		x"85a90400",
		x"8fa20004",
		x"aee50000",
		x"ac480000",
		x"afc90000",
		x"8fa3000c",
		x"8fa80008",
		x"24630001",
		x"8fa20004",
		x"afa3000c",
		x"25080004",
		x"8fa30000",
		x"24420004",
		x"afa80008",
		x"8fa8000c",
		x"afa20004",
		x"24630004",
		x"24020008",
		x"26b50004",
		x"afa30000",
		x"27de0004",
		x"26f70004",
		x"26d60004",
		x"1502ff28",
		x"27390004",
		x"8fbe0038",
		x"8fb70034",
		x"8fb60030",
		x"8fb5002c",
		x"8fb40028",
		x"8fb30024",
		x"8fb20020",
		x"8fb1001c",
		x"8fb00018",
		x"03e00008",
		x"27bd0040",
		x"3c050000",
		x"27bdfee0",
		x"24a50c98",
		x"24040004",
		x"00003021",
		x"00003821",
		x"afbf011c",
		x"afb10114",
		x"afb20118",
		x"0c000008",
		x"afb00110",
		x"00002821",
		x"00003021",
		x"00003821",
		x"0c000008",
		x"24040003",
		x"0c00000c",
		x"00402021",
		x"00402821",
		x"24040004",
		x"00003021",
		x"0c000008",
		x"00003821",
		x"00008821",
		x"3c100000",
		x"26121510",
		x"24040002",
		x"02402821",
		x"24060001",
		x"0c000008",
		x"00003821",
		x"1040fff8",
		x"3c020000",
		x"8e061510",
		x"24451514",
		x"00002021",
		x"080002e5",
		x"27a30010",
		x"8ca2fffc",
		x"00000000",
		x"ac62fffc",
		x"0086102a",
		x"24a50004",
		x"24840001",
		x"1440fff9",
		x"24630004",
		x"27b00010",
		x"02002021",
		x"0c000116",
		x"24050008",
		x"3c020000",
		x"24030040",
		x"ac431510",
		x"3c020000",
		x"24451514",
		x"00002021",
		x"24060040",
		x"8e020000",
		x"24840001",
		x"0086182a",
		x"aca20000",
		x"26100004",
		x"1460fffa",
		x"24a50004",
		x"24040001",
		x"02402821",
		x"24060003",
		x"0c000008",
		x"00003821",
		x"1040fffb",
		x"24040001",
		x"26310001",
		x"2a220014",
		x"1440ffce",
		x"00002821",
		x"00003021",
		x"00003821",
		x"0c000008",
		x"24040003",
		x"0c00000c",
		x"00402021",
		x"00402821",
		x"24040004",
		x"00003021",
		x"0c000008",
		x"00003821",
		x"3c050000",
		x"24a50cb4",
		x"24040004",
		x"00003021",
		x"0c000008",
		x"00003821",
		x"00002021",
		x"00002821",
		x"00003021",
		x"0c000008",
		x"00003821",
		x"1040fffb",
		x"00002021",
		x"8fbf011c",
		x"8fb20118",
		x"8fb10114",
		x"8fb00110",
		x"00001021",
		x"03e00008",
		x"27bd0120",
		x"4d504547",
		x"20546173",
		x"6b204420",
		x"73746172",
		x"743a2069",
		x"44435420",
		x"00000000",
		x"456e6420",
		x"5461736b",
		x"2044202d",
		x"204d5045",
		x"47000000",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff00",
		x"ff00ff01",
		x"ff02ff03",
		x"ff04ff05",
		x"ff06ff07",
		x"ff08ff09",
		x"ff0aff0b",
		x"ff0cff0d",
		x"ff0eff0f",
		x"ff10ff11",
		x"ff12ff13",
		x"ff14ff15",
		x"ff16ff17",
		x"ff18ff19",
		x"ff1aff1b",
		x"ff1cff1d",
		x"ff1eff1f",
		x"ff20ff21",
		x"ff22ff23",
		x"ff24ff25",
		x"ff26ff27",
		x"ff28ff29",
		x"ff2aff2b",
		x"ff2cff2d",
		x"ff2eff2f",
		x"ff30ff31",
		x"ff32ff33",
		x"ff34ff35",
		x"ff36ff37",
		x"ff38ff39",
		x"ff3aff3b",
		x"ff3cff3d",
		x"ff3eff3f",
		x"ff40ff41",
		x"ff42ff43",
		x"ff44ff45",
		x"ff46ff47",
		x"ff48ff49",
		x"ff4aff4b",
		x"ff4cff4d",
		x"ff4eff4f",
		x"ff50ff51",
		x"ff52ff53",
		x"ff54ff55",
		x"ff56ff57",
		x"ff58ff59",
		x"ff5aff5b",
		x"ff5cff5d",
		x"ff5eff5f",
		x"ff60ff61",
		x"ff62ff63",
		x"ff64ff65",
		x"ff66ff67",
		x"ff68ff69",
		x"ff6aff6b",
		x"ff6cff6d",
		x"ff6eff6f",
		x"ff70ff71",
		x"ff72ff73",
		x"ff74ff75",
		x"ff76ff77",
		x"ff78ff79",
		x"ff7aff7b",
		x"ff7cff7d",
		x"ff7eff7f",
		x"ff80ff81",
		x"ff82ff83",
		x"ff84ff85",
		x"ff86ff87",
		x"ff88ff89",
		x"ff8aff8b",
		x"ff8cff8d",
		x"ff8eff8f",
		x"ff90ff91",
		x"ff92ff93",
		x"ff94ff95",
		x"ff96ff97",
		x"ff98ff99",
		x"ff9aff9b",
		x"ff9cff9d",
		x"ff9eff9f",
		x"ffa0ffa1",
		x"ffa2ffa3",
		x"ffa4ffa5",
		x"ffa6ffa7",
		x"ffa8ffa9",
		x"ffaaffab",
		x"ffacffad",
		x"ffaeffaf",
		x"ffb0ffb1",
		x"ffb2ffb3",
		x"ffb4ffb5",
		x"ffb6ffb7",
		x"ffb8ffb9",
		x"ffbaffbb",
		x"ffbcffbd",
		x"ffbeffbf",
		x"ffc0ffc1",
		x"ffc2ffc3",
		x"ffc4ffc5",
		x"ffc6ffc7",
		x"ffc8ffc9",
		x"ffcaffcb",
		x"ffccffcd",
		x"ffceffcf",
		x"ffd0ffd1",
		x"ffd2ffd3",
		x"ffd4ffd5",
		x"ffd6ffd7",
		x"ffd8ffd9",
		x"ffdaffdb",
		x"ffdcffdd",
		x"ffdeffdf",
		x"ffe0ffe1",
		x"ffe2ffe3",
		x"ffe4ffe5",
		x"ffe6ffe7",
		x"ffe8ffe9",
		x"ffeaffeb",
		x"ffecffed",
		x"ffeeffef",
		x"fff0fff1",
		x"fff2fff3",
		x"fff4fff5",
		x"fff6fff7",
		x"fff8fff9",
		x"fffafffb",
		x"fffcfffd",
		x"fffeffff",
		x"00000001",
		x"00020003",
		x"00040005",
		x"00060007",
		x"00080009",
		x"000a000b",
		x"000c000d",
		x"000e000f",
		x"00100011",
		x"00120013",
		x"00140015",
		x"00160017",
		x"00180019",
		x"001a001b",
		x"001c001d",
		x"001e001f",
		x"00200021",
		x"00220023",
		x"00240025",
		x"00260027",
		x"00280029",
		x"002a002b",
		x"002c002d",
		x"002e002f",
		x"00300031",
		x"00320033",
		x"00340035",
		x"00360037",
		x"00380039",
		x"003a003b",
		x"003c003d",
		x"003e003f",
		x"00400041",
		x"00420043",
		x"00440045",
		x"00460047",
		x"00480049",
		x"004a004b",
		x"004c004d",
		x"004e004f",
		x"00500051",
		x"00520053",
		x"00540055",
		x"00560057",
		x"00580059",
		x"005a005b",
		x"005c005d",
		x"005e005f",
		x"00600061",
		x"00620063",
		x"00640065",
		x"00660067",
		x"00680069",
		x"006a006b",
		x"006c006d",
		x"006e006f",
		x"00700071",
		x"00720073",
		x"00740075",
		x"00760077",
		x"00780079",
		x"007a007b",
		x"007c007d",
		x"007e007f",
		x"00800081",
		x"00820083",
		x"00840085",
		x"00860087",
		x"00880089",
		x"008a008b",
		x"008c008d",
		x"008e008f",
		x"00900091",
		x"00920093",
		x"00940095",
		x"00960097",
		x"00980099",
		x"009a009b",
		x"009c009d",
		x"009e009f",
		x"00a000a1",
		x"00a200a3",
		x"00a400a5",
		x"00a600a7",
		x"00a800a9",
		x"00aa00ab",
		x"00ac00ad",
		x"00ae00af",
		x"00b000b1",
		x"00b200b3",
		x"00b400b5",
		x"00b600b7",
		x"00b800b9",
		x"00ba00bb",
		x"00bc00bd",
		x"00be00bf",
		x"00c000c1",
		x"00c200c3",
		x"00c400c5",
		x"00c600c7",
		x"00c800c9",
		x"00ca00cb",
		x"00cc00cd",
		x"00ce00cf",
		x"00d000d1",
		x"00d200d3",
		x"00d400d5",
		x"00d600d7",
		x"00d800d9",
		x"00da00db",
		x"00dc00dd",
		x"00de00df",
		x"00e000e1",
		x"00e200e3",
		x"00e400e5",
		x"00e600e7",
		x"00e800e9",
		x"00ea00eb",
		x"00ec00ed",
		x"00ee00ef",
		x"00f000f1",
		x"00f200f3",
		x"00f400f5",
		x"00f600f7",
		x"00f800f9",
		x"00fa00fb",
		x"00fc00fd",
		x"00fe00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"00ff00ff",
		x"241d3fff",	 --iquant.c
		x"0c00014f",
		x"00000000",
		x"00002021",
		x"0000000c",
		x"00000000",
		x"08000006",
		x"00000000",
		x"0000000c",
		x"00000000",
		x"03e00008",
		x"00000000",
		x"14800007",
		x"3c050000",
		x"24a30794",
		x"24020030",
		x"00602021",
		x"a0a20794",
		x"08000045",
		x"a0600001",
		x"3c02cccc",
		x"3442cccd",
		x"00820019",
		x"00404021",
		x"24a70794",
		x"24060001",
		x"2409000b",
		x"00001810",
		x"000318c2",
		x"000310c0",
		x"00031840",
		x"00621821",
		x"00831823",
		x"24630030",
		x"0800002f",
		x"a0a30794",
		x"00880019",
		x"24c60001",
		x"00001010",
		x"000210c2",
		x"000218c0",
		x"00021040",
		x"00431021",
		x"00821023",
		x"24420030",
		x"10c90006",
		x"a0e20000",
		x"00880019",
		x"00001010",
		x"000220c2",
		x"1480fff1",
		x"24e70001",
		x"3c020000",
		x"24420788",
		x"24c4ffff",
		x"3c030000",
		x"00822821",
		x"24630794",
		x"00c21021",
		x"08000040",
		x"a0400000",
		x"9062ffff",
		x"2484ffff",
		x"a0a20001",
		x"24630001",
		x"0481fffb",
		x"24a5ffff",
		x"3c020000",
		x"24440788",
		x"03e00008",
		x"00801021",
		x"3c020000",
		x"24050030",
		x"2443077c",
		x"a045077c",
		x"24020078",
		x"a0620001",
		x"1480000a",
		x"a060000a",
		x"a0650009",
		x"a0650002",
		x"a0650003",
		x"a0650004",
		x"a0650005",
		x"a0650006",
		x"a0650007",
		x"08000068",
		x"a0650008",
		x"3c020000",
		x"24450785",
		x"3c020000",
		x"2447077d",
		x"3082000f",
		x"24460030",
		x"24430057",
		x"2c42000a",
		x"10400003",
		x"00000000",
		x"08000065",
		x"a0a60000",
		x"a0a30000",
		x"24a5ffff",
		x"14a7fff5",
		x"00042102",
		x"3c020000",
		x"03e00008",
		x"2442077c",
		x"04810002",
		x"00801021",
		x"00041023",
		x"03e00008",
		x"00000000",
		x"30820001",
		x"00021023",
		x"3042b400",
		x"00042043",
		x"00822026",
		x"14c00002",
		x"0086001a",
		x"0007000d",
		x"00001010",
		x"03e00008",
		x"00451021",
		x"03e00008",
		x"00851021",
		x"03e00008",
		x"00851023",
		x"00801021",
		x"08000084",
		x"00801821",
		x"a0650000",
		x"24630001",
		x"1cc0fffd",
		x"24c6ffff",
		x"03e00008",
		x"00000000",
		x"0481003c",
		x"00801021",
		x"3c020000",
		x"2447076c",
		x"3c026666",
		x"00042823",
		x"344a6667",
		x"00003021",
		x"24090030",
		x"080000a3",
		x"2408000c",
		x"080000a0",
		x"a0e90000",
		x"00aa0018",
		x"00001010",
		x"00021083",
		x"00431023",
		x"00021840",
		x"000220c0",
		x"00641821",
		x"00a31823",
		x"24630030",
		x"00402821",
		x"a0e30000",
		x"24c60001",
		x"10c80006",
		x"24e70001",
		x"00051fc3",
		x"14a0fff0",
		x"28c20005",
		x"1440ffec",
		x"00000000",
		x"3c030000",
		x"2463075c",
		x"3c020000",
		x"24c40001",
		x"00604021",
		x"2447076c",
		x"00c31821",
		x"00002821",
		x"24090004",
		x"2406002e",
		x"080000be",
		x"a0600002",
		x"14a90003",
		x"00000000",
		x"a0460000",
		x"2484ffff",
		x"90e30000",
		x"00881021",
		x"24a50001",
		x"a0430000",
		x"2484ffff",
		x"24e70001",
		x"0481fff5",
		x"00881021",
		x"3c030000",
		x"2402002d",
		x"2465075c",
		x"08000104",
		x"a062075c",
		x"10400005",
		x"3c040000",
		x"00402821",
		x"2487076c",
		x"080000e5",
		x"00003021",
		x"2483076c",
		x"24020030",
		x"00602821",
		x"a082076c",
		x"08000104",
		x"a0600001",
		x"24020030",
		x"080000e1",
		x"a0e20000",
		x"3c026666",
		x"34426667",
		x"00a20018",
		x"00001010",
		x"00021083",
		x"00431023",
		x"00021840",
		x"000220c0",
		x"00641821",
		x"00a31823",
		x"24630030",
		x"00402821",
		x"a0e30000",
		x"24c60001",
		x"2402000c",
		x"10c20006",
		x"24e70001",
		x"00051fc3",
		x"14a0ffed",
		x"28c20005",
		x"1440ffe8",
		x"00000000",
		x"3c030000",
		x"2463075c",
		x"3c020000",
		x"00c02021",
		x"00604021",
		x"2447076c",
		x"00c31821",
		x"00002821",
		x"24090004",
		x"2406002e",
		x"08000100",
		x"a0600001",
		x"14a90003",
		x"00000000",
		x"a0460000",
		x"2484ffff",
		x"90e30000",
		x"00881021",
		x"24a50001",
		x"a0430000",
		x"2484ffff",
		x"24e70001",
		x"0481fff5",
		x"00881021",
		x"3c020000",
		x"2445075c",
		x"03e00008",
		x"00a01021",
		x"00801821",
		x"80a20000",
		x"24a50001",
		x"a0620000",
		x"1440fffc",
		x"24630001",
		x"03e00008",
		x"00801021",
		x"00801821",
		x"80620000",
		x"00000000",
		x"1440fffd",
		x"24630001",
		x"00641023",
		x"03e00008",
		x"2442ffff",
		x"8c820000",
		x"24030003",
		x"00661823",
		x"00625804",
		x"3c020000",
		x"ac8b0000",
		x"2459071c",
		x"00057080",
		x"00805021",
		x"00006821",
		x"24180008",
		x"240f0008",
		x"000d10c0",
		x"00594821",
		x"01404021",
		x"00006021",
		x"01ac1025",
		x"10400014",
		x"00000000",
		x"91220000",
		x"8d030000",
		x"00e20018",
		x"00001012",
		x"00000000",
		x"00000000",
		x"00430018",
		x"00001012",
		x"00021903",
		x"2862f800",
		x"10400003",
		x"28660800",
		x"0800013a",
		x"2403f800",
		x"14c00002",
		x"00000000",
		x"240307ff",
		x"01635821",
		x"ad030000",
		x"258c0001",
		x"25080004",
		x"1598ffe7",
		x"25290001",
		x"25ad0001",
		x"15afffe0",
		x"014e5021",
		x"000510c0",
		x"31630001",
		x"14600007",
		x"00451023",
		x"00021880",
		x"00831821",
		x"8c62001c",
		x"00000000",
		x"38420001",
		x"ac62001c",
		x"03e00008",
		x"00000000",
		x"3c050000",
		x"27bdfee0",
		x"24a506ec",
		x"24040004",
		x"00003021",
		x"00003821",
		x"afbf011c",
		x"afb10114",
		x"afb20118",
		x"0c000008",
		x"afb00110",
		x"00002821",
		x"00003021",
		x"00003821",
		x"0c000008",
		x"24040003",
		x"0c00000c",
		x"00402021",
		x"00402821",
		x"24040004",
		x"00003021",
		x"0c000008",
		x"00003821",
		x"00008821",
		x"3c100000",
		x"261207a0",
		x"24040002",
		x"02402821",
		x"24060002",
		x"0c000008",
		x"00003821",
		x"1040fff8",
		x"3c020000",
		x"8e0607a0",
		x"244507a4",
		x"00002021",
		x"08000178",
		x"27a30010",
		x"8ca2fffc",
		x"00000000",
		x"ac62fffc",
		x"0086102a",
		x"24a50004",
		x"24840001",
		x"1440fff9",
		x"24630004",
		x"27b00010",
		x"02002021",
		x"24050008",
		x"00003021",
		x"0c000116",
		x"24070001",
		x"3c020000",
		x"24030040",
		x"ac4307a0",
		x"3c020000",
		x"244507a4",
		x"00002021",
		x"24060040",
		x"8e020000",
		x"24840001",
		x"0086182a",
		x"aca20000",
		x"26100004",
		x"1460fffa",
		x"24a50004",
		x"24040001",
		x"02402821",
		x"00003021",
		x"0c000008",
		x"00003821",
		x"1040fffb",
		x"24040001",
		x"26310001",
		x"2a220014",
		x"1440ffcc",
		x"00002821",
		x"00003021",
		x"00003821",
		x"0c000008",
		x"24040003",
		x"0c00000c",
		x"00402021",
		x"00402821",
		x"24040004",
		x"00003021",
		x"0c000008",
		x"00003821",
		x"3c050000",
		x"24a50708",
		x"24040004",
		x"00003021",
		x"0c000008",
		x"00003821",
		x"00002021",
		x"00002821",
		x"00003021",
		x"0c000008",
		x"00003821",
		x"1040fffb",
		x"00002021",
		x"8fbf011c",
		x"8fb20118",
		x"8fb10114",
		x"8fb00110",
		x"00001021",
		x"03e00008",
		x"27bd0120",
		x"4d504547",
		x"20546173",
		x"6b204320",
		x"73746172",
		x"743a2069",
		x"7175616e",
		x"74200000",
		x"456e6420",
		x"5461736b",
		x"20432d20",
		x"4d504547",
		x"00000000",
		x"08101316",
		x"1a1b1d22",
		x"10101618",
		x"1b1d2225",
		x"13161a1b",
		x"1d222226",
		x"16161a1b",
		x"1d222528",
		x"161a1b1d",
		x"20232830",
		x"1a1b1d20",
		x"2328303a",
		x"1a1b1d22",
		x"262e3845",
		x"1b1d2326",
		x"2e384553",
		x"241d3fff",	 --ivlc.c
		x"0c000247",
		x"00000000",
		x"00002021",
		x"0000000c",
		x"00000000",
		x"08000006",
		x"00000000",
		x"0000000c",
		x"00000000",
		x"03e00008",
		x"00000000",
		x"14800007",
		x"3c050000",
		x"24a3106c",
		x"24020030",
		x"00602021",
		x"a0a2106c",
		x"08000045",
		x"a0600001",
		x"3c02cccc",
		x"3442cccd",
		x"00820019",
		x"00404021",
		x"24a7106c",
		x"24060001",
		x"2409000b",
		x"00001810",
		x"000318c2",
		x"000310c0",
		x"00031840",
		x"00621821",
		x"00831823",
		x"24630030",
		x"0800002f",
		x"a0a3106c",
		x"00880019",
		x"24c60001",
		x"00001010",
		x"000210c2",
		x"000218c0",
		x"00021040",
		x"00431021",
		x"00821023",
		x"24420030",
		x"10c90006",
		x"a0e20000",
		x"00880019",
		x"00001010",
		x"000220c2",
		x"1480fff1",
		x"24e70001",
		x"3c020000",
		x"24421060",
		x"24c4ffff",
		x"3c030000",
		x"00822821",
		x"2463106c",
		x"00c21021",
		x"08000040",
		x"a0400000",
		x"9062ffff",
		x"2484ffff",
		x"a0a20001",
		x"24630001",
		x"0481fffb",
		x"24a5ffff",
		x"3c020000",
		x"24441060",
		x"03e00008",
		x"00801021",
		x"3c020000",
		x"24050030",
		x"24431054",
		x"a0451054",
		x"24020078",
		x"a0620001",
		x"1480000a",
		x"a060000a",
		x"a0650009",
		x"a0650002",
		x"a0650003",
		x"a0650004",
		x"a0650005",
		x"a0650006",
		x"a0650007",
		x"08000068",
		x"a0650008",
		x"3c020000",
		x"2445105d",
		x"3c020000",
		x"24471055",
		x"3082000f",
		x"24460030",
		x"24430057",
		x"2c42000a",
		x"10400003",
		x"00000000",
		x"08000065",
		x"a0a60000",
		x"a0a30000",
		x"24a5ffff",
		x"14a7fff5",
		x"00042102",
		x"3c020000",
		x"03e00008",
		x"24421054",
		x"04810002",
		x"00801021",
		x"00041023",
		x"03e00008",
		x"00000000",
		x"30820001",
		x"00021023",
		x"3042b400",
		x"00042043",
		x"00822026",
		x"14c00002",
		x"0086001a",
		x"0007000d",
		x"00001010",
		x"03e00008",
		x"00451021",
		x"03e00008",
		x"00851021",
		x"03e00008",
		x"00851023",
		x"00801021",
		x"08000084",
		x"00801821",
		x"a0650000",
		x"24630001",
		x"1cc0fffd",
		x"24c6ffff",
		x"03e00008",
		x"00000000",
		x"0481003c",
		x"00801021",
		x"3c020000",
		x"24471044",
		x"3c026666",
		x"00042823",
		x"344a6667",
		x"00003021",
		x"24090030",
		x"080000a3",
		x"2408000c",
		x"080000a0",
		x"a0e90000",
		x"00aa0018",
		x"00001010",
		x"00021083",
		x"00431023",
		x"00021840",
		x"000220c0",
		x"00641821",
		x"00a31823",
		x"24630030",
		x"00402821",
		x"a0e30000",
		x"24c60001",
		x"10c80006",
		x"24e70001",
		x"00051fc3",
		x"14a0fff0",
		x"28c20005",
		x"1440ffec",
		x"00000000",
		x"3c030000",
		x"24631034",
		x"3c020000",
		x"24c40001",
		x"00604021",
		x"24471044",
		x"00c31821",
		x"00002821",
		x"24090004",
		x"2406002e",
		x"080000be",
		x"a0600002",
		x"14a90003",
		x"00000000",
		x"a0460000",
		x"2484ffff",
		x"90e30000",
		x"00881021",
		x"24a50001",
		x"a0430000",
		x"2484ffff",
		x"24e70001",
		x"0481fff5",
		x"00881021",
		x"3c030000",
		x"2402002d",
		x"24651034",
		x"08000104",
		x"a0621034",
		x"10400005",
		x"3c040000",
		x"00402821",
		x"24871044",
		x"080000e5",
		x"00003021",
		x"24831044",
		x"24020030",
		x"00602821",
		x"a0821044",
		x"08000104",
		x"a0600001",
		x"24020030",
		x"080000e1",
		x"a0e20000",
		x"3c026666",
		x"34426667",
		x"00a20018",
		x"00001010",
		x"00021083",
		x"00431023",
		x"00021840",
		x"000220c0",
		x"00641821",
		x"00a31823",
		x"24630030",
		x"00402821",
		x"a0e30000",
		x"24c60001",
		x"2402000c",
		x"10c20006",
		x"24e70001",
		x"00051fc3",
		x"14a0ffed",
		x"28c20005",
		x"1440ffe8",
		x"00000000",
		x"3c030000",
		x"24631034",
		x"3c020000",
		x"00c02021",
		x"00604021",
		x"24471044",
		x"00c31821",
		x"00002821",
		x"24090004",
		x"2406002e",
		x"08000100",
		x"a0600001",
		x"14a90003",
		x"00000000",
		x"a0460000",
		x"2484ffff",
		x"90e30000",
		x"00881021",
		x"24a50001",
		x"a0430000",
		x"2484ffff",
		x"24e70001",
		x"0481fff5",
		x"00881021",
		x"3c020000",
		x"24451034",
		x"03e00008",
		x"00a01021",
		x"00801821",
		x"80a20000",
		x"24a50001",
		x"a0620000",
		x"1440fffc",
		x"24630001",
		x"03e00008",
		x"00801021",
		x"00801821",
		x"80620000",
		x"00000000",
		x"1440fffd",
		x"24630001",
		x"00641023",
		x"03e00008",
		x"2442ffff",
		x"00073c00",
		x"00047400",
		x"3c0b0000",
		x"3c030000",
		x"3c090000",
		x"00052c00",
		x"00073c03",
		x"000e7403",
		x"856a1030",
		x"84681028",
		x"8524102a",
		x"14e0002c",
		x"00052c03",
		x"000a1080",
		x"00463021",
		x"308700ff",
		x"00006821",
		x"00006021",
		x"0800013b",
		x"240fffff",
		x"8cc20000",
		x"152f0006",
		x"00000000",
		x"000b5400",
		x"000a5403",
		x"24c60004",
		x"24090007",
		x"24040080",
		x"00471024",
		x"01021007",
		x"00021400",
		x"000d1840",
		x"00021403",
		x"258c0001",
		x"00626821",
		x"01204021",
		x"00803821",
		x"000c1400",
		x"00021403",
		x"2503ffff",
		x"00072042",
		x"00034c00",
		x"004e102a",
		x"254b0001",
		x"00094c03",
		x"1440ffe6",
		x"308400ff",
		x"10a0000e",
		x"00000000",
		x"3c020000",
		x"a44a1030",
		x"3c020000",
		x"a4481028",
		x"3c020000",
		x"08000154",
		x"a447102a",
		x"24020007",
		x"a4621028",
		x"24020080",
		x"a522102a",
		x"a5601030",
		x"00006821",
		x"03e00008",
		x"01a01021",
		x"27bdffe0",
		x"afb10014",
		x"00a08821",
		x"afb00010",
		x"00002821",
		x"00048400",
		x"02203021",
		x"24040005",
		x"afbf0018",
		x"0c000116",
		x"00003821",
		x"00021c00",
		x"00031c03",
		x"2862001f",
		x"10400009",
		x"00108403",
		x"12000004",
		x"00031840",
		x"3c020000",
		x"0800017a",
		x"24420b0c",
		x"3c020000",
		x"0800017a",
		x"24420b4c",
		x"12000012",
		x"02203021",
		x"2404000a",
		x"00002821",
		x"0c000116",
		x"00003821",
		x"2442fc20",
		x"00021400",
		x"00021403",
		x"3c030000",
		x"00021040",
		x"24630b8c",
		x"00431021",
		x"80440001",
		x"80500000",
		x"24050001",
		x"02203021",
		x"08000191",
		x"00003821",
		x"24040009",
		x"00002821",
		x"0c000116",
		x"00003821",
		x"2442fe10",
		x"00021400",
		x"00021403",
		x"3c030000",
		x"00021040",
		x"24630bcc",
		x"00431021",
		x"80440001",
		x"80500000",
		x"24050001",
		x"02203021",
		x"00003821",
		x"0c000116",
		x"00000000",
		x"12000012",
		x"00002021",
		x"02002021",
		x"02203021",
		x"24050001",
		x"0c000116",
		x"00003821",
		x"00022400",
		x"00042403",
		x"2602ffff",
		x"00441007",
		x"30420001",
		x"14400006",
		x"24020001",
		x"02021004",
		x"00821023",
		x"24420001",
		x"00022400",
		x"00042403",
		x"8fbf0018",
		x"8fb10014",
		x"8fb00010",
		x"00801021",
		x"03e00008",
		x"27bd0020",
		x"27bdffd8",
		x"afb00010",
		x"00058400",
		x"afb40020",
		x"afb3001c",
		x"0006a400",
		x"afb20018",
		x"00108403",
		x"00809821",
		x"00e09021",
		x"00002021",
		x"00002821",
		x"00003021",
		x"24070001",
		x"afbf0024",
		x"afb10014",
		x"0c000116",
		x"0014a403",
		x"12000002",
		x"00002021",
		x"24040001",
		x"0c000156",
		x"02402821",
		x"ae620000",
		x"24110001",
		x"24040010",
		x"00002821",
		x"02403021",
		x"0c000116",
		x"00003821",
		x"00402021",
		x"2c420400",
		x"14400007",
		x"00041202",
		x"00021840",
		x"00621821",
		x"3c020000",
		x"24420c2c",
		x"08000204",
		x"2442fff4",
		x"2c820200",
		x"14400007",
		x"00041182",
		x"00021840",
		x"00621821",
		x"3c020000",
		x"24420f20",
		x"08000204",
		x"2442ffe8",
		x"2c820100",
		x"14400006",
		x"00041102",
		x"00021840",
		x"00621821",
		x"3c020000",
		x"08000203",
		x"24420f38",
		x"2c820080",
		x"14400006",
		x"000410c2",
		x"00021840",
		x"00621821",
		x"3c020000",
		x"08000203",
		x"24420f68",
		x"2c820040",
		x"14400006",
		x"00041082",
		x"00021840",
		x"00621821",
		x"3c020000",
		x"08000203",
		x"24420f98",
		x"2c820020",
		x"14400006",
		x"00041042",
		x"00021840",
		x"00621821",
		x"3c020000",
		x"08000203",
		x"24420fc8",
		x"2c820010",
		x"14400040",
		x"00041840",
		x"3c020000",
		x"00641821",
		x"24420ff8",
		x"2442ffd0",
		x"00628021",
		x"82040002",
		x"24050001",
		x"02403021",
		x"0c000116",
		x"00003821",
		x"82030000",
		x"24020040",
		x"10620032",
		x"24020041",
		x"14620016",
		x"24040001",
		x"24040006",
		x"24050001",
		x"02403021",
		x"0c000116",
		x"00003821",
		x"2404000c",
		x"24050001",
		x"02403021",
		x"00003821",
		x"0c000116",
		x"02228821",
		x"00408021",
		x"304207ff",
		x"10400021",
		x"2a020800",
		x"38440001",
		x"1080000c",
		x"2a220040",
		x"24021000",
		x"0800022c",
		x"00508023",
		x"24050001",
		x"02403021",
		x"00003821",
		x"82100001",
		x"0c000116",
		x"02238821",
		x"00402021",
		x"2a220040",
		x"10400011",
		x"3c020000",
		x"24420bec",
		x"02221021",
		x"90450000",
		x"10800002",
		x"000518c2",
		x"00108023",
		x"00740018",
		x"000318c0",
		x"00a31823",
		x"26310001",
		x"00001012",
		x"00431021",
		x"00021080",
		x"00531021",
		x"080001c5",
		x"ac500000",
		x"8fbf0024",
		x"8fb40020",
		x"8fb3001c",
		x"8fb20018",
		x"8fb10014",
		x"8fb00010",
		x"03e00008",
		x"27bd0028",
		x"3c050000",
		x"27bdfce0",
		x"24a50adc",
		x"24040004",
		x"00003021",
		x"00003821",
		x"afbf031c",
		x"afb10314",
		x"afb20318",
		x"0c000008",
		x"afb00310",
		x"00002821",
		x"00003021",
		x"00003821",
		x"0c000008",
		x"24040003",
		x"0c00000c",
		x"00402021",
		x"00402821",
		x"24040004",
		x"00003021",
		x"0c000008",
		x"00003821",
		x"00008821",
		x"3c100000",
		x"26121078",
		x"24040002",
		x"02402821",
		x"24060004",
		x"0c000008",
		x"00003821",
		x"1040fff8",
		x"3c020000",
		x"8e061078",
		x"2445107c",
		x"00002021",
		x"08000270",
		x"27a30110",
		x"8ca2fffc",
		x"00000000",
		x"ac62fffc",
		x"0086102a",
		x"24a50004",
		x"24840001",
		x"1440fff9",
		x"24630004",
		x"27a70010",
		x"27a20110",
		x"ace00000",
		x"24e70004",
		x"14e2fffd",
		x"27b00010",
		x"02002021",
		x"00002821",
		x"0c0001ac",
		x"24060008",
		x"3c020000",
		x"24030040",
		x"ac431078",
		x"3c020000",
		x"2445107c",
		x"00002021",
		x"24060040",
		x"8e020000",
		x"24840001",
		x"0086182a",
		x"aca20000",
		x"26100004",
		x"1460fffa",
		x"24a50004",
		x"24040001",
		x"02402821",
		x"24060001",
		x"0c000008",
		x"00003821",
		x"1040fffb",
		x"24040001",
		x"26310001",
		x"2a220014",
		x"1440ffc8",
		x"00002821",
		x"00003021",
		x"00003821",
		x"0c000008",
		x"24040003",
		x"0c00000c",
		x"00402021",
		x"00402821",
		x"24040004",
		x"00003021",
		x"0c000008",
		x"00003821",
		x"3c050000",
		x"24a50af8",
		x"24040004",
		x"00003021",
		x"0c000008",
		x"00003821",
		x"00002021",
		x"00002821",
		x"00003021",
		x"0c000008",
		x"00003821",
		x"1040fffb",
		x"00002021",
		x"8fbf031c",
		x"8fb20318",
		x"8fb10314",
		x"8fb00310",
		x"00001021",
		x"03e00008",
		x"27bd0320",
		x"4d504547",
		x"20546173",
		x"6b204220",
		x"73746172",
		x"743a2069",
		x"564c4320",
		x"00000000",
		x"456e6420",
		x"5461736b",
		x"2042202d",
		x"204d5045",
		x"47000000",
		x"00020002",
		x"00020002",
		x"00020002",
		x"00020002",
		x"01020102",
		x"01020102",
		x"01020102",
		x"01020102",
		x"02020202",
		x"02020202",
		x"02020202",
		x"02020202",
		x"03030303",
		x"03030303",
		x"04040404",
		x"05050000",
		x"01020102",
		x"01020102",
		x"01020102",
		x"01020102",
		x"02020202",
		x"02020202",
		x"02020202",
		x"02020202",
		x"00030003",
		x"00030003",
		x"03030303",
		x"03030303",
		x"04030403",
		x"04030403",
		x"05040504",
		x"06050000",
		x"06060606",
		x"06060606",
		x"06060606",
		x"06060606",
		x"06060606",
		x"06060606",
		x"06060606",
		x"06060606",
		x"07070707",
		x"07070707",
		x"07070707",
		x"07070707",
		x"08080808",
		x"08080808",
		x"09090909",
		x"0a0a0b0a",
		x"07060706",
		x"07060706",
		x"07060706",
		x"07060706",
		x"08070807",
		x"08070807",
		x"09080908",
		x"0a090b09",
		x"00010810",
		x"0902030a",
		x"11182019",
		x"120b0405",
		x"0c131a21",
		x"28302922",
		x"1b140d06",
		x"070e151c",
		x"232a3138",
		x"39322b24",
		x"1d160f17",
		x"1e252c33",
		x"3a3b342d",
		x"261f272e",
		x"353c3d36",
		x"2f373e3f",
		x"41000641",
		x"00064100",
		x"06410006",
		x"07010707",
		x"01070801",
		x"07080107",
		x"06010706",
		x"01070202",
		x"07020207",
		x"00070600",
		x"07060007",
		x"06000706",
		x"00060600",
		x"06060006",
		x"06000606",
		x"04010604",
		x"01060401",
		x"06040106",
		x"05010605",
		x"01060501",
		x"06050106",
		x"0105080b",
		x"0108000b",
		x"08000a08",
		x"0d01080c",
		x"01080302",
		x"08010408",
		x"02010502",
		x"01050201",
		x"05020105",
		x"02010502",
		x"01050201",
		x"05020105",
		x"01020501",
		x"02050102",
		x"05010205",
		x"01020501",
		x"02050102",
		x"05010205",
		x"03010503",
		x"01050301",
		x"05030105",
		x"03010503",
		x"01050301",
		x"05030105",
		x"01010301",
		x"01030101",
		x"03010103",
		x"01010301",
		x"01030101",
		x"03010103",
		x"01010301",
		x"01030101",
		x"03010103",
		x"01010301",
		x"01030101",
		x"03010103",
		x"01010301",
		x"01030101",
		x"03010103",
		x"01010301",
		x"01030101",
		x"03010103",
		x"01010301",
		x"01030101",
		x"03010103",
		x"01010301",
		x"01030101",
		x"03010103",
		x"40000440",
		x"00044000",
		x"04400004",
		x"40000440",
		x"00044000",
		x"04400004",
		x"40000440",
		x"00044000",
		x"04400004",
		x"40000440",
		x"00044000",
		x"04400004",
		x"00030400",
		x"03040003",
		x"04000304",
		x"00030400",
		x"03040003",
		x"04000304",
		x"00030400",
		x"03040003",
		x"04000304",
		x"00030400",
		x"03040003",
		x"04000304",
		x"00010200",
		x"01020001",
		x"02000102",
		x"00010200",
		x"01020001",
		x"02000102",
		x"00010200",
		x"01020001",
		x"02000102",
		x"00010200",
		x"01020001",
		x"02000102",
		x"00010200",
		x"01020001",
		x"02000102",
		x"00010200",
		x"01020001",
		x"02000102",
		x"00010200",
		x"01020001",
		x"02000102",
		x"00010200",
		x"01020001",
		x"02000102",
		x"00010200",
		x"01020001",
		x"02000102",
		x"00010200",
		x"01020001",
		x"02000102",
		x"00010200",
		x"01020001",
		x"02000102",
		x"00010200",
		x"01020001",
		x"02000102",
		x"00010200",
		x"01020001",
		x"02000102",
		x"00010200",
		x"01020001",
		x"02000102",
		x"00010200",
		x"01020001",
		x"02000102",
		x"00010200",
		x"01020001",
		x"02000102",
		x"00020300",
		x"02030002",
		x"03000203",
		x"00020300",
		x"02030002",
		x"03000203",
		x"00020300",
		x"02030002",
		x"03000203",
		x"00020300",
		x"02030002",
		x"03000203",
		x"00020300",
		x"02030002",
		x"03000203",
		x"00020300",
		x"02030002",
		x"03000203",
		x"00020300",
		x"02030002",
		x"03000203",
		x"00020300",
		x"02030002",
		x"03000203",
		x"00040500",
		x"04050004",
		x"05000405",
		x"00040500",
		x"04050004",
		x"05000405",
		x"00050500",
		x"05050005",
		x"05000505",
		x"00050500",
		x"05050005",
		x"05000505",
		x"09010709",
		x"01070103",
		x"07010307",
		x"0a01070a",
		x"01070008",
		x"07000807",
		x"00090700",
		x"0907000c",
		x"08000d08",
		x"02030804",
		x"0208000e",
		x"08000f08",
		x"05020905",
		x"02090e01",
		x"090e0109",
		x"02040a10",
		x"010a0f01",
		x"090f0109",
		x"000b0c08",
		x"020c0403",
		x"0c000a0c",
		x"02040c07",
		x"020c1501",
		x"0c14010c",
		x"00090c13",
		x"010c1201",
		x"0c01050c",
		x"03030c00",
		x"080c0602",
		x"0c11010c",
		x"0a020d09",
		x"020d0503",
		x"0d03040d",
		x"02050d01",
		x"070d0106",
		x"0d000f0d",
		x"000e0d00",
		x"0d0d000c",
		x"0d1a010d",
		x"19010d18",
		x"010d1701",
		x"0d16010d",
		x"001f0e00",
		x"1e0e001d",
		x"0e001c0e",
		x"001b0e00",
		x"1a0e0019",
		x"0e00180e",
		x"00170e00",
		x"160e0015",
		x"0e00140e",
		x"00130e00",
		x"120e0011",
		x"0e00100e",
		x"00280f00",
		x"270f0026",
		x"0f00250f",
		x"00240f00",
		x"230f0022",
		x"0f00210f",
		x"00200f01",
		x"0e0f010d",
		x"0f010c0f",
		x"010b0f01",
		x"0a0f0109",
		x"0f01080f",
		x"01121001",
		x"11100110",
		x"10010f10",
		x"06031010",
		x"02100f02",
		x"100e0210",
		x"0d02100c",
		x"02100b02",
		x"101f0110",
		x"1e01101d",
		x"01101c01",
		x"101b0110",
		x"00070080",
		x"241d3fff",	 --print.c
		x"0c000116",
		x"00000000",
		x"00002021",
		x"0000000c",
		x"00000000",
		x"08000006",
		x"00000000",
		x"0000000c",
		x"00000000",
		x"03e00008",
		x"00000000",
		x"14800007",
		x"3c050000",
		x"24a30584",
		x"24020030",
		x"00602021",
		x"a0a20584",
		x"08000045",
		x"a0600001",
		x"3c02cccc",
		x"3442cccd",
		x"00820019",
		x"00404021",
		x"24a70584",
		x"24060001",
		x"2409000b",
		x"00001810",
		x"000318c2",
		x"000310c0",
		x"00031840",
		x"00621821",
		x"00831823",
		x"24630030",
		x"0800002f",
		x"a0a30584",
		x"00880019",
		x"24c60001",
		x"00001010",
		x"000210c2",
		x"000218c0",
		x"00021040",
		x"00431021",
		x"00821023",
		x"24420030",
		x"10c90006",
		x"a0e20000",
		x"00880019",
		x"00001010",
		x"000220c2",
		x"1480fff1",
		x"24e70001",
		x"3c020000",
		x"24420578",
		x"24c4ffff",
		x"3c030000",
		x"00822821",
		x"24630584",
		x"00c21021",
		x"08000040",
		x"a0400000",
		x"9062ffff",
		x"2484ffff",
		x"a0a20001",
		x"24630001",
		x"0481fffb",
		x"24a5ffff",
		x"3c020000",
		x"24440578",
		x"03e00008",
		x"00801021",
		x"3c020000",
		x"24050030",
		x"2443056c",
		x"a045056c",
		x"24020078",
		x"a0620001",
		x"1480000a",
		x"a060000a",
		x"a0650009",
		x"a0650002",
		x"a0650003",
		x"a0650004",
		x"a0650005",
		x"a0650006",
		x"a0650007",
		x"08000068",
		x"a0650008",
		x"3c020000",
		x"24450575",
		x"3c020000",
		x"2447056d",
		x"3082000f",
		x"24460030",
		x"24430057",
		x"2c42000a",
		x"10400003",
		x"00000000",
		x"08000065",
		x"a0a60000",
		x"a0a30000",
		x"24a5ffff",
		x"14a7fff5",
		x"00042102",
		x"3c020000",
		x"03e00008",
		x"2442056c",
		x"04810002",
		x"00801021",
		x"00041023",
		x"03e00008",
		x"00000000",
		x"30820001",
		x"00021023",
		x"3042b400",
		x"00042043",
		x"00822026",
		x"14c00002",
		x"0086001a",
		x"0007000d",
		x"00001010",
		x"03e00008",
		x"00451021",
		x"03e00008",
		x"00851021",
		x"03e00008",
		x"00851023",
		x"00801021",
		x"08000084",
		x"00801821",
		x"a0650000",
		x"24630001",
		x"1cc0fffd",
		x"24c6ffff",
		x"03e00008",
		x"00000000",
		x"0481003c",
		x"00801021",
		x"3c020000",
		x"2447055c",
		x"3c026666",
		x"00042823",
		x"344a6667",
		x"00003021",
		x"24090030",
		x"080000a3",
		x"2408000c",
		x"080000a0",
		x"a0e90000",
		x"00aa0018",
		x"00001010",
		x"00021083",
		x"00431023",
		x"00021840",
		x"000220c0",
		x"00641821",
		x"00a31823",
		x"24630030",
		x"00402821",
		x"a0e30000",
		x"24c60001",
		x"10c80006",
		x"24e70001",
		x"00051fc3",
		x"14a0fff0",
		x"28c20005",
		x"1440ffec",
		x"00000000",
		x"3c030000",
		x"2463054c",
		x"3c020000",
		x"24c40001",
		x"00604021",
		x"2447055c",
		x"00c31821",
		x"00002821",
		x"24090004",
		x"2406002e",
		x"080000be",
		x"a0600002",
		x"14a90003",
		x"00000000",
		x"a0460000",
		x"2484ffff",
		x"90e30000",
		x"00881021",
		x"24a50001",
		x"a0430000",
		x"2484ffff",
		x"24e70001",
		x"0481fff5",
		x"00881021",
		x"3c030000",
		x"2402002d",
		x"2465054c",
		x"08000104",
		x"a062054c",
		x"10400005",
		x"3c040000",
		x"00402821",
		x"2487055c",
		x"080000e5",
		x"00003021",
		x"2483055c",
		x"24020030",
		x"00602821",
		x"a082055c",
		x"08000104",
		x"a0600001",
		x"24020030",
		x"080000e1",
		x"a0e20000",
		x"3c026666",
		x"34426667",
		x"00a20018",
		x"00001010",
		x"00021083",
		x"00431023",
		x"00021840",
		x"000220c0",
		x"00641821",
		x"00a31823",
		x"24630030",
		x"00402821",
		x"a0e30000",
		x"24c60001",
		x"2402000c",
		x"10c20006",
		x"24e70001",
		x"00051fc3",
		x"14a0ffed",
		x"28c20005",
		x"1440ffe8",
		x"00000000",
		x"3c030000",
		x"2463054c",
		x"3c020000",
		x"00c02021",
		x"00604021",
		x"2447055c",
		x"00c31821",
		x"00002821",
		x"24090004",
		x"2406002e",
		x"08000100",
		x"a0600001",
		x"14a90003",
		x"00000000",
		x"a0460000",
		x"2484ffff",
		x"90e30000",
		x"00881021",
		x"24a50001",
		x"a0430000",
		x"2484ffff",
		x"24e70001",
		x"0481fff5",
		x"00881021",
		x"3c020000",
		x"2445054c",
		x"03e00008",
		x"00a01021",
		x"00801821",
		x"80a20000",
		x"24a50001",
		x"a0620000",
		x"1440fffc",
		x"24630001",
		x"03e00008",
		x"00801021",
		x"00801821",
		x"80620000",
		x"00000000",
		x"1440fffd",
		x"24630001",
		x"00641023",
		x"03e00008",
		x"2442ffff",
		x"3c050000",
		x"27bdffe8",
		x"24a50520",
		x"24040004",
		x"00003021",
		x"00003821",
		x"afb00010",
		x"afbf0014",
		x"0c000008",
		x"24100013",
		x"3c050000",
		x"24a50590",
		x"24040002",
		x"00003021",
		x"0c000008",
		x"00003821",
		x"00002821",
		x"00003021",
		x"00003821",
		x"1040fff6",
		x"24040003",
		x"0c000008",
		x"2610ffff",
		x"0c00000c",
		x"00402021",
		x"00402821",
		x"24040004",
		x"00003021",
		x"0c000008",
		x"00003821",
		x"0601ffec",
		x"3c050000",
		x"3c050000",
		x"24a50538",
		x"24040004",
		x"00003021",
		x"0c000008",
		x"00003821",
		x"00002021",
		x"00002821",
		x"00003021",
		x"0c000008",
		x"00003821",
		x"1040fffb",
		x"00002021",
		x"8fbf0014",
		x"8fb00010",
		x"00001021",
		x"03e00008",
		x"27bd0018",
		x"4d504547",
		x"20546173",
		x"6b205052",
		x"494e5420",
		x"73746172",
		x"743a0000",
		x"456e6420",
		x"5461736b",
		x"2045202d",
		x"204d5045",
		x"47000000",
		x"241d3fff",	 --start.c
		x"0c000116",
		x"00000000",
		x"00002021",
		x"0000000c",
		x"00000000",
		x"08000006",
		x"00000000",
		x"0000000c",
		x"00000000",
		x"03e00008",
		x"00000000",
		x"14800007",
		x"3c050000",
		x"24a308a4",
		x"24020030",
		x"00602021",
		x"a0a208a4",
		x"08000045",
		x"a0600001",
		x"3c02cccc",
		x"3442cccd",
		x"00820019",
		x"00404021",
		x"24a708a4",
		x"24060001",
		x"2409000b",
		x"00001810",
		x"000318c2",
		x"000310c0",
		x"00031840",
		x"00621821",
		x"00831823",
		x"24630030",
		x"0800002f",
		x"a0a308a4",
		x"00880019",
		x"24c60001",
		x"00001010",
		x"000210c2",
		x"000218c0",
		x"00021040",
		x"00431021",
		x"00821023",
		x"24420030",
		x"10c90006",
		x"a0e20000",
		x"00880019",
		x"00001010",
		x"000220c2",
		x"1480fff1",
		x"24e70001",
		x"3c020000",
		x"24420898",
		x"24c4ffff",
		x"3c030000",
		x"00822821",
		x"246308a4",
		x"00c21021",
		x"08000040",
		x"a0400000",
		x"9062ffff",
		x"2484ffff",
		x"a0a20001",
		x"24630001",
		x"0481fffb",
		x"24a5ffff",
		x"3c020000",
		x"24440898",
		x"03e00008",
		x"00801021",
		x"3c020000",
		x"24050030",
		x"2443088c",
		x"a045088c",
		x"24020078",
		x"a0620001",
		x"1480000a",
		x"a060000a",
		x"a0650009",
		x"a0650002",
		x"a0650003",
		x"a0650004",
		x"a0650005",
		x"a0650006",
		x"a0650007",
		x"08000068",
		x"a0650008",
		x"3c020000",
		x"24450895",
		x"3c020000",
		x"2447088d",
		x"3082000f",
		x"24460030",
		x"24430057",
		x"2c42000a",
		x"10400003",
		x"00000000",
		x"08000065",
		x"a0a60000",
		x"a0a30000",
		x"24a5ffff",
		x"14a7fff5",
		x"00042102",
		x"3c020000",
		x"03e00008",
		x"2442088c",
		x"04810002",
		x"00801021",
		x"00041023",
		x"03e00008",
		x"00000000",
		x"30820001",
		x"00021023",
		x"3042b400",
		x"00042043",
		x"00822026",
		x"14c00002",
		x"0086001a",
		x"0007000d",
		x"00001010",
		x"03e00008",
		x"00451021",
		x"03e00008",
		x"00851021",
		x"03e00008",
		x"00851023",
		x"00801021",
		x"08000084",
		x"00801821",
		x"a0650000",
		x"24630001",
		x"1cc0fffd",
		x"24c6ffff",
		x"03e00008",
		x"00000000",
		x"0481003c",
		x"00801021",
		x"3c020000",
		x"2447087c",
		x"3c026666",
		x"00042823",
		x"344a6667",
		x"00003021",
		x"24090030",
		x"080000a3",
		x"2408000c",
		x"080000a0",
		x"a0e90000",
		x"00aa0018",
		x"00001010",
		x"00021083",
		x"00431023",
		x"00021840",
		x"000220c0",
		x"00641821",
		x"00a31823",
		x"24630030",
		x"00402821",
		x"a0e30000",
		x"24c60001",
		x"10c80006",
		x"24e70001",
		x"00051fc3",
		x"14a0fff0",
		x"28c20005",
		x"1440ffec",
		x"00000000",
		x"3c030000",
		x"2463086c",
		x"3c020000",
		x"24c40001",
		x"00604021",
		x"2447087c",
		x"00c31821",
		x"00002821",
		x"24090004",
		x"2406002e",
		x"080000be",
		x"a0600002",
		x"14a90003",
		x"00000000",
		x"a0460000",
		x"2484ffff",
		x"90e30000",
		x"00881021",
		x"24a50001",
		x"a0430000",
		x"2484ffff",
		x"24e70001",
		x"0481fff5",
		x"00881021",
		x"3c030000",
		x"2402002d",
		x"2465086c",
		x"08000104",
		x"a062086c",
		x"10400005",
		x"3c040000",
		x"00402821",
		x"2487087c",
		x"080000e5",
		x"00003021",
		x"2483087c",
		x"24020030",
		x"00602821",
		x"a082087c",
		x"08000104",
		x"a0600001",
		x"24020030",
		x"080000e1",
		x"a0e20000",
		x"3c026666",
		x"34426667",
		x"00a20018",
		x"00001010",
		x"00021083",
		x"00431023",
		x"00021840",
		x"000220c0",
		x"00641821",
		x"00a31823",
		x"24630030",
		x"00402821",
		x"a0e30000",
		x"24c60001",
		x"2402000c",
		x"10c20006",
		x"24e70001",
		x"00051fc3",
		x"14a0ffed",
		x"28c20005",
		x"1440ffe8",
		x"00000000",
		x"3c030000",
		x"2463086c",
		x"3c020000",
		x"00c02021",
		x"00604021",
		x"2447087c",
		x"00c31821",
		x"00002821",
		x"24090004",
		x"2406002e",
		x"08000100",
		x"a0600001",
		x"14a90003",
		x"00000000",
		x"a0460000",
		x"2484ffff",
		x"90e30000",
		x"00881021",
		x"24a50001",
		x"a0430000",
		x"2484ffff",
		x"24e70001",
		x"0481fff5",
		x"00881021",
		x"3c020000",
		x"2445086c",
		x"03e00008",
		x"00a01021",
		x"00801821",
		x"80a20000",
		x"24a50001",
		x"a0620000",
		x"1440fffc",
		x"24630001",
		x"03e00008",
		x"00801021",
		x"00801821",
		x"80620000",
		x"00000000",
		x"1440fffd",
		x"24630001",
		x"00641023",
		x"03e00008",
		x"2442ffff",
		x"3c050000",
		x"27bdffe0",
		x"24a50638",
		x"24040004",
		x"00003021",
		x"00003821",
		x"afbf001c",
		x"afb20018",
		x"afb10014",
		x"0c000008",
		x"afb00010",
		x"00002821",
		x"00003021",
		x"00003821",
		x"0c000008",
		x"24040003",
		x"0c00000c",
		x"00402021",
		x"00402821",
		x"24040004",
		x"00003021",
		x"0c000008",
		x"00003821",
		x"3c020000",
		x"2443066c",
		x"3c020000",
		x"244408b4",
		x"3c020000",
		x"2445086c",
		x"8c620000",
		x"24630004",
		x"ac820000",
		x"1465fffc",
		x"24840004",
		x"24030080",
		x"3c020000",
		x"ac4308b0",
		x"00009021",
		x"24040003",
		x"00002821",
		x"00003021",
		x"0c000008",
		x"00003821",
		x"00408821",
		x"3c050000",
		x"24a508b0",
		x"24040001",
		x"24060002",
		x"0c000008",
		x"00003821",
		x"1040fffa",
		x"3c050000",
		x"24040003",
		x"00002821",
		x"00003021",
		x"0c000008",
		x"00003821",
		x"3c050000",
		x"24a50650",
		x"00003021",
		x"00003821",
		x"24040004",
		x"0c000008",
		x"00408021",
		x"0c00000c",
		x"02202021",
		x"00402821",
		x"24040004",
		x"00003021",
		x"0c000008",
		x"00003821",
		x"3c050000",
		x"24a50654",
		x"00003021",
		x"00003821",
		x"0c000008",
		x"24040004",
		x"0c00000c",
		x"02002021",
		x"00402821",
		x"24040004",
		x"00003021",
		x"0c000008",
		x"00003821",
		x"26520001",
		x"24020014",
		x"1642ffd0",
		x"24040003",
		x"00002821",
		x"00003021",
		x"00003821",
		x"0c000008",
		x"24040003",
		x"0c00000c",
		x"00402021",
		x"00402821",
		x"24040004",
		x"00003021",
		x"0c000008",
		x"00003821",
		x"3c050000",
		x"24a50658",
		x"24040004",
		x"00003021",
		x"0c000008",
		x"00003821",
		x"00002021",
		x"00002821",
		x"00003021",
		x"0c000008",
		x"00003821",
		x"1040fffb",
		x"00002021",
		x"8fbf001c",
		x"8fb20018",
		x"8fb10014",
		x"8fb00010",
		x"00001021",
		x"03e00008",
		x"27bd0020",
		x"4d504547",
		x"20546173",
		x"6b204120",
		x"73746172",
		x"743a2020",
		x"00000000",
		x"54310000",
		x"54320000",
		x"456e6420",
		x"5461736b",
		x"2041202d",
		x"204d5045",
		x"47000000",
		x"000000fa",
		x"000000b8",
		x"00000020",
		x"00000005",
		x"00000020",
		x"00000020",
		x"00000002",
		x"00000038",
		x"00000020",
		x"0000007e",
		x"0000007f",
		x"000000f0",
		x"00000010",
		x"0000003f",
		x"00000054",
		x"0000008a",
		x"00000008",
		x"0000001f",
		x"000000a8",
		x"00000000",
		x"00000042",
		x"00000000",
		x"000000d2",
		x"00000080",
		x"0000003e",
		x"000000f6",
		x"000000a0",
		x"0000000e",
		x"0000003e",
		x"00000045",
		x"00000080",
		x"0000003e",
		x"000000c0",
		x"00000007",
		x"000000bc",
		x"00000079",
		x"00000000",
		x"0000003f",
		x"000000c2",
		x"00000028",
		x"000000b2",
		x"0000003f",
		x"0000000e",
		x"00000078",
		x"000000be",
		x"00000088",
		x"0000009c",
		x"00000082",
		x"00000017",
		x"000000fc",
		x"00000011",
		x"000000bc",
		x"00000085",
		x"00000074",
		x"00000027",
		x"000000a7",
		x"000000f2",
		x"00000024",
		x"00000002",
		x"000000ce",
		x"0000005f",
		x"000000c7",
		x"000000ce",
		x"0000004e",
		x"000000a7",
		x"0000003c",
		x"00000073",
		x"000000b6",
		x"00000031",
		x"00000001",
		x"00000001",
		x"00000001",
		x"00000001",
		x"00000001",
		x"00000001",
		x"00000001",
		x"00000001",
		x"00000001",
		x"00000001",
		x"00000001",
		x"00000001",
		x"00000001",
		x"00000001",
		x"00000001",
		x"00000001",
		x"00000001",
		x"00000001",
		x"00000001",
		x"00000001",
		x"00000001",
		x"00000001",
		x"00000001",
		x"00000001",
		x"00000001",
		x"00000001",
		x"00000001",
		x"00000001",
		x"00000001",
		x"00000001",
		x"00000001",
		x"00000001",
		x"00000001",
		x"00000001",
		x"00000001",
		x"00000001",
		x"00000001",
		x"00000001",
		x"00000001",
		x"00000001",
		x"00000001",
		x"00000001",
		x"00000001",
		x"00000001",
		x"00000001",
		x"00000001",
		x"00000001",
		x"00000001",
		x"00000001",
		x"00000001",
		x"00000001",
		x"00000001",
		x"00000001",
		x"00000001",
		x"00000001",
		x"00000001",
		x"00000001",
		x"00000001",
		x"00000001",
		(others=>'0'));
end memory_pack;
