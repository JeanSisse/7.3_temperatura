library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_misc.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library UNISIM;
use UNISIM.vcomponents.all;

entity ram_master is
	port(clk             : in  std_logic;
        address_a       : in  std_logic_vector(31 downto 2);
        enable_a        : in  std_logic;
        wbe_a           : in  std_logic_vector(3 downto 0);
        data_write_a    : in  std_logic_vector(31 downto 0);
        data_read_a     : out std_logic_vector(31 downto 0);

        address_b       : in  std_logic_vector(31 downto 2);
        enable_b        : in  std_logic;
        wbe_b           : in  std_logic_vector(3 downto 0);
        data_write_b    : in  std_logic_vector(31 downto 0);
        data_read_b     : out std_logic_vector(31 downto 0));
end; --entity ram     

architecture ram_master of ram_master is
signal enable_a_lo       : std_logic;
signal wbe_a_lo          : std_logic_vector(3 downto 0);
signal data_write_a_lo   : std_logic_vector(31 downto 0);
signal data_read_a_lo    : std_logic_vector(31 downto 0);
signal enable_b_lo       : std_logic;
signal wbe_b_lo          : std_logic_vector(3 downto 0);
signal data_read_b_lo    : std_logic_vector(31 downto 0);
signal enable_a_hi       : std_logic;
signal wbe_a_hi          : std_logic_vector(3 downto 0);
signal data_read_a_hi   : std_logic_vector(31 downto 0);
signal enable_b_hi       : std_logic;
signal wbe_b_hi          : std_logic_vector(3 downto 0);
signal data_read_b_hi    : std_logic_vector(31 downto 0);
signal address_a_reg     : std_logic_vector(31 downto 2);
signal address_b_reg     : std_logic_vector(31 downto 2);
signal enable_a_lo_256       : std_logic;
signal wbe_a_lo_256          : std_logic_vector(3 downto 0);
signal data_write_a_lo_256   : std_logic_vector(31 downto 0);
signal data_read_a_lo_256    : std_logic_vector(31 downto 0);
signal enable_b_lo_256       : std_logic;
signal wbe_b_lo_256          : std_logic_vector(3 downto 0);
signal data_read_b_lo_256    : std_logic_vector(31 downto 0);
signal enable_a_hi_256       : std_logic;
signal wbe_a_hi_256          : std_logic_vector(3 downto 0);
signal data_read_a_hi_256   : std_logic_vector(31 downto 0);
signal enable_b_hi_256       : std_logic;
signal wbe_b_hi_256          : std_logic_vector(3 downto 0);
signal data_read_b_hi_256    : std_logic_vector(31 downto 0);
signal enable_a_lo_512       : std_logic;
signal wbe_a_lo_512          : std_logic_vector(3 downto 0);
signal data_write_a_lo_512   : std_logic_vector(31 downto 0);
signal data_read_a_lo_512    : std_logic_vector(31 downto 0);
signal enable_b_lo_512       : std_logic;
signal wbe_b_lo_512          : std_logic_vector(3 downto 0);
signal data_read_b_lo_512    : std_logic_vector(31 downto 0);
signal enable_a_hi_512       : std_logic;
signal wbe_a_hi_512          : std_logic_vector(3 downto 0);
signal data_read_a_hi_512   : std_logic_vector(31 downto 0);
signal enable_b_hi_512       : std_logic;
signal wbe_b_hi_512          : std_logic_vector(3 downto 0);
signal data_read_b_hi_512    : std_logic_vector(31 downto 0);
signal enable_a_lo_512_2       : std_logic;
signal wbe_a_lo_512_2          : std_logic_vector(3 downto 0);
signal data_write_a_lo_512_2   : std_logic_vector(31 downto 0);
signal data_read_a_lo_512_2    : std_logic_vector(31 downto 0);
signal enable_b_lo_512_2       : std_logic;
signal wbe_b_lo_512_2          : std_logic_vector(3 downto 0);
signal data_read_b_lo_512_2    : std_logic_vector(31 downto 0);
signal enable_a_hi_512_2       : std_logic;
signal wbe_a_hi_512_2          : std_logic_vector(3 downto 0);
signal data_read_a_hi_512_2   : std_logic_vector(31 downto 0);
signal enable_b_hi_512_2       : std_logic;
signal wbe_b_hi_512_2          : std_logic_vector(3 downto 0);
signal data_read_b_hi_512_2    : std_logic_vector(31 downto 0);
begin
process(clk)
begin
if rising_edge(clk) then
	address_a_reg <= address_a;
	address_b_reg <= address_b;
	end if;
end process;
data_read_a <= data_read_a_lo when (address_a_reg < x"0001000"&"00") else
data_read_a_hi when ((address_a_reg >= x"0001000"&"00") and (address_a_reg < x"0002000"&"00")) else 
data_read_a_lo_256 when ((address_a_reg >= x"0002000"&"00") and (address_a_reg < x"0003000"&"00")) else 
data_read_a_hi_256 when ((address_a_reg >= x"0003000"&"00") and (address_a_reg < x"0004000"&"00")) else 
data_read_a_lo_512 when ((address_a_reg >= x"0004000"&"00") and (address_a_reg < x"0005000"&"00")) else 
data_read_a_hi_512 when ((address_a_reg >= x"0005000"&"00") and (address_a_reg < x"0006000"&"00")) else 
data_read_a_lo_512_2 when ((address_a_reg >= x"0006000"&"00") and (address_a_reg < x"0007000"&"00")) else 
data_read_a_hi_512_2 when ((address_a_reg >= x"0007000"&"00") and (address_a_reg < x"0008000"&"00")); 
data_read_b <= data_read_b_lo when (address_b_reg < x"0001000"&"00") else
data_read_b_hi when ((address_b_reg >= x"0001000"&"00") and (address_b_reg < x"0002000"&"00")) else
data_read_b_lo_256 when ((address_b_reg >= x"0002000"&"00") and (address_a_reg < x"0003000"&"00")) else 
data_read_b_hi_256 when ((address_b_reg >= x"0003000"&"00") and (address_b_reg< x"0004000"&"00")) else 
data_read_b_lo_512 when ((address_b_reg >= x"0004000"&"00") and (address_b_reg< x"0005000"&"00")) else 
data_read_b_hi_512 when ((address_b_reg >= x"0005000"&"00") and (address_b_reg< x"0006000"&"00")) else 
data_read_b_lo_512_2 when ((address_b_reg >= x"0006000"&"00") and (address_b_reg< x"0007000"&"00")) else 
data_read_b_hi_512_2 when ((address_b_reg >= x"0007000"&"00") and (address_b_reg< x"0008000"&"00")); 
enable_a_lo <= enable_a when (address_a < x"0001000"&"00") else '0';
enable_b_lo <= enable_b when (address_b < x"0001000"&"00") else '0';
enable_a_hi <= enable_a when ((address_a >= x"0001000"&"00") and (address_a < x"0002000"&"00")) else '0';
enable_b_hi <= enable_b when ((address_b >= x"0001000"&"00") and (address_b < x"0002000"&"00")) else '0';
enable_a_lo_256 <= enable_a when ((address_a >= x"0002000"&"00") and (address_a < x"0003000"&"00")) else '0';
enable_b_lo_256 <= enable_b when ((address_b >= x"0002000"&"00") and (address_b < x"0003000"&"00")) else '0';
enable_a_hi_256 <= enable_a when ((address_a >= x"0003000"&"00") and (address_a < x"0004000"&"00")) else '0';
enable_b_hi_256 <= enable_b when ((address_b >= x"0003000"&"00") and (address_b < x"0004000"&"00")) else '0';
enable_a_lo_512 <= enable_a when ((address_a >= x"0004000"&"00") and (address_a < x"0005000"&"00")) else '0';
enable_b_lo_512 <= enable_b when ((address_b >= x"0004000"&"00") and (address_b < x"0005000"&"00")) else '0';
enable_a_hi_512 <= enable_a when ((address_a >= x"0005000"&"00") and (address_a < x"0006000"&"00")) else '0';
enable_b_hi_512 <= enable_b when ((address_b >= x"0005000"&"00") and (address_b < x"0006000"&"00")) else '0';
enable_a_lo_512_2 <= enable_a when ((address_a >= x"0006000"&"00") and (address_a < x"0007000"&"00")) else '0';
enable_b_lo_512_2 <= enable_b when ((address_b >= x"0006000"&"00") and (address_b < x"0007000"&"00")) else '0';
enable_a_hi_512_2 <= enable_a when ((address_a >= x"0007000"&"00") and (address_a < x"0008000"&"00")) else '0';
enable_b_hi_512_2 <= enable_b when ((address_b >= x"0007000"&"00") and (address_b < x"0008000"&"00")) else '0';
wbe_a_lo <= wbe_a when  enable_a_lo='1' else x"0";
wbe_a_hi <= wbe_a when  enable_a_hi='1' else x"0";
wbe_b_lo <= wbe_b when  enable_b_lo='1' else x"0";
wbe_b_hi <= wbe_b when  enable_b_hi='1' else x"0";
wbe_a_lo_256 <= wbe_a when  enable_a_lo_256='1' else x"0";
wbe_a_hi_256 <= wbe_a when  enable_a_hi_256='1' else x"0";
wbe_b_lo_256 <= wbe_b when  enable_b_lo_256='1' else x"0";
wbe_b_hi_256 <= wbe_b when  enable_b_hi_256='1' else x"0";
wbe_a_lo_512 <= wbe_a when  enable_a_lo_512='1' else x"0";
wbe_a_hi_512 <= wbe_a when  enable_a_hi_512='1' else x"0";
wbe_b_lo_512 <= wbe_b when  enable_b_lo_512='1' else x"0";
wbe_b_hi_512 <= wbe_b when  enable_b_hi_512='1' else x"0";
wbe_a_lo_512_2 <= wbe_a when  enable_a_lo_512_2='1' else x"0";
wbe_a_hi_512_2 <= wbe_a when  enable_a_hi_512_2='1' else x"0";
wbe_b_lo_512_2 <= wbe_b when  enable_b_lo_512_2='1' else x"0";
wbe_b_hi_512_2 <= wbe_b when  enable_b_hi_512_2='1' else x"0";



ram_bit_0_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"ED39BA795990D275FB4A6E96ACC4731DEA4598B0AFB54867F6EE4618C3749807",
INIT_01 => X"58A0047D8607944AC7DA180001ECA2444042106208408208C20022E9173734B3",
INIT_02 => X"8B1E49562021F8051500147A0E162923024F28000415F5787B09FBF999BB1EFC",
INIT_03 => X"1013BF028A959403C06A23A147723C01E140088280C4CF6996088862C7922221",
INIT_04 => X"781A003802015D9078011DE20340699198600000B08694916434804825241311",
INIT_05 => X"2CA000587E10C880036A3103C00F2000E1E0383C00730002B4409845E4425171",
INIT_06 => X"179B48CFF95DCF9EF730E1C3BB731138AF7B888025340C0888430047040FEE18",
INIT_07 => X"AF155113160400185F87C1F05707D415E664A6E7C5551EBE783060CEB164833F",
INIT_08 => X"4D7E40002B7AE005FDB47600208229010C6101001EFE198C96B0528202C0DCB4",
INIT_09 => X"062400608234D864444081048A80CC00062D42D30222108091C107A1DA040267",
INIT_0A => X"204A21008E514844EB5145000255DA599581D3A9583C24351240B58298011308",
INIT_0B => X"E08C4830F81380CE0F89E07A9E0789E07A9E0789E07A9E0789E070CF0184F038",
INIT_0C => X"3A4E9D63EA180EB150CA1CA45C254D4AF4AA414568729139F2A12C0000016110",
INIT_0D => X"F0009E0FC048211E9C11C31F82E4A000890022B827EB52F52347F174E93A749D",
INIT_0E => X"F0009E0FCC42EFDFBF0AE03080E2AEB2E0F1F80FA97FE0F0009E0FC40FA97FE0",
INIT_0F => X"0231F0BD9E3FC08FEBD6F661C0E008C3CB5F040FAB3FE0F0009E0FC40FAB3FE0",
INIT_10 => X"20180309A0F83BE2B87C7C42EFDFBF187806013879BA878FE807F65FBF12E038",
INIT_11 => X"0BE9F01FC8B38C2098DAE007F323A0C83136B248831ACBFC8BBDCAB779BC699F",
INIT_12 => X"004C72BEC800FE7464290626D7003F9947184131B59003FFEC07F00003F01FB9",
INIT_13 => X"A0FFDA2A3C0202B8776A2FA7F023F7D065703080E29F1B2BE9F8A27E6E915C0E",
INIT_14 => X"016C2D25E52630BB1AE49C2BA7F98D6F846DFC0C2352A0024B83F07F198BE9F8",
INIT_15 => X"749D2749D2749D2749D2749D2749F285F25D2C500815A5522CB5A4B400000CD4",
INIT_16 => X"49D2749D2749D2749D2749D2749D2749D2749D2749D2749D2749D2749D2749D2",
INIT_17 => X"9D2749D2749D2749D2749D2749D2749D2749D2749D2749D2749D2749D2749D27",
INIT_18 => X"31C136AD8E9B562BA39E2600654BA800000000000000000749D2749D2749D274",
INIT_19 => X"4104104104104104104104104104104104104104104104109C83B8E38E2ABE71",
INIT_1A => X"0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0410410410",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000007C3E1F0F87C3E1F0F87C3E1F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000187FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"BAF7FFD55EF007FD75EFFFAE97555557BD75EF5D000000000000000000000000",
INIT_1F => X"000AA843FE00AAFBE8B45AA803DFEFA28428B455D0017410A28428AAAA2FBD54",
INIT_20 => X"FEBAA2D5401450051401555D7FC0145F7AEBFFFF08002AA10A2AABFEAAA2FFC0",
INIT_21 => X"D755555517FFEFA280021FF082E974AA5D7BFFE000804000BAAAAAAAB45557FF",
INIT_22 => X"EA8B45005168A10AA8028A10087FD7410557FC21555D51574AAA2FFE8B455D7B",
INIT_23 => X"AE95410AA80000005D003FEAAFFAEBFE00A2803FEBA002A820AA0800174BA5D2",
INIT_24 => X"2AEA8A10000417410A2FFE8BEFF7FFE8B45FFFBC00005D003FF45557FC01FFFF",
INIT_25 => X"00000000000000000000000000000000000000557DF5500003DFEFFF84175EFA",
INIT_26 => X"5F524AFE38B780154BAFFF1D54AF0075D75EFEBAE9554540754717F1F8000000",
INIT_27 => X"50B6AABDE12BEA0AF010B7D1F8F47E00A2DB45AA8A3AFD7B68E2AB78550E1255",
INIT_28 => X"E9257F1E816D557095EAAA2D1401D500002A150038038E285D7F78FD7000B6AB",
INIT_29 => X"5A87AAD178A8002D1D21C5E8257D5C7AA854008700249243A412EBFF5542A43F",
INIT_2A => X"52A82000E3A5D2150AB8F401471EDBC0B680900AAF52B474385D75C502D15754",
INIT_2B => X"FD7E9541242FE920AD082E10A28F6A150012A2F02AFFDF40E85F475451D502D1",
INIT_2C => X"0550E87B7A405B52AAD152BD00151EAFEDB52E3F1EFFFF485A2DA3D5D24BD417",
INIT_2D => X"57F40545850000000000000000000000000000000000000000000005AAF55508",
INIT_2E => X"F7AEAABFF5D2A81151FB8635A02FA69574BAF7D5555AF0D79D55FFA2AC974450",
INIT_2F => X"8D46F6ABE7082AAAAF2FAC77FE00FF16565B2FA9075F4F7B3EBDF50FEAEAAB55",
INIT_30 => X"56803CE3AEB038662E5D81406014D5D51F5E08A394003A908B8410E707EF34A0",
INIT_31 => X"4AF0151555AF58794040077D774FAE8C798A11A0EAEF75F7AA84001A7052C952",
INIT_32 => X"4E1870108B11020AD4AA05542A0A05051023F9A9D57B63BFBF906CB45FABC095",
INIT_33 => X"F5F0DA6BC9525688C1A2A0C06E9FEE5555BE48AB2A2AE0A0F20C43EAC562245B",
INIT_34 => X"000000FF80F55E25C00A0BA7FBED407A97F6F35F498B96BEB12DAAB77558ABD5",
INIT_35 => X"8000000FF8000000FF8000000FF8000000FF8000000FF8000000FF8000000FF8",
INIT_36 => X"00000000000000000000000000FF8000000FF8000000FF8000000FF8000000FF",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000008000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(0),        -- Port A data input
DOA(0)   => data_read_a_lo(0),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(0),        -- Port B data input
DOB(0)   => data_read_b_lo(0),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_1_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"212C001411984004084D000508C53810A03D1450E839B003342114428A000803",
INIT_01 => X"08000010400A0008010600000084005000400002000000000000000000140000",
INIT_02 => X"C084484000002014400205851002007030450E0000A606C8C44CB4C6666C00E0",
INIT_03 => X"CCF7CE0002058001000000800240200001018CA1800001091408463061120118",
INIT_04 => X"082800100000000040000900010000100040000000008411600401C02100000C",
INIT_05 => X"10800202080422000020012200000000810000200000000004020C00200011A0",
INIT_06 => X"56BDBFBC48C315A8660C18305750C008940D8000011000820001000104050004",
INIT_07 => X"8B4344400004000150248912154404C6060A2FE24555013E13060C158AC97F01",
INIT_08 => X"00082080087A000559102400200281000469000008B000000090108000400430",
INIT_09 => X"0000000000001004140545402820020000010010208000008041060008200001",
INIT_0A => X"2102210182004840007845004044020000200080080844200000048088000000",
INIT_0B => X"48800000190191064620646A06468064680646A0646A06468064690321503234",
INIT_0C => X"02008100200800A1100707040101E20BE0B002605C1C110848200C0000000800",
INIT_0D => X"F000A000C0000012187087010AE4B00000000810010040108104100408020401",
INIT_0E => X"F000A000CC4200002F08E03080000010F18058000003C0F000A000C4000003C0",
INIT_0F => X"000000078808C00000023461C0E00000012704000003C0F000A000C4000003C0",
INIT_10 => X"201803000000240218C0044200001E1878060000000AAC00680000001F10E038",
INIT_11 => X"2100B00048230C200009A0001303204800025200040A00D000000202090C281F",
INIT_12 => X"00000002C9000260640900004D0000904618400012900001EC03F00000000039",
INIT_13 => X"80025A0A3C020000002A8400B00007806070308000000961002880204A901C0E",
INIT_14 => X"000801046004308A185000020128000904285C0C0312A0020000000838810028",
INIT_15 => X"0401004010040100401004010040100010410C002000040280100000000008D0",
INIT_16 => X"4010040100401004010040100401004010040100401004010040100401004010",
INIT_17 => X"0100401004010040100401004010040100401004010040100401004010040100",
INIT_18 => X"48D757DF8A9410218E8A56085142020000000000000000004010040100401004",
INIT_19 => X"555555555555555555555555555554514514514514550431A581924924B02651",
INIT_1A => X"4BA5D2E974BA5D2E974BA5D2E974BA5D2EB75BADD6EB75BADD6EB75555555555",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800005D2E974BA5D2E974BA5D2E97",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000607FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"10AAAABFFFFFF803FE10F7D17FEBA55556AAAAAA800000000000000000000000",
INIT_1F => X"EBAFFD555400557BD54BA5D7FFDF45A2FBD75EFA2AE97555F7FBFFF45FFAE800",
INIT_20 => X"ABEFA2D568A005D5157400AA8028AAAF7FBD54AA002A955555D7FE8ABA082EBF",
INIT_21 => X"FDF55AAFBC0010555540010550417555AA8028BEFAAAE97555082A80000AA802",
INIT_22 => X"BD7410550428ABA5D5168ABA552EBDFEF5D7FEAA00AAAABFEAA007BC0145FFFF",
INIT_23 => X"FFEAB55557FFFEBAAAD568B45A2D5575555D7FC2155F7AEA8BEFAAAA954BA557",
INIT_24 => X"D7BD74000804154BA082ABFF55FFD57DF45F7D568ABAF7AABFFFF082ABFFFFFF",
INIT_25 => X"000000000000000000000000000000000000002EBFFEFA280021FF082E974AA5",
INIT_26 => X"5E175EFF57BF8FC2000BEA4BAE97F78A3FE28E3D17DEAA485FE8E02B50000000",
INIT_27 => X"455571E8A2A087BF8EAAEB8E0016D5D75D54BA5D7BFFF7DA2FFD55EFAAA49554",
INIT_28 => X"157428145A00AA8A2FBD7B6DF6AA28550E10405F7A4AFE38EAA0924921C2FD55",
INIT_29 => X"8E971471C7010B7D168F47400A07A28415A001684104155C5B6DF6DBEFBFAA07",
INIT_2A => X"BFBD7B6A0BF492415FC20105D24AAABF1FFBC7010FF8A38FEF557FEAB78B6AAB",
INIT_2B => X"017EBA4A8EB8F6FFD5FE8B7D557495EAAA2D16D1FDBED56A55557A43DE385FD4",
INIT_2C => X"854008700249243A417FFF41542F5D717FE2AAAA56DEBD17FE3DF7FB7FEBFE38",
INIT_2D => X"07DFCA127B8000000000000000000000000000000000000000000002A3D5C7AA",
INIT_2E => X"AAFBD55FFAA8416545A6FB60F47AF2A00010F78028B15F7823FEAAA2D57DFBA0",
INIT_2F => X"22A38C20B2552E975F758516AAAA0869AAAB8A7C19C55550E8574BA557BFFFEF",
INIT_30 => X"55FFEFBCEE5FBAACB10085EE5DE10A2AEBFF55F7BAAA8565DBAC1112FFAC21A0",
INIT_31 => X"BEA097BEAAFAF2863FA00DD574201E7AD1FFF5575841DE08007FC20480028957",
INIT_32 => X"54FF57EFBFA18D4FBFFF40FF809D4000D7FC00FC5D062BBA05ED5034472A02EA",
INIT_33 => X"7DFBFF6963FCAAA2283CF14050062B0A2F7AE8B5D5D51F5E18ABD5EAFFF2AF95",
INIT_34 => X"000000002CB75F7AA84001A7052C95256807DC31AA8114DE55F5BED201FFFED1",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000008000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(1),        -- Port A data input
DOA(0)   => data_read_a_lo(1),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(1),        -- Port B data input
DOB(0)   => data_read_b_lo(1),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_2_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10E44660018259B2843913100062C98004802322D3E030235201006009B2813",
INIT_01 => X"000AC188084900481C8024A542400340404000720885800802000906E4910204",
INIT_02 => X"82040072AC248C31010204880000007401044C0550200000480E0080001300E0",
INIT_03 => X"0080812C130D0A0D1193088802182142494D218220021100001A8020C1004A00",
INIT_04 => X"090D0AD62824A44A428408540D1610020C6E510818923441A4908B0503404201",
INIT_05 => X"5000A004081122242420480A14A99C428908122144244150906124248C002168",
INIT_06 => X"1400088400450000460000001308890094082015800011012D41D518044C1100",
INIT_07 => X"26731111491C1541324C1114BD880004002040204050413F1400100480000201",
INIT_08 => X"02410582881E0C1511D02082AAAB016A2463288549B044605201D10AE11B0020",
INIT_09 => X"E80394280E40158020B591000800481051241A4A404B5035C60904502054E000",
INIT_0A => X"0102C9E12202EA6014D027C418428E220A5500024808922801A0900A84454458",
INIT_0B => X"4600070110C10D04340043400434A043420434A04342043480434102184021A0",
INIT_0C => X"E9CA34328E44CA1401306100A246000402100C088104010AC8005C5681812B04",
INIT_0D => X"0000A0000801487334E34C1A980001550055481204090A4C01351253A728D194",
INIT_0E => X"0000A000013800004000080000000000500000B01480010000A0000150148001",
INIT_0F => X"0000000608000A500409000800000000012001501480010000A00000B0148001",
INIT_10 => X"1000000000002400000001A100004002000000000000A0000360018040001000",
INIT_11 => X"380001C01048000000090298040440000002400008C400022042004080028000",
INIT_12 => X"0000000009530080880000004813802090000000120C94000200000000000001",
INIT_13 => X"4C000100000000000002E0000950002018000000000001580002508010440000",
INIT_14 => X"7120642000000400015020500004221018000082008000000000000820180002",
INIT_15 => X"5094A5294A5294A52942509425094209461468000822241A03835D88482AB001",
INIT_16 => X"09465094A5294A5294A5294250942509425094A5294A5294A529425094250942",
INIT_17 => X"94650946509465294E5294E5294E5094650946509465294E5294E5294E509465",
INIT_18 => X"080271AE180616A38A18FA204452A7F03F03F07E07E07E05294E5294E5294E50",
INIT_19 => X"20820820820820820820820820820820820820820820490C04102CB2CB2EB2C0",
INIT_1A => X"8944A25128944A25128944A25128944A25128944A25128944A25128208208208",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF1F804A25128944A25128944A2512",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000787FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"AAAA843DFFFAAD1554005D7FD74AA00040015500000000000000000000000000",
INIT_1F => X"F45AAAAA8A10A2AE80010A2AA975FF5D003FE10F7D17FEBAF7D5420AA0855420",
INIT_20 => X"FF45A2AA975EFA2FFD7555FFFBFFF45AAFBC20AAF7D1575EF55517DF555D2EBF",
INIT_21 => X"95555552E974105D517DF55AAAAAABEFAAD1575EFAAAE974AA5D51554BA5D7FF",
INIT_22 => X"E82010F7AABFE10FFD542145FFD5554AA555555555557FE8ABA082EBFFFFAAAE",
INIT_23 => X"FBC0010AA802ABEFAAD540000FFD540000AA802AABAF7FFC2010AAAE821EF552",
INIT_24 => X"A8028BEFAAAE821550851420AA002E800AA08042AB45007FC00BAFFD168BEFF7",
INIT_25 => X"000000000000000000000000000000000000002E80010555540010550417555A",
INIT_26 => X"AE95F40002157F470AABE803AE97A2DF55400557FD54AA1D04001C5150000000",
INIT_27 => X"EF55517DFC5552ABDF45B6AEAFFD5F7A482000BEAE905C755003FE28E3D17DEA",
INIT_28 => X"0BA5FD0154BA5D7BFAF7DA2AE955EFAAA495545E3F5EFF57F7FE80082FFDE105",
INIT_29 => X"8AAF082AB8EAAEB8E0016D5D2A924105D5B7FF7DB6AAAABC7BEDB505EFBEA407",
INIT_2A => X"95038AAAEAF1D7410E80000FF8438E00B6DF68FEF4871D24BA495B5556D5571E",
INIT_2B => X"1ED1EFEAF1EFFFDEAD1C5010AA8E2FBD7B6DF47A00EBDB50000A380AAE28E804",
INIT_2C => X"5A001684104155C5B68E2DBEFBFFBC703AE2DF42AAA002A851C214003FF68007",
INIT_2D => X"50002155510000000000000000000000000000000000000000000002087A2841",
INIT_2E => X"55003FEAAAAD57DEBAA2FDDC01051FBD74BAF7802AB05AAFBD5400557BD54AA5",
INIT_2F => X"7AF7FC20B2F7FBC015D58517FF555D2ABDF55F782BEB47AFAD00010F7AA82155",
INIT_30 => X"55FFFFC20FFF3AE544108410174BA557BEABEFAAEBD55FFAA1456547A2D360F4",
INIT_31 => X"0BA547FD75FF58516AAAA0828AAAB4A78016545540400010557BFDFFFF7822A9",
INIT_32 => X"550AAFACAAA122AA8954BAA2AE9D545002A800A8FF862BA00F2F9E8F0050D442",
INIT_33 => X"954505C417FFFF08555555BAAD335B57AB5155400A2AEBFF45FFFB404007FFBD",
INIT_34 => X"00000000061DE08007FC2048002895755FFAEBCFE57BBA57002DF3C4AAAA002E",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000010000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(2),        -- Port A data input
DOA(0)   => data_read_a_lo(2),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(2),        -- Port B data input
DOB(0)   => data_read_b_lo(2),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_3_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"210C44A20020248B08431120001604B8156023104C40771B3430400A02380206",
INIT_01 => X"015A2A4050B009683C0422C992000B61404040028804A0080A000C16A8990A0C",
INIT_02 => X"C0A406500CE0A95011000D1501005274B5041AB330860281CC08008222170060",
INIT_03 => X"AB488054270F08E1289084C8020420E005A48DA16C021100003A46B06900C91A",
INIT_04 => X"848966150DA0A02941A4080C612A104201C689044382FD403C17E491829B259B",
INIT_05 => X"D006620608843116942508120A208D18A5050160C600D4C894600094B49CA068",
INIT_06 => X"12002D9401C70008060408141788E2C094887033080071913209CC8004640100",
INIT_07 => X"221111454874CCC4122C0932155400C2023940284000003E15020525CE805E11",
INIT_08 => X"020103C9984A0AC511102029869D974214EDBA132891000052C1750B48290020",
INIT_09 => X"60808C8A2E41351020004148A289428730A51E5E644C8233A0090E1020208100",
INIT_0A => X"A4000041A600417914506F955D6422000934000A090A94A020229603A414144D",
INIT_0B => X"469100841001000406D04065040650406D0406D04065040670406C8201782032",
INIT_0C => X"6A4AF532A8040AF821042D01F14084030070262810340402C0000CCE4CC12520",
INIT_0D => X"000800000401C333494594532980733302CCC81300094E5C91200257AD2AD795",
INIT_0E => X"00080000051C0000400000000000000800000190148000000800000450148000",
INIT_0F => X"0000010000000B100409000000000004000005101480000008000004F0148000",
INIT_10 => X"0000000002000000000001B00000400000000000000400000168018040000000",
INIT_11 => X"1000034010480000010002D804044000004000812E4400002440014080028000",
INIT_12 => X"0000000100570080880000080015C02090000002000CCC000200000000000040",
INIT_13 => X"1C0001000000000000104000094C002018000000000040100006418010440000",
INIT_14 => X"4128652000004404010E20500004208018800082008000000000010000100006",
INIT_15 => X"5795A5595A5595A5595A5595A5595E1152556D008028341B13924D80C2E67009",
INIT_16 => X"69565795A5595A5595A5595A5595A5595A559525795257952579525795257952",
INIT_17 => X"95256956579525495E5595A5495E5595A5495E5595A569565795256956579525",
INIT_18 => X"7818F18E0C8514298B0C52A0115009AA9556AAD552AAD5556956579525695657",
INIT_19 => X"24924924924924924924924924924820820820820825042C0000249249202A60",
INIT_1A => X"8D46A351A8D46A351A8D46A351A8D46A353A9D4EA753A9D4EA753A9249249249",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF248086A351A8D46A351A8D46A351A",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"EFAAFFD54AAF7D168B45AAAABDF5500002AA1000000000000000000000000000",
INIT_1F => X"F45FFD168AAA0855420AAAA843DFFFAAD1554005D7FD74AAA284001550055421",
INIT_20 => X"55FF5D003FE10F7803FEBAFFD5420AA080400155AAD5554AAF7802AB4500043D",
INIT_21 => X"28B45A2AE82155A2FBFFEBA0800021550855555FFAA84001FFAAAE80010A2AA9",
INIT_22 => X"168ABAFFFBD54BAAAAE97400A2FBC20AAA284175EF55517DF555D2EBFE00AA80",
INIT_23 => X"AA954AA5D7FFFF45AAAA975EF007BD7555FFFBFDF55AAFBD55EF5D2EBFE10085",
INIT_24 => X"AD1575EFAAAE974AA5D00175555D0015410F7AAAAAAA55043DE00FFFFD5555AA",
INIT_25 => X"0000000000000000000000000000000000000004174105D517DF55AAAAAABEFA",
INIT_26 => X"ABC04001C51551471D7AAF1D05D2EBD56DB7DBEAEBFF551C042AA101D0000000",
INIT_27 => X"92EB842FB5508043FF55EBD56ABD75D5B470AABE8A3AFD7A2DF55400557FD54A",
INIT_28 => X"557FD2082000BEAE905C755003FE28E3D17DEAAEBDF40002550F47155AADB504",
INIT_29 => X"DF40552ABDF45B6AEAFFD5F7A48017DAAFFFAE821C0A0717D1C5B575FFB68E82",
INIT_2A => X"C55D7492E90E3808756DA92EBFFD74BAE3AE85480FFFFC00AABE8E105C755517",
INIT_2B => X"43AE10EAF5C5547FF80954AA5D7FFAF7DA2AE905EF0075D5545E3F5EFF57F7D5",
INIT_2C => X"5B7FF7DB6AAAABC7BEDB505EFBEF5C7092FF801756D490A10438EBA4B8E92410",
INIT_2D => X"D0028A00510000000000000000000000000000000000000000000000E124105D",
INIT_2E => X"AAFBD54005D7BD54AAF78002155515157555AAD142040A2D57FFFFFFAEBFF555",
INIT_2F => X"051AE955F7AAFBC0000AF843FF5500003FF55AAFD6AB455157D74BAF7AAA8B45",
INIT_30 => X"FF557BD74EFFBACD41577B8400010F7AA8215555003FEAAAAC53DEB8A2FDDC01",
INIT_31 => X"0BAF7AA8015558517FF555D2ABDF51F782BCB47ABAE801FFAAFBEAA105D2E955",
INIT_32 => X"214FA2D3EAF57AFFDD7555082AA0AAA00557FEA8A2FDD64BAAF8282012AFFEC2",
INIT_33 => X"820AAAB842AA00000028AB0AAFF48547AE04174BA557BEABEFA2AA951FF88554",
INIT_34 => X"000000002A80010557BFDFFFF7822A955FFFFC21FFF3BE40412DE02955FF082A",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000008000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(3),        -- Port A data input
DOA(0)   => data_read_a_lo(3),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(3),        -- Port B data input
DOB(0)   => data_read_b_lo(3),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_4_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"A108400020612C80284210081034849800A000303100048B3432C82904204006",
INIT_01 => X"210668000008004C1C20250E12100368403008418984014902030906A8910200",
INIT_02 => X"120404C0024C0600000206100008402404040C00F104008040080080001310E0",
INIT_03 => X"7728805052470B5C1B873C04121D03845D0020CA0822018000080084C1000002",
INIT_04 => X"0B899E43891686690790485D5C3E02000E9892201D306D03A9835C16029AC186",
INIT_05 => X"C001E080005030767434C0003C8A01D6B81C5703C82CDBC000072400089C8120",
INIT_06 => X"1000088100410000460002041300004084080070D00030032009700024641102",
INIT_07 => X"4261950408CCBC2012048310951000000003402A4000143E1008912480000211",
INIT_08 => X"00811007AC0A1EB5131120C79E7D176251E53E80E8B361604041340838452020",
INIT_09 => X"C08360820C0912800035F1801630A8260900180C00C8021C800FEE522020A108",
INIT_0A => X"8400F88C166262E940D00D410D62AD02091704024D0A02882192020DA0544043",
INIT_0B => X"4011078510C90D143142430C243042430C24304243042430C24305121A612186",
INIT_0C => X"C08060101000C00401008800F004140009400E4002A0010240000DC3C080002C",
INIT_0D => X"000800100001C07261C51C42390240F050C3C000950008088130040100018000",
INIT_0E => X"00080010003510004000000000000048010002E0100000000800100220100000",
INIT_0F => X"0000014008001550000800000000000400800280100000000800100360100000",
INIT_10 => X"00000000020000080080009410004000000000000044080000D8008000000000",
INIT_11 => X"000005800008000001040168000040000041000100EC00004002214000008000",
INIT_12 => X"00000041003C000008000008200D00001000000208050C000200000000002040",
INIT_13 => X"17000100000000000090000002C8000008000000000060000004480000400000",
INIT_14 => X"8400C00208004844C00800000000528008000000008000000000010040000000",
INIT_15 => X"0100800004030080000C010000A00D1804404912802A261B53104810DB1E0028",
INIT_16 => X"000C030000200C01000020040300800004030000000C03000000040100802004",
INIT_17 => X"008020040100C010000200800004010040300800000020040100C03000020000",
INIT_18 => X"40C700FC0A000280C68A08A950520E964C3269B2C9864D30000C030040100800",
INIT_19 => X"555555555555555555555555555554514514514514526991A199A28A28981451",
INIT_1A => X"41A0D068341A0D068341A0D068341A0D06A351A8D46A351A8D46A35555555555",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF771F60D068341A0D068341A0D0683",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FF087FFDF5508003FEBA087FD54BAAA841540055000000000000000000000000",
INIT_1F => X"F5500003DF455555421EFAAFFD54AAF7D168B45AAAABDF55A2802AA1000002AB",
INIT_20 => X"DFFFAAD1554005D7FD74AAAA840015500002AABA082E954005500021FF5D2EBF",
INIT_21 => X"68BEF080028BFF0855555455500174BAA2AABDE0055517FF555555420AAAA843",
INIT_22 => X"168ABA0055574BA5555554BA5D0400155AAD1554AAF7802AB4500043DF45FFD1",
INIT_23 => X"0400010A2AA955FF55003FE10F7803FEBAFFD5420BA085168A00007BFDE10085",
INIT_24 => X"855555FFAA84001FFAAFBEAB45002A97545F7D1555EF55043DF5555517DEAA5D",
INIT_25 => X"000000000000000000000000000000000000002A82155A2FBFFEBA0800021550",
INIT_26 => X"5BC042AA101D0A28BC7007FFDF45080A3AEAA007BD2482BE84124285C0000000",
INIT_27 => X"004100021FF492AB8F7D1C0438E381451471D7AAFBD0492EBD56DB7DBEAEBFF5",
INIT_28 => X"FED1C5F470AABE8A3AFD7A2DF55400557FD54AABE84001C5550A28ABA1424974",
INIT_29 => X"FB5508043FF55EBD56ABD75D0428BEF005557545490012482B6A0BAE2849557A",
INIT_2A => X"6DA101475FDE10145F68A921C55504924955524AA140E0717DAADB50492EB842",
INIT_2B => X"43AF6D405F78E3A1C2002000BEAA905C755003FE28E3803DEAAEBDF40002557F",
INIT_2C => X"FFFAE821C0A0717D1C5B575FFB6DF425575D7BEFB55002097555FFD5401EF5D0",
INIT_2D => X"784000AA59000000000000000000000000000000000000000000000208017DAA",
INIT_2E => X"A2D57FFFFF7AEBFF55FF8028A00512EAAB45007FFFF55082EA8AAA087FC2010F",
INIT_2F => X"5512AAAA085D04174100800021FF002EA8BEF5D0428ABA595557555AAFBC2000",
INIT_30 => X"00FF802ABAA04552ABFF597FD74BAF7AAA8B45AAFBD54005D7BD54AAF7800215",
INIT_31 => X"5FFAAFBC0000AF843FF5500003FF55AAFD6AB4551002ABEF0055555550004020",
INIT_32 => X"DEB0A2FD5600051537DE005D557DE005D7BE8AA85555400100879560AA592F95",
INIT_33 => X"17545FFD5421FF5D0428BEF0079FCABA598400010F7AA8215555003FEAAAA843",
INIT_34 => X"0000000004001FFAAFBEAA105D2E955FF557BD75EFFBBCD415521FBFDF450004",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000010000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(4),        -- Port A data input
DOA(0)   => data_read_a_lo(4),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(4),        -- Port B data input
DOB(0)   => data_read_b_lo(4),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_5_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50DB0A0791B1B41694368283C81F9996A091A32152007AB36B20E03C040C002",
INIT_01 => X"880015C49830884C446A40000C34C24841280A00084000C8C212892EEA953231",
INIT_02 => X"408F417400B1D9100002171C1FA20171124E6AA00D8633F8CD09DBFBBB972F7C",
INIT_03 => X"88538F0182058082D800C3314722DC08A34084A100C4D7C99208521063D00148",
INIT_04 => X"F45E41AFAF420996B8411CA282F80A9091224800A2C61490363080C8A4000308",
INIT_05 => X"0EA416069640420901A01505C4410020C6E228DC30532839B043289D9C005031",
INIT_06 => X"13992D9AF8C74E92B7B568D19708C038AFFA89F0B9348C9204C389672407EF12",
INIT_07 => X"6255000016053C18162589725146F442222CE6AF844012BE795224458BA4DE0F",
INIT_08 => X"4F3F00503B4AE104B5347230418190420821006016FC18843630D285FC416CB4",
INIT_09 => X"EEA33E700340902C4424C442B0344724066C56C2248130A2D9C185B24A24832B",
INIT_0A => X"315325008348CC40AB570500204462508135D5AA593E043731E9B18A98440137",
INIT_0B => X"E0CD463C5813804E0258E0358E02D8E03D8E0258E03D8E02D8E03447012C701E",
INIT_0C => X"F8DE3C27CA181E5D710664A5F140C14BD32A2E281992940AFAA15C3FC0836310",
INIT_0D => X"F000BE0FC80020130841840308653FF0313FE92C23FB1EECB367C0F3E378F0BC",
INIT_0E => X"F000BE0FCD806FFFAF0AE83080E2AEB2F0F1E01BE53FE1F000BE0FC41BE53FE1",
INIT_0F => X"0231F0BF9E3F02A7FFD63669C0E008C3CB7F041BE1BFE1F000BE0FC41BE1BFE1",
INIT_10 => X"30180309A0F83FE2B87C7D006FFF9F1A7806013879BAA78FC103FF5F1F12F038",
INIT_11 => X"39E9C1DBF8A30C2098DBE2FF7F2320483136F200A822CBACAB9DDEB7F9BC291F",
INIT_12 => X"004C72BEC95FEF64E4090626DF15B7D1C6184131B7980DFFFC03F00003F01FB9",
INIT_13 => X"1DFFFA0A3C0202B8776AE7A7C9CBFFF060703080E29F1B79E9F6427EFE901C0E",
INIT_14 => X"2B716CA5C56620590350ACD3A7D5B7EFAC6DFC8C0312A0024B83F07F3999E9F2",
INIT_15 => X"F0BCAF3BC2F3BC6F0BCEF2BC2F3BC6DBC67C251104A2261253904580207E1C81",
INIT_16 => X"1BCEF0BC2F3BC2F1BCEF0BC6F2BC2F1BCAF1BC6F2BC6F2BCAF1BC2F3BC6F2BCE",
INIT_17 => X"BCEF0BC2F3BC2F1BCAF1BCAF3BC6F0BCEF0BCEF2BC6F2BCAF1BCAF1BC2F3BCAF",
INIT_18 => X"69CFEF73B6FFE7436DB6FD0831518424965B4D2492CB69AF1BCEF0BC6F2BC6F0",
INIT_19 => X"F7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF3EF9FBFBB9E79E7BEBCB7",
INIT_1A => X"DEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDF7DF7DF7D",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF29FDAF77BBDDEEF77BBDDEEF77BBD",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"AAA2802AA10FFFFFDE0008556AABA5D2ABFFEFFF800000000000000000000000",
INIT_1F => X"ABAF7AAA8BFFAA802ABFF087FFDF5508003FEBA087FD54BA0804154005555574",
INIT_20 => X"54AAF7D168B45AAAABDF55AA802AA1000003FEBA00002AABA5D2EBFEBAAAD16A",
INIT_21 => X"3DE005555575EFA2D142145A2FFE8B45FF80001555D2E955FFFFD5421EFAAFFD",
INIT_22 => X"FC00BA5D5568AAAF7AAAAAAAAA802AABA082E954005500021FF5D2EBFF550000",
INIT_23 => X"D5420AAAA843DFFFAAD1554005D7FD74AAAA840014500517FFEF007BEABFF5D7",
INIT_24 => X"2AABDE0055517FF555504154BAA2FBEAA105D2E97410FFD16AAAA5D2ABDEBAFF",
INIT_25 => X"000000000000000000000000000000000000000028BFF0855555455500174BAA",
INIT_26 => X"21E84124285C51574BAB68A2DA00FFFFFFE38085F6FA92552AB8FEFF78000000",
INIT_27 => X"925D2AB8EBABEDB6AA92F7AAA8BC7B68A28BC70075FDF45080A3AEAA007BD248",
INIT_28 => X"5FFFFD1471D7AAFBD0492EBD56DB7DBEAEBFF55BE842AA105D0A38EBA1C0428A",
INIT_29 => X"21FF492AB8F7D1C0438E38145B575EFA2DB45145B6F5EFB6DF78E05145552A92",
INIT_2A => X"7DFC70875EABC7557FC20AA415F68AAAF7AAAAA82BE8A28A9214249740041000",
INIT_2B => X"B6FABA542ABAE2AF7DF470AABE8A3AFD7A2DF55400557FD54AABE84001C55551",
INIT_2C => X"5557545490012482B6A0BAE2849043AFED1C0E10492B6FFEFA105D2A95410FFD",
INIT_2D => X"D2AAABEFFB8000000000000000000000000000000000000000000000428BEF00",
INIT_2E => X"082EA8AAA087FC20105504000AA5955554BAFFAEBDE10F7FBFDEBA007BFDE005",
INIT_2F => X"0512AA8AAA5D0028A005D2AA8ABAF7FBE8A00FFAEAAB45F3AAAAB4500557FF55",
INIT_30 => X"EFFFAA97545552A821EFFBD557555AAFBC2000A2D57FFFFF7AEBFF55FF8028A0",
INIT_31 => X"A005D04174100800021FF002EA8BEF5D0428ABA597FD55FFA2FFD5555FFD57FF",
INIT_32 => X"54AAF7800015551517DF45005168B55557FC0012087FEAABAF7AAAAA10F3AAAA",
INIT_33 => X"FFE005D2A95410F7FFFFEBA5D2EA8ABAFBFFD74BAF7AAA8B45AAFBD54005D7BD",
INIT_34 => X"00000000002ABEF005555555000402000FF802AAAA04452ABFF592E80010FFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000060000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(5),        -- Port A data input
DOA(0)   => data_read_a_lo(5),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(5),        -- Port B data input
DOB(0)   => data_read_b_lo(5),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_6_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10800B0061A01002840002C030028180004003220200403312301C4389B2082",
INIT_01 => X"060009C838394848188160000C42426041000000090800090210090000510200",
INIT_02 => X"00043040009001100000061000018070002408000000000648080000001210E0",
INIT_03 => X"0000800002054081020080801200A0000300008000201184681A0000410C4800",
INIT_04 => X"0808801040000001401048008100022401400002024024053200020089000100",
INIT_05 => X"0240040408402202002000C200400020A50000A0000010010001260808000520",
INIT_06 => X"44000881064500004600000013088002840C240F5048011200010000440C0146",
INIT_07 => X"0241914041FE83E010040110110003040020402A0000003E1000000488000201",
INIT_08 => X"8001BF002C4A01041B112020200110024029006FE09081002004902000012068",
INIT_09 => X"0083FE38A040100281353150ACB645AEF8C01404448000008011061204200108",
INIT_0A => X"3103AD0413424E4014D627C470462200011504420C0A962A2189002881404060",
INIT_0B => X"46C1060C16C96D15B0425B0425B1425B1425B0C25B0C25B1C25B1512D8212D82",
INIT_0C => X"009000140401100601016600A040220203A004480598010248000D0010420C0C",
INIT_0D => X"0000A01033A00013000000000018800F2400091081100C0090A5008200410020",
INIT_0E => X"0000A0103142000000000000000000455D0018100000000000A0103410000000",
INIT_0F => X"000000466800C200000000000000000001A0F4100000000000A0103410000000",
INIT_10 => X"00000000000024094680014200000000000000000041E8002900000000000000",
INIT_11 => X"F000322000000000000D1A000000000000034D240C2000502000000000000000",
INIT_12 => X"000000403F4000000000000068D24000000000001A60F0000000000000002007",
INIT_13 => X"C0000000000000000087C0003014000000000000000025D00008958000000000",
INIT_14 => X"02000000000814C219500150002800101280000000000000000000086670000C",
INIT_15 => X"8120C82208812048120882208892055A0060011280222413130449010301F051",
INIT_16 => X"3200802008320C82200802048320C82200812048320880200812048220880204",
INIT_17 => X"20C83208812048020883204802048120882204812008220C8220081204822088",
INIT_18 => X"79CFF1FE1E9F52ABEF9EFE8150120EC718638E38E30C71C812088220C8120080",
INIT_19 => X"71C71C71C71C71C71C71C71C71C71C71C71C71C71C736D9DBD9BBEFBEFBEBEF1",
INIT_1A => X"CFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FC71C71C71C",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCF29A7F3F9FCFE7F3F9FCFE7F3F9F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000607FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"EFA2FBD54BA5555554BAAAFBC20BA5D7BEAAAAFF800000000000000000000000",
INIT_1F => X"EBA0855421455555574AAA2802AA10FFFFFDE0008556AABA5D2ABFFEFFF843DF",
INIT_20 => X"DF5508003FEBA087FD54BA000415400550428AAAAA84021FF007BD54BAAAD17D",
INIT_21 => X"A8BFFAAD1554BA002A95555A28417400AAFBE8ABAF7FFD54AAAA802ABFF087FF",
INIT_22 => X"BD5545080417555A2D17FE1000003FEBA00002AABA5D2EBFEBAAAD16AABAF7AA",
INIT_23 => X"D5421EFAAFFD54AAF7D168B45AAAABDF55AA802AA100000001EF087FEAA00FFF",
INIT_24 => X"F80001555D2E955FFFF843DEAAA2803DFEF0855401FF082EA8B555D7FC21FFFF",
INIT_25 => X"0000000000000000000000000000000000000055575EFA2D142145A2FFE8B45F",
INIT_26 => X"2552AB8FEFF78E3DFFFAAFFD04AA415B52492B6F5C20825D7FE8A92FF8000000",
INIT_27 => X"EF147BD2482BED57AE921451421555551574BAB68A2DA00FFFFFFE38085F6FA9",
INIT_28 => X"4BAB68A28BC70075FDF45080A3AEAA007BD24821C04124281C0E2DA82BE8E001",
INIT_29 => X"8EBABEDB6AA92F7AAA8BC7B6D5524AA14209557DA28E15400BEF1EFA92FFFFD2",
INIT_2A => X"071FF0071EDA38F7F1D5555000417545B6D178E281C0A38EBA1C0428A925D2AB",
INIT_2B => X"4A8B555C7FC2147F7D1471D7AAFBD0492EBD56DB7DBEAEBFF55BE842AA105D0E",
INIT_2C => X"DB45145B6F5EFB6DF78E05145552A925FFFF8E3DE82BE8E38FFF0851401C7082",
INIT_2D => X"57FE8A00F38000000000000000000000000000000000000000000005B575EFA2",
INIT_2E => X"F7FBFDEBA007BFDE005D2AAABEFFBAABDFEFAAFBC00BA007BC0000FFD5420005",
INIT_2F => X"A592ABFE00F7AA821FF557FC0010F7D168A105D55421455155554BAFFAEBDE10",
INIT_30 => X"10F7D57DE00FFFBC00AAFBAAAAB4500557FF55082EA8AAA087FC20105504000A",
INIT_31 => X"AAA5D0028A005D2AA8ABAF7FBE8A00FFAEAAB45F3D5400BA5504155EFAAAE954",
INIT_32 => X"FF55FF8028A00512E975FF08557FEAAF7D157545080417545F7D56AAAA592AA8",
INIT_33 => X"AABEF005542155000028B555D7FC2145F3D557555AAFBC2000A2D57FFFFF7AEB",
INIT_34 => X"000000007FD55FFA2FFD5555FFD57FFEFFFAA97545552A821EFFBAABDE00F7AA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000048000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(6),        -- Port A data input
DOA(0)   => data_read_a_lo(6),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(6),        -- Port B data input
DOB(0)   => data_read_b_lo(6),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_7_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10844B00482258A2842112C02450418800002300500030B313300C418992002",
INIT_01 => X"020009C23838684D1C20E0000E11424840000000080000080200000000110204",
INIT_02 => X"000520700CA08910000206101180803081144880010400044808000000122160",
INIT_03 => X"000080040305208000008000328080040304008020303194289A000041484800",
INIT_04 => X"08088000000000010000CA008008060441000000028234493410820191000000",
INIT_05 => X"03500404000022020020044000000C208400408000001000984005949C002928",
INIT_06 => X"54000881044500004680000013008002940C24001A4A010200018920646410C7",
INIT_07 => X"22510040400500011204813015012204002040280000013E1000000488000201",
INIT_08 => X"9001A0602C4A01051B132820208001024069004008908002120851420001226A",
INIT_09 => X"01100020A2401008A20404E08200A05000A4264640800022C8198C4E05200018",
INIT_0A => X"20002000024040400050450440C48A0041140C420B0904208800904286000008",
INIT_0B => X"50822002120D2134800648006480064800648106481064810648193240432404",
INIT_0C => X"284A142288042A5C24202451505E00A621A5220A8091444040188C001B41210A",
INIT_0D => X"00F001F021141A12004104020810B000100000000109064C80010050A3285194",
INIT_0E => X"00F001F027420000400004C3201C514408081C1014800000F001F02810148000",
INIT_0F => X"E00E0E404100E200040900000B0380383480C81014800000F001F02810148000",
INIT_10 => X"4160C0301D07001D0402034200004000019860078641004039000180400002C0",
INIT_11 => X"08103BA0104810C8462416E8040446120C890814600010512000000080028400",
INIT_12 => X"98038D4030DD008088C2419120B740209021908C4846FC000200030F000FE006",
INIT_13 => X"DD000100411C81078884204035DC00201804C3201C60A408100DD58010440130",
INIT_14 => X"412024202211148019064200402A32901A8000B2048902C0807C0E00C448100D",
INIT_15 => X"50942509425194651946519465894619421421102000269243854D8002000250",
INIT_16 => X"19465194E50942509425094E51946519465094A50942509425194E5194651942",
INIT_17 => X"9425094251946539465094250946539465194250942509465194650942509425",
INIT_18 => X"0000000000000000000000080150890820800041041000052942509465194653",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF21E6C000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"AAF7D5575455D557DFEF002AAAB55002E820AAAA800000000000000000000000",
INIT_1F => X"B55007FD74AAAA843DFEFA2FBD54BA5555554BAAAFBC20BA5D7BEAAAAFFFBC00",
INIT_20 => X"AA10FFFFFDE0008556AABA5D2ABFFEFFFAAAAAAAF7D57FFEFF7D555555A2AEAA",
INIT_21 => X"42145552ABDFEFFFAA801EFFFFBFDF550000175555504175450055574AAA2802",
INIT_22 => X"A975EF00003DF55555168A00000428AAAAA84021FF007BD54BAAAD17DEBA0855",
INIT_23 => X"802ABFF087FFDF5508003FEBA087FD54BA000415400557BD74BAFFD140000082",
INIT_24 => X"AFBE8ABAF7FFD54AAAAAEA8ABA55557FEAAA2843FF55A2AEA8B55AAAABDEAAFF",
INIT_25 => X"0000000000000000000000000000000000000051554BA002A95555A28417400A",
INIT_26 => X"25D7FE8A92FFFFC70BAE3D155555415178FD7082EAAB550820870BAAA8000000",
INIT_27 => X"FFEBD55557DBEA4AFB550871D7482AA8E3DFFFAAFFD04AA415B52492B6F5C208",
INIT_28 => X"5550051574BAB68A2DA00FFFFFFE38085F6FA92552AB8FEFF7A0ADABAEBD578F",
INIT_29 => X"2482BED57AE921451421555524BDFD7FFA4801D7F7F5FDF55000E17545410E17",
INIT_2A => X"D2482E3D1450381C20905EF08003AF55415F6DA38080E2DA82BE8E001EF147BD",
INIT_2B => X"AAFB55ABA0BDE02EB8A28BC70075FDF45080A3AEAA007BD24821C04124281C7B",
INIT_2C => X"209557DA28E15400BEF1EFA92FFFFD24BAB6A4A8A82495F78E92AA843DF45BEA",
INIT_2D => X"800174BAA680000000000000000000000000000000000000000000055524AA14",
INIT_2E => X"007BC0000FFD542000557FE8A00F3FFD54BAAAD15754508556AB45002AA8B450",
INIT_2F => X"FFB803DEAAAAD56ABEFAAD5575EFF7803DF45085557410AEAABDFEFAAFBC00BA",
INIT_30 => X"55082E97555002E955550C55554BAFFAEBDE10F7FBFDEBA007BFDE005D2AAABE",
INIT_31 => X"E00F7AA821FF557FC0010F7D168A105D554214551003FF45FF8400145FFD57FF",
INIT_32 => X"20105504000AA597FC2010A2D1554AA5500021EF000028B55087BFDEBA042ABF",
INIT_33 => X"E8A00A2803FF45F7AABDF55AA843FE10AEAAAAB4500557FF55082EA8AAA087FC",
INIT_34 => X"0000000055400BA5504155EFAAAE95410F7D57DE00FFFBC00AAFB8028A00007F",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000007FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(7),        -- Port A data input
DOA(0)   => data_read_a_lo(7),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(7),        -- Port B data input
DOB(0)   => data_read_b_lo(7),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_8_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000B0000040042840002C0000001800000070000000033022000000000086",
INIT_01 => X"000009C21838284D1C2160000E12426840000000180800080200080040510200",
INIT_02 => X"0001004000900110000006100080003000240800014400004808000000122160",
INIT_03 => X"00008000020440810002A0801010A0044300000000200086011A000040404800",
INIT_04 => X"8000801000020401400040408108022029400000124004041200000089000100",
INIT_05 => X"02080424085022020000040200480020850010A0002010010120060800040400",
INIT_06 => X"50000880006500000680000011008006840C200018C1010200018920E0640102",
INIT_07 => X"426000404005000112048130150120240020400A0000013E1000000488000010",
INIT_08 => X"220100402C42010413110020200100024029004000A200002004902200012141",
INIT_09 => X"0000000080400008010410A2940A45240040140440800022C8388E1200A00008",
INIT_0A => X"00420100020048405000070440C0000001140412090000000021002081000048",
INIT_0B => X"0000000800000100011000010000100001000010000100001000010000880008",
INIT_0C => X"001000040001100008012008004020102180800804802000C0080D00100A0008",
INIT_0D => X"0FF0000002200A1200410402080080003000091085100C008124008000400020",
INIT_0E => X"0FF000000140000040F517CF600000000104081010001E0FF00000001010001E",
INIT_0F => X"E000000000804200000809963F1F80000000001010001E0FF00000001010001E",
INIT_10 => X"CFE7C0F00000000000810140000040E587F9E000000008100900008000ED0FC7",
INIT_11 => X"00021040030C73D80000021000585F3600000020240020102000000802419660",
INIT_12 => X"F80000000042000B0BD6C0000010800618E7B000000C000003F80FFF00000000",
INIT_13 => X"800005D5C3FD800000000008180000078A8FCF600000000002028001006AA3F1",
INIT_14 => X"020000000008808219002100100C000041120370DCAD1FC18000000000000202",
INIT_15 => X"8020080200812048120481204812055A04604930A02026934215410102000110",
INIT_16 => X"0200802008020080200802048120481204812048120481204802008020080200",
INIT_17 => X"2008020081204812048120481200802008020080200802048120481204812048",
INIT_18 => X"414A87D78AF42143CEBAC88151120A0000000000000000081204812008020080",
INIT_19 => X"F3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF7E799B1BEB65B65948051",
INIT_1A => X"C3E9F0FA7C3E9F0FA7C3E9F0FA7C3E9F0F87C3E1F0F87C3E1F0F87CF3CF3CF3C",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF1B5DA9F0FA7C3E9F0FA7C3E9F0FA7",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"0000043DF55087BC01EF007FD75FFFF84000AAFF800000000000000000000000",
INIT_1F => X"E10A28028AAAAAFBC00AAF7D5575455D557DFEF002AAAB55002E820AAAA84000",
INIT_20 => X"54BA5555554BAAAFBC20BA5D7BEAAAAFFAA95545552ABFE00087BC00AA082EBF",
INIT_21 => X"D74AAAAD57FF45002A975FF007BE8BFFA2FBFFFFFAAD5400AAFF843DFEFA2FBD",
INIT_22 => X"BE8A00082A97410F7D5555EFAAAAAAAAAF7D57FFEFF7D555555A2AEAAB55007F",
INIT_23 => X"55574AAA2802AA10FFFFFDE0008556AABA5D2ABFFEFFFAA82000555555545AAF",
INIT_24 => X"00017555550417545000015545087BC2010AAD54014500516ABFFA2AABDF4500",
INIT_25 => X"000000000000000000000000000000000000002ABDFEFFFAA801EFFFFBFDF550",
INIT_26 => X"50820870BAAA8407000140038F450075C71FF087BD75D7FF84050BAEB8000000",
INIT_27 => X"10007FC50BA002ABFE00AA8A2AABABEFFC70BAE3D155555415178FD7082EAAB5",
INIT_28 => X"082EB8E3DFFFAAFFD04AA415B52492B6F5C20825D7FE8A92FFA497545552AB8E",
INIT_29 => X"557DBEA4AFB550871D7482AAD17DF451C24955EF0875EFBD7B6F1FFFC7BEDB45",
INIT_2A => X"87000415B5057DAAFBE8A10082092410EBD5505EFB6A0ADABAEBD578FFFEBD55",
INIT_2B => X"B6ABC7B6AABFFED0051574BAB68A2DA00FFFFFFE38085F6FA92552AB8FEFF7AA",
INIT_2C => X"A4801D7F7F5FDF55000E17545410E17555000E17545007BC0000BED14217D005",
INIT_2D => X"784174AAA280000000000000000000000000000000000000000000024BDFD7FF",
INIT_2E => X"08556AB45002AA8B450800174BAA684174105D042AB550055555FF007BD7555F",
INIT_2F => X"0F384175555D2EA8A00087BD74BA082EBDE10AAAEA8ABAF7FFD54BAAAD157545",
INIT_30 => X"55FFD57DF55FFFBD5400A2AABDFEFAAFBC00BA007BC0000FFD542000557FE8A0",
INIT_31 => X"EAAAAD56ABEFAAD5575EFF7803DF45085557410AED17FF455D04155FF00557DF",
INIT_32 => X"DE005D2AAABEFFBAE97410087BC21EFA2FFEAA00000002010A2D5421FFFF803D",
INIT_33 => X"C0010FFD1401EF087FE8B55FFAEBDFEF0855554BAFFAEBDE10F7FBFDEBA007BF",
INIT_34 => X"00000000003FF45FF8400145FFD57FF55082E97555002E955550C2E95555087B",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000020000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(8),        -- Port A data input
DOA(0)   => data_read_a_lo(8),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(8),        -- Port B data input
DOB(0)   => data_read_b_lo(8),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_9_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00018248A2840112C00002C18000002300500030B3132000400812002",
INIT_01 => X"A140098218302849180060000C004240413C0A61590001D90213C90008510204",
INIT_02 => X"102008700CB089100002061031285074810448800104008048080080001210E2",
INIT_03 => X"00008015074608840390A0040040800203140000A00010800408108448020042",
INIT_04 => X"082080400004A00100000100840602020100000002C2344156108201811801C0",
INIT_05 => X"0200048480011502049500280020CC2084000080008010019161249C9C002188",
INIT_06 => X"70000881004500004E01020411D08000940C00001800010200018B20206C0102",
INIT_07 => X"EA70C0040005000312048130150100040020404A0000017E10408104C8000110",
INIT_08 => X"000000402C220104131004202081120050A5104000A204617201D10801002000",
INIT_09 => X"000800002F4924003085E51420A0100400641E4E40800022C8088C1220200908",
INIT_0A => X"20102000024040484028450001648C2229150400080244000401900284000440",
INIT_0B => X"0880110901081110411204112040120411204012041120401204111020090208",
INIT_0C => X"685B34A688841A5C21200101A01A0004009024028004044248404D00104B2100",
INIT_0D => X"0000A01000000213000000000000B0001000010000190E44802002D1A168D0B4",
INIT_0E => X"0000A010014000000000000000000040500008100400000000A0100410040000",
INIT_0F => X"0000004608004200040000000000000001A004100080000000A0100410008000",
INIT_10 => X"00000000000024080000014000000000000000000040A0000900010000000000",
INIT_11 => X"300013E010000000000D00F804000000000340000C0000102000000080000000",
INIT_12 => X"00000040091F0000800000006807C000800000001A0CFC000000000000002001",
INIT_13 => X"DD000000000000000082C00019DC002000000000000021500006D58010000000",
INIT_14 => X"03206420000000C019502050000C32901A800080000000000000000860100006",
INIT_15 => X"D1B46D1B46D0B42D0B42D0B42D8B424342342832002A24921082158802001011",
INIT_16 => X"0B42D0B42D0B42D0B42D0B46D1B46D1B46D1B46D1B46D1B46D1B46D1B46D1B46",
INIT_17 => X"B42D0B42D1B46D1B46D1B46D1B46D1B46D1B46D1B46D1B42D0B42D0B42D0B42D",
INIT_18 => X"89999E91BCD1512B871C4A0100000000000000000000000D0B42D0B42D0B42D0",
INIT_19 => X"A28A28A28A28A28A28A28A28A28A29A69A69A69A69A51C200807249041202AE6",
INIT_1A => X"8349A4D068341A0D269341A0D269341A0D068341A0D068341A0D068A28A28A28",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF2DA921A0D269341A0D068349A4D06",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"45A280154BA5555401EFFFD5421EFA2FFFFF555D000000000000000000000000",
INIT_1F => X"5EF00557DF555D040000000043DF55087BC01EF007FD75FFFF84000AAFFD57DF",
INIT_20 => X"75455D557DFEF002AAAB55002E820AAAA843DFEF00517DEBA007BFDFEFFFD157",
INIT_21 => X"28AAAAAAABDF45F7803FFEF555568AAAF7802AA00FFFBD7555087BC00AAF7D55",
INIT_22 => X"BD54BA550417400085155555082A95545552ABFE00087BC00AA082EBFE10A280",
INIT_23 => X"043DFEFA2FBD54BA5555554BAAAFBC20BA5D7BEAAAAFFFBC00AA552E95545087",
INIT_24 => X"2FBFFFFFAAD5400AAFF8402000A2FFFDF555D7BE8BFF5D51575EFA280175555D",
INIT_25 => X"00000000000000000000000000000000000000557FF45002A975FF007BE8BFFA",
INIT_26 => X"7FF84050BAEBDF78F45B68010482415B471C7E3DF451EFBEFBFAF45490000000",
INIT_27 => X"82007FFAFEFE3DB505EF1C5B7AF45490407000140038F450075C71FF087BD75D",
INIT_28 => X"5451C7FC70BAE3D155555415178FD7082EAAB550820870BAAA8438FFF00517DE",
INIT_29 => X"50BA002ABFE00AA8A2AABABEAEB8F45F78A3DFD741516DAAAE38E2DA28EBFFD5",
INIT_2A => X"C20BA5D2E905550071D54825D0A1543808515756D1C2497545552AB8E10007FC",
INIT_2B => X"5505FFBE801256D490E3DFFFAAFFD04AA415B52492B6F5C20825D7FE8A92FFFF",
INIT_2C => X"24955EF0875EFBD7B6F1FFFC7BEDB45082EB8002000AAFFFDF6D417FEABEF5D5",
INIT_2D => X"7FBE8B5500000000000000000000000000000000000000000000000517DF451C",
INIT_2E => X"0055555FF007BD7555F784174AAA2FBEAB45F78402010007BD5545AAFFD55EFF",
INIT_2F => X"AA68028BEF00517FE10007BE8BFFAAFFC01FF557FE8B550004174105D042AB55",
INIT_30 => X"AAAAAEBFEAAAAFFD5545557FD54BAAAD15754508556AB45002AA8B450800174B",
INIT_31 => X"5555D2EA8A00087BD74BA082EBDE10AAAEA8ABAF7AAAAB45F7AEBFF4508557FE",
INIT_32 => X"2000557FE8A00F3FFC00BA552E80145005557400552A954BA0051575EF550417",
INIT_33 => X"FDFFF007FE8BFF5551401EFF784021FF002ABDFEFAAFBC00BA007BC0000FFD54",
INIT_34 => X"00000000517FF455D04155FF00557DF55FFD57DF55FFFBD5400A28400010A2FB",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000040000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(9),        -- Port A data input
DOA(0)   => data_read_a_lo(9),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(9),        -- Port B data input
DOB(0)   => data_read_b_lo(9),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_10_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00018248A2840112C00002C18000202300500030B3132000400992006",
INIT_01 => X"A140098218302849180060000C00424040000000080000080200090008510204",
INIT_02 => X"102100400C8001100000061000A8503401044880010400004808000000122160",
INIT_03 => X"000080150746088401908000100080020304000020201080001A108448404842",
INIT_04 => X"800080400004A001000040008406020201000000020004401000000180180080",
INIT_05 => X"02000484800133020495040800208C20A4000080000010000001249010042008",
INIT_06 => X"50000881004500004681020411808000940C20001800010200018920206C0102",
INIT_07 => X"024084044005000112048130150120040020400A0000013E10408104C8000010",
INIT_08 => X"000100402C020105131100200000124250A51040088084614001110801012000",
INIT_09 => X"00080082CD09240820800000000000040000180840800022C8088C1220200108",
INIT_0A => X"841201000200484910000F050560262229140402080200A00402000484140400",
INIT_0B => X"0010118900080010000200102001020000200002001020010200001000010008",
INIT_0C => X"408120900404004821202001F05E00040180260A8080044240004C0010800228",
INIT_0D => X"0000A01000000813004104020800800030000800010008088124020102008100",
INIT_0E => X"0000A010014000004000000000000040500008101480000000A0100410148000",
INIT_0F => X"0000004608004200040900000000000001A004101480000000A0100410148000",
INIT_10 => X"00000000000024080000014000004000000000000040A0000900018040000000",
INIT_11 => X"3800100010480000000D00000404400000034000282000102000000080028000",
INIT_12 => X"00000040090000808800000068000020900000001A0000000200000000002001",
INIT_13 => X"80000100000000000082E0001000002018000000000021580000800010440000",
INIT_14 => X"00004000000004C0195000500008000000000082008000000000000860180000",
INIT_15 => X"0100401004010040100401004090055804404110802A24921317580802001011",
INIT_16 => X"0000000000000000000000040100401004010040100401004010040100401004",
INIT_17 => X"0040100400000000000000000000000000000000000000000000000000000000",
INIT_18 => X"215281FC1A72E2486AAA40A85052020000000000000000001004010040100401",
INIT_19 => X"51451451451451451451451451451451451451451452AA83330A8A28A29EA8D1",
INIT_1A => X"5CA6532994CA6532B95CAE572994CA6532994CA6532994CA6532994514514514",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF31CE2E572994CA6532994CAE572B9",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"10AAFBE8AAAA2D540000F7D57DF55A2AABFFEF08000000000000000000000000",
INIT_1F => X"F45FFFBC2010AAD57DF45A280154BA5555401EFFFD5421EFA2FFFFF555D003FE",
INIT_20 => X"DF55087BC01EF007FD75FFFF84000AAFF8002155AAFFE8B45AAD540000087FFD",
INIT_21 => X"7DF555D517FEBA082A801EFF7FBD5400FFD568B555D00155EF08040000000043",
INIT_22 => X"BFDE00A2FBC0145005168A10AA843DFEF00517DEBA007BFDFEFFFD1575EF0055",
INIT_23 => X"7BC00AAF7D5575455D557DFEF002AAAB55002E820AAAA803FEBA082AAAAAAF7F",
INIT_24 => X"7802AA00FFFBD7555082E82155FFAEAAB55AAD568B455D00154BAFFFBD75EF5D",
INIT_25 => X"000000000000000000000000000000000000002ABDF45F7803FFEF555568AAAF",
INIT_26 => X"FBEFBFAF4549003DE10BEF5EDAAAAAD547038EBD57DF7DA2AEB8FC7000000000",
INIT_27 => X"6DAADF470280075FFF45E3F1C7038A2DF78F45B68010482415B471C7E3DF451E",
INIT_28 => X"5C7000407000140038F450075C71FF087BD75D7FF84050BAEB8002155BEF5EDB",
INIT_29 => X"AFEFE3DB505EF1C5B7AF45495B7DEAA0824851EFEBFBD2410EBD168B7D410A17",
INIT_2A => X"38EAA0824A8AAAEBF5FAE28AAF1C2155005F68A10A28438FFF00517DE82007FF",
INIT_2B => X"4104AAF7F1D75EF557FC70BAE3D155555415178FD7082EAAB550820870BAAA80",
INIT_2C => X"8A3DFD741516DAAAE38E2DA28EBFFD55451C2087155EBA4A8B7DAADF68B7D410",
INIT_2D => X"2AEAAB55000000000000000000000000000000000000000000000002EB8F45F7",
INIT_2E => X"007BD5545AAFFD55EFF7FBE8B5500043FE00F7D17FEBAA2D5574BAAAD17DFEFA",
INIT_2F => X"AA28002155FFD17FFFFA2FBD74BA00557FF45A2D5554AAA2FBEAB45F78402010",
INIT_30 => X"00AAD16ABFF002A975450004174105D042AB550055555FF007BD7555F784174A",
INIT_31 => X"BEF00517FE10007BE8BFFAAFFC01FF557FE8B55007FFDEAA0004175FFA2FBC20",
INIT_32 => X"8B450800174BAA68428AAA08042AABAAAD56AABAAAD140155087FEAA10A28028",
INIT_33 => X"2ABEFAAFBE8BFF0004020AAFFD5555EF557FD54BAAAD15754508556AB45002AA",
INIT_34 => X"000000002AAAB45F7AEBFF4508557FEAAAAAEBFEAAAAFFD5545550015555A284",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000047FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(10),        -- Port A data input
DOA(0)   => data_read_a_lo(10),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(10),        -- Port B data input
DOB(0)   => data_read_b_lo(10),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_11_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10180B05A0010402840602C2D001019000000300000000330A20080EC180002",
INIT_01 => X"AB400984B830084C1820E0000C36424840000000080000088200000802112220",
INIT_02 => X"102A68440080011000000618062AD03502640800010410424908136019920868",
INIT_03 => X"001282118644C88481908001106088022300000080F4925CDC9A10844A9A4842",
INIT_04 => X"401280480004A1011000418084460002E12000000200040010000040A8000000",
INIT_05 => X"0FC8048484011502059511488020802084400888001110000000050000005400",
INIT_06 => X"1011088AE24500001631024511C08004A70AA40008B90D0200018B60A0650D45",
INIT_07 => X"020011005405000910040150110041040024400D800002BE18408104C9205908",
INIT_08 => X"89390040280241041D175820000001020061004004800567403512A801014C46",
INIT_09 => X"050800E20D09A424C5840400808000040680180840800022D8288E946CA00833",
INIT_0A => X"85002000024040410A000D0504408C32E915D9C208050084840201A099100400",
INIT_0B => X"B01011934A005101431CA821CA831CA821CA831CA831CA821CA83165410E5410",
INIT_0C => X"00010080028000010402214850444091019B02080885200042A9CC001000003A",
INIT_0D => X"5A5018C5A0A00812004104020808B00030000808024008008325820000000000",
INIT_0E => X"5A5018C5AB0062C38A4DB680A0D8241500D5761B011986695014A96E1A811986",
INIT_0F => X"42056A289A1BB2078A922DA2A8B180A2600AAE1A811986695014A96E1B011986",
INIT_10 => X"05AA429189B60AC43C6C7F0272C3841DB528802CAB18468F4101621B1BAC8455",
INIT_11 => X"C003104289A668B8CAB270106338317A3D94392020224ACDE215883078681B5C",
INIT_12 => X"804B020A06020C67061BC785938085134CD551BCA1C90006C0C2958502861120",
INIT_13 => X"80819A5539D503336D61056ABA006282806CA64090B89E015AAA880E48382EB8",
INIT_14 => X"40000000E808989003066E03513E41470126C6284B2D20410AB4503089C00A82",
INIT_15 => X"0000000000000000000000000000041800400110200026124202500802000800",
INIT_16 => X"1004010040100401004010000000000000000000000000000000000000000000",
INIT_17 => X"0040100401004010040100401004010040100401004010040100401004010040",
INIT_18 => X"C110083018162148420840280050800000000000000000001004010040100401",
INIT_19 => X"000000000000000000000000000001041041041041003882928E0000000AA0C4",
INIT_1A => X"0000000000008040000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3E0FC000000000000020100000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"EFAA842ABEFA280155EFFFFBC01EF08554000055000000000000000000000000",
INIT_1F => X"F4508514000000003FE10AAFBE8AAAA2D540000F7D57DF55A2AABFFEF0804155",
INIT_20 => X"54BA5555401EFFFD5421EFA2FFFFF555D51575FFA2FFD75FF550015400FFFBFF",
INIT_21 => X"C2010AAD568AAAAAD142145FF80155EF0051555FF0804155FFF7D57DF45A2801",
INIT_22 => X"01540008514215555003DFFFA28002155AAFFE8B45AAD540000087FFDF45FFFB",
INIT_23 => X"040000000043DF55087BC01EF007FD75FFFF84000AAFF802ABFFA2AABFE10080",
INIT_24 => X"FD568B555D00155EF085168B45085142010FFAE800AA5D7BFDF45F7FFEAA0000",
INIT_25 => X"00000000000000000000000000000000000000517FEBA082A801EFF7FBD5400F",
INIT_26 => X"DA2AEB8FC70000175EFB6802DBC7BE8A155EFE3FBC71FF145B42038550000000",
INIT_27 => X"EF550E15400E3F1FFF7D085B420381C003DE10BEF5EDAAAAAD547038EBD57DF7",
INIT_28 => X"5C7F7DF78F45B68010482415B471C7E3DF451EFBEFBFAF45495F575FFBEF5D05",
INIT_29 => X"70280075FFF45E3F1C7038A2DB68ABAB6D145145FF84155D7085B555C7140410",
INIT_2A => X"28BEFBEA4BDE28140A1543800514515549003FFC7BE8002155BEF5EDB6DAADF4",
INIT_2B => X"FFFF7DE3F1EFA10140407000140038F450075C71FF087BD75D7FF84050BAEB84",
INIT_2C => X"24851EFEBFBD2410EBD168B7D410A175C7005B6DB55145140000FFAE85082417",
INIT_2D => X"57BC20AA5D0000000000000000000000000000000000000000000005B7DEAA08",
INIT_2E => X"A2D5574BAAAD17DFEFA2AEAAB550004175FFF7803DF45FFAE955EFAAFBD55EF5",
INIT_2F => X"5007FD75FFF7D5401EF5D2E97410AAD17DFEF007FC20AA5D043FE00F7D17FEBA",
INIT_30 => X"55007FD5545550400145FFFBEAB45F78402010007BD5545AAFFD55EFF7FBE8B5",
INIT_31 => X"155FFD17FFFFA2FBD74BA00557FF45A2D5554AAA2FBEAAAAFFD555545FF80155",
INIT_32 => X"7555F784174AAA2842ABEFFF803DEAA5D2E974AA00515754500003FF55FF8002",
INIT_33 => X"40000FFAE97410007BFFFFFA2D57FE105D04174105D042AB550055555FF007BD",
INIT_34 => X"000000007FFDEAA0004175FFA2FBC2000AAD16ABFF002A97545007FFFF455555",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000040000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(11),        -- Port A data input
DOA(0)   => data_read_a_lo(11),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(11),        -- Port B data input
DOB(0)   => data_read_b_lo(11),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_12_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50080B01BC002006940202C0DE041196A83183000000023322287E0FC000006",
INIT_01 => X"0E000C068000E04D40238000001702484000000008000008820009280A553231",
INIT_02 => X"400B71440C8001100000171C0283813013766A800586235ECC09C8423B962966",
INIT_03 => X"CC618E048306E082000081000040900003548421A080025EDF08421042DC0108",
INIT_04 => X"00028020000000812000012080080000E100001002000448100000C1BC18008C",
INIT_05 => X"0FF8060610000402010015E100004C2084800090000310000000079010007C19",
INIT_06 => X"33992D98DEC74A003EA468D01510C03E8F580C800A3F018200418927E0668645",
INIT_07 => X"0204000406050013142409121142F746222EE2498000007E111204058B84C50C",
INIT_08 => X"E826A0602902A10491165C200000820018A5104010C01086003C13E000004EDF",
INIT_09 => X"023000000000000867000000000000040000600060801022C9F88D244FA40133",
INIT_0A => X"00100000820040482B28050001600010C13499F01B334015980001E09F000000",
INIT_0B => X"B80460124F16F06BC20CBC30CBC20CBC20CBC30CBC20CBC20CBC3065E1865E10",
INIT_0C => X"00000000029D204B7C0382FD0100F3F9F80FA0200E0BF40063F99C0010000012",
INIT_0D => X"93900F6EE230301208008001007A80001100002002801000A042000000000000",
INIT_0E => X"93900F6EEC421392C96B1237E0D8BD9629F97E0B348EDAC3900F6EFA0B158EDA",
INIT_0F => X"622DBC31D73F6006A5891533EF9500EAE64BCA0B158EDAC3900F6EFA0B348EDA",
INIT_10 => X"C2B083798D341B10DEFE14400392C74CAEAD412EDD2B4FCFF812A383430C669E",
INIT_11 => X"49FAB442994B3238D4E2FB104636652E19B8BA30C022DAD8C100CA39E8CEBE66",
INIT_12 => X"30469392526208C6CC95C33717D88532966471A9C5DD00B12728D5360234D62A",
INIT_13 => X"828C4999AF580395542D27CDBA0020F0FABAC800DA550C29F36A8A2554E48A64",
INIT_14 => X"40000000873FB80B8A00EF03F56CC12B416A51B60585A5C28895962502E9F36A",
INIT_15 => X"0000000000000000000000000000008000000410802A26924010000002000EE0",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"28C1111026C152A121960A884042020000000000000000000000000000000000",
INIT_19 => X"2082082082082082082082082082092492492492492400200005A8A28A200A37",
INIT_1A => X"964B2592C964B2592C964B2592C964B2590C86432190C86432190C8208208208",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF400FEB2592C964B2592C964B2592C",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FF00042ABEFFF8400010082EAABFF55002ABEF08000000000000000000000000",
INIT_1F => X"BEFFFFBD54000004155EFAA842ABEFA280155EFFFFBC01EF0855400005555421",
INIT_20 => X"8AAAA2D540000F7D57DF55A2AABFFEF08556AA10000028AAAFFD15541000002A",
INIT_21 => X"40000005168AAA087BFFFFF5D04001FF00041554555557FE005D003FE10AAFBE",
INIT_22 => X"1555FF082AA8B55F7AEA8BEF5551575FFA2FFD75FF550015400FFFBFFF450851",
INIT_23 => X"D57DF45A280154BA5555401EFFFD5421EFA2FFFFF555D0000145082E955FF085",
INIT_24 => X"051555FF0804155FFF7842AA100000020BAAA801541055042ABEFFFFBD5410AA",
INIT_25 => X"000000000000000000000000000000000000005568AAAAAD142145FF80155EF0",
INIT_26 => X"F145B42038555F401D71C0A2DBC7EB80000280824ADBD7490E28BEF080000000",
INIT_27 => X"82FFDB5243800002FBD7EBFBD24101C00175EFB6802DBC7BE8A155EFE3FBC71F",
INIT_28 => X"E1041003DE10BEF5EDAAAAAD547038EBD57DF7DA2AEB8FC7005F6AA381C0A2DA",
INIT_29 => X"5400E3F1FFF7D085B420381C5B6AA82147FF8FEF410E001FF000E17555555B7A",
INIT_2A => X"0017D142E905EF1451525C7082AADB45F7AEA8BEF555F575FFBEF5D05EF550E1",
INIT_2B => X"02FBEFEBFBD2410AADF78F45B68010482415B471C7E3DF451EFBEFBFAF454900",
INIT_2C => X"D145145FF84155D7085B555C71404105C7F7842FA381C0A00082AA8A10410410",
INIT_2D => X"02AA8BEF000000000000000000000000000000000000000000000005B68ABAB6",
INIT_2E => X"FFAE955EFAAFBD55EF557BC20AA5D7BC01555D2EBFF55A284000AA08003FF550",
INIT_2F => X"5007BE8AAA5D2EBDE00FFFFC00AA08003FF55A2FBC00105D04175FFF7803DF45",
INIT_30 => X"FF082A97555557FE8A0000043FE00F7D17FEBAA2D5574BAAAD17DFEFA2AEAAB5",
INIT_31 => X"5FFF7D5401EF5D2E97410AAD17DFEF007FC20AA5D7BE8A005D7FEABFF002E821",
INIT_32 => X"55EFF7FBE8B550004001FF5D2A801EF5D5142145082EBFF55F7AAAABEF5D7FD7",
INIT_33 => X"82010A2AA8000008043FFFFA2FBC2010A2FBEAB45F78402010007BD5545AAFFD",
INIT_34 => X"000000007BEAAAAFFD555545FF8015555007FD5545550400145FF843DEAA552A",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000007FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(12),        -- Port A data input
DOA(0)   => data_read_a_lo(12),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(12),        -- Port B data input
DOB(0)   => data_read_b_lo(12),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_13_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10110A0441812402840402822007818000E00700000000330A3000000008042",
INIT_01 => X"A1400986B830E84D182260000C1042484001000008220008A20019080A510200",
INIT_02 => X"10A108600C9141100000C6180CA85035010E4880010431004908135980122D60",
INIT_03 => X"0013881507460886C190832175809C02030400002020124C441A108468424842",
INIT_04 => X"203080680204A0113801D600864E0C96C12000008244244052200201801802C0",
INIT_05 => X"030004849601110204950409C0208C2084E0009C0000100120A00C9918002098",
INIT_06 => X"10000882804544921681428591908000AF28A8002BC00D020003896020658FC4",
INIT_07 => X"CA20400450050009100501501102E0042020448D0000023E10408144C800D800",
INIT_08 => X"1D2B00402B220104B53100200001020218A5104016CC1C616401910801010100",
INIT_09 => X"050800404D49A42EB08000000000000406481C8C408000A2D8088D1820200B00",
INIT_0A => X"0010000002004048AA08050401604462E9144002090740148441200484000500",
INIT_0B => X"000A112100000000010000000001000000000000001000000000000000800000",
INIT_0C => X"509528954404144C200425010040000001B020081094040072005C0030864208",
INIT_0D => X"1C10B3831034081200000000000430003000206822F20CA8826AC2A14250A128",
INIT_0E => X"1C10B383110218CB0E54C2EA404A4F03D404A41AA5B7344C10B383081BA4B734",
INIT_0F => X"8001CE3E20A5B284ED1132909C72885A2B2C381BA4B7344C10B383081AA5B734",
INIT_10 => X"AC3CC0C0B8182597A801610218CB0C3548B3A008E730A01AB113A5524E6ACA67",
INIT_11 => X"A151EC5952E44128CA194517354C180A3C066430202021252991C22C99731014",
INIT_12 => X"1804C8A0ADA2E6A983014780CA28B2A5C8825194332B018A444AEA2701288A15",
INIT_13 => X"02D09852745F80112C428562EE0353635232D50048A411C158BB0A7910142C77",
INIT_14 => X"4240480068001C9B9150A0000297046E4023F8BE8E3E1E0109472C3EB50158BB",
INIT_15 => X"A1284A1284A1284A1284A1284A12851A84284110406A26924302590806000110",
INIT_16 => X"1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284",
INIT_17 => X"284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A",
INIT_18 => X"7DDFE7EFBEFFE7D3EFBEFC48A0550000000000000000000A1284A1284A1284A1",
INIT_19 => X"D75D75D75D75D75D75D75D75D75D75D75D75D75D75D7EFBFBFBBAAAAAABEFDF7",
INIT_1A => X"5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5D75D75D75",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000FEFD7EBF5FAFD7EBF5FAFD7EBF",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"AA5D043FFFFAAAABDEAA557BFDE00FFD140155F7800000000000000000000000",
INIT_1F => X"400AAD540155A2D5421FF00042ABEFFF8400010082EAABFF55002ABEF08556AA",
INIT_20 => X"ABEFA280155EFFFFBC01EF08554000055043DEBAF7843FFFFF7AABDF55A2AA97",
INIT_21 => X"D5400005568A1055043DEBAAAFFE8B45557FD7410552EAAABAAA84155EFAA842",
INIT_22 => X"FE8ABAAA8428A00087BD7555FFD56AA10000028AAAFFD15541000002ABEFFFFB",
INIT_23 => X"803FE10AAFBE8AAAA2D540000F7D57DF55A2AABFFEF085557545FFD17DEBAA2F",
INIT_24 => X"0041554555557FE005D0000155557BEAABA5D2ABDF450851420AA5D7FD5555A2",
INIT_25 => X"000000000000000000000000000000000000005168AAA087BFFFFF5D04001FF0",
INIT_26 => X"7490E28BEF08516DA82410A3FFD7AAA4B8E824971F8E38E3DF45155EB8000000",
INIT_27 => X"D7EBA4BDF45AAAA90410BEDF45155A2DF401D71C0A2DBC7EB80000280824ADBD",
INIT_28 => X"A82B680175EFB6802DBC7BE8A155EFE3FBC71FF145B42038550E38E92EB803FF",
INIT_29 => X"243800002FBD7EBFBD24101C556FA38490A3FE92BEFFEAB45417FD24385D2AAF",
INIT_2A => X"5056DE3D17FE92BEF1EFA92AA8428A10007FD557DFFDF6AA381C0A2DA82FFDB5",
INIT_2B => X"B400925D7FD557DA2803DE10BEF5EDAAAAAD547038EBD57DF7DA2AEB8FC70051",
INIT_2C => X"7FF8FEF410E001FF000E17555555B7AE10410E00155497FEFABA4120B8F55085",
INIT_2D => X"2FBD7545AA8000000000000000000000000000000000000000000005B6AA8214",
INIT_2E => X"A284000AA08003FF55002AA8BEF00517FE00082EBDF45AA8428A10085568ABAA",
INIT_2F => X"A5D2EA8A00A2803DF45AA843DF55AAAE82000F7FBD5545AAFBC01555D2EBFF55",
INIT_30 => X"55087FC00BA552ABFE10F784175FFF7803DF45FFAE955EFAAFBD55EF557BC20A",
INIT_31 => X"AAA5D2EBDE00FFFFC00AA08003FF55A2FBC00105D517FEAA082EBFE10F7FFE8B",
INIT_32 => X"DFEFA2AEAAB550051401FFA2D57FE10F7D57DE00AA842AA00007FD75FFF7FBE8",
INIT_33 => X"FDEAA08042AB45087FC0010557FD55FFAA843FE00F7D17FEBAA2D5574BAAAD17",
INIT_34 => X"000000007BE8A005D7FEABFF002E821FF082A97555557FE8A00002E82155007B",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000067FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(13),        -- Port A data input
DOA(0)   => data_read_a_lo(13),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(13),        -- Port B data input
DOB(0)   => data_read_b_lo(13),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_14_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10020A000180000284008280000281800000030000000033022000000580002",
INIT_01 => X"A14009821830284D186860000C30C24840000000084000084200090008510200",
INIT_02 => X"102100600C9001100000061020A8503401044880010400204908012018122F64",
INIT_03 => X"00008015074608840190800010008002030400002074F401209A108448404842",
INIT_04 => X"000080400004A00100004000840E000201000000024024401200020180180080",
INIT_05 => X"0A000484800111020495040800208C2084000080000010010020049818002008",
INIT_06 => X"1000088020450402B6A1420511C080008468A80008000D0200018B202067AF10",
INIT_07 => X"422000044005000910040110510260040024400C800000BE3850A144C924080E",
INIT_08 => X"000B004028020104111100200001020210A51040008004616001910801010000",
INIT_09 => X"000800004D492408208000000000000406401C0C40800022C8088DB420200900",
INIT_0A => X"0010000002004048000005040160042229140002090200000401000484000400",
INIT_0B => X"0000110100000000010000100000000000000100000000000000100000000000",
INIT_0C => X"409120940404104C2000210100400000011020080084040040005C0010820208",
INIT_0D => X"E0E0A0000190081200000000000000003000000000100C088020028102408120",
INIT_0E => X"E0E0A0000B02740421A0E5D1A024002050805210040000B0E0A0000210040000",
INIT_0F => X"E01200860008920106460D4501CB000111300210008000B0E0A0000210008000",
INIT_10 => X"0ABBC00905C33C6000400F02740412C0715C40110080A4006110510C14D18178",
INIT_11 => X"20000041DB011CC000090012565306500002411420220080220C0093C3892324",
INIT_12 => X"5809240C09024A4AE0CA00004800839682398000120800658992F3C700C30181",
INIT_13 => X"002B46867DBC002A830280000800F7B7A0B1E240240A8340000200067EAA8CB6",
INIT_14 => X"42004005800004801150A00341244000845C7DB0D0200900422ACA4B28000002",
INIT_15 => X"8120481204812048120481204812051A04204110002A26924302590802000000",
INIT_16 => X"1204812048120481204812048120481204812048120481204812048120481204",
INIT_17 => X"2048120481204812048120481204812048120481204812048120481204812048",
INIT_18 => X"69CB91FE1EF7D3ABEFBECA080050000000000000000000081204812048120481",
INIT_19 => X"F3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF7EFBBBBBF9E79E7BEAAF3",
INIT_1A => X"CFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCF3CF3CF3C",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FF007F3F9FCFE7F3F9FCFE7F3F9F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"45AAD157400007BEAAAAAAAE955555D5568A105D000000000000000000000000",
INIT_1F => X"0AAF784020AAF7D56AAAA5D043FFFFAAAABDEAA557BFDE00FFD140155F7D17DF",
INIT_20 => X"ABEFFF8400010082EAABFF55002ABEF085155400FFD1420100055574AAA2AA80",
INIT_21 => X"40155A28028B550051574005D7FFFE105D7BD7545A284020BA0055421FF00042",
INIT_22 => X"1421FF5D7FFDEBA085168B45FF843DEBAF7843FFFFF7AABDF55A2AA97400AAD5",
INIT_23 => X"04155EFAA842ABEFA280155EFFFFBC01EF08554000055002AB455D5142010085",
INIT_24 => X"57FD7410552EAAABAAA8017400AAD140000002EBFFEFA2AAA8BEFF780021FF55",
INIT_25 => X"000000000000000000000000000000000000005568A1055043DEBAAAFFE8B455",
INIT_26 => X"8E3DF45155EBD17FF6DAADB504001C71EDA82AAA0955455D556DA00490000000",
INIT_27 => X"101C55554AAAAA480082FF84000BAEBD16DA82410A3FFD7AAA4B8E824971F8E3",
INIT_28 => X"092085F401D71C0A2DBC7EB80000280824ADBD7490E28BEF085157428FFDB420",
INIT_29 => X"DF45AAAA90410BEDF45155A28E2AB7D0051504005D71F8E004975D556DB68405",
INIT_2A => X"28B6D5D51420101C5B401EF417BFAEAA08516AB45E38E38E92EB803FFD7EBA4B",
INIT_2B => X"EAFBC7EB80071FF5500175EFB6802DBC7BE8A155EFE3FBC71FF145B420385500",
INIT_2C => X"0A3FE92BEFFEAB45417FD24385D2AAFA82B68015400AADB40000082EBFFC7A2A",
INIT_2D => X"5557FE1000000000000000000000000000000000000000000000000556FA3849",
INIT_2E => X"AA8428A10085568ABAA2FBD7545AAD17DFFFAAFFC200055557DE00A280155455",
INIT_2F => X"F0051554AAFFFFC00105D55554BAA28400000F784020BAAAD17FE00082EBDF45",
INIT_30 => X"000051575FFF78415410087BC01555D2EBFF55A284000AA08003FF55002AA8BE",
INIT_31 => X"A00A2803DF45AA843DF55AAAE82000F7FBD5545AAAEAABFF0051400105D5568A",
INIT_32 => X"55EF557BC20AA5D042ABFF555142000557FC01EF007FEAABA00556AB55A2AEA8",
INIT_33 => X"C0010082EBDF55A2AABDF45A284175FF5D04175FFF7803DF45FFAE955EFAAFBD",
INIT_34 => X"00000000517FEAA082EBFE10F7FFE8B55087FC00BA552ABFE10F78415400A2FB",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000007FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(14),        -- Port A data input
DOA(0)   => data_read_a_lo(14),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(14),        -- Port B data input
DOB(0)   => data_read_b_lo(14),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_15_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000A000000000284000280000001800020030000000033022000000180002",
INIT_01 => X"A140098018300848180060000C00426040000000080000080200000000110200",
INIT_02 => X"1020004000801110000006100028503400040800010430004808000180120278",
INIT_03 => X"00008011064408840190800000228002A3000000000010000008108448000042",
INIT_04 => X"701280400004A991000000A28406000211000000220004941000000880000000",
INIT_05 => X"02000484800155020495000800218020C4002880005310000000040000000001",
INIT_06 => X"10000880004540000711224491C08000850A880008000D020001892020656300",
INIT_07 => X"8A04000016050009140501505100000420204008000000BE70408104C8000000",
INIT_08 => X"001F004028026104111002200000000200210040008004614001100801010000",
INIT_09 => X"000800000D09240000800000000000040600180840800022C8088C1020200000",
INIT_0A => X"0000000002004040000105000040042229140002080000000400000080000400",
INIT_0B => X"0000110100000000010000100001000010000000000000000000100000800008",
INIT_0C => X"0001008000000000000025000040000001300008009400006200580010000000",
INIT_0D => X"0000000002300012000000000004200030000000000008008020020000000000",
INIT_0E => X"0000000001000000400000000000000000000010108000000000000010108000",
INIT_0F => X"0000000000000200000900000000000000000010140000000000000010140000",
INIT_10 => X"0140000000000000000001000000400000000000000000000100008040000000",
INIT_11 => X"0000004000480000000000100004400000000030002000406000000000068409",
INIT_12 => X"8000000000020080080000000000802010000000000800000201000800000000",
INIT_13 => X"00000100000000000000000008000000184400A0000000000002000000441108",
INIT_14 => X"4000000000000000010620000004000000000242038B82800000000000000002",
INIT_15 => X"0000000000000000000000000000041800000110000024130202500802000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000080050000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"000804154AA5D00001EFF78428AAA007BC2145F7800000000000000000000000",
INIT_1F => X"0AA007FC2000F7D17DF45AAD157400007BEAAAAAAAE955555D5568A105D7FC00",
INIT_20 => X"FFFFAAAABDEAA557BFDE00FFD140155F7FBD74AAAAD17DF45F7D1421EF005540",
INIT_21 => X"020AAF7FFFDF45FF84000BA552ABDFEF08517DF55A2FBEAB555D556AAAA5D043",
INIT_22 => X"FEAB45F7843FF45082A801FF005155400FFD1420100055574AAA2AA800AAF784",
INIT_23 => X"D5421FF00042ABEFFF8400010082EAABFF55002ABEF087BE8ABA555168B55AAF",
INIT_24 => X"D7BD7545A284020BA007FFFE10A284000AA0055401550055574005D2E800AAA2",
INIT_25 => X"000000000000000000000000000000000000000028B550051574005D7FFFE105",
INIT_26 => X"55D556DA004971C7038140012482550E021C7EB8028A821C7BC516DFF8000000",
INIT_27 => X"45E3DF471C70851400BA0071C5028FFD17FF6DAADB504001C71EDA82AAA09554",
INIT_28 => X"B555D516DA82410A3FFD7AAA4B8E824971F8E38E3DF45155EBF1D5492BED17FF",
INIT_29 => X"54AAAAA480082FF84000BAEBF1FFF7DEB8000092552ABFFEF08517DF6DB6FBE8",
INIT_2A => X"EFA8241516DB55A2FFEAB6DEB843DF551C20801C71C5157428FFDB420101C555",
INIT_2B => X"550428412A85082BEDF401D71C0A2DBC7EB80000280824ADBD7490E28BEF087F",
INIT_2C => X"51504005D71F8E004975D556DB68405092087FF8E00BE8A02082005F47145085",
INIT_2D => X"57BD75EFF78000000000000000000000000000000000000000000000E2AB7D00",
INIT_2E => X"55557DE00A2801554555557FE100055554BA5504000105D2A80145AA842AA005",
INIT_2F => X"5AAD557410F7D57DF55AAFBD55450055420BA0055574BAF7D17DFFFAAFFC2000",
INIT_30 => X"FF08517FFFFF7FBEAB455D517FE00082EBDF45AA8428A10085568ABAA2FBD754",
INIT_31 => X"4AAFFFFC00105D55554BAA28400000F784020BAAAD57FFEFA28402010552ABDF",
INIT_32 => X"FF55002AA8BEF007FFDE1000557DF45AAFBE8BEFA2803FF45550400155555155",
INIT_33 => X"80000087BD55450855400BA002A95400F7FBC01555D2EBFF55A284000AA08003",
INIT_34 => X"000000002EAABFF0051400105D5568A000051575FFF78415410087FEAA10F7AE",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000060000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(15),        -- Port A data input
DOA(0)   => data_read_a_lo(15),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(15),        -- Port B data input
DOB(0)   => data_read_b_lo(15),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_16_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"DA22C618B1000482B688B186588884862A400438255FC38381441205BA803003",
INIT_01 => X"264AC80028404C211203A952A90341080B173340412000E1005D628000820484",
INIT_02 => X"400034C206C405000001A48202084004003008255040826EE008B440200E2042",
INIT_03 => X"2916704900606AC82B49CC56DF8CC1E50E4800202115005760010010000C0400",
INIT_04 => X"052DCA856DC7504B82BF6614C86D2B7F85AAD17F4B100000B88148C4804A428A",
INIT_05 => X"373CB02A00C0502F301180141A42A5720E0F43C17A8479580001AC20000000E2",
INIT_06 => X"303E2094282B85242C85001038D5710E8410D5959BC4800015001219D0550077",
INIT_07 => X"880100000159954501280B0080146F7112D949A0015018220540000382805001",
INIT_08 => X"30015452880C8D90409A05B2CB2CA400200209E5601044A24000000462A60018",
INIT_09 => X"452D54000C0907000330000000000096480050000685400005FC014743E0DC92",
INIT_0A => X"00014808A02004200E540480212000A448C0080024AEA00C9688000000000005",
INIT_0B => X"000D58460018F6D3D84400044000440004400044000440004400042000220002",
INIT_0C => X"0001004010A8812831605DA0000A054052E40000817680220040025699200002",
INIT_0D => X"AAADA0C343F1AC1B01040A002024895514554485D00000012400240000000000",
INIT_0E => X"AAADA0CC421CA003B694B68018FAAA708E2CB5320018CAC99BA0A3B9320018CA",
INIT_0F => X"B1443A1891E4A928C29020E6A8524CE7A3EE59320018CAC99BA0ACB9320018CA",
INIT_10 => X"04B2A5A40B1E6644AF0F021EA003AC24352AB2449A3FF2FA04E5E09B128834AD",
INIT_11 => X"60ED838E890B703C6260D8E3A21275714C902375B801324301AB0067622E5E54",
INIT_12 => X"064F70DBDB1C74424E91E1C194C71D1216F50A8C241815FEB6A9158863F638FB",
INIT_13 => X"45FDF9D364DBD9435A6D45C9E81BED555E4C15F11133D171727A2550EE2F1BA0",
INIT_14 => X"08150013F162119014204373517700ACCC59432A2B2D001F803471A9A960E572",
INIT_15 => X"000000000000000000000000000000880002054000229088542210206B2AB015",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"2A898D21B4C98389ED146C080000000000000000000000000000000000000000",
INIT_19 => X"A29A29A29A29A29A29A29A29A29A28A28A28A28A28A53CBF0F0D3CF3CF0AB1A2",
INIT_1A => X"8F47A3D1E8F4FA7D3E9F4FA7D3E9F4FA7D3E8F4FA3D3E8F4FA3D3E9A29A29A29",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000FA7D3E9F4FA7D1E8F47A3D1E",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFF7FBE8B45AAD568BFFFFAA975FF00003FE0055000000000000000000000000",
INIT_1F => X"0005D2A95410FFFFC00000804154AA5D00001EFF78428AAA007BC2145F7843FF",
INIT_20 => X"7400007BEAAAAAAAE955555D5568A105D2E974BAF7FBEAB45FFFFC00BAF78002",
INIT_21 => X"C2000F78000010552E800AA002E821FFA2AAAAA00000417555FFD17DF45AAD15",
INIT_22 => X"43FEBA5D55575FFF7AABFE00557BD74AAAAD17DF45F7D1421EF0055400AA007F",
INIT_23 => X"D56AAAA5D043FFFFAAAABDEAA557BFDE00FFD140155F7AABDF55F7AE820AA080",
INIT_24 => X"8517DF55A2FBEAB555D04154BAA2FBE8B55FFFFD55FF557FC2000FF8015410FF",
INIT_25 => X"000000000000000000000000000000000000007FFDF45FF84000BA552ABDFEF0",
INIT_26 => X"21C7BC516DFF8438FC7E3F1EAB55B6DF6DBFFF7AA955C71C043FE10490000000",
INIT_27 => X"55FFF1C70BAF78A000005D2097438FFF1C7038140012482550E021C7EB8028A8",
INIT_28 => X"57DEBD17FF6DAADB504001C71EDA82AAA0955455D556DA00492490492F7FBE8B",
INIT_29 => X"71C70851400BA0071C5028FF84020285D2085092002A801FFB6AAA8A10080E17",
INIT_2A => X"BAF6DE3AA8709208043FEBA555B555FFE3AABFE005D71D5492BED17FF45E3DF4",
INIT_2B => X"BC0028E38412428EBD16DA82410A3FFD7AAA4B8E824971F8E38E3DF45155EBA4",
INIT_2C => X"8000092552ABFFEF08517DF6DB6FBE8B555D04124BAB6FBE8B45E3FBD55D7557",
INIT_2D => X"5003DE000000000000000000000000000000000000000000000000071FFF7DEB",
INIT_2E => X"5D2A80145AA842AA00557BD75EFF78428B55AAD168B55F7FFFDFEFFFAA955555",
INIT_2F => X"0000000010F7FBEAB45FFD1554AAFFAE820105500154AAF7D5554BA550400010",
INIT_30 => X"EFF7AEA8A10002E955FFA2D17DFFFAAFFC200055557DE00A2801554555557FE1",
INIT_31 => X"410F7D57DF55AAFBD55450055420BA0055574BAF784000BA5D0017410082E801",
INIT_32 => X"8ABAA2FBD7545AA802ABEFA2AA9541000003DEBA557BD75EFA2AEBDE105D5557",
INIT_33 => X"EAB45AAFFD55555D7FC20AAA280000AAAAD17FE00082EBDF45AA8428A1008556",
INIT_34 => X"00000000557FFEFA28402010552ABDFFF08517FFFFF7FBEAB455D04020AAFFFB",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000020000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(16),        -- Port A data input
DOA(0)   => data_read_a_lo(16),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(16),        -- Port B data input
DOB(0)   => data_read_b_lo(16),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_17_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"5284CE4FB7BD2C8994A13392DBD02E14006B82AC7E800D44D3DD2FD5F9B961C0",
INIT_01 => X"F9BA301F7E03FC6793F2199B39FC233C11D93AE6F3BB92B32091DBC339B24542",
INIT_02 => X"1D5FC0C08F040404446965C0607FB8A217C400C33A908078551BD04222186338",
INIT_03 => X"A14124C28DFD960832C90446DF8400A5055C25295B695FF97E1B5AC757F06D6B",
INIT_04 => X"04A106866DA3D02A01FB660C08A4AB7F840EDB6F48100DFC8081081D78AC7402",
INIT_05 => X"51E072F0C0C58D9C125EBFC00A46CF0388054100F680E0CE0107B8D040DAFCDA",
INIT_06 => X"019A4D00786B048112C58B16307F15DE8408B233661C10BBA5DAAFA9DDA1194D",
INIT_07 => X"8E00001660700CE170284A00891C7C03D29DE26814515835902AC089A2801540",
INIT_08 => X"C009F3A1B0120A1C51DFF881861CBE0305A12A0321810217C01D34EDC98FFA1C",
INIT_09 => X"747E6610052CDEE97FF1F9F63E3EF790380078002CE976AB6BF769769E4D437D",
INIT_0A => X"00185C44B91BC1740B7605040BE0018CFC7429F326B9D045FF8000E9AB415606",
INIT_0B => X"3A28FC1AAF5CF6F3D3EF3D3EF3D3EF3D3EF3D3EF3D3EF3D3EF3D3EF9E9F79E9E",
INIT_0C => X"0000020012E9E10A31EB5FF9296A67F5B4FFBD2FAD7FE653C3FBFF33E10C001B",
INIT_0D => X"333EA16031F2BD47BDA2CA5D8164FCCFE833C5C3D00018006C68170000000000",
INIT_0E => X"333EA160391BEFF2C32FB695F919110D5ECE542A6FEEB2533EA160782A6FEEB2",
INIT_0F => X"D18C0D06638A207CFDE1F7DDAD76D5282400F82A6FEEB2533EA160782A6FEEB2",
INIT_10 => X"E6E43E59AFE4A59B57679D19EFF2C7573FAD5A86840354D1706FFFA3EF6E24B6",
INIT_11 => X"F7D7A0ABD6DAAAB96529382B74E4E1FE4ACA4D77FAAB77CE3AF3EE78F58DB737",
INIT_12 => X"2D1281017F056E9C9C3FC95949C157ADB55572CA52606DFED6CA55334C04C04F",
INIT_13 => X"59FDEB974F486905001FDF5FA0D719F9956EAA1A184045D5D7A870D2F5A5D752",
INIT_14 => X"60158015177F916A039EF41FDB34A91F432EA58949D5B5C85F97871876F7D7E8",
INIT_15 => X"000000000000000000000000000004DC200005E705B7B3D9FC22F00BE419FB55",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"06013DB9880A5D22E229F3030018000000000000000000000000000000000000",
INIT_19 => X"D35D74D35D74D34D35D74D35D74D34D34D34D34D34D0D30D0D303AEBAE886E40",
INIT_1A => X"51A8D46A351A0D068341A0D068341A0D068341A8D468341A8D46834D35D74D34",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000008D46A351A8D46A351A8D46A3",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFF7FBFDF55A28402000F7D56ABFF55000000000000000000000000",
INIT_1F => X"A00F7843FEBA55043FFFFF7FBE8B45AAD568BFFFFAA975FF00003FE0055043FF",
INIT_20 => X"54AA5D00001EFF78428AAA007BC2145F7D568B45000002010552EBDF45A28028",
INIT_21 => X"95410FFAE800105D2A95410002A95410AAAEBFF55AAFFC00BAF7FFC000008041",
INIT_22 => X"57DE00F7AE800AAAAAABDFEF5D2E974BAF7FBEAB45FFFFC00BAF780020005D2A",
INIT_23 => X"517DF45AAD157400007BEAAAAAAAE955555D5568A105D7FFFFEFA2D568BFFFFD",
INIT_24 => X"2AAAAA00000417555FF8028B55082A974105D003FF55F7802AAAAAAD168AAA5D",
INIT_25 => X"000000000000000000000000000000000000000000010552E800AA002E821FFA",
INIT_26 => X"71C043FE10490A3FFFFFFFFFDFEFE3F5FAF45AA8000038F7DB6FBD7490000000",
INIT_27 => X"384124BFF7DB68A28A38F7803DE82490438FC7E3F1EAB55B6DF6DBFFF7AA955C",
INIT_28 => X"0BAFFF1C7038140012482550E021C7EB8028A821C7BC516DFFDF68B551C0E050",
INIT_29 => X"70BAF78A000005D2097438FFAA85000492495428082E95400AAA0BDF7DB6F5C7",
INIT_2A => X"FAFFFB6D56FBFFEBDB78E38F7AA800BAB6AEBDFD75D2490492F7FBE8B55FFF1C",
INIT_2B => X"028AAAB6D16FA8249517FF6DAADB504001C71EDA82AAA0955455D556DA00497F",
INIT_2C => X"2085092002A801FFB6AAA8A10080E1757DEB8A2DB5514249243841003FF6DEB8",
INIT_2D => X"7FFFDF550000000000000000000000000000000000000000000000004020285D",
INIT_2E => X"F7FFFDFEFFFAA9555555003DE00002ABFFEFF7FBFDFFFAAD168B55AA80000BAF",
INIT_2F => X"FF7FBEAB45552E954BA08003DFFFFFAAA8AAAF7843FE10000428B55AAD168B55",
INIT_30 => X"10AA843FFFFF7D5554BAF7D5554BA5504000105D2A80145AA842AA00557BD75E",
INIT_31 => X"010F7FBEAB45FFD1554AAFFAE820105500154AAF7AE974000800154AA002E954",
INIT_32 => X"554555557FE10007FEABEFFFD57FFEFAAFFE8ABAFFAA820BAF7AEBFF55550000",
INIT_33 => X"020AA08003DFFFA28028AAAF7D17DE0000517DFFFAAFFC200055557DE00A2801",
INIT_34 => X"0000000004000BA5D0017410082E801EFF7AEA8A10002E955FFA2AABFF455500",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000067FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(17),        -- Port A data input
DOA(0)   => data_read_a_lo(17),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(17),        -- Port B data input
DOB(0)   => data_read_b_lo(17),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_18_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"69844019080000A21A611406840014122A641074155FC28A2024001001801003",
INIT_01 => X"01067920034004180005E9E3C90360C0041C0181002001602025800008440084",
INIT_02 => X"40AC3CAA22D605200000856E2481902400344A20F802C22054001000021E2379",
INIT_03 => X"A95308ECD3207AC81D91C4002004C08A06008080BA868007E58040102B0E0100",
INIT_04 => X"044CC183800CA00780808004C8DB841405A80A100B586200FAC24AE4805242CA",
INIT_05 => X"771C10000000000B1135883C08A115320E0401C0200038394230070A19000020",
INIT_06 => X"3001499C602A8A003E800A042D8132A00098408F79E3901218050018024110D6",
INIT_07 => X"5029401000C983E60004010030400353C05806800104004E0000042E52800E20",
INIT_08 => X"0000117088080990419005B0C309402030060860E01004A828408800440405E3",
INIT_09 => X"6B8186185C42900693A002004040001E1950850C848601008708114A2030B480",
INIT_0A => X"100180A8062026000DC425C0301311324AA237108857220BA089420440000030",
INIT_0B => X"C44703657083080C2800C2000C2000C2000C2000C2000C2000C2000610006100",
INIT_0C => X"C1B0609C05013065CC042004040808084001E000108010230400800FD9B286C4",
INIT_0D => X"CCC15F9CBA45505640000A402019003F140FC2060014250B9080008306C18360",
INIT_0E => X"CCC15F9FB1962FCB69E08AAAEAEBCDDF7C728582081483ACC15F9C3982081483",
INIT_0F => X"EBF1CFFF7670ACC3811A28AB57523CDFEBFBF982081483ACC15F9F3982081483",
INIT_10 => X"C9002BF05800D875E63CC9962FCB52CAA02FE3F8E7F5E3AC3620805298B15A3F",
INIT_11 => X"F1B72A8A800B7546DB9F1CA320037F01BD67DC4041D4CF03138DD865103EFEEA",
INIT_12 => X"81CCFAFDBF9464006FD037AEFAE5150016EA8DB7BFE25208E8F46A228BF8A757",
INIT_13 => X"641256EC844B8AF92FD7CEDC24A9E181A8A29509EAAE7FD3B749471C48F8A459",
INIT_14 => X"0297D086E00036D2440E0880AAD62BEFF5778802A3AF8E8FB0440CE78773B709",
INIT_15 => X"8360D8360D8360D8360D8360D83609220D20D00000080C0601400B402307E480",
INIT_16 => X"360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D",
INIT_17 => X"60D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8",
INIT_18 => X"D9D701DC2E784601EFBE2C00000000000000000000000008360D8360D8360D83",
INIT_19 => X"5155555545145145155555545145145145145145145220B22A0B820820965177",
INIT_1A => X"44A25128944A25128944A25128944A25128944AA552A954A2512895554514514",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000025128944A25128944A251289",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFEFF7AE954BA5D04174AA00000000000000000000000000",
INIT_1F => X"145AA801741000043FFFFFFFFFFFFFF7FBFDF55A28402000F7D56ABFF55043FF",
INIT_20 => X"8B45AAD568BFFFFAA975FF00003FE0055043FFFFFFFFFDFEFA2D56AB45AA8400",
INIT_21 => X"3FEBA55557FFEFA2D168B55AAFBFFFFFFF80021EF0855421EF00043FFFFF7FBE",
INIT_22 => X"A82155F7AEBFEBAFFD56AA00A2D568B45000002010552EBDF45A28028A00F784",
INIT_23 => X"FFC00000804154AA5D00001EFF78428AAA007BC2145F7D5400000004020AA5D2",
INIT_24 => X"AAEBFF55AAFFC00BAF7AE80010082E954BA0004174AAAA8428B45082ABFEBAA2",
INIT_25 => X"000000000000000000000000000000000000002E800105D2A95410002A95410A",
INIT_26 => X"8F7DB6FBD7490E3FFFFFFFFFFFFFFFFBFDFEFFFAE954AA550415492140000000",
INIT_27 => X"D7AAD16FB6DBE8E00155BE8015410140A3FFFFFFFFFDFEFE3F5FAF45AA800003",
INIT_28 => X"1C7140438FC7E3F1EAB55B6DF6DBFFF7AA955C71C043FE1049043FFEFE3F1F8F",
INIT_29 => X"FF7DB68A28A38F7803DE82495B78FC7AAD56FB6DBEF1FAFD7E384001EF145B47",
INIT_2A => X"420381C0A02082492A85155E3A4BDE92FFD56FA28B6DF68B551C0E050384124B",
INIT_2B => X"E28B7D1420BDEAAA2F1C7038140012482550E021C7EB8028A821C7BC516DFFD1",
INIT_2C => X"2495428082E95400AAA0BDF7DB6F5C70BAFFAE870280024904BA1400174AABE8",
INIT_2D => X"50415410550000000000000000000000000000000000000000000002A8500049",
INIT_2E => X"AAD168B55AA80000BAF7FFFDF55002ABFFFFFFFFFFFEFF7FBFDFFFF7AA974BA5",
INIT_2F => X"000043DFEFA2D56AB45AAD57DFEFF7AA82155F78015400552ABFFEFF7FBFDFFF",
INIT_30 => X"55A280021EF557FD7555550428B55AAD168B55F7FFFDFEFFFAA9555555003DE0",
INIT_31 => X"B45552E954BA08003DFFFFFAAA8AAAF7843FE10007FEAB55A2D17FFEFFFD568B",
INIT_32 => X"AA00557BD75EFF7D1400AA5D2A82000002A95545A2843FE00F7D17FEAAF7FBEA",
INIT_33 => X"020AA5D04154BAF7AEA8BEF55003DEAAA2D5554BA5504000105D2A80145AA842",
INIT_34 => X"000000002E974000800154AA002E95410AA843FFFFF7D5554BAF7AE974BA0004",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000020000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(18),        -- Port A data input
DOA(0)   => data_read_a_lo(18),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(18),        -- Port B data input
DOB(0)   => data_read_b_lo(18),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_19_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"042200000000000041088001001AA00000000000000000000000500802000003",
INIT_01 => X"074018000024000000000404000000000A22000800000800004A200000000001",
INIT_02 => X"0000048002C405000000000006A84000000000200893C246A20000000020031A",
INIT_03 => X"020A9639044012C80001C4000004C08006000000001025000000000000000000",
INIT_04 => X"0400C0800000000380800004C8000000058800000B1000009880480480024200",
INIT_05 => X"420410000000000B10804004080001320E0401C0200038080000000000000000",
INIT_06 => X"2002409006F00A8428050A000280493104004500480090080A01120220140020",
INIT_07 => X"0000000000418026090240923240002190400000000000C0054A912054004021",
INIT_08 => X"0000115080000990000000B0C308000000000860200160000000000038380000",
INIT_09 => X"8000F80001012590001000000000001618000000020280008180810200000000",
INIT_0A => X"0000000000000000000000000000000100008000110000000000000000000017",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000840007600000000000000000800259000000",
INIT_0D => X"0008A0034078104B41A41000000000031400C002000000000000000000000000",
INIT_0E => X"0008A0004263C0343EDD414004042228DC0D385598035D0008A003B05598035D",
INIT_0F => X"040231068187C39F5A4F985C008902041124505598035D0008A000B05598035D",
INIT_10 => X"1BFBD406451B02000E033263C0343CB740500401180DE053A98F6ECC739D8140",
INIT_11 => X"420851546B2400000040D8549B5800000010227848D4303807FC8CC5508AEAED",
INIT_12 => X"52210402120A936B0000000004C2A8D6480000000018A700FCF980CC300318A2",
INIT_13 => X"B1427ED430B41402D025082359700181C21140E40511802208D6B30C48F8A8A4",
INIT_14 => X"9C000018440021011821B35254E99AF9E9410006362A2B6424287B08286208D6",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000023006000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"7747E18E0218CC18E88324000000000000000000000000000000000000000000",
INIT_19 => X"34C30C30C30C30D34C30C30C30C30C30C30C30C30C3504118982A69A6980E411",
INIT_1A => X"C26130984C26130984C26130984C261309A4D26130984C26130984C30C30C30D",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000130984C26130984C26130984",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAA954BA5500020BA5D000000000000000000000000",
INIT_1F => X"4BA5D517FFFF08043FFFFFFFFFFFFFFFFFFFFEFF7AE954BA5D04174AA007BFFF",
INIT_20 => X"FFFFF7FBFDF55A28402000F7D56ABFF557BFFFFFFFFFFFFFFFFFBFDFEFFFAA97",
INIT_21 => X"17410007BFFFFFFFFFFFFEFF7D16AB45AA8002000F7D5575455D043FFFFFFFFF",
INIT_22 => X"568B55F7AE955FFAA840201008043FFFFFFFFFDFEFA2D56AB45AA8400145AA80",
INIT_23 => X"043FFFFF7FBE8B45AAD568BFFFFAA975FF00003FE00557BFFFFFFFFBFDF45AAD",
INIT_24 => X"F80021EF0855421EF002ABFFEFF7D168B55AAD17FFEFF7AE975FF00557FFFF5D",
INIT_25 => X"00000000000000000000000000000000000000557FFEFA2D168B55AAFBFFFFFF",
INIT_26 => X"A5504154921471FFFFFFFFFFFFFFFFFFFFFFFF7AA954BA550000082550000000",
INIT_27 => X"EFF7FBFAFD7E3A4954BA555B7AFC7080E3FFFFFFFFFFFFFFFFBFDFEFFFAE954A",
INIT_28 => X"545550A3FFFFFFFFFDFEFE3F5FAF45AA8000038F7DB6FBD74975FFFFFFFFFFFF",
INIT_29 => X"FB6DBE8E00155BE8015410147FFFFFFF7FBF8FC7EBD568B55A28000000FFDF52",
INIT_2A => X"FDFC7E3F1FAF55A2DB6FB7DF7AE955C7BE800000008043FFEFE3F1F8FD7AAD16",
INIT_2B => X"0955FF145B7AFC7410438FC7E3F1EAB55B6DF6DBFFF7AA955C71C043FE10497B",
INIT_2C => X"D56FB6DBEF1FAFD7E384001EF145B471C71424B8FC7E3D56AB6DB6DF7AFC7EBA",
INIT_2D => X"50002000550000000000000000000000000000000000000000000005B78FC7AA",
INIT_2E => X"F7FBFDFFFF7AA974BA55041541055517FFFFFFFFFFFFFFFFFFFFEFF7AA974AA5",
INIT_2F => X"500517FFFFFFFBFDFEFFFFFEAB45AA80154AA557BEAB45002ABFFFFFFFFFFFEF",
INIT_30 => X"55A28002000F7FFC2155552ABFFEFF7FBFDFFFAAD168B55AA80000BAF7FFFDF5",
INIT_31 => X"FEFA2D56AB45AAD57DFEFF7AA82155F78015400557BFDFEFF7FBEAB55A2D56AB",
INIT_32 => X"555555003DE00007FFDF45AAD568B45AAFBFFFFFFFAA95545F7840201000043D",
INIT_33 => X"6ABFFFFFBEAB45A280155EF557FE8B55000428B55AAD168B55F7FFFDFEFFFAA9",
INIT_34 => X"000000007FEAB55A2D17FFEFFFD568B55A280021EF557FD755555042AB55AAD1",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000040000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(19),        -- Port A data input
DOA(0)   => data_read_a_lo(19),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(19),        -- Port B data input
DOB(0)   => data_read_b_lo(19),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_20_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000003",
INIT_01 => X"A65FF80000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000048002CC070000000000000000000000002FF86100200000000220002362",
INIT_03 => X"00000000000203D80025DC18004DC3D01E000000000000000000000000000000",
INIT_04 => X"07E5DF808071026F87C4191DD8005080679800000F300002998058068002C000",
INIT_05 => X"C205F23A2100557F70000004390021F61E1E87C3FD0CFBF80880072042000044",
INIT_06 => X"1209244C2000100006800000020010000008407FC800B0000000100600040000",
INIT_07 => X"8802000009FFBFE51886018002040020000800000554003E0000000002800000",
INIT_08 => X"30801F5780259FB0000000F7DF78020004011FEFE00000000020031502000083",
INIT_09 => X"00000000001000000000000000000056F8000001000000040000040141800802",
INIT_0A => X"0000000000000008000800000000000000000000000000000010010014800000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"00010240001721214E000004000000080000008000001000040080FFDB000000",
INIT_0D => X"0000000F3008001E00000000001803FF14FFC006000000008010200000000000",
INIT_0E => X"0000000F3040200000020000000026A70C0008020000200000000F3002000020",
INIT_0F => X"000030B86000400080000200000000004A58F0020000200000000F3002000020",
INIT_10 => X"0000000002183E61E6000040200001000000000019B140000800800000020000",
INIT_11 => X"C00010080000000000525801000000000014AC08000000508001030A0A400100",
INIT_12 => X"000002BC360020000000000292C0100000000000A56000090100000000001F86",
INIT_13 => X"8010000000000000574500001001060600000000001716800000803102020000",
INIT_14 => X"00000000000040040040002000080506049CDF70C08040100000706707600000",
INIT_15 => X"00000000000000000000000000802040200200604040000000000024FB7FE008",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"060070400020112240209A408004000000000000000000000000000000000000",
INIT_19 => X"65965965965965965965965965965861861861861860D30424343CF3CF340E00",
INIT_1A => X"90C86432190C86432190C86432190C86432190C86432190C8643219659659659",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000086432190C86432190C864321",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974AA55040201008000000000000000000000000",
INIT_1F => X"4AA550002000007BFFFFFFFFFFFFFFFFFFFFFFFFFAA954BA5500020BA5D7FFFF",
INIT_20 => X"FFFFFFFFFFFEFF7AE954BA5D04174AA00003FFFFFFFFFFFFFFFFFFFFFFF7AA97",
INIT_21 => X"7FFFF087FFFFFFFFFFFFFFFFFFFFDFEFFFAE974AA5D003FE005D043FFFFFFFFF",
INIT_22 => X"BFDFFFAA84000105D556AB55557BFFFFFFFFFFFFFFFFFBFDFEFFFAA974BA5D51",
INIT_23 => X"043FFFFFFFFFFFFFF7FBFDF55A28402000F7D56ABFF55003FFFFFFFFFFFFFF7F",
INIT_24 => X"A8002000F7D5575455D2EBFFFFFFFFFFFEFF7FBEAB55A28000010F7D16ABEF08",
INIT_25 => X"000000000000000000000000000000000000007BFFFFFFFFFFFFEFF7D16AB45A",
INIT_26 => X"A550000082557FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550400028000000000",
INIT_27 => X"FFFFFFFDFEFF7AE974BA5500050380071FFFFFFFFFFFFFFFFFFFFFFFF7AA954B",
INIT_28 => X"E285D0E3FFFFFFFFFFFFFFFFBFDFEFFFAE954AA55041549214043FFFFFFFFFFF",
INIT_29 => X"AFD7E3A4954BA555B7AFC70871FFFFFFFFFFFFFFF7FBFDFFFFFAA974BA550038",
INIT_2A => X"3FFFFFFFFFDFEFF7F1FAFC7A28002028555F6FB7D5D75FFFFFFFFFFFFEFF7FBF",
INIT_2B => X"402010FFDB6ABEF140A3FFFFFFFFFDFEFE3F5FAF45AA8000038F7DB6FBD7490E",
INIT_2C => X"FBF8FC7EBD568B55A28000000FFDF525455524BFFFFFFFBFDFC7E3F5E8B45A28",
INIT_2D => X"504000BA080000000000000000000000000000000000000000000007FFFFFFF7",
INIT_2E => X"FFFFFFFEFF7AA974AA550002000557FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5",
INIT_2F => X"055043FFFFFFFFFFFFFF7FBFDFEFFFAE954BA5500174AA08517FFFFFFFFFFFFF",
INIT_30 => X"EFF7AE974AA550028AAA5D2ABFFFFFFFFFFFEFF7FBFDFFFF7AA974BA55041541",
INIT_31 => X"FFFFFFBFDFEFFFFFEAB45AA80154AA557BEAB4500557FFFFFFFFFDFEFF7FFFFF",
INIT_32 => X"00BAF7FFFDF55002EBFFFFF7FBFDFEFFFD568B55A284020BA557FFFFFF5D517F",
INIT_33 => X"FFF55A2D16AB45AA8402000F7FBEABEF5D2ABFFEFF7FBFDFFFAAD168B55AA800",
INIT_34 => X"000000007BFDFEFF7FBEAB55A2D56AB55A28002000F7FFC215555043DFEFF7FB",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000007FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(20),        -- Port A data input
DOA(0)   => data_read_a_lo(20),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(20),        -- Port B data input
DOB(0)   => data_read_b_lo(20),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_21_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"4A302428B824900A128C090A5C1800261500213C005FE812D10420054085A202",
INIT_01 => X"081FFE3440B609703B0427F801A40B8115BC4F655300340288A40D30040E4DD8",
INIT_02 => X"04CA478082CC1740002019824E0203100640303FF8C0B31061096E21A1840814",
INIT_03 => X"230CA7A4810083F80095DE00102DC3823EA821094EC68248923200013290C800",
INIT_04 => X"07CFFFC04904AA7F8780409DF84A0202879800000F3000029980780EA2C3C002",
INIT_05 => X"DE87F0280000407FF900D914382091FE1E1C0FC3E01EFFF8000480200008D062",
INIT_06 => X"010E2182002BC107A03448808F0D7C002822987FC830F40134CC74D002016612",
INIT_07 => X"0401000011FBFFE00520000200422033025C4209104500000012004C004D8C0B",
INIT_08 => X"00EF1F5FA0041FF080AC70FFDF78220010841EFFE7116E144071268DFD3E4C24",
INIT_09 => X"FC8BFE18008083B4443151462A28C6DFF80010002605302248088950484550A3",
INIT_0A => X"10018C241102068006C620C03882019480E631A0855E924E2598038938404037",
INIT_0B => X"A641165448C80C103648A3648A3648A3648A3648A3648A3648A366451B2451B2",
INIT_0C => X"011100841200D001000624000100C002804A08221890004806A310FFDF000454",
INIT_0D => X"5004D8158809C86065941840B1014FFF56FFC0281280080180B2948004400220",
INIT_0E => X"5004D815810D42E04A08A80098C02450025360694101816002D41A4068C10181",
INIT_0F => X"134160C8125B0B271802242880A04482418A0068C101816002D41A4069410181",
INIT_10 => X"10080E05C0B06AA8B12CFD0D42E0441A300012682960828F05C96A001B029010",
INIT_11 => X"00010362A8A20826A88660D86B202049F115100920C54E8EA256ECF078BA081C",
INIT_12 => X"064802C0081B0D64040936443306C55144104F30A8801406D002900062803201",
INIT_13 => X"4581BA0038005A706680012280506A8010602011819E290048A2118EC8140C08",
INIT_14 => X"CC158092C044600466208CC5091011C322A4C40A0300600C0A80509F41800880",
INIT_15 => X"80200802008020080200802008020412002001000000381C02004000FBFFF80D",
INIT_16 => X"0200802008020080200802008020080200802008020080200802008020080200",
INIT_17 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_18 => X"FDDFEFFFBEFFE7C7BFBEFC000000000000000000000000080200802008020080",
INIT_19 => X"F7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7FFBFBFFF9E79E7FFFDF3",
INIT_1A => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFDFEFF7FBFDFEFF7FBFDF7DF7DF7D",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00001FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D000200008000000000000000000000000",
INIT_1F => X"4AA5D00020AA5D7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550402010087FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAA954BA5500020BA5D7FFFFFFFFFFFFFFFFFFFFFFFFFFAE95",
INIT_21 => X"0200000003FFFFFFFFFFFFFFFFFFFFFFF7AA974BA5D0402000557BFFFFFFFFFF",
INIT_22 => X"FFFFEFF7AE974BA5D00174BA00003FFFFFFFFFFFFFFFFFFFFFFF7AA974AA5500",
INIT_23 => X"043FFFFFFFFFFFFFFFFFFFFEFF7AE954BA5D04174AA00003FFFFFFFFFFFFFFFF",
INIT_24 => X"FAE974AA5D003FE005D2EBFFFFFFFFFFFFFFFFFFDFEFF7AE954AA5500174BA5D",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFDFEFF",
INIT_26 => X"A550400028007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0000010000000000",
INIT_27 => X"FFFFFFFFFFFFFAA954BA5D00000BA557FFFFFFFFFFFFFFFFFFFFFFFFFFAE974A",
INIT_28 => X"0005571FFFFFFFFFFFFFFFFFFFFFFFF7AA954BA550000082557BFFFFFFFFFFFF",
INIT_29 => X"DFEFF7AE974BA55000503800003FFFFFFFFFFFFFFFFFFFFEFF7AA974AA5D0405",
INIT_2A => X"3FFFFFFFFFFFFFFFFFFDFEFF7AE954BA5D00154AA00043FFFFFFFFFFFFFFFFFF",
INIT_2B => X"A974BA5D00104925D0E3FFFFFFFFFFFFFFFFBFDFEFFFAE954AA550415492140E",
INIT_2C => X"FFFFFFFF7FBFDFFFFFAA974BA550038E285D2ABFFFFFFFFFFFFFFFFBFDFEFFFA",
INIT_2D => X"D00000100000000000000000000000000000000000000000000000071FFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE954AA5504000BA087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0557BFFFFFFFFFFFFFFFFFFFFFFFF7AA954BA5D00000BA5D7FFFFFFFFFFFFFFF",
INIT_30 => X"EFF7AE954AA5D041740055517FFFFFFFFFFFFFFFFFFFFEFF7AA974AA55000200",
INIT_31 => X"FFFFFFFFFFFFF7FBFDFEFFFAE954BA5500174AA08043FFFFFFFFFFFFFFFFBFDF",
INIT_32 => X"74BA550415410552ABFFFFFFFFFFFFFF7FBFDFFFFFAA974AA5D00174BA08043F",
INIT_33 => X"FDFEFF7FBFFFFFF7AE954BA5D0000010552ABFFFFFFFFFFFEFF7FBFDFFFF7AA9",
INIT_34 => X"00000000557FFFFFFFFFDFEFF7FFFFFEFF7AE974AA550028AAA5D2EBFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(21),        -- Port A data input
DOA(0)   => data_read_a_lo(21),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(21),        -- Port B data input
DOB(0)   => data_read_b_lo(21),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_22_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"5290F4CDE914905A14A43D33F488243E17122300F55FEB189B343A1140548380",
INIT_01 => X"A94007B259F6A975386262000C344BA9573C6FF57B18A5FB0ABFCD3C2C5F4F0C",
INIT_02 => X"D56B4302AC01005111011BD506AA5205274056900596A539584E2E6DFE4B2418",
INIT_03 => X"9AC0FCBD854688207C90007A1000047A00E588632CA213C8903AD6B55AD0EB5A",
INIT_04 => X"30002047A6FCA110086C402022F2124A8022492580040440002021C922D9109B",
INIT_05 => X"14A206B6838151008D95DD1847811C08002380041F1104002205AC4140DAD060",
INIT_06 => X"1727FF2EB9EF113A10BD32F44289D1F840C1710010344DB9A808FDFF3DE03130",
INIT_07 => X"050700154A00401D00495A06A8D464C5F6B54AA8551040818F4C997AC80CBE05",
INIT_08 => X"0141008801018040E48D50080002B00A0C00801014541E9504703680017F6CB4",
INIT_09 => X"02680000010937986481514E2A29CE010708C0804C6A033F7FCFF9426A41F1AB",
INIT_0A => X"00500001840000C80B410014088040F4A944B1AA313C004554002381B8000500",
INIT_0B => X"A004D1594832824A070AA070AA070AA070AA070AA070AA070AA0725503855038",
INIT_0C => X"501428054278142151262CA50343854E506A2C6898B2950AA6A35B0004284058",
INIT_0D => X"90078E1F840A2B0114020104022460002200050F60E220A06880D2A14050A028",
INIT_0E => X"90078E1F891C239F8908003099C1ACF06273612B3482C0C0078E1F412B1582C0",
INIT_0F => X"1BA1B0FD16770236A4091621C08055C2C0DB012B1582C0C0078E1F412B3482C0",
INIT_10 => X"00101F09C030AB28B03C111C239F870828041BA859F213AFC14AA38043006018",
INIT_11 => X"10E8822A984B0025B0DE6089462660095337B08AA600CA88B143AB11880C2806",
INIT_12 => X"055412D4481128C4CC012A66F304553096004B61BD8068B92400D0004E303689",
INIT_13 => X"589C48082C006A9057CA4385809520F07830001AC2173B00E162563454C40804",
INIT_14 => X"00460848952220592745AC11A544B1BF006850840180A00E1C81900C4190E160",
INIT_15 => X"22088220882208822088220882208CD888088D940D2A3A9D5002001300800C8C",
INIT_16 => X"0080200882208822088220882208822088220882208822088220882208822088",
INIT_17 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_18 => X"FBDFD1FE3EFBD7BBEFBEFA0A245120000000007FFFFFFFF20080200802008020",
INIT_19 => X"F3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF7FFBFAFBBBEFBEFBEFBF7",
INIT_1A => X"CFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCF3CF3CF3C",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000007F3F9FCFE7F3F9FCFE7F3F9F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040000000000000000000000000000000",
INIT_1F => X"4BA550000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0002000087FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974AA550402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"020AA5D7FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5D00000AA007FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAA954BA5504000AA557FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5D00",
INIT_23 => X"7BFFFFFFFFFFFFFFFFFFFFFFFFFAA954BA5500020BA5D7FFFFFFFFFFFFFFFFFF",
INIT_24 => X"7AA974BA5D040200055517FFFFFFFFFFFFFFFFFFFFFFFFAA954BA5500000BA5D",
INIT_25 => X"00000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000080000000",
INIT_27 => X"FFFFFFFFFFFFFAE974AA550002010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"0BA087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550400028007FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAA954BA5D00000BA557FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5D0002",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAA954BA5504020AA5D7BFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"A974AA5D00070925D71FFFFFFFFFFFFFFFFFFFFFFFF7AA954BA5500000825571",
INIT_2C => X"FFFFFFFFFFFFFFEFF7AA974AA5D040500055517FFFFFFFFFFFFFFFFFFFFFFF7A",
INIT_2D => X"D040200008000000000000000000000000000000000000000000000003FFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"A087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550002000087FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAA954AA5D00020AA007FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5504000B",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFF7AA954BA5D00000BA5D7BFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"74AA55000200055517FFFFFFFFFFFFFFFFFFFFEFF7AA974BA5504020BA557BFF",
INIT_33 => X"FFFFFFFFFFDFEFF7AE974AA5D00154105D517FFFFFFFFFFFFFFFFFFFFEFF7AA9",
INIT_34 => X"00000000043FFFFFFFFFFFFFFFFBFDFEFF7AE954AA5D041740055557FFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000007FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(22),        -- Port A data input
DOA(0)   => data_read_a_lo(22),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(22),        -- Port B data input
DOB(0)   => data_read_b_lo(22),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_23_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"EF20906D902424807BC8241BC81801B97D38AD3C0800103362A6741C80A12A02",
INIT_01 => X"001FFF8409F089003B4422000D80C80106804A7951C5B9D1C828043EA28838F9",
INIT_02 => X"028406A002DC176444683862400003111001303FFC00F240D50146013B300500",
INIT_03 => X"0006C90C010203F80005DC00C52FC380BEAC25886C02034800200200A1008008",
INIT_04 => X"17DFFF8049000BFF878314BFF8488890979800002F702002BB807A068403C280",
INIT_05 => X"DA07F0000000007FF020C814380011FE5E1C2FC3E05FFFF90020000808900010",
INIT_06 => X"10004C9690A8CA008024685184097E81E872C8FFE900FC31348EFDF03BE15E22",
INIT_07 => X"402000001FFBFFFD00080200B8140011F0D8C108155542018D1A302193E94004",
INIT_08 => X"41BE1F5F80003FF0002023FFDF79000000000EFFE309606020008005FC000000",
INIT_09 => X"FC83FE1840C0902400300000000000DFFD4004040C4D32BF7C0EE860003CE680",
INIT_0A => X"10018C24110A860006C620C0312241C482B20420CC56924E2199000C00415037",
INIT_0B => X"4669070510C90C14304043040430404304043040430404304043040218202182",
INIT_0C => X"008000105400C00400100000A018000801000C024000004A940000FFDF820604",
INIT_0D => X"100152100801C17E61841950B1C10FFF57FFC02812F00429DC92C40002000100",
INIT_0E => X"10015210088528E00E02C8200A430A424202A1CAF13F214001521001CBF03F21",
INIT_0F => X"01C1C044006D0C94FB94320880603C420B8001CBF03F214001521001CAF13F21",
INIT_10 => X"30182800A018D9CA8000648528E00D12480202C86040902AC60BACDF0E02D020",
INIT_11 => X"0445C19960A00026880C006739000009B00300010AF5052419D1964419028014",
INIT_12 => X"01844068880CE72000013600600332C140004D101808458A5602E00089202911",
INIT_13 => X"41D0B9023402085020825132C8CB5B4040301009408021144CB042F880100C06",
INIT_14 => X"8E17C0D240406519400500840A9524EE38A1F80E02120018390320F050144CB2",
INIT_15 => X"01004010040100401004010040100100040040000000000001000900FBFFE000",
INIT_16 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_17 => X"0040100401004010040100401004010040100401004010040100401004010040",
INIT_18 => X"0000000000000000000000000000000000000000000000001004010040100401",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000000000000000000000000",
INIT_1F => X"4BA5D0400010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000007FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974BA5D0002000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"00010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA550002000007FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAE974AA550400000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5500",
INIT_23 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550402010087FFFFFFFFFFFFFFFFFF",
INIT_24 => X"FAE954AA5D00000AA007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA55040200008",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010000000000",
INIT_27 => X"FFFFFFFFFFFFFAE974BA5D0400010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0000010007FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAE974AA550002010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA550002",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550400010087FFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"E954AA5D0402038007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550400028007F",
INIT_2C => X"FFFFFFFFFFFFFFFFFFAE954AA5D00020BA087FFFFFFFFFFFFFFFFFFFFFFFFFFA",
INIT_2D => X"D0402010000000000000000000000000000000000000000000000007FFFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000087FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAE974BA550002010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D000001",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFFFAE974AA550002000087FFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"54AA5504000BA087FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA550400010007FFF",
INIT_33 => X"FFFFFFFFFFFFFFFFAA954AA5D04000AA087FFFFFFFFFFFFFFFFFFFFFFFFFFAE9",
INIT_34 => X"000000007BFFFFFFFFFFFFFFFFFFFFFFFFFAA954AA5D00020AA007BFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000007FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(23),        -- Port A data input
DOA(0)   => data_read_a_lo(23),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(23),        -- Port B data input
DOB(0)   => data_read_b_lo(23),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_24_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100600007FFF000080108004000800020000840041000080808",
INIT_02 => X"0000068002CC07400000090C080002000000103FF811F150231000520ABE4404",
INIT_03 => X"210A0600000203F80005DC00000DC3801EA000000745C4010220000000008000",
INIT_04 => X"07C5FF804900026F8780001DF8000000079800000F300002998078068003C080",
INIT_05 => X"C207F0000000007FF0000004380001FE1E1C07C3E00CFFF80000000000000000",
INIT_06 => X"0002648240F20035A0102000BD0000002802C87FC800FCAA035400001B918600",
INIT_07 => X"0000000001FBFFEC4D2B4AD0B8129063B2CC0000100042018408142F16C01848",
INIT_08 => X"008E1F5F80001FF0000000FFDF78000000000EFFE001600000000005FC000000",
INIT_09 => X"E883FE180000000000300000000000DFFD0000002A80D500000671000004A000",
INIT_0A => X"10018C0411020600048620C030020502000200000400920A2198000800404037",
INIT_0B => X"0641060400C00C00304003040030400304003040030400304003040018200182",
INIT_0C => X"000000001000C00000000000000240058000000000000000000000FFDF000404",
INIT_0D => X"E00880104809C1666594584031010FFF56FFC000104000000010440000000000",
INIT_0E => X"E0088010492064206100E81084200048C0804012500021B00880108012500021",
INIT_0F => X"04100144800803419043064900C0020501840012500021B00880108012500021",
INIT_10 => X"1018140F02C0000809408D206420530270040410004C840041A0D80054109038",
INIT_11 => X"110002C9E8010C00010480B35A0300400041020902F60002260D65B361BAA104",
INIT_12 => X"0228204300166B4060080008240593D0021800020818B06D9802F00030C02060",
INIT_13 => X"143B62023C00142800B04400095DFF90203020042108603100061516EE800C06",
INIT_14 => X"DC1180C7804400044029208301040214AE4C7C02000040206602C10B48110006",
INIT_15 => X"00000000000000000000000000000000000000000000000000000000FBFFE000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"DD5EDCF9822659B6888332000000000000000000000000000000000000000000",
INIT_19 => X"F3CF3CF3CF3CF3DF7DF7DF7DF7DF7DF3DF3DF3DF3DF4D30C2432AEBAEBFE5A15",
INIT_1A => X"C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783DF7DF7DF7C",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000F0783C1E0F0783C1E0F0783",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201008000000000000000000000000",
INIT_1F => X"4BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974BA5D0400000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"00010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000007FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAE974BA5D0000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_23 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0002000087FFFFFFFFFFFFFFFFFF",
INIT_24 => X"FAE974BA550002000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D000200000",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010080000000",
INIT_27 => X"FFFFFFFFFFFFFAE974BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000087FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAE974BA5D0400010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0000010007FFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"E974BA550002000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0000010007F",
INIT_2C => X"FFFFFFFFFFFFFFFFFFAE974BA550002000007FFFFFFFFFFFFFFFFFFFFFFFFFFA",
INIT_2D => X"D0402010080000000000000000000000000000000000000000000007FFFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAE974BA5D0400000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040200",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000087FFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"74BA5D0000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0000010087FFF",
INIT_33 => X"FFFFFFFFFFFFFFFFAE974BA550000010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE9",
INIT_34 => X"000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA550002010087FFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(24),        -- Port A data input
DOA(0)   => data_read_a_lo(24),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(24),        -- Port B data input
DOB(0)   => data_read_b_lo(24),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_25_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100200002000000080100004000000020000800041000080808",
INIT_02 => X"0000068002CC474000000800000002000000103FFCE302008000000880844A04",
INIT_03 => X"00000040700803FC0105DE00020DC3801EA00000040000000020000000008000",
INIT_04 => X"47C5FFC04904026F8780081DFC040000079C92484F30499299837C168003E400",
INIT_05 => X"C207F0382004407FF0000004382281FF1E1C07C3E00CFFFC090004B05000200A",
INIT_06 => X"1009015C4000000020000000390C10002802C87FC800F8000000000019810600",
INIT_07 => X"0501000001FBFFFD480A0280A816002010800001000054018408102000000002",
INIT_08 => X"0C8E1F5FA21C9FF8004000FFDF7C062031863EFFF75D78004001010DFC000020",
INIT_09 => X"E883FE180C00000000300000000000DFFF00180800000000000660100000A000",
INIT_0A => X"1001DCCC31222730A49620C030020100000200000400921A21D8000804404037",
INIT_0B => X"0641062400C00C00304003040030400304003040030400304003040018200182",
INIT_0C => X"C11160845004D04820000000000000000000000000000000940000FFDF000404",
INIT_0D => X"000800000801C0786184185031810FFF56FFC02812E0182000F2C48304418220",
INIT_0E => X"0008000000002020000008000000000800800002400001000800000002400001",
INIT_0F => X"0000010000000000900000080000000400000002400001000800000002400001",
INIT_10 => X"1000000002002000004000002020000200000000000404000000880000001000",
INIT_11 => X"010000082000000001000001080000000040000100C600800001040000040009",
INIT_12 => X"0000000100002100000000080000104000000002000000081001000000000040",
INIT_13 => X"0010200000000000001004000001080000400080000040010000001080001008",
INIT_14 => X"8C11808200400000400000C20000000420000000030280000000010000010000",
INIT_15 => X"82208822088220882208822088A20C52082081A30080000002005008FBFFF001",
INIT_16 => X"2208822088220882208822088220882208822088220882208822088220882208",
INIT_17 => X"2088220882208822088220882208822088220882208822088220882208822088",
INIT_18 => X"29432D518B45265D82BB4101000005FFFFFFFFFFFFFFFFF82208822088220882",
INIT_19 => X"24924924924924820820820820820820924820924824000A6242B4D34D7F7451",
INIT_1A => X"AC562B158AC562B158AC562B158AC562B1188C46231188C46231189249249249",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000162B158AC562B158AC562B158",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000000000000000000000000",
INIT_1F => X"4BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"02000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAE974BA5D0402000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_23 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000007FFFFFFFFFFFFFFFFFF",
INIT_24 => X"FAE974BA5D0400000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040000008",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010000000000",
INIT_27 => X"FFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAE974BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000007FFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"E974BA5D0400000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000087F",
INIT_2C => X"FFFFFFFFFFFFFFFFFFAE974BA5D0400000007FFFFFFFFFFFFFFFFFFFFFFFFFFA",
INIT_2D => X"D0402010000000000000000000000000000000000000000000000007FFFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"74BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000007FFF",
INIT_33 => X"FFFFFFFFFFFFFFFFAE974BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE9",
INIT_34 => X"000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000007FFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000007FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(25),        -- Port A data input
DOA(0)   => data_read_a_lo(25),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(25),        -- Port B data input
DOB(0)   => data_read_b_lo(25),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_26_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"E9264EAB20190CA3BA4997AA9002AE9C001006B0778015CFA17E0811039879C7",
INIT_01 => X"F1FFF9BB1F773C7F9BB07DFFFDD863FC5FFF3FEFFBBF9FFB22FFFBC7B9F30686",
INIT_02 => X"9B3184F8AFDEAF300029E4E300FC78A6258548EFFA71C00172082400003A2161",
INIT_03 => X"0084F0FF7FFF1FDD3FEFDCDE981DC3FF5F0D294A7B2B18A0001B9CE6CC606E73",
INIT_04 => X"0FC5DFD7EDFFD66F87FE605DDDBFF3690F9EDB7F5F7AFF639BD7DE37C2FEF591",
INIT_05 => X"F205F0F8E9D199FF76DFEE1C3FCC3FF7BE1FD7C3FFACFBFFDFF7B4FEFFDAA10E",
INIT_06 => X"042648C40179912406C1830639AFBEC14489737FDC00B13BB79DFDB83BF4112A",
INIT_07 => X"763A844769FFBFE4398E4390BB9C28B1D0F049080414583F9468D1AEFC000060",
INIT_08 => X"02C05FD7BC471FBD13D981F7DF7D7E6171AF3FEFE8A3E679FAC1FD1FFFBEB000",
INIT_09 => X"F8CFFE38FF7F6BD928F1ABB47476B5FEF9F59F5FCEEDE73FEE0EFC53B079F5CC",
INIT_0A => X"315BDDCC3B336F7C548667D47B7737AF3FD62601EDC2B66A67B9D60FE4C4427F",
INIT_0B => X"06E19F4DA0E80E903DE3035E3035E3035E3035E3035E3035E3035E981AF181AE",
INIT_0C => X"EBFBF7FEBD66DBFCA3F87501AE7B080607307DCFE1D4077B4D026FFFFBFFAFCD",
INIT_0D => X"0007E010084BCD7FF1B61B5C33813FFFFCFFC7D7D51D6F5FDCB935D7AFEBD7F5",
INIT_0E => X"0007E01001BD8020500008001F010040520201F45EC0010007E01001F45EC001",
INIT_0F => X"1DC0004600400F781429C0080000770001A001F45EC0010007E01001F45EC001",
INIT_10 => X"10003C064000E408010081BD8020600200001EC00040B02007EC09A0E0001000",
INIT_11 => X"360403E434588007200D00F88C84C081C203404B3BFD0402346235408402C080",
INIT_12 => X"07B00040091F1190982038406807C868B1000E401A08FE0012040000FC002001",
INIT_13 => X"7D00212000007C400082D81009FC08281D00001F010021560406758091454000",
INIT_14 => X"FFBFF5FA1040076065F730FC08043A903A80008320C0403C3400008860160406",
INIT_15 => X"D7F5FD7F5FD7F5FD7F5FD7F5FDFF7F7F7F77F9F761FFBFDFFDE5BFFFFF7FF005",
INIT_16 => X"7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5F",
INIT_17 => X"F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD",
INIT_18 => X"B79E923C2CD990AA7F0DDB6B910C8DFFFFFFFFFFFFFFFFFD7F5FD7F5FD7F5FD7",
INIT_19 => X"30C30C30C30C30C30C30C30C30C30C30D34D34C30C35F7AA9ABF0E38E3A8EB62",
INIT_1A => X"C26130984C26130984C26130984C26130984C26130984C26130984C30C30C30C",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000130984C26130984C26130984",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000000000000000000000000",
INIT_1F => X"4BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"02010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_23 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFF",
INIT_24 => X"FAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010000000000",
INIT_27 => X"FFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"E974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007F",
INIT_2C => X"FFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFA",
INIT_2D => X"D0402010000000000000000000000000000000000000000000000007FFFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"74BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFF",
INIT_33 => X"FFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE9",
INIT_34 => X"000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(26),        -- Port A data input
DOA(0)   => data_read_a_lo(26),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(26),        -- Port B data input
DOB(0)   => data_read_b_lo(26),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_27_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"00080A40000A41248002029000050A088000008242A0004404480002000A1155",
INIT_01 => X"F1FFF1C11F781C129C107DFFFE0860941E81258CA2B71C2220EC1B86E1A00002",
INIT_02 => X"183080988B2EAE00002BE001117C78C6848140CFFA0000800042008000011081",
INIT_03 => X"000000FF7CF91F1D3DEF3CDA881D23FB5C0C21085B0B0820001318C60C204C63",
INIT_04 => X"8FC51FD7EDFDD66E47EE205D1DB7F1490E5EDB7D5CBADB2385D79C3643D4E580",
INIT_05 => X"E001F0C0C991BBFC76DFEA1A3F8C3BC7391F9723FF2CE3FCD6D13096B79C8106",
INIT_06 => X"40000001000000084041830600A40C415004637FC4003021259CFDB01BF80028",
INIT_07 => X"3158954761FA3FE402088220AC1108001080400A400041018468D1A060000050",
INIT_08 => X"02005F0784411E390A4881C7BEFC5F6171CE2F8FE823E778DAC16C1FFBBC9000",
INIT_09 => X"F0C7FEBABF3F6BD108F40E04C0C084F0F8B58B5B8849673F6C0E7A01B00914C4",
INIT_0A => X"B51BFDCC39732F3554866AD57C37BEAF1C152201A4C0B6EA63AAD60B60D4427F",
INIT_0B => X"06F18FC5A0E00F0038D1030D1030D1030D1030D1030D1030D1030F0818688186",
INIT_0C => X"AB6AD7EAB962CBD8A3A83101F47E08040510768EA0C406630D0226FFE375ADE5",
INIT_0D => X"000760000843C561E5C55C42B9011FFF48FFCC57550D63564D1D2556ADAB56D5",
INIT_0E => X"0007600004BD8020100008001F010000130201E44A40010007600005E44A4001",
INIT_0F => X"1DC0000208400D781020C00800007700002005E44A40010007600005E44A4001",
INIT_10 => X"10003C064000C400018080BD8020200200001EC00000382006EC0820A0001000",
INIT_11 => X"3E0403A424108007200102E888808081C20040431BC504021462354004004080",
INIT_12 => X"07B00000015D1110102038400817484821000E400204FE0010040000FC000000",
INIT_13 => X"7D00202000007C400000F81001FC08080500001F0100005E0404758081014000",
INIT_14 => X"8DBBB5FA10400360649310FC08003A903A8000012040403C34000080201E0404",
INIT_15 => X"56D5B56D5B56D5B56D5B56D5B56D7E3D7B57B1C4E17F0944B8D596EEFC7FF001",
INIT_16 => X"6D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B",
INIT_17 => X"D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B5",
INIT_18 => X"2D0200903950C080420948E2D10E8FFFFFFFFFFFFFFFFFF56D5B56D5B56D5B56",
INIT_19 => X"00000000000000000000000000000104000000000004000E5E420000002921C4",
INIT_1A => X"28140A05028140A05028140A05028140A0100804020100804020100000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000140A05028140A05028140A050",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000000000000000000000000",
INIT_1F => X"4BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_23 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFF",
INIT_24 => X"FAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201008",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010000000000",
INIT_27 => X"FFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"E974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087F",
INIT_2C => X"FFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFA",
INIT_2D => X"D0402010000000000000000000000000000000000000000000000007FFFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"74BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFF",
INIT_33 => X"FFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE9",
INIT_34 => X"000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000007FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(27),        -- Port A data input
DOA(0)   => data_read_a_lo(27),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(27),        -- Port B data input
DOB(0)   => data_read_b_lo(27),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_28_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"02200AA400180030808802A900002A08001280A08A801044104A1000001818C3",
INIT_01 => X"50A00011460214428114180000882214413D0A71592A01D92213D28005210202",
INIT_02 => X"8A54800A210200111100C2110054289220810440030404010844000444410001",
INIT_03 => X"1080010208B51400007800000A000001000108C21008092000018C6295200631",
INIT_04 => X"0008000000017000000028000001610300000010000802202040012040040011",
INIT_05 => X"2000044440048880026A22000026A20000000000000000004994140203000064",
INIT_06 => X"1400922401041008004891224228810080010200040001020800000004000008",
INIT_07 => X"150B001328000001404010040084088404200020455514000224489028492201",
INIT_08 => X"00414000201800004080A0000002480B04008100011000088800081002C19020",
INIT_09 => X"000400001036584108415B4A6A694A0000100101C08200000001000190200044",
INIT_0A => X"004800210C19808400500010009110091500020B408820000200400040811600",
INIT_0B => X"40000800B00100040D8140581405814058140581405814058140580A02C0A02C",
INIT_0C => X"00200248010201008298150006210802043058C46054032981002D00201C8081",
INIT_0D => X"0000A00000400600841041108280300008000140000401028008330000800040",
INIT_0E => X"0000A000000080001000000000000000500000040A40000000A00000040A4000",
INIT_0F => X"00000006000000080020C00000000000012000040A40000000A00000040A4000",
INIT_10 => X"00000000000024000000000080002000000000000000A00000040020A0000000",
INIT_11 => X"2200000404108000000900008080808000024040152000000020000004004080",
INIT_12 => X"0000000009001010102000004800080821000000120002000004000000000001",
INIT_13 => X"2000002000000000000288000020000805000000000001420000200001014000",
INIT_14 => X"408010000000022000D610280000080000000001204000000000000820020000",
INIT_15 => X"00401004010040100401004010042024210218734CD52150A840827504000000",
INIT_16 => X"0401004010040100401004010040100401004010040100401004010040100401",
INIT_17 => X"4010040100401004010040100401004010040100401004010040100401004010",
INIT_18 => X"05822140048D2E57B1348141845C200000000000000000000401004010040100",
INIT_19 => X"04104104104104104104104104104104104104104101A6A0A0EB1861863BC422",
INIT_1A => X"2C160B0582C160B0582C160B0582C160B0180C06030180C06030181041041041",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000160B0582C160B0582C160B058",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000000000000000000000000",
INIT_1F => X"4BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_23 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFF",
INIT_24 => X"FAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010000000000",
INIT_27 => X"FFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"E974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007F",
INIT_2C => X"FFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFA",
INIT_2D => X"D0402010000000000000000000000000000000000000000000000007FFFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"74BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFF",
INIT_33 => X"FFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE9",
INIT_34 => X"000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000007FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(28),        -- Port A data input
DOA(0)   => data_read_a_lo(28),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(28),        -- Port B data input
DOB(0)   => data_read_b_lo(28),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_29_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"79964E4BA01DACAB9E659792D00AAE160002829C7FDFEFCEE97C2815039D70C3",
INIT_01 => X"50BFF9AB0775343F9AB01DF80D5821FC0FFF3FEFD1AF9FF1207FFBC7B9720586",
INIT_02 => X"0D15846807D207200021C4E200D428A2018408600271C000720A0000003A2161",
INIT_03 => X"0000B0027BBF17C43E6DC05E1A0DC07D1F0000803B2819A00019084345606421",
INIT_04 => X"07CDC047A4FB526F807C681DC4B97369078249370F482E62BA414627C2FE3000",
INIT_05 => X"F204007861C088FF0EFF260407C427F19E03C7C01F8CF80749B390EA4BCA202C",
INIT_06 => X"000248C00079800406C081023B233E804488527FDC008019968D74982C94110A",
INIT_07 => X"5229000221FF8000398641903B082831D05000200000083F942850AEB4000221",
INIT_08 => X"00805FD0180E1F8C1111A0F041056A0100A11FE000916249A800B915FE82B020",
INIT_09 => X"F80C000055FF7C492840AAB45456B55E015015058665A31DA603A4539058F54C",
INIT_0A => X"000850400A11414C005005000B51158936D20601A98A204006114005C4800217",
INIT_0B => X"40201948B029029409A3401A3401A3401A3401A3401A3401A3401A9A00D1A00C",
INIT_0C => X"40B1225C1506512C83E85500AC3A080406305587A154023141006DFFF89E82C9",
INIT_0D => X"0000A01008480D3EB4A24A0C910037FFFC0007C7C0140D0B50A8218102C08160",
INIT_0E => X"0000A010010080005000000000000040520000141EC0000000A01000141EC000",
INIT_0F => X"00000046000002080429C0000000000001A000141EC0000000A01000141EC000",
INIT_10 => X"00000000000024080100010080006000000000000040B000010401A0E0000000",
INIT_11 => X"3600004414588000000D00108484C080000340483B590000202000008402C080",
INIT_12 => X"00000040090210909820000068008828B10000001A0802000204000000002001",
INIT_13 => X"20000120000000000082D800082000281D000000000021560002200011454000",
INIT_14 => X"B29450580000066021F6303C000408000000008320C000000000000860160002",
INIT_15 => X"816058160581605816058160589625662522506344FF9FCFFF62EB6DFF001004",
INIT_16 => X"1605816058160581605816058160581605816058160581605816058160581605",
INIT_17 => X"6058160581605816058160581605816058160581605816058160581605816058",
INIT_18 => X"F2DDCFFFBEFFCF07FFBFFD41800C05FFFFFFFFFFFFFFFFF81605816058160581",
INIT_19 => X"7DF7DF7DF7DF7DF7DF7DF7DF7DF7DD75D75D75D75D77FFBF3F7DFFFFFFD779F3",
INIT_1A => X"FEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDF7DF7DF7DF",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00001F7FBFDFEFF7FBFDFEFF7FBFD",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000000000000000000000000",
INIT_1F => X"4BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_23 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFF",
INIT_24 => X"FAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010000000000",
INIT_27 => X"FFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"E974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007F",
INIT_2C => X"FFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFA",
INIT_2D => X"D0402010000000000000000000000000000000000000000000000007FFFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"74BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFF",
INIT_33 => X"FFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE9",
INIT_34 => X"000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(29),        -- Port A data input
DOA(0)   => data_read_a_lo(29),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(29),        -- Port B data input
DOB(0)   => data_read_b_lo(29),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_30_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"FFDFF3FC3EFFF7FFFFBFFA000000000000000000000000000000000000000000",
INIT_19 => X"F3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF5F7AEBEBFBEFBEFFEFFF7",
INIT_1A => X"CFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCF3CF3CF3C",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000007F3F9FCFE7F3F9FCFE7F3F9F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000000000000000000000000",
INIT_1F => X"4BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_23 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFF",
INIT_24 => X"FAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010000000000",
INIT_27 => X"FFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"E974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007F",
INIT_2C => X"FFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFA",
INIT_2D => X"D0402010000000000000000000000000000000000000000000000007FFFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"74BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFF",
INIT_33 => X"FFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE9",
INIT_34 => X"000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(30),        -- Port A data input
DOA(0)   => data_read_a_lo(30),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(30),        -- Port B data input
DOB(0)   => data_read_b_lo(30),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_31_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"129000008004A00804A40000400800020000000C005FEA005800200400050100",
INIT_01 => X"A15FF18019700810180065FFFC0040801E80258CA2951C2200EC0906A0804140",
INIT_02 => X"146000808A0C060444692000402850040400408FF80000000010000000004000",
INIT_03 => X"000000FD74480B1C3D951C5A800D03FA1C0C21084B0300000012108518004842",
INIT_04 => X"07C51FC7EDFCA26E07EE001D1CB6904A061EDB6D4C30490281831C1602D0E480",
INIT_05 => X"C001F0808181117C7C95C8183FA099C7181F8703FF0CE3FC0201209010988002",
INIT_06 => X"00000000000000010001020400840C41C000617FC0003021259CFDB01BF00020",
INIT_07 => X"0000000441FA3FE400080200A810000010804008100040018448912040000040",
INIT_08 => X"00011F0780011E38004801C79E7C162231862E8FE00166704041240DF93D0000",
INIT_09 => X"F0C3FE180D89279000B00000000000D0F80088080849673F6C0E780020091480",
INIT_0A => X"1011DCCC31222730048620C4382204A608142002A440924A6188020920404437",
INIT_0B => X"0661874500E00E00304003040030400304003040030400304003060018200182",
INIT_0C => X"810040801060C04821202001A05A00040100240A80800442040202FFC3200444",
INIT_0D => X"000740000803C0616184184031010FFF40FFC407500020004C10060204010200",
INIT_0E => X"0007400000BD0020000008001F010000020201E04000010007400001E0400001",
INIT_0F => X"1DC0000000400D701000000800007700000001E04000010007400001E0400001",
INIT_10 => X"10003C064000C000010080BD0020000200001EC00000102006E8080000001000",
INIT_11 => X"140403A020000007200000E808000001C200000308C504021442354000000000",
INIT_12 => X"07B00000001D0100000038400007404000000E400000FC0010000000FC000000",
INIT_13 => X"5D00200000007C400000501001DC08000000001F010000140404558080000000",
INIT_14 => X"8C1380DA10400140640100D4080032903A8000000000403C3400008000140404",
INIT_15 => X"02008020080200802008020080200C1808008184012A08041202500AF87FF001",
INIT_16 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_17 => X"0080200802008020080200802008020080200802008020080200802008020080",
INIT_18 => X"000000000000000000000002001005FFFFFFFFFFFFFFFFF02008020080200802",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000000000000000000000000",
INIT_1F => X"4BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_23 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFF",
INIT_24 => X"FAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010000000000",
INIT_27 => X"FFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"E974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007F",
INIT_2C => X"FFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFA",
INIT_2D => X"D0402010000000000000000000000000000000000000000000000007FFFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"74BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFF",
INIT_33 => X"FFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE9",
INIT_34 => X"000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(31),        -- Port A data input
DOA(0)   => data_read_a_lo(31),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(31),        -- Port B data input
DOB(0)   => data_read_b_lo(31),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_0_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"ED39BA795990D275FB4A6E96ACC4731DEA4598B0AFB54867F6EE4618C3749807",
INIT_01 => X"58A0047D8607944AC7DA180001ECA2444042106208408208C20022E9173734B3",
INIT_02 => X"8B1E49562021F8051500147A0E162923024F28000415F5787B09FBF999BB1EFC",
INIT_03 => X"1013BF028A959403C06A23A147723C01E140088280C4CF6996088862C7922221",
INIT_04 => X"781A003802015D9078011DE20340699198600000B08694916434804825241311",
INIT_05 => X"2CA000587E10C880036A3103C00F2000E1E0383C00730002B4409845E4425171",
INIT_06 => X"179B48CFF95DCF9EF730E1C3BB731138AF7B888025340C0888430047040FEE18",
INIT_07 => X"AF155113160400185F87C1F05707D415E664A6E7C5551EBE783060CEB164833F",
INIT_08 => X"4D7E40002B7AE005FDB47600208229010C6101001EFE198C96B0528202C0DCB4",
INIT_09 => X"062400608234D864444081048A80CC00062D42D30222108091C107A1DA040267",
INIT_0A => X"204A21008E514844EB5145000255DA599581D3A9583C24351240B58298011308",
INIT_0B => X"E08C4830F81380CE0F89E07A9E0789E07A9E0789E07A9E0789E070CF0184F038",
INIT_0C => X"3A4E9D63EA180EB150CA1CA45C254D4AF4AA414568729139F2A12C0000016110",
INIT_0D => X"F0009E0FC048211E9C11C31F82E4A000890022B827EB52F52347F174E93A749D",
INIT_0E => X"F0009E0FCC42EFDFBF0AE03080E2AEB2E0F1F80FA97FE0F0009E0FC40FA97FE0",
INIT_0F => X"0231F0BD9E3FC08FEBD6F661C0E008C3CB5F040FAB3FE0F0009E0FC40FAB3FE0",
INIT_10 => X"20180309A0F83BE2B87C7C42EFDFBF187806013879BA878FE807F65FBF12E038",
INIT_11 => X"0BE9F01FC8B38C2098DAE007F323A0C83136B248831ACBFC8BBDCAB779BC699F",
INIT_12 => X"004C72BEC800FE7464290626D7003F9947184131B59003FFEC07F00003F01FB9",
INIT_13 => X"A0FFDA2A3C0202B8776A2FA7F023F7D065703080E29F1B2BE9F8A27E6E915C0E",
INIT_14 => X"016C2D25E52630BB1AE49C2BA7F98D6F846DFC0C2352A0024B83F07F198BE9F8",
INIT_15 => X"749D2749D2749D2749D2749D2749F285F25D2C500815A5522CB5A4B400000CD4",
INIT_16 => X"49D2749D2749D2749D2749D2749D2749D2749D2749D2749D2749D2749D2749D2",
INIT_17 => X"9D2749D2749D2749D2749D2749D2749D2749D2749D2749D2749D2749D2749D27",
INIT_18 => X"31C136AD8E9B562BA39E2600654BA800000000000000000749D2749D2749D274",
INIT_19 => X"4104104104104104104104104104104104104104104104109C83B8E38E2ABE71",
INIT_1A => X"0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0410410410",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000007C3E1F0F87C3E1F0F87C3E1F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000187FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"BAF7FFD55EF007FD75EFFFAE97555557BD75EF5D000000000000000000000000",
INIT_1F => X"000AA843FE00AAFBE8B45AA803DFEFA28428B455D0017410A28428AAAA2FBD54",
INIT_20 => X"FEBAA2D5401450051401555D7FC0145F7AEBFFFF08002AA10A2AABFEAAA2FFC0",
INIT_21 => X"D755555517FFEFA280021FF082E974AA5D7BFFE000804000BAAAAAAAB45557FF",
INIT_22 => X"EA8B45005168A10AA8028A10087FD7410557FC21555D51574AAA2FFE8B455D7B",
INIT_23 => X"AE95410AA80000005D003FEAAFFAEBFE00A2803FEBA002A820AA0800174BA5D2",
INIT_24 => X"2AEA8A10000417410A2FFE8BEFF7FFE8B45FFFBC00005D003FF45557FC01FFFF",
INIT_25 => X"00000000000000000000000000000000000000557DF5500003DFEFFF84175EFA",
INIT_26 => X"5F524AFE38B780154BAFFF1D54AF0075D75EFEBAE9554540754717F1F8000000",
INIT_27 => X"50B6AABDE12BEA0AF010B7D1F8F47E00A2DB45AA8A3AFD7B68E2AB78550E1255",
INIT_28 => X"E9257F1E816D557095EAAA2D1401D500002A150038038E285D7F78FD7000B6AB",
INIT_29 => X"5A87AAD178A8002D1D21C5E8257D5C7AA854008700249243A412EBFF5542A43F",
INIT_2A => X"52A82000E3A5D2150AB8F401471EDBC0B680900AAF52B474385D75C502D15754",
INIT_2B => X"FD7E9541242FE920AD082E10A28F6A150012A2F02AFFDF40E85F475451D502D1",
INIT_2C => X"0550E87B7A405B52AAD152BD00151EAFEDB52E3F1EFFFF485A2DA3D5D24BD417",
INIT_2D => X"57F40545850000000000000000000000000000000000000000000005AAF55508",
INIT_2E => X"F7AEAABFF5D2A81151FB8635A02FA69574BAF7D5555AF0D79D55FFA2AC974450",
INIT_2F => X"8D46F6ABE7082AAAAF2FAC77FE00FF16565B2FA9075F4F7B3EBDF50FEAEAAB55",
INIT_30 => X"56803CE3AEB038662E5D81406014D5D51F5E08A394003A908B8410E707EF34A0",
INIT_31 => X"4AF0151555AF58794040077D774FAE8C798A11A0EAEF75F7AA84001A7052C952",
INIT_32 => X"4E1870108B11020AD4AA05542A0A05051023F9A9D57B63BFBF906CB45FABC095",
INIT_33 => X"F5F0DA6BC9525688C1A2A0C06E9FEE5555BE48AB2A2AE0A0F20C43EAC562245B",
INIT_34 => X"000000FF80F55E25C00A0BA7FBED407A97F6F35F498B96BEB12DAAB77558ABD5",
INIT_35 => X"8000000FF8000000FF8000000FF8000000FF8000000FF8000000FF8000000FF8",
INIT_36 => X"00000000000000000000000000FF8000000FF8000000FF8000000FF8000000FF",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000008000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(0),        -- Port A data input
DOA(0)   => data_read_a_hi(0),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(0),        -- Port B data input
DOB(0)   => data_read_b_hi(0),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_1_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"212C001411984004084D000508C53810A03D1450E839B003342114428A000803",
INIT_01 => X"08000010400A0008010600000084005000400002000000000000000000140000",
INIT_02 => X"C084484000002014400205851002007030450E0000A606C8C44CB4C6666C00E0",
INIT_03 => X"CCF7CE0002058001000000800240200001018CA1800001091408463061120118",
INIT_04 => X"082800100000000040000900010000100040000000008411600401C02100000C",
INIT_05 => X"10800202080422000020012200000000810000200000000004020C00200011A0",
INIT_06 => X"56BDBFBC48C315A8660C18305750C008940D8000011000820001000104050004",
INIT_07 => X"8B4344400004000150248912154404C6060A2FE24555013E13060C158AC97F01",
INIT_08 => X"00082080087A000559102400200281000469000008B000000090108000400430",
INIT_09 => X"0000000000001004140545402820020000010010208000008041060008200001",
INIT_0A => X"2102210182004840007845004044020000200080080844200000048088000000",
INIT_0B => X"48800000190191064620646A06468064680646A0646A06468064690321503234",
INIT_0C => X"02008100200800A1100707040101E20BE0B002605C1C110848200C0000000800",
INIT_0D => X"F000A000C0000012187087010AE4B00000000810010040108104100408020401",
INIT_0E => X"F000A000CC4200002F08E03080000010F18058000003C0F000A000C4000003C0",
INIT_0F => X"000000078808C00000023461C0E00000012704000003C0F000A000C4000003C0",
INIT_10 => X"201803000000240218C0044200001E1878060000000AAC00680000001F10E038",
INIT_11 => X"2100B00048230C200009A0001303204800025200040A00D000000202090C281F",
INIT_12 => X"00000002C9000260640900004D0000904618400012900001EC03F00000000039",
INIT_13 => X"80025A0A3C020000002A8400B00007806070308000000961002880204A901C0E",
INIT_14 => X"000801046004308A185000020128000904285C0C0312A0020000000838810028",
INIT_15 => X"0401004010040100401004010040100010410C002000040280100000000008D0",
INIT_16 => X"4010040100401004010040100401004010040100401004010040100401004010",
INIT_17 => X"0100401004010040100401004010040100401004010040100401004010040100",
INIT_18 => X"48D757DF8A9410218E8A56085142020000000000000000004010040100401004",
INIT_19 => X"555555555555555555555555555554514514514514550431A581924924B02651",
INIT_1A => X"4BA5D2E974BA5D2E974BA5D2E974BA5D2EB75BADD6EB75BADD6EB75555555555",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800005D2E974BA5D2E974BA5D2E97",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000607FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"10AAAABFFFFFF803FE10F7D17FEBA55556AAAAAA800000000000000000000000",
INIT_1F => X"EBAFFD555400557BD54BA5D7FFDF45A2FBD75EFA2AE97555F7FBFFF45FFAE800",
INIT_20 => X"ABEFA2D568A005D5157400AA8028AAAF7FBD54AA002A955555D7FE8ABA082EBF",
INIT_21 => X"FDF55AAFBC0010555540010550417555AA8028BEFAAAE97555082A80000AA802",
INIT_22 => X"BD7410550428ABA5D5168ABA552EBDFEF5D7FEAA00AAAABFEAA007BC0145FFFF",
INIT_23 => X"FFEAB55557FFFEBAAAD568B45A2D5575555D7FC2155F7AEA8BEFAAAA954BA557",
INIT_24 => X"D7BD74000804154BA082ABFF55FFD57DF45F7D568ABAF7AABFFFF082ABFFFFFF",
INIT_25 => X"000000000000000000000000000000000000002EBFFEFA280021FF082E974AA5",
INIT_26 => X"5E175EFF57BF8FC2000BEA4BAE97F78A3FE28E3D17DEAA485FE8E02B50000000",
INIT_27 => X"455571E8A2A087BF8EAAEB8E0016D5D75D54BA5D7BFFF7DA2FFD55EFAAA49554",
INIT_28 => X"157428145A00AA8A2FBD7B6DF6AA28550E10405F7A4AFE38EAA0924921C2FD55",
INIT_29 => X"8E971471C7010B7D168F47400A07A28415A001684104155C5B6DF6DBEFBFAA07",
INIT_2A => X"BFBD7B6A0BF492415FC20105D24AAABF1FFBC7010FF8A38FEF557FEAB78B6AAB",
INIT_2B => X"017EBA4A8EB8F6FFD5FE8B7D557495EAAA2D16D1FDBED56A55557A43DE385FD4",
INIT_2C => X"854008700249243A417FFF41542F5D717FE2AAAA56DEBD17FE3DF7FB7FEBFE38",
INIT_2D => X"07DFCA127B8000000000000000000000000000000000000000000002A3D5C7AA",
INIT_2E => X"AAFBD55FFAA8416545A6FB60F47AF2A00010F78028B15F7823FEAAA2D57DFBA0",
INIT_2F => X"22A38C20B2552E975F758516AAAA0869AAAB8A7C19C55550E8574BA557BFFFEF",
INIT_30 => X"55FFEFBCEE5FBAACB10085EE5DE10A2AEBFF55F7BAAA8565DBAC1112FFAC21A0",
INIT_31 => X"BEA097BEAAFAF2863FA00DD574201E7AD1FFF5575841DE08007FC20480028957",
INIT_32 => X"54FF57EFBFA18D4FBFFF40FF809D4000D7FC00FC5D062BBA05ED5034472A02EA",
INIT_33 => X"7DFBFF6963FCAAA2283CF14050062B0A2F7AE8B5D5D51F5E18ABD5EAFFF2AF95",
INIT_34 => X"000000002CB75F7AA84001A7052C95256807DC31AA8114DE55F5BED201FFFED1",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000008000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(1),        -- Port A data input
DOA(0)   => data_read_a_hi(1),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(1),        -- Port B data input
DOB(0)   => data_read_b_hi(1),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_2_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10E44660018259B2843913100062C98004802322D3E030235201006009B2813",
INIT_01 => X"000AC188084900481C8024A542400340404000720885800802000906E4910204",
INIT_02 => X"82040072AC248C31010204880000007401044C0550200000480E0080001300E0",
INIT_03 => X"0080812C130D0A0D1193088802182142494D218220021100001A8020C1004A00",
INIT_04 => X"090D0AD62824A44A428408540D1610020C6E510818923441A4908B0503404201",
INIT_05 => X"5000A004081122242420480A14A99C428908122144244150906124248C002168",
INIT_06 => X"1400088400450000460000001308890094082015800011012D41D518044C1100",
INIT_07 => X"26731111491C1541324C1114BD880004002040204050413F1400100480000201",
INIT_08 => X"02410582881E0C1511D02082AAAB016A2463288549B044605201D10AE11B0020",
INIT_09 => X"E80394280E40158020B591000800481051241A4A404B5035C60904502054E000",
INIT_0A => X"0102C9E12202EA6014D027C418428E220A5500024808922801A0900A84454458",
INIT_0B => X"4600070110C10D04340043400434A043420434A04342043480434102184021A0",
INIT_0C => X"E9CA34328E44CA1401306100A246000402100C088104010AC8005C5681812B04",
INIT_0D => X"0000A0000801487334E34C1A980001550055481204090A4C01351253A728D194",
INIT_0E => X"0000A000013800004000080000000000500000B01480010000A0000150148001",
INIT_0F => X"0000000608000A500409000800000000012001501480010000A00000B0148001",
INIT_10 => X"1000000000002400000001A100004002000000000000A0000360018040001000",
INIT_11 => X"380001C01048000000090298040440000002400008C400022042004080028000",
INIT_12 => X"0000000009530080880000004813802090000000120C94000200000000000001",
INIT_13 => X"4C000100000000000002E0000950002018000000000001580002508010440000",
INIT_14 => X"7120642000000400015020500004221018000082008000000000000820180002",
INIT_15 => X"5094A5294A5294A52942509425094209461468000822241A03835D88482AB001",
INIT_16 => X"09465094A5294A5294A5294250942509425094A5294A5294A529425094250942",
INIT_17 => X"94650946509465294E5294E5294E5094650946509465294E5294E5294E509465",
INIT_18 => X"080271AE180616A38A18FA204452A7F03F03F07E07E07E05294E5294E5294E50",
INIT_19 => X"20820820820820820820820820820820820820820820490C04102CB2CB2EB2C0",
INIT_1A => X"8944A25128944A25128944A25128944A25128944A25128944A25128208208208",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF1F804A25128944A25128944A2512",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000787FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"AAAA843DFFFAAD1554005D7FD74AA00040015500000000000000000000000000",
INIT_1F => X"F45AAAAA8A10A2AE80010A2AA975FF5D003FE10F7D17FEBAF7D5420AA0855420",
INIT_20 => X"FF45A2AA975EFA2FFD7555FFFBFFF45AAFBC20AAF7D1575EF55517DF555D2EBF",
INIT_21 => X"95555552E974105D517DF55AAAAAABEFAAD1575EFAAAE974AA5D51554BA5D7FF",
INIT_22 => X"E82010F7AABFE10FFD542145FFD5554AA555555555557FE8ABA082EBFFFFAAAE",
INIT_23 => X"FBC0010AA802ABEFAAD540000FFD540000AA802AABAF7FFC2010AAAE821EF552",
INIT_24 => X"A8028BEFAAAE821550851420AA002E800AA08042AB45007FC00BAFFD168BEFF7",
INIT_25 => X"000000000000000000000000000000000000002E80010555540010550417555A",
INIT_26 => X"AE95F40002157F470AABE803AE97A2DF55400557FD54AA1D04001C5150000000",
INIT_27 => X"EF55517DFC5552ABDF45B6AEAFFD5F7A482000BEAE905C755003FE28E3D17DEA",
INIT_28 => X"0BA5FD0154BA5D7BFAF7DA2AE955EFAAA495545E3F5EFF57F7FE80082FFDE105",
INIT_29 => X"8AAF082AB8EAAEB8E0016D5D2A924105D5B7FF7DB6AAAABC7BEDB505EFBEA407",
INIT_2A => X"95038AAAEAF1D7410E80000FF8438E00B6DF68FEF4871D24BA495B5556D5571E",
INIT_2B => X"1ED1EFEAF1EFFFDEAD1C5010AA8E2FBD7B6DF47A00EBDB50000A380AAE28E804",
INIT_2C => X"5A001684104155C5B68E2DBEFBFFBC703AE2DF42AAA002A851C214003FF68007",
INIT_2D => X"50002155510000000000000000000000000000000000000000000002087A2841",
INIT_2E => X"55003FEAAAAD57DEBAA2FDDC01051FBD74BAF7802AB05AAFBD5400557BD54AA5",
INIT_2F => X"7AF7FC20B2F7FBC015D58517FF555D2ABDF55F782BEB47AFAD00010F7AA82155",
INIT_30 => X"55FFFFC20FFF3AE544108410174BA557BEABEFAAEBD55FFAA1456547A2D360F4",
INIT_31 => X"0BA547FD75FF58516AAAA0828AAAB4A78016545540400010557BFDFFFF7822A9",
INIT_32 => X"550AAFACAAA122AA8954BAA2AE9D545002A800A8FF862BA00F2F9E8F0050D442",
INIT_33 => X"954505C417FFFF08555555BAAD335B57AB5155400A2AEBFF45FFFB404007FFBD",
INIT_34 => X"00000000061DE08007FC2048002895755FFAEBCFE57BBA57002DF3C4AAAA002E",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000010000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(2),        -- Port A data input
DOA(0)   => data_read_a_hi(2),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(2),        -- Port B data input
DOB(0)   => data_read_b_hi(2),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_3_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"210C44A20020248B08431120001604B8156023104C40771B3430400A02380206",
INIT_01 => X"015A2A4050B009683C0422C992000B61404040028804A0080A000C16A8990A0C",
INIT_02 => X"C0A406500CE0A95011000D1501005274B5041AB330860281CC08008222170060",
INIT_03 => X"AB488054270F08E1289084C8020420E005A48DA16C021100003A46B06900C91A",
INIT_04 => X"848966150DA0A02941A4080C612A104201C689044382FD403C17E491829B259B",
INIT_05 => X"D006620608843116942508120A208D18A5050160C600D4C894600094B49CA068",
INIT_06 => X"12002D9401C70008060408141788E2C094887033080071913209CC8004640100",
INIT_07 => X"221111454874CCC4122C0932155400C2023940284000003E15020525CE805E11",
INIT_08 => X"020103C9984A0AC511102029869D974214EDBA132891000052C1750B48290020",
INIT_09 => X"60808C8A2E41351020004148A289428730A51E5E644C8233A0090E1020208100",
INIT_0A => X"A4000041A600417914506F955D6422000934000A090A94A020229603A414144D",
INIT_0B => X"469100841001000406D04065040650406D0406D04065040670406C8201782032",
INIT_0C => X"6A4AF532A8040AF821042D01F14084030070262810340402C0000CCE4CC12520",
INIT_0D => X"000800000401C333494594532980733302CCC81300094E5C91200257AD2AD795",
INIT_0E => X"00080000051C0000400000000000000800000190148000000800000450148000",
INIT_0F => X"0000010000000B100409000000000004000005101480000008000004F0148000",
INIT_10 => X"0000000002000000000001B00000400000000000000400000168018040000000",
INIT_11 => X"1000034010480000010002D804044000004000812E4400002440014080028000",
INIT_12 => X"0000000100570080880000080015C02090000002000CCC000200000000000040",
INIT_13 => X"1C0001000000000000104000094C002018000000000040100006418010440000",
INIT_14 => X"4128652000004404010E20500004208018800082008000000000010000100006",
INIT_15 => X"5795A5595A5595A5595A5595A5595E1152556D008028341B13924D80C2E67009",
INIT_16 => X"69565795A5595A5595A5595A5595A5595A559525795257952579525795257952",
INIT_17 => X"95256956579525495E5595A5495E5595A5495E5595A569565795256956579525",
INIT_18 => X"7818F18E0C8514298B0C52A0115009AA9556AAD552AAD5556956579525695657",
INIT_19 => X"24924924924924924924924924924820820820820825042C0000249249202A60",
INIT_1A => X"8D46A351A8D46A351A8D46A351A8D46A353A9D4EA753A9D4EA753A9249249249",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF248086A351A8D46A351A8D46A351A",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"EFAAFFD54AAF7D168B45AAAABDF5500002AA1000000000000000000000000000",
INIT_1F => X"F45FFD168AAA0855420AAAA843DFFFAAD1554005D7FD74AAA284001550055421",
INIT_20 => X"55FF5D003FE10F7803FEBAFFD5420AA080400155AAD5554AAF7802AB4500043D",
INIT_21 => X"28B45A2AE82155A2FBFFEBA0800021550855555FFAA84001FFAAAE80010A2AA9",
INIT_22 => X"168ABAFFFBD54BAAAAE97400A2FBC20AAA284175EF55517DF555D2EBFE00AA80",
INIT_23 => X"AA954AA5D7FFFF45AAAA975EF007BD7555FFFBFDF55AAFBD55EF5D2EBFE10085",
INIT_24 => X"AD1575EFAAAE974AA5D00175555D0015410F7AAAAAAA55043DE00FFFFD5555AA",
INIT_25 => X"0000000000000000000000000000000000000004174105D517DF55AAAAAABEFA",
INIT_26 => X"ABC04001C51551471D7AAF1D05D2EBD56DB7DBEAEBFF551C042AA101D0000000",
INIT_27 => X"92EB842FB5508043FF55EBD56ABD75D5B470AABE8A3AFD7A2DF55400557FD54A",
INIT_28 => X"557FD2082000BEAE905C755003FE28E3D17DEAAEBDF40002550F47155AADB504",
INIT_29 => X"DF40552ABDF45B6AEAFFD5F7A48017DAAFFFAE821C0A0717D1C5B575FFB68E82",
INIT_2A => X"C55D7492E90E3808756DA92EBFFD74BAE3AE85480FFFFC00AABE8E105C755517",
INIT_2B => X"43AE10EAF5C5547FF80954AA5D7FFAF7DA2AE905EF0075D5545E3F5EFF57F7D5",
INIT_2C => X"5B7FF7DB6AAAABC7BEDB505EFBEF5C7092FF801756D490A10438EBA4B8E92410",
INIT_2D => X"D0028A00510000000000000000000000000000000000000000000000E124105D",
INIT_2E => X"AAFBD54005D7BD54AAF78002155515157555AAD142040A2D57FFFFFFAEBFF555",
INIT_2F => X"051AE955F7AAFBC0000AF843FF5500003FF55AAFD6AB455157D74BAF7AAA8B45",
INIT_30 => X"FF557BD74EFFBACD41577B8400010F7AA8215555003FEAAAAC53DEB8A2FDDC01",
INIT_31 => X"0BAF7AA8015558517FF555D2ABDF51F782BCB47ABAE801FFAAFBEAA105D2E955",
INIT_32 => X"214FA2D3EAF57AFFDD7555082AA0AAA00557FEA8A2FDD64BAAF8282012AFFEC2",
INIT_33 => X"820AAAB842AA00000028AB0AAFF48547AE04174BA557BEABEFA2AA951FF88554",
INIT_34 => X"000000002A80010557BFDFFFF7822A955FFFFC21FFF3BE40412DE02955FF082A",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000008000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(3),        -- Port A data input
DOA(0)   => data_read_a_hi(3),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(3),        -- Port B data input
DOB(0)   => data_read_b_hi(3),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_4_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"A108400020612C80284210081034849800A000303100048B3432C82904204006",
INIT_01 => X"210668000008004C1C20250E12100368403008418984014902030906A8910200",
INIT_02 => X"120404C0024C0600000206100008402404040C00F104008040080080001310E0",
INIT_03 => X"7728805052470B5C1B873C04121D03845D0020CA0822018000080084C1000002",
INIT_04 => X"0B899E43891686690790485D5C3E02000E9892201D306D03A9835C16029AC186",
INIT_05 => X"C001E080005030767434C0003C8A01D6B81C5703C82CDBC000072400089C8120",
INIT_06 => X"1000088100410000460002041300004084080070D00030032009700024641102",
INIT_07 => X"4261950408CCBC2012048310951000000003402A4000143E1008912480000211",
INIT_08 => X"00811007AC0A1EB5131120C79E7D176251E53E80E8B361604041340838452020",
INIT_09 => X"C08360820C0912800035F1801630A8260900180C00C8021C800FEE522020A108",
INIT_0A => X"8400F88C166262E940D00D410D62AD02091704024D0A02882192020DA0544043",
INIT_0B => X"4011078510C90D143142430C243042430C24304243042430C24305121A612186",
INIT_0C => X"C08060101000C00401008800F004140009400E4002A0010240000DC3C080002C",
INIT_0D => X"000800100001C07261C51C42390240F050C3C000950008088130040100018000",
INIT_0E => X"00080010003510004000000000000048010002E0100000000800100220100000",
INIT_0F => X"0000014008001550000800000000000400800280100000000800100360100000",
INIT_10 => X"00000000020000080080009410004000000000000044080000D8008000000000",
INIT_11 => X"000005800008000001040168000040000041000100EC00004002214000008000",
INIT_12 => X"00000041003C000008000008200D00001000000208050C000200000000002040",
INIT_13 => X"17000100000000000090000002C8000008000000000060000004480000400000",
INIT_14 => X"8400C00208004844C00800000000528008000000008000000000010040000000",
INIT_15 => X"0100800004030080000C010000A00D1804404912802A261B53104810DB1E0028",
INIT_16 => X"000C030000200C01000020040300800004030000000C03000000040100802004",
INIT_17 => X"008020040100C010000200800004010040300800000020040100C03000020000",
INIT_18 => X"40C700FC0A000280C68A08A950520E964C3269B2C9864D30000C030040100800",
INIT_19 => X"555555555555555555555555555554514514514514526991A199A28A28981451",
INIT_1A => X"41A0D068341A0D068341A0D068341A0D06A351A8D46A351A8D46A35555555555",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF771F60D068341A0D068341A0D0683",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FF087FFDF5508003FEBA087FD54BAAA841540055000000000000000000000000",
INIT_1F => X"F5500003DF455555421EFAAFFD54AAF7D168B45AAAABDF55A2802AA1000002AB",
INIT_20 => X"DFFFAAD1554005D7FD74AAAA840015500002AABA082E954005500021FF5D2EBF",
INIT_21 => X"68BEF080028BFF0855555455500174BAA2AABDE0055517FF555555420AAAA843",
INIT_22 => X"168ABA0055574BA5555554BA5D0400155AAD1554AAF7802AB4500043DF45FFD1",
INIT_23 => X"0400010A2AA955FF55003FE10F7803FEBAFFD5420BA085168A00007BFDE10085",
INIT_24 => X"855555FFAA84001FFAAFBEAB45002A97545F7D1555EF55043DF5555517DEAA5D",
INIT_25 => X"000000000000000000000000000000000000002A82155A2FBFFEBA0800021550",
INIT_26 => X"5BC042AA101D0A28BC7007FFDF45080A3AEAA007BD2482BE84124285C0000000",
INIT_27 => X"004100021FF492AB8F7D1C0438E381451471D7AAFBD0492EBD56DB7DBEAEBFF5",
INIT_28 => X"FED1C5F470AABE8A3AFD7A2DF55400557FD54AABE84001C5550A28ABA1424974",
INIT_29 => X"FB5508043FF55EBD56ABD75D0428BEF005557545490012482B6A0BAE2849557A",
INIT_2A => X"6DA101475FDE10145F68A921C55504924955524AA140E0717DAADB50492EB842",
INIT_2B => X"43AF6D405F78E3A1C2002000BEAA905C755003FE28E3803DEAAEBDF40002557F",
INIT_2C => X"FFFAE821C0A0717D1C5B575FFB6DF425575D7BEFB55002097555FFD5401EF5D0",
INIT_2D => X"784000AA59000000000000000000000000000000000000000000000208017DAA",
INIT_2E => X"A2D57FFFFF7AEBFF55FF8028A00512EAAB45007FFFF55082EA8AAA087FC2010F",
INIT_2F => X"5512AAAA085D04174100800021FF002EA8BEF5D0428ABA595557555AAFBC2000",
INIT_30 => X"00FF802ABAA04552ABFF597FD74BAF7AAA8B45AAFBD54005D7BD54AAF7800215",
INIT_31 => X"5FFAAFBC0000AF843FF5500003FF55AAFD6AB4551002ABEF0055555550004020",
INIT_32 => X"DEB0A2FD5600051537DE005D557DE005D7BE8AA85555400100879560AA592F95",
INIT_33 => X"17545FFD5421FF5D0428BEF0079FCABA598400010F7AA8215555003FEAAAA843",
INIT_34 => X"0000000004001FFAAFBEAA105D2E955FF557BD75EFFBBCD415521FBFDF450004",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000010000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(4),        -- Port A data input
DOA(0)   => data_read_a_hi(4),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(4),        -- Port B data input
DOB(0)   => data_read_b_hi(4),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_5_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50DB0A0791B1B41694368283C81F9996A091A32152007AB36B20E03C040C002",
INIT_01 => X"880015C49830884C446A40000C34C24841280A00084000C8C212892EEA953231",
INIT_02 => X"408F417400B1D9100002171C1FA20171124E6AA00D8633F8CD09DBFBBB972F7C",
INIT_03 => X"88538F0182058082D800C3314722DC08A34084A100C4D7C99208521063D00148",
INIT_04 => X"F45E41AFAF420996B8411CA282F80A9091224800A2C61490363080C8A4000308",
INIT_05 => X"0EA416069640420901A01505C4410020C6E228DC30532839B043289D9C005031",
INIT_06 => X"13992D9AF8C74E92B7B568D19708C038AFFA89F0B9348C9204C389672407EF12",
INIT_07 => X"6255000016053C18162589725146F442222CE6AF844012BE795224458BA4DE0F",
INIT_08 => X"4F3F00503B4AE104B5347230418190420821006016FC18843630D285FC416CB4",
INIT_09 => X"EEA33E700340902C4424C442B0344724066C56C2248130A2D9C185B24A24832B",
INIT_0A => X"315325008348CC40AB570500204462508135D5AA593E043731E9B18A98440137",
INIT_0B => X"E0CD463C5813804E0258E0358E02D8E03D8E0258E03D8E02D8E03447012C701E",
INIT_0C => X"F8DE3C27CA181E5D710664A5F140C14BD32A2E281992940AFAA15C3FC0836310",
INIT_0D => X"F000BE0FC80020130841840308653FF0313FE92C23FB1EECB367C0F3E378F0BC",
INIT_0E => X"F000BE0FCD806FFFAF0AE83080E2AEB2F0F1E01BE53FE1F000BE0FC41BE53FE1",
INIT_0F => X"0231F0BF9E3F02A7FFD63669C0E008C3CB7F041BE1BFE1F000BE0FC41BE1BFE1",
INIT_10 => X"30180309A0F83FE2B87C7D006FFF9F1A7806013879BAA78FC103FF5F1F12F038",
INIT_11 => X"39E9C1DBF8A30C2098DBE2FF7F2320483136F200A822CBACAB9DDEB7F9BC291F",
INIT_12 => X"004C72BEC95FEF64E4090626DF15B7D1C6184131B7980DFFFC03F00003F01FB9",
INIT_13 => X"1DFFFA0A3C0202B8776AE7A7C9CBFFF060703080E29F1B79E9F6427EFE901C0E",
INIT_14 => X"2B716CA5C56620590350ACD3A7D5B7EFAC6DFC8C0312A0024B83F07F3999E9F2",
INIT_15 => X"F0BCAF3BC2F3BC6F0BCEF2BC2F3BC6DBC67C251104A2261253904580207E1C81",
INIT_16 => X"1BCEF0BC2F3BC2F1BCEF0BC6F2BC2F1BCAF1BC6F2BC6F2BCAF1BC2F3BC6F2BCE",
INIT_17 => X"BCEF0BC2F3BC2F1BCAF1BCAF3BC6F0BCEF0BCEF2BC6F2BCAF1BCAF1BC2F3BCAF",
INIT_18 => X"69CFEF73B6FFE7436DB6FD0831518424965B4D2492CB69AF1BCEF0BC6F2BC6F0",
INIT_19 => X"F7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF3EF9FBFBB9E79E7BEBCB7",
INIT_1A => X"DEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDF7DF7DF7D",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF29FDAF77BBDDEEF77BBDDEEF77BBD",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"AAA2802AA10FFFFFDE0008556AABA5D2ABFFEFFF800000000000000000000000",
INIT_1F => X"ABAF7AAA8BFFAA802ABFF087FFDF5508003FEBA087FD54BA0804154005555574",
INIT_20 => X"54AAF7D168B45AAAABDF55AA802AA1000003FEBA00002AABA5D2EBFEBAAAD16A",
INIT_21 => X"3DE005555575EFA2D142145A2FFE8B45FF80001555D2E955FFFFD5421EFAAFFD",
INIT_22 => X"FC00BA5D5568AAAF7AAAAAAAAA802AABA082E954005500021FF5D2EBFF550000",
INIT_23 => X"D5420AAAA843DFFFAAD1554005D7FD74AAAA840014500517FFEF007BEABFF5D7",
INIT_24 => X"2AABDE0055517FF555504154BAA2FBEAA105D2E97410FFD16AAAA5D2ABDEBAFF",
INIT_25 => X"000000000000000000000000000000000000000028BFF0855555455500174BAA",
INIT_26 => X"21E84124285C51574BAB68A2DA00FFFFFFE38085F6FA92552AB8FEFF78000000",
INIT_27 => X"925D2AB8EBABEDB6AA92F7AAA8BC7B68A28BC70075FDF45080A3AEAA007BD248",
INIT_28 => X"5FFFFD1471D7AAFBD0492EBD56DB7DBEAEBFF55BE842AA105D0A38EBA1C0428A",
INIT_29 => X"21FF492AB8F7D1C0438E38145B575EFA2DB45145B6F5EFB6DF78E05145552A92",
INIT_2A => X"7DFC70875EABC7557FC20AA415F68AAAF7AAAAA82BE8A28A9214249740041000",
INIT_2B => X"B6FABA542ABAE2AF7DF470AABE8A3AFD7A2DF55400557FD54AABE84001C55551",
INIT_2C => X"5557545490012482B6A0BAE2849043AFED1C0E10492B6FFEFA105D2A95410FFD",
INIT_2D => X"D2AAABEFFB8000000000000000000000000000000000000000000000428BEF00",
INIT_2E => X"082EA8AAA087FC20105504000AA5955554BAFFAEBDE10F7FBFDEBA007BFDE005",
INIT_2F => X"0512AA8AAA5D0028A005D2AA8ABAF7FBE8A00FFAEAAB45F3AAAAB4500557FF55",
INIT_30 => X"EFFFAA97545552A821EFFBD557555AAFBC2000A2D57FFFFF7AEBFF55FF8028A0",
INIT_31 => X"A005D04174100800021FF002EA8BEF5D0428ABA597FD55FFA2FFD5555FFD57FF",
INIT_32 => X"54AAF7800015551517DF45005168B55557FC0012087FEAABAF7AAAAA10F3AAAA",
INIT_33 => X"FFE005D2A95410F7FFFFEBA5D2EA8ABAFBFFD74BAF7AAA8B45AAFBD54005D7BD",
INIT_34 => X"00000000002ABEF005555555000402000FF802AAAA04452ABFF592E80010FFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000060000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(5),        -- Port A data input
DOA(0)   => data_read_a_hi(5),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(5),        -- Port B data input
DOB(0)   => data_read_b_hi(5),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_6_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10800B0061A01002840002C030028180004003220200403312301C4389B2082",
INIT_01 => X"060009C838394848188160000C42426041000000090800090210090000510200",
INIT_02 => X"00043040009001100000061000018070002408000000000648080000001210E0",
INIT_03 => X"0000800002054081020080801200A0000300008000201184681A0000410C4800",
INIT_04 => X"0808801040000001401048008100022401400002024024053200020089000100",
INIT_05 => X"0240040408402202002000C200400020A50000A0000010010001260808000520",
INIT_06 => X"44000881064500004600000013088002840C240F5048011200010000440C0146",
INIT_07 => X"0241914041FE83E010040110110003040020402A0000003E1000000488000201",
INIT_08 => X"8001BF002C4A01041B112020200110024029006FE09081002004902000012068",
INIT_09 => X"0083FE38A040100281353150ACB645AEF8C01404448000008011061204200108",
INIT_0A => X"3103AD0413424E4014D627C470462200011504420C0A962A2189002881404060",
INIT_0B => X"46C1060C16C96D15B0425B0425B1425B1425B0C25B0C25B1C25B1512D8212D82",
INIT_0C => X"009000140401100601016600A040220203A004480598010248000D0010420C0C",
INIT_0D => X"0000A01033A00013000000000018800F2400091081100C0090A5008200410020",
INIT_0E => X"0000A0103142000000000000000000455D0018100000000000A0103410000000",
INIT_0F => X"000000466800C200000000000000000001A0F4100000000000A0103410000000",
INIT_10 => X"00000000000024094680014200000000000000000041E8002900000000000000",
INIT_11 => X"F000322000000000000D1A000000000000034D240C2000502000000000000000",
INIT_12 => X"000000403F4000000000000068D24000000000001A60F0000000000000002007",
INIT_13 => X"C0000000000000000087C0003014000000000000000025D00008958000000000",
INIT_14 => X"02000000000814C219500150002800101280000000000000000000086670000C",
INIT_15 => X"8120C82208812048120882208892055A0060011280222413130449010301F051",
INIT_16 => X"3200802008320C82200802048320C82200812048320880200812048220880204",
INIT_17 => X"20C83208812048020883204802048120882204812008220C8220081204822088",
INIT_18 => X"79CFF1FE1E9F52ABEF9EFE8150120EC718638E38E30C71C812088220C8120080",
INIT_19 => X"71C71C71C71C71C71C71C71C71C71C71C71C71C71C736D9DBD9BBEFBEFBEBEF1",
INIT_1A => X"CFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FC71C71C71C",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCF29A7F3F9FCFE7F3F9FCFE7F3F9F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000607FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"EFA2FBD54BA5555554BAAAFBC20BA5D7BEAAAAFF800000000000000000000000",
INIT_1F => X"EBA0855421455555574AAA2802AA10FFFFFDE0008556AABA5D2ABFFEFFF843DF",
INIT_20 => X"DF5508003FEBA087FD54BA000415400550428AAAAA84021FF007BD54BAAAD17D",
INIT_21 => X"A8BFFAAD1554BA002A95555A28417400AAFBE8ABAF7FFD54AAAA802ABFF087FF",
INIT_22 => X"BD5545080417555A2D17FE1000003FEBA00002AABA5D2EBFEBAAAD16AABAF7AA",
INIT_23 => X"D5421EFAAFFD54AAF7D168B45AAAABDF55AA802AA100000001EF087FEAA00FFF",
INIT_24 => X"F80001555D2E955FFFF843DEAAA2803DFEF0855401FF082EA8B555D7FC21FFFF",
INIT_25 => X"0000000000000000000000000000000000000055575EFA2D142145A2FFE8B45F",
INIT_26 => X"2552AB8FEFF78E3DFFFAAFFD04AA415B52492B6F5C20825D7FE8A92FF8000000",
INIT_27 => X"EF147BD2482BED57AE921451421555551574BAB68A2DA00FFFFFFE38085F6FA9",
INIT_28 => X"4BAB68A28BC70075FDF45080A3AEAA007BD24821C04124281C0E2DA82BE8E001",
INIT_29 => X"8EBABEDB6AA92F7AAA8BC7B6D5524AA14209557DA28E15400BEF1EFA92FFFFD2",
INIT_2A => X"071FF0071EDA38F7F1D5555000417545B6D178E281C0A38EBA1C0428A925D2AB",
INIT_2B => X"4A8B555C7FC2147F7D1471D7AAFBD0492EBD56DB7DBEAEBFF55BE842AA105D0E",
INIT_2C => X"DB45145B6F5EFB6DF78E05145552A925FFFF8E3DE82BE8E38FFF0851401C7082",
INIT_2D => X"57FE8A00F38000000000000000000000000000000000000000000005B575EFA2",
INIT_2E => X"F7FBFDEBA007BFDE005D2AAABEFFBAABDFEFAAFBC00BA007BC0000FFD5420005",
INIT_2F => X"A592ABFE00F7AA821FF557FC0010F7D168A105D55421455155554BAFFAEBDE10",
INIT_30 => X"10F7D57DE00FFFBC00AAFBAAAAB4500557FF55082EA8AAA087FC20105504000A",
INIT_31 => X"AAA5D0028A005D2AA8ABAF7FBE8A00FFAEAAB45F3D5400BA5504155EFAAAE954",
INIT_32 => X"FF55FF8028A00512E975FF08557FEAAF7D157545080417545F7D56AAAA592AA8",
INIT_33 => X"AABEF005542155000028B555D7FC2145F3D557555AAFBC2000A2D57FFFFF7AEB",
INIT_34 => X"000000007FD55FFA2FFD5555FFD57FFEFFFAA97545552A821EFFBAABDE00F7AA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000048000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(6),        -- Port A data input
DOA(0)   => data_read_a_hi(6),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(6),        -- Port B data input
DOB(0)   => data_read_b_hi(6),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_7_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10844B00482258A2842112C02450418800002300500030B313300C418992002",
INIT_01 => X"020009C23838684D1C20E0000E11424840000000080000080200000000110204",
INIT_02 => X"000520700CA08910000206101180803081144880010400044808000000122160",
INIT_03 => X"000080040305208000008000328080040304008020303194289A000041484800",
INIT_04 => X"08088000000000010000CA008008060441000000028234493410820191000000",
INIT_05 => X"03500404000022020020044000000C208400408000001000984005949C002928",
INIT_06 => X"54000881044500004680000013008002940C24001A4A010200018920646410C7",
INIT_07 => X"22510040400500011204813015012204002040280000013E1000000488000201",
INIT_08 => X"9001A0602C4A01051B132820208001024069004008908002120851420001226A",
INIT_09 => X"01100020A2401008A20404E08200A05000A4264640800022C8198C4E05200018",
INIT_0A => X"20002000024040400050450440C48A0041140C420B0904208800904286000008",
INIT_0B => X"50822002120D2134800648006480064800648106481064810648193240432404",
INIT_0C => X"284A142288042A5C24202451505E00A621A5220A8091444040188C001B41210A",
INIT_0D => X"00F001F021141A12004104020810B000100000000109064C80010050A3285194",
INIT_0E => X"00F001F027420000400004C3201C514408081C1014800000F001F02810148000",
INIT_0F => X"E00E0E404100E200040900000B0380383480C81014800000F001F02810148000",
INIT_10 => X"4160C0301D07001D0402034200004000019860078641004039000180400002C0",
INIT_11 => X"08103BA0104810C8462416E8040446120C890814600010512000000080028400",
INIT_12 => X"98038D4030DD008088C2419120B740209021908C4846FC000200030F000FE006",
INIT_13 => X"DD000100411C81078884204035DC00201804C3201C60A408100DD58010440130",
INIT_14 => X"412024202211148019064200402A32901A8000B2048902C0807C0E00C448100D",
INIT_15 => X"50942509425194651946519465894619421421102000269243854D8002000250",
INIT_16 => X"19465194E50942509425094E51946519465094A50942509425194E5194651942",
INIT_17 => X"9425094251946539465094250946539465194250942509465194650942509425",
INIT_18 => X"0000000000000000000000080150890820800041041000052942509465194653",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF21E6C000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"AAF7D5575455D557DFEF002AAAB55002E820AAAA800000000000000000000000",
INIT_1F => X"B55007FD74AAAA843DFEFA2FBD54BA5555554BAAAFBC20BA5D7BEAAAAFFFBC00",
INIT_20 => X"AA10FFFFFDE0008556AABA5D2ABFFEFFFAAAAAAAF7D57FFEFF7D555555A2AEAA",
INIT_21 => X"42145552ABDFEFFFAA801EFFFFBFDF550000175555504175450055574AAA2802",
INIT_22 => X"A975EF00003DF55555168A00000428AAAAA84021FF007BD54BAAAD17DEBA0855",
INIT_23 => X"802ABFF087FFDF5508003FEBA087FD54BA000415400557BD74BAFFD140000082",
INIT_24 => X"AFBE8ABAF7FFD54AAAAAEA8ABA55557FEAAA2843FF55A2AEA8B55AAAABDEAAFF",
INIT_25 => X"0000000000000000000000000000000000000051554BA002A95555A28417400A",
INIT_26 => X"25D7FE8A92FFFFC70BAE3D155555415178FD7082EAAB550820870BAAA8000000",
INIT_27 => X"FFEBD55557DBEA4AFB550871D7482AA8E3DFFFAAFFD04AA415B52492B6F5C208",
INIT_28 => X"5550051574BAB68A2DA00FFFFFFE38085F6FA92552AB8FEFF7A0ADABAEBD578F",
INIT_29 => X"2482BED57AE921451421555524BDFD7FFA4801D7F7F5FDF55000E17545410E17",
INIT_2A => X"D2482E3D1450381C20905EF08003AF55415F6DA38080E2DA82BE8E001EF147BD",
INIT_2B => X"AAFB55ABA0BDE02EB8A28BC70075FDF45080A3AEAA007BD24821C04124281C7B",
INIT_2C => X"209557DA28E15400BEF1EFA92FFFFD24BAB6A4A8A82495F78E92AA843DF45BEA",
INIT_2D => X"800174BAA680000000000000000000000000000000000000000000055524AA14",
INIT_2E => X"007BC0000FFD542000557FE8A00F3FFD54BAAAD15754508556AB45002AA8B450",
INIT_2F => X"FFB803DEAAAAD56ABEFAAD5575EFF7803DF45085557410AEAABDFEFAAFBC00BA",
INIT_30 => X"55082E97555002E955550C55554BAFFAEBDE10F7FBFDEBA007BFDE005D2AAABE",
INIT_31 => X"E00F7AA821FF557FC0010F7D168A105D554214551003FF45FF8400145FFD57FF",
INIT_32 => X"20105504000AA597FC2010A2D1554AA5500021EF000028B55087BFDEBA042ABF",
INIT_33 => X"E8A00A2803FF45F7AABDF55AA843FE10AEAAAAB4500557FF55082EA8AAA087FC",
INIT_34 => X"0000000055400BA5504155EFAAAE95410F7D57DE00FFFBC00AAFB8028A00007F",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000007FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(7),        -- Port A data input
DOA(0)   => data_read_a_hi(7),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(7),        -- Port B data input
DOB(0)   => data_read_b_hi(7),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_8_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000B0000040042840002C0000001800000070000000033022000000000086",
INIT_01 => X"000009C21838284D1C2160000E12426840000000180800080200080040510200",
INIT_02 => X"0001004000900110000006100080003000240800014400004808000000122160",
INIT_03 => X"00008000020440810002A0801010A0044300000000200086011A000040404800",
INIT_04 => X"8000801000020401400040408108022029400000124004041200000089000100",
INIT_05 => X"02080424085022020000040200480020850010A0002010010120060800040400",
INIT_06 => X"50000880006500000680000011008006840C200018C1010200018920E0640102",
INIT_07 => X"426000404005000112048130150120240020400A0000013E1000000488000010",
INIT_08 => X"220100402C42010413110020200100024029004000A200002004902200012141",
INIT_09 => X"0000000080400008010410A2940A45240040140440800022C8388E1200A00008",
INIT_0A => X"00420100020048405000070440C0000001140412090000000021002081000048",
INIT_0B => X"0000000800000100011000010000100001000010000100001000010000880008",
INIT_0C => X"001000040001100008012008004020102180800804802000C0080D00100A0008",
INIT_0D => X"0FF0000002200A1200410402080080003000091085100C008124008000400020",
INIT_0E => X"0FF000000140000040F517CF600000000104081010001E0FF00000001010001E",
INIT_0F => X"E000000000804200000809963F1F80000000001010001E0FF00000001010001E",
INIT_10 => X"CFE7C0F00000000000810140000040E587F9E000000008100900008000ED0FC7",
INIT_11 => X"00021040030C73D80000021000585F3600000020240020102000000802419660",
INIT_12 => X"F80000000042000B0BD6C0000010800618E7B000000C000003F80FFF00000000",
INIT_13 => X"800005D5C3FD800000000008180000078A8FCF600000000002028001006AA3F1",
INIT_14 => X"020000000008808219002100100C000041120370DCAD1FC18000000000000202",
INIT_15 => X"8020080200812048120481204812055A04604930A02026934215410102000110",
INIT_16 => X"0200802008020080200802048120481204812048120481204802008020080200",
INIT_17 => X"2008020081204812048120481200802008020080200802048120481204812048",
INIT_18 => X"414A87D78AF42143CEBAC88151120A0000000000000000081204812008020080",
INIT_19 => X"F3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF7E799B1BEB65B65948051",
INIT_1A => X"C3E9F0FA7C3E9F0FA7C3E9F0FA7C3E9F0F87C3E1F0F87C3E1F0F87CF3CF3CF3C",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF1B5DA9F0FA7C3E9F0FA7C3E9F0FA7",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"0000043DF55087BC01EF007FD75FFFF84000AAFF800000000000000000000000",
INIT_1F => X"E10A28028AAAAAFBC00AAF7D5575455D557DFEF002AAAB55002E820AAAA84000",
INIT_20 => X"54BA5555554BAAAFBC20BA5D7BEAAAAFFAA95545552ABFE00087BC00AA082EBF",
INIT_21 => X"D74AAAAD57FF45002A975FF007BE8BFFA2FBFFFFFAAD5400AAFF843DFEFA2FBD",
INIT_22 => X"BE8A00082A97410F7D5555EFAAAAAAAAAF7D57FFEFF7D555555A2AEAAB55007F",
INIT_23 => X"55574AAA2802AA10FFFFFDE0008556AABA5D2ABFFEFFFAA82000555555545AAF",
INIT_24 => X"00017555550417545000015545087BC2010AAD54014500516ABFFA2AABDF4500",
INIT_25 => X"000000000000000000000000000000000000002ABDFEFFFAA801EFFFFBFDF550",
INIT_26 => X"50820870BAAA8407000140038F450075C71FF087BD75D7FF84050BAEB8000000",
INIT_27 => X"10007FC50BA002ABFE00AA8A2AABABEFFC70BAE3D155555415178FD7082EAAB5",
INIT_28 => X"082EB8E3DFFFAAFFD04AA415B52492B6F5C20825D7FE8A92FFA497545552AB8E",
INIT_29 => X"557DBEA4AFB550871D7482AAD17DF451C24955EF0875EFBD7B6F1FFFC7BEDB45",
INIT_2A => X"87000415B5057DAAFBE8A10082092410EBD5505EFB6A0ADABAEBD578FFFEBD55",
INIT_2B => X"B6ABC7B6AABFFED0051574BAB68A2DA00FFFFFFE38085F6FA92552AB8FEFF7AA",
INIT_2C => X"A4801D7F7F5FDF55000E17545410E17555000E17545007BC0000BED14217D005",
INIT_2D => X"784174AAA280000000000000000000000000000000000000000000024BDFD7FF",
INIT_2E => X"08556AB45002AA8B450800174BAA684174105D042AB550055555FF007BD7555F",
INIT_2F => X"0F384175555D2EA8A00087BD74BA082EBDE10AAAEA8ABAF7FFD54BAAAD157545",
INIT_30 => X"55FFD57DF55FFFBD5400A2AABDFEFAAFBC00BA007BC0000FFD542000557FE8A0",
INIT_31 => X"EAAAAD56ABEFAAD5575EFF7803DF45085557410AED17FF455D04155FF00557DF",
INIT_32 => X"DE005D2AAABEFFBAE97410087BC21EFA2FFEAA00000002010A2D5421FFFF803D",
INIT_33 => X"C0010FFD1401EF087FE8B55FFAEBDFEF0855554BAFFAEBDE10F7FBFDEBA007BF",
INIT_34 => X"00000000003FF45FF8400145FFD57FF55082E97555002E955550C2E95555087B",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000020000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(8),        -- Port A data input
DOA(0)   => data_read_a_hi(8),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(8),        -- Port B data input
DOB(0)   => data_read_b_hi(8),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_9_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00018248A2840112C00002C18000002300500030B3132000400812002",
INIT_01 => X"A140098218302849180060000C004240413C0A61590001D90213C90008510204",
INIT_02 => X"102008700CB089100002061031285074810448800104008048080080001210E2",
INIT_03 => X"00008015074608840390A0040040800203140000A00010800408108448020042",
INIT_04 => X"082080400004A00100000100840602020100000002C2344156108201811801C0",
INIT_05 => X"0200048480011502049500280020CC2084000080008010019161249C9C002188",
INIT_06 => X"70000881004500004E01020411D08000940C00001800010200018B20206C0102",
INIT_07 => X"EA70C0040005000312048130150100040020404A0000017E10408104C8000110",
INIT_08 => X"000000402C220104131004202081120050A5104000A204617201D10801002000",
INIT_09 => X"000800002F4924003085E51420A0100400641E4E40800022C8088C1220200908",
INIT_0A => X"20102000024040484028450001648C2229150400080244000401900284000440",
INIT_0B => X"0880110901081110411204112040120411204012041120401204111020090208",
INIT_0C => X"685B34A688841A5C21200101A01A0004009024028004044248404D00104B2100",
INIT_0D => X"0000A01000000213000000000000B0001000010000190E44802002D1A168D0B4",
INIT_0E => X"0000A010014000000000000000000040500008100400000000A0100410040000",
INIT_0F => X"0000004608004200040000000000000001A004100080000000A0100410008000",
INIT_10 => X"00000000000024080000014000000000000000000040A0000900010000000000",
INIT_11 => X"300013E010000000000D00F804000000000340000C0000102000000080000000",
INIT_12 => X"00000040091F0000800000006807C000800000001A0CFC000000000000002001",
INIT_13 => X"DD000000000000000082C00019DC002000000000000021500006D58010000000",
INIT_14 => X"03206420000000C019502050000C32901A800080000000000000000860100006",
INIT_15 => X"D1B46D1B46D0B42D0B42D0B42D8B424342342832002A24921082158802001011",
INIT_16 => X"0B42D0B42D0B42D0B42D0B46D1B46D1B46D1B46D1B46D1B46D1B46D1B46D1B46",
INIT_17 => X"B42D0B42D1B46D1B46D1B46D1B46D1B46D1B46D1B46D1B42D0B42D0B42D0B42D",
INIT_18 => X"89999E91BCD1512B871C4A0100000000000000000000000D0B42D0B42D0B42D0",
INIT_19 => X"A28A28A28A28A28A28A28A28A28A29A69A69A69A69A51C200807249041202AE6",
INIT_1A => X"8349A4D068341A0D269341A0D269341A0D068341A0D068341A0D068A28A28A28",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF2DA921A0D269341A0D068349A4D06",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"45A280154BA5555401EFFFD5421EFA2FFFFF555D000000000000000000000000",
INIT_1F => X"5EF00557DF555D040000000043DF55087BC01EF007FD75FFFF84000AAFFD57DF",
INIT_20 => X"75455D557DFEF002AAAB55002E820AAAA843DFEF00517DEBA007BFDFEFFFD157",
INIT_21 => X"28AAAAAAABDF45F7803FFEF555568AAAF7802AA00FFFBD7555087BC00AAF7D55",
INIT_22 => X"BD54BA550417400085155555082A95545552ABFE00087BC00AA082EBFE10A280",
INIT_23 => X"043DFEFA2FBD54BA5555554BAAAFBC20BA5D7BEAAAAFFFBC00AA552E95545087",
INIT_24 => X"2FBFFFFFAAD5400AAFF8402000A2FFFDF555D7BE8BFF5D51575EFA280175555D",
INIT_25 => X"00000000000000000000000000000000000000557FF45002A975FF007BE8BFFA",
INIT_26 => X"7FF84050BAEBDF78F45B68010482415B471C7E3DF451EFBEFBFAF45490000000",
INIT_27 => X"82007FFAFEFE3DB505EF1C5B7AF45490407000140038F450075C71FF087BD75D",
INIT_28 => X"5451C7FC70BAE3D155555415178FD7082EAAB550820870BAAA8438FFF00517DE",
INIT_29 => X"50BA002ABFE00AA8A2AABABEAEB8F45F78A3DFD741516DAAAE38E2DA28EBFFD5",
INIT_2A => X"C20BA5D2E905550071D54825D0A1543808515756D1C2497545552AB8E10007FC",
INIT_2B => X"5505FFBE801256D490E3DFFFAAFFD04AA415B52492B6F5C20825D7FE8A92FFFF",
INIT_2C => X"24955EF0875EFBD7B6F1FFFC7BEDB45082EB8002000AAFFFDF6D417FEABEF5D5",
INIT_2D => X"7FBE8B5500000000000000000000000000000000000000000000000517DF451C",
INIT_2E => X"0055555FF007BD7555F784174AAA2FBEAB45F78402010007BD5545AAFFD55EFF",
INIT_2F => X"AA68028BEF00517FE10007BE8BFFAAFFC01FF557FE8B550004174105D042AB55",
INIT_30 => X"AAAAAEBFEAAAAFFD5545557FD54BAAAD15754508556AB45002AA8B450800174B",
INIT_31 => X"5555D2EA8A00087BD74BA082EBDE10AAAEA8ABAF7AAAAB45F7AEBFF4508557FE",
INIT_32 => X"2000557FE8A00F3FFC00BA552E80145005557400552A954BA0051575EF550417",
INIT_33 => X"FDFFF007FE8BFF5551401EFF784021FF002ABDFEFAAFBC00BA007BC0000FFD54",
INIT_34 => X"00000000517FF455D04155FF00557DF55FFD57DF55FFFBD5400A28400010A2FB",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000040000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(9),        -- Port A data input
DOA(0)   => data_read_a_hi(9),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(9),        -- Port B data input
DOB(0)   => data_read_b_hi(9),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_10_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00018248A2840112C00002C18000202300500030B3132000400992006",
INIT_01 => X"A140098218302849180060000C00424040000000080000080200090008510204",
INIT_02 => X"102100400C8001100000061000A8503401044880010400004808000000122160",
INIT_03 => X"000080150746088401908000100080020304000020201080001A108448404842",
INIT_04 => X"800080400004A001000040008406020201000000020004401000000180180080",
INIT_05 => X"02000484800133020495040800208C20A4000080000010000001249010042008",
INIT_06 => X"50000881004500004681020411808000940C20001800010200018920206C0102",
INIT_07 => X"024084044005000112048130150120040020400A0000013E10408104C8000010",
INIT_08 => X"000100402C020105131100200000124250A51040088084614001110801012000",
INIT_09 => X"00080082CD09240820800000000000040000180840800022C8088C1220200108",
INIT_0A => X"841201000200484910000F050560262229140402080200A00402000484140400",
INIT_0B => X"0010118900080010000200102001020000200002001020010200001000010008",
INIT_0C => X"408120900404004821202001F05E00040180260A8080044240004C0010800228",
INIT_0D => X"0000A01000000813004104020800800030000800010008088124020102008100",
INIT_0E => X"0000A010014000004000000000000040500008101480000000A0100410148000",
INIT_0F => X"0000004608004200040900000000000001A004101480000000A0100410148000",
INIT_10 => X"00000000000024080000014000004000000000000040A0000900018040000000",
INIT_11 => X"3800100010480000000D00000404400000034000282000102000000080028000",
INIT_12 => X"00000040090000808800000068000020900000001A0000000200000000002001",
INIT_13 => X"80000100000000000082E0001000002018000000000021580000800010440000",
INIT_14 => X"00004000000004C0195000500008000000000082008000000000000860180000",
INIT_15 => X"0100401004010040100401004090055804404110802A24921317580802001011",
INIT_16 => X"0000000000000000000000040100401004010040100401004010040100401004",
INIT_17 => X"0040100400000000000000000000000000000000000000000000000000000000",
INIT_18 => X"215281FC1A72E2486AAA40A85052020000000000000000001004010040100401",
INIT_19 => X"51451451451451451451451451451451451451451452AA83330A8A28A29EA8D1",
INIT_1A => X"5CA6532994CA6532B95CAE572994CA6532994CA6532994CA6532994514514514",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF31CE2E572994CA6532994CAE572B9",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"10AAFBE8AAAA2D540000F7D57DF55A2AABFFEF08000000000000000000000000",
INIT_1F => X"F45FFFBC2010AAD57DF45A280154BA5555401EFFFD5421EFA2FFFFF555D003FE",
INIT_20 => X"DF55087BC01EF007FD75FFFF84000AAFF8002155AAFFE8B45AAD540000087FFD",
INIT_21 => X"7DF555D517FEBA082A801EFF7FBD5400FFD568B555D00155EF08040000000043",
INIT_22 => X"BFDE00A2FBC0145005168A10AA843DFEF00517DEBA007BFDFEFFFD1575EF0055",
INIT_23 => X"7BC00AAF7D5575455D557DFEF002AAAB55002E820AAAA803FEBA082AAAAAAF7F",
INIT_24 => X"7802AA00FFFBD7555082E82155FFAEAAB55AAD568B455D00154BAFFFBD75EF5D",
INIT_25 => X"000000000000000000000000000000000000002ABDF45F7803FFEF555568AAAF",
INIT_26 => X"FBEFBFAF4549003DE10BEF5EDAAAAAD547038EBD57DF7DA2AEB8FC7000000000",
INIT_27 => X"6DAADF470280075FFF45E3F1C7038A2DF78F45B68010482415B471C7E3DF451E",
INIT_28 => X"5C7000407000140038F450075C71FF087BD75D7FF84050BAEB8002155BEF5EDB",
INIT_29 => X"AFEFE3DB505EF1C5B7AF45495B7DEAA0824851EFEBFBD2410EBD168B7D410A17",
INIT_2A => X"38EAA0824A8AAAEBF5FAE28AAF1C2155005F68A10A28438FFF00517DE82007FF",
INIT_2B => X"4104AAF7F1D75EF557FC70BAE3D155555415178FD7082EAAB550820870BAAA80",
INIT_2C => X"8A3DFD741516DAAAE38E2DA28EBFFD55451C2087155EBA4A8B7DAADF68B7D410",
INIT_2D => X"2AEAAB55000000000000000000000000000000000000000000000002EB8F45F7",
INIT_2E => X"007BD5545AAFFD55EFF7FBE8B5500043FE00F7D17FEBAA2D5574BAAAD17DFEFA",
INIT_2F => X"AA28002155FFD17FFFFA2FBD74BA00557FF45A2D5554AAA2FBEAB45F78402010",
INIT_30 => X"00AAD16ABFF002A975450004174105D042AB550055555FF007BD7555F784174A",
INIT_31 => X"BEF00517FE10007BE8BFFAAFFC01FF557FE8B55007FFDEAA0004175FFA2FBC20",
INIT_32 => X"8B450800174BAA68428AAA08042AABAAAD56AABAAAD140155087FEAA10A28028",
INIT_33 => X"2ABEFAAFBE8BFF0004020AAFFD5555EF557FD54BAAAD15754508556AB45002AA",
INIT_34 => X"000000002AAAB45F7AEBFF4508557FEAAAAAEBFEAAAAFFD5545550015555A284",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000047FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(10),        -- Port A data input
DOA(0)   => data_read_a_hi(10),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(10),        -- Port B data input
DOB(0)   => data_read_b_hi(10),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_11_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10180B05A0010402840602C2D001019000000300000000330A20080EC180002",
INIT_01 => X"AB400984B830084C1820E0000C36424840000000080000088200000802112220",
INIT_02 => X"102A68440080011000000618062AD03502640800010410424908136019920868",
INIT_03 => X"001282118644C88481908001106088022300000080F4925CDC9A10844A9A4842",
INIT_04 => X"401280480004A1011000418084460002E12000000200040010000040A8000000",
INIT_05 => X"0FC8048484011502059511488020802084400888001110000000050000005400",
INIT_06 => X"1011088AE24500001631024511C08004A70AA40008B90D0200018B60A0650D45",
INIT_07 => X"020011005405000910040150110041040024400D800002BE18408104C9205908",
INIT_08 => X"89390040280241041D175820000001020061004004800567403512A801014C46",
INIT_09 => X"050800E20D09A424C5840400808000040680180840800022D8288E946CA00833",
INIT_0A => X"85002000024040410A000D0504408C32E915D9C208050084840201A099100400",
INIT_0B => X"B01011934A005101431CA821CA831CA821CA831CA831CA821CA83165410E5410",
INIT_0C => X"00010080028000010402214850444091019B02080885200042A9CC001000003A",
INIT_0D => X"5A5018C5A0A00812004104020808B00030000808024008008325820000000000",
INIT_0E => X"5A5018C5AB0062C38A4DB680A0D8241500D5761B011986695014A96E1A811986",
INIT_0F => X"42056A289A1BB2078A922DA2A8B180A2600AAE1A811986695014A96E1B011986",
INIT_10 => X"05AA429189B60AC43C6C7F0272C3841DB528802CAB18468F4101621B1BAC8455",
INIT_11 => X"C003104289A668B8CAB270106338317A3D94392020224ACDE215883078681B5C",
INIT_12 => X"804B020A06020C67061BC785938085134CD551BCA1C90006C0C2958502861120",
INIT_13 => X"80819A5539D503336D61056ABA006282806CA64090B89E015AAA880E48382EB8",
INIT_14 => X"40000000E808989003066E03513E41470126C6284B2D20410AB4503089C00A82",
INIT_15 => X"0000000000000000000000000000041800400110200026124202500802000800",
INIT_16 => X"1004010040100401004010000000000000000000000000000000000000000000",
INIT_17 => X"0040100401004010040100401004010040100401004010040100401004010040",
INIT_18 => X"C110083018162148420840280050800000000000000000001004010040100401",
INIT_19 => X"000000000000000000000000000001041041041041003882928E0000000AA0C4",
INIT_1A => X"0000000000008040000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3E0FC000000000000020100000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"EFAA842ABEFA280155EFFFFBC01EF08554000055000000000000000000000000",
INIT_1F => X"F4508514000000003FE10AAFBE8AAAA2D540000F7D57DF55A2AABFFEF0804155",
INIT_20 => X"54BA5555401EFFFD5421EFA2FFFFF555D51575FFA2FFD75FF550015400FFFBFF",
INIT_21 => X"C2010AAD568AAAAAD142145FF80155EF0051555FF0804155FFF7D57DF45A2801",
INIT_22 => X"01540008514215555003DFFFA28002155AAFFE8B45AAD540000087FFDF45FFFB",
INIT_23 => X"040000000043DF55087BC01EF007FD75FFFF84000AAFF802ABFFA2AABFE10080",
INIT_24 => X"FD568B555D00155EF085168B45085142010FFAE800AA5D7BFDF45F7FFEAA0000",
INIT_25 => X"00000000000000000000000000000000000000517FEBA082A801EFF7FBD5400F",
INIT_26 => X"DA2AEB8FC70000175EFB6802DBC7BE8A155EFE3FBC71FF145B42038550000000",
INIT_27 => X"EF550E15400E3F1FFF7D085B420381C003DE10BEF5EDAAAAAD547038EBD57DF7",
INIT_28 => X"5C7F7DF78F45B68010482415B471C7E3DF451EFBEFBFAF45495F575FFBEF5D05",
INIT_29 => X"70280075FFF45E3F1C7038A2DB68ABAB6D145145FF84155D7085B555C7140410",
INIT_2A => X"28BEFBEA4BDE28140A1543800514515549003FFC7BE8002155BEF5EDB6DAADF4",
INIT_2B => X"FFFF7DE3F1EFA10140407000140038F450075C71FF087BD75D7FF84050BAEB84",
INIT_2C => X"24851EFEBFBD2410EBD168B7D410A175C7005B6DB55145140000FFAE85082417",
INIT_2D => X"57BC20AA5D0000000000000000000000000000000000000000000005B7DEAA08",
INIT_2E => X"A2D5574BAAAD17DFEFA2AEAAB550004175FFF7803DF45FFAE955EFAAFBD55EF5",
INIT_2F => X"5007FD75FFF7D5401EF5D2E97410AAD17DFEF007FC20AA5D043FE00F7D17FEBA",
INIT_30 => X"55007FD5545550400145FFFBEAB45F78402010007BD5545AAFFD55EFF7FBE8B5",
INIT_31 => X"155FFD17FFFFA2FBD74BA00557FF45A2D5554AAA2FBEAAAAFFD555545FF80155",
INIT_32 => X"7555F784174AAA2842ABEFFF803DEAA5D2E974AA00515754500003FF55FF8002",
INIT_33 => X"40000FFAE97410007BFFFFFA2D57FE105D04174105D042AB550055555FF007BD",
INIT_34 => X"000000007FFDEAA0004175FFA2FBC2000AAD16ABFF002A97545007FFFF455555",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000040000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(11),        -- Port A data input
DOA(0)   => data_read_a_hi(11),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(11),        -- Port B data input
DOB(0)   => data_read_b_hi(11),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_12_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50080B01BC002006940202C0DE041196A83183000000023322287E0FC000006",
INIT_01 => X"0E000C068000E04D40238000001702484000000008000008820009280A553231",
INIT_02 => X"400B71440C8001100000171C0283813013766A800586235ECC09C8423B962966",
INIT_03 => X"CC618E048306E082000081000040900003548421A080025EDF08421042DC0108",
INIT_04 => X"00028020000000812000012080080000E100001002000448100000C1BC18008C",
INIT_05 => X"0FF8060610000402010015E100004C2084800090000310000000079010007C19",
INIT_06 => X"33992D98DEC74A003EA468D01510C03E8F580C800A3F018200418927E0668645",
INIT_07 => X"0204000406050013142409121142F746222EE2498000007E111204058B84C50C",
INIT_08 => X"E826A0602902A10491165C200000820018A5104010C01086003C13E000004EDF",
INIT_09 => X"023000000000000867000000000000040000600060801022C9F88D244FA40133",
INIT_0A => X"00100000820040482B28050001600010C13499F01B334015980001E09F000000",
INIT_0B => X"B80460124F16F06BC20CBC30CBC20CBC20CBC30CBC20CBC20CBC3065E1865E10",
INIT_0C => X"00000000029D204B7C0382FD0100F3F9F80FA0200E0BF40063F99C0010000012",
INIT_0D => X"93900F6EE230301208008001007A80001100002002801000A042000000000000",
INIT_0E => X"93900F6EEC421392C96B1237E0D8BD9629F97E0B348EDAC3900F6EFA0B158EDA",
INIT_0F => X"622DBC31D73F6006A5891533EF9500EAE64BCA0B158EDAC3900F6EFA0B348EDA",
INIT_10 => X"C2B083798D341B10DEFE14400392C74CAEAD412EDD2B4FCFF812A383430C669E",
INIT_11 => X"49FAB442994B3238D4E2FB104636652E19B8BA30C022DAD8C100CA39E8CEBE66",
INIT_12 => X"30469392526208C6CC95C33717D88532966471A9C5DD00B12728D5360234D62A",
INIT_13 => X"828C4999AF580395542D27CDBA0020F0FABAC800DA550C29F36A8A2554E48A64",
INIT_14 => X"40000000873FB80B8A00EF03F56CC12B416A51B60585A5C28895962502E9F36A",
INIT_15 => X"0000000000000000000000000000008000000410802A26924010000002000EE0",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"28C1111026C152A121960A884042020000000000000000000000000000000000",
INIT_19 => X"2082082082082082082082082082092492492492492400200005A8A28A200A37",
INIT_1A => X"964B2592C964B2592C964B2592C964B2590C86432190C86432190C8208208208",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF400FEB2592C964B2592C964B2592C",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FF00042ABEFFF8400010082EAABFF55002ABEF08000000000000000000000000",
INIT_1F => X"BEFFFFBD54000004155EFAA842ABEFA280155EFFFFBC01EF0855400005555421",
INIT_20 => X"8AAAA2D540000F7D57DF55A2AABFFEF08556AA10000028AAAFFD15541000002A",
INIT_21 => X"40000005168AAA087BFFFFF5D04001FF00041554555557FE005D003FE10AAFBE",
INIT_22 => X"1555FF082AA8B55F7AEA8BEF5551575FFA2FFD75FF550015400FFFBFFF450851",
INIT_23 => X"D57DF45A280154BA5555401EFFFD5421EFA2FFFFF555D0000145082E955FF085",
INIT_24 => X"051555FF0804155FFF7842AA100000020BAAA801541055042ABEFFFFBD5410AA",
INIT_25 => X"000000000000000000000000000000000000005568AAAAAD142145FF80155EF0",
INIT_26 => X"F145B42038555F401D71C0A2DBC7EB80000280824ADBD7490E28BEF080000000",
INIT_27 => X"82FFDB5243800002FBD7EBFBD24101C00175EFB6802DBC7BE8A155EFE3FBC71F",
INIT_28 => X"E1041003DE10BEF5EDAAAAAD547038EBD57DF7DA2AEB8FC7005F6AA381C0A2DA",
INIT_29 => X"5400E3F1FFF7D085B420381C5B6AA82147FF8FEF410E001FF000E17555555B7A",
INIT_2A => X"0017D142E905EF1451525C7082AADB45F7AEA8BEF555F575FFBEF5D05EF550E1",
INIT_2B => X"02FBEFEBFBD2410AADF78F45B68010482415B471C7E3DF451EFBEFBFAF454900",
INIT_2C => X"D145145FF84155D7085B555C71404105C7F7842FA381C0A00082AA8A10410410",
INIT_2D => X"02AA8BEF000000000000000000000000000000000000000000000005B68ABAB6",
INIT_2E => X"FFAE955EFAAFBD55EF557BC20AA5D7BC01555D2EBFF55A284000AA08003FF550",
INIT_2F => X"5007BE8AAA5D2EBDE00FFFFC00AA08003FF55A2FBC00105D04175FFF7803DF45",
INIT_30 => X"FF082A97555557FE8A0000043FE00F7D17FEBAA2D5574BAAAD17DFEFA2AEAAB5",
INIT_31 => X"5FFF7D5401EF5D2E97410AAD17DFEF007FC20AA5D7BE8A005D7FEABFF002E821",
INIT_32 => X"55EFF7FBE8B550004001FF5D2A801EF5D5142145082EBFF55F7AAAABEF5D7FD7",
INIT_33 => X"82010A2AA8000008043FFFFA2FBC2010A2FBEAB45F78402010007BD5545AAFFD",
INIT_34 => X"000000007BEAAAAFFD555545FF8015555007FD5545550400145FF843DEAA552A",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000007FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(12),        -- Port A data input
DOA(0)   => data_read_a_hi(12),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(12),        -- Port B data input
DOB(0)   => data_read_b_hi(12),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_13_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10110A0441812402840402822007818000E00700000000330A3000000008042",
INIT_01 => X"A1400986B830E84D182260000C1042484001000008220008A20019080A510200",
INIT_02 => X"10A108600C9141100000C6180CA85035010E4880010431004908135980122D60",
INIT_03 => X"0013881507460886C190832175809C02030400002020124C441A108468424842",
INIT_04 => X"203080680204A0113801D600864E0C96C12000008244244052200201801802C0",
INIT_05 => X"030004849601110204950409C0208C2084E0009C0000100120A00C9918002098",
INIT_06 => X"10000882804544921681428591908000AF28A8002BC00D020003896020658FC4",
INIT_07 => X"CA20400450050009100501501102E0042020448D0000023E10408144C800D800",
INIT_08 => X"1D2B00402B220104B53100200001020218A5104016CC1C616401910801010100",
INIT_09 => X"050800404D49A42EB08000000000000406481C8C408000A2D8088D1820200B00",
INIT_0A => X"0010000002004048AA08050401604462E9144002090740148441200484000500",
INIT_0B => X"000A112100000000010000000001000000000000001000000000000000800000",
INIT_0C => X"509528954404144C200425010040000001B020081094040072005C0030864208",
INIT_0D => X"1C10B3831034081200000000000430003000206822F20CA8826AC2A14250A128",
INIT_0E => X"1C10B383110218CB0E54C2EA404A4F03D404A41AA5B7344C10B383081BA4B734",
INIT_0F => X"8001CE3E20A5B284ED1132909C72885A2B2C381BA4B7344C10B383081AA5B734",
INIT_10 => X"AC3CC0C0B8182597A801610218CB0C3548B3A008E730A01AB113A5524E6ACA67",
INIT_11 => X"A151EC5952E44128CA194517354C180A3C066430202021252991C22C99731014",
INIT_12 => X"1804C8A0ADA2E6A983014780CA28B2A5C8825194332B018A444AEA2701288A15",
INIT_13 => X"02D09852745F80112C428562EE0353635232D50048A411C158BB0A7910142C77",
INIT_14 => X"4240480068001C9B9150A0000297046E4023F8BE8E3E1E0109472C3EB50158BB",
INIT_15 => X"A1284A1284A1284A1284A1284A12851A84284110406A26924302590806000110",
INIT_16 => X"1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284",
INIT_17 => X"284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A",
INIT_18 => X"7DDFE7EFBEFFE7D3EFBEFC48A0550000000000000000000A1284A1284A1284A1",
INIT_19 => X"D75D75D75D75D75D75D75D75D75D75D75D75D75D75D7EFBFBFBBAAAAAABEFDF7",
INIT_1A => X"5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5D75D75D75",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000FEFD7EBF5FAFD7EBF5FAFD7EBF",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"AA5D043FFFFAAAABDEAA557BFDE00FFD140155F7800000000000000000000000",
INIT_1F => X"400AAD540155A2D5421FF00042ABEFFF8400010082EAABFF55002ABEF08556AA",
INIT_20 => X"ABEFA280155EFFFFBC01EF08554000055043DEBAF7843FFFFF7AABDF55A2AA97",
INIT_21 => X"D5400005568A1055043DEBAAAFFE8B45557FD7410552EAAABAAA84155EFAA842",
INIT_22 => X"FE8ABAAA8428A00087BD7555FFD56AA10000028AAAFFD15541000002ABEFFFFB",
INIT_23 => X"803FE10AAFBE8AAAA2D540000F7D57DF55A2AABFFEF085557545FFD17DEBAA2F",
INIT_24 => X"0041554555557FE005D0000155557BEAABA5D2ABDF450851420AA5D7FD5555A2",
INIT_25 => X"000000000000000000000000000000000000005168AAA087BFFFFF5D04001FF0",
INIT_26 => X"7490E28BEF08516DA82410A3FFD7AAA4B8E824971F8E38E3DF45155EB8000000",
INIT_27 => X"D7EBA4BDF45AAAA90410BEDF45155A2DF401D71C0A2DBC7EB80000280824ADBD",
INIT_28 => X"A82B680175EFB6802DBC7BE8A155EFE3FBC71FF145B42038550E38E92EB803FF",
INIT_29 => X"243800002FBD7EBFBD24101C556FA38490A3FE92BEFFEAB45417FD24385D2AAF",
INIT_2A => X"5056DE3D17FE92BEF1EFA92AA8428A10007FD557DFFDF6AA381C0A2DA82FFDB5",
INIT_2B => X"B400925D7FD557DA2803DE10BEF5EDAAAAAD547038EBD57DF7DA2AEB8FC70051",
INIT_2C => X"7FF8FEF410E001FF000E17555555B7AE10410E00155497FEFABA4120B8F55085",
INIT_2D => X"2FBD7545AA8000000000000000000000000000000000000000000005B6AA8214",
INIT_2E => X"A284000AA08003FF55002AA8BEF00517FE00082EBDF45AA8428A10085568ABAA",
INIT_2F => X"A5D2EA8A00A2803DF45AA843DF55AAAE82000F7FBD5545AAFBC01555D2EBFF55",
INIT_30 => X"55087FC00BA552ABFE10F784175FFF7803DF45FFAE955EFAAFBD55EF557BC20A",
INIT_31 => X"AAA5D2EBDE00FFFFC00AA08003FF55A2FBC00105D517FEAA082EBFE10F7FFE8B",
INIT_32 => X"DFEFA2AEAAB550051401FFA2D57FE10F7D57DE00AA842AA00007FD75FFF7FBE8",
INIT_33 => X"FDEAA08042AB45087FC0010557FD55FFAA843FE00F7D17FEBAA2D5574BAAAD17",
INIT_34 => X"000000007BE8A005D7FEABFF002E821FF082A97555557FE8A00002E82155007B",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000067FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(13),        -- Port A data input
DOA(0)   => data_read_a_hi(13),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(13),        -- Port B data input
DOB(0)   => data_read_b_hi(13),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_14_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10020A000180000284008280000281800000030000000033022000000580002",
INIT_01 => X"A14009821830284D186860000C30C24840000000084000084200090008510200",
INIT_02 => X"102100600C9001100000061020A8503401044880010400204908012018122F64",
INIT_03 => X"00008015074608840190800010008002030400002074F401209A108448404842",
INIT_04 => X"000080400004A00100004000840E000201000000024024401200020180180080",
INIT_05 => X"0A000484800111020495040800208C2084000080000010010020049818002008",
INIT_06 => X"1000088020450402B6A1420511C080008468A80008000D0200018B202067AF10",
INIT_07 => X"422000044005000910040110510260040024400C800000BE3850A144C924080E",
INIT_08 => X"000B004028020104111100200001020210A51040008004616001910801010000",
INIT_09 => X"000800004D492408208000000000000406401C0C40800022C8088DB420200900",
INIT_0A => X"0010000002004048000005040160042229140002090200000401000484000400",
INIT_0B => X"0000110100000000010000100000000000000100000000000000100000000000",
INIT_0C => X"409120940404104C2000210100400000011020080084040040005C0010820208",
INIT_0D => X"E0E0A0000190081200000000000000003000000000100C088020028102408120",
INIT_0E => X"E0E0A0000B02740421A0E5D1A024002050805210040000B0E0A0000210040000",
INIT_0F => X"E01200860008920106460D4501CB000111300210008000B0E0A0000210008000",
INIT_10 => X"0ABBC00905C33C6000400F02740412C0715C40110080A4006110510C14D18178",
INIT_11 => X"20000041DB011CC000090012565306500002411420220080220C0093C3892324",
INIT_12 => X"5809240C09024A4AE0CA00004800839682398000120800658992F3C700C30181",
INIT_13 => X"002B46867DBC002A830280000800F7B7A0B1E240240A8340000200067EAA8CB6",
INIT_14 => X"42004005800004801150A00341244000845C7DB0D0200900422ACA4B28000002",
INIT_15 => X"8120481204812048120481204812051A04204110002A26924302590802000000",
INIT_16 => X"1204812048120481204812048120481204812048120481204812048120481204",
INIT_17 => X"2048120481204812048120481204812048120481204812048120481204812048",
INIT_18 => X"69CB91FE1EF7D3ABEFBECA080050000000000000000000081204812048120481",
INIT_19 => X"F3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF7EFBBBBBF9E79E7BEAAF3",
INIT_1A => X"CFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCF3CF3CF3C",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FF007F3F9FCFE7F3F9FCFE7F3F9F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"45AAD157400007BEAAAAAAAE955555D5568A105D000000000000000000000000",
INIT_1F => X"0AAF784020AAF7D56AAAA5D043FFFFAAAABDEAA557BFDE00FFD140155F7D17DF",
INIT_20 => X"ABEFFF8400010082EAABFF55002ABEF085155400FFD1420100055574AAA2AA80",
INIT_21 => X"40155A28028B550051574005D7FFFE105D7BD7545A284020BA0055421FF00042",
INIT_22 => X"1421FF5D7FFDEBA085168B45FF843DEBAF7843FFFFF7AABDF55A2AA97400AAD5",
INIT_23 => X"04155EFAA842ABEFA280155EFFFFBC01EF08554000055002AB455D5142010085",
INIT_24 => X"57FD7410552EAAABAAA8017400AAD140000002EBFFEFA2AAA8BEFF780021FF55",
INIT_25 => X"000000000000000000000000000000000000005568A1055043DEBAAAFFE8B455",
INIT_26 => X"8E3DF45155EBD17FF6DAADB504001C71EDA82AAA0955455D556DA00490000000",
INIT_27 => X"101C55554AAAAA480082FF84000BAEBD16DA82410A3FFD7AAA4B8E824971F8E3",
INIT_28 => X"092085F401D71C0A2DBC7EB80000280824ADBD7490E28BEF085157428FFDB420",
INIT_29 => X"DF45AAAA90410BEDF45155A28E2AB7D0051504005D71F8E004975D556DB68405",
INIT_2A => X"28B6D5D51420101C5B401EF417BFAEAA08516AB45E38E38E92EB803FFD7EBA4B",
INIT_2B => X"EAFBC7EB80071FF5500175EFB6802DBC7BE8A155EFE3FBC71FF145B420385500",
INIT_2C => X"0A3FE92BEFFEAB45417FD24385D2AAFA82B68015400AADB40000082EBFFC7A2A",
INIT_2D => X"5557FE1000000000000000000000000000000000000000000000000556FA3849",
INIT_2E => X"AA8428A10085568ABAA2FBD7545AAD17DFFFAAFFC200055557DE00A280155455",
INIT_2F => X"F0051554AAFFFFC00105D55554BAA28400000F784020BAAAD17FE00082EBDF45",
INIT_30 => X"000051575FFF78415410087BC01555D2EBFF55A284000AA08003FF55002AA8BE",
INIT_31 => X"A00A2803DF45AA843DF55AAAE82000F7FBD5545AAAEAABFF0051400105D5568A",
INIT_32 => X"55EF557BC20AA5D042ABFF555142000557FC01EF007FEAABA00556AB55A2AEA8",
INIT_33 => X"C0010082EBDF55A2AABDF45A284175FF5D04175FFF7803DF45FFAE955EFAAFBD",
INIT_34 => X"00000000517FEAA082EBFE10F7FFE8B55087FC00BA552ABFE10F78415400A2FB",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000007FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(14),        -- Port A data input
DOA(0)   => data_read_a_hi(14),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(14),        -- Port B data input
DOB(0)   => data_read_b_hi(14),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_15_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000A000000000284000280000001800020030000000033022000000180002",
INIT_01 => X"A140098018300848180060000C00426040000000080000080200000000110200",
INIT_02 => X"1020004000801110000006100028503400040800010430004808000180120278",
INIT_03 => X"00008011064408840190800000228002A3000000000010000008108448000042",
INIT_04 => X"701280400004A991000000A28406000211000000220004941000000880000000",
INIT_05 => X"02000484800155020495000800218020C4002880005310000000040000000001",
INIT_06 => X"10000880004540000711224491C08000850A880008000D020001892020656300",
INIT_07 => X"8A04000016050009140501505100000420204008000000BE70408104C8000000",
INIT_08 => X"001F004028026104111002200000000200210040008004614001100801010000",
INIT_09 => X"000800000D09240000800000000000040600180840800022C8088C1020200000",
INIT_0A => X"0000000002004040000105000040042229140002080000000400000080000400",
INIT_0B => X"0000110100000000010000100001000010000000000000000000100000800008",
INIT_0C => X"0001008000000000000025000040000001300008009400006200580010000000",
INIT_0D => X"0000000002300012000000000004200030000000000008008020020000000000",
INIT_0E => X"0000000001000000400000000000000000000010108000000000000010108000",
INIT_0F => X"0000000000000200000900000000000000000010140000000000000010140000",
INIT_10 => X"0140000000000000000001000000400000000000000000000100008040000000",
INIT_11 => X"0000004000480000000000100004400000000030002000406000000000068409",
INIT_12 => X"8000000000020080080000000000802010000000000800000201000800000000",
INIT_13 => X"00000100000000000000000008000000184400A0000000000002000000441108",
INIT_14 => X"4000000000000000010620000004000000000242038B82800000000000000002",
INIT_15 => X"0000000000000000000000000000041800000110000024130202500802000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000080050000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"000804154AA5D00001EFF78428AAA007BC2145F7800000000000000000000000",
INIT_1F => X"0AA007FC2000F7D17DF45AAD157400007BEAAAAAAAE955555D5568A105D7FC00",
INIT_20 => X"FFFFAAAABDEAA557BFDE00FFD140155F7FBD74AAAAD17DF45F7D1421EF005540",
INIT_21 => X"020AAF7FFFDF45FF84000BA552ABDFEF08517DF55A2FBEAB555D556AAAA5D043",
INIT_22 => X"FEAB45F7843FF45082A801FF005155400FFD1420100055574AAA2AA800AAF784",
INIT_23 => X"D5421FF00042ABEFFF8400010082EAABFF55002ABEF087BE8ABA555168B55AAF",
INIT_24 => X"D7BD7545A284020BA007FFFE10A284000AA0055401550055574005D2E800AAA2",
INIT_25 => X"000000000000000000000000000000000000000028B550051574005D7FFFE105",
INIT_26 => X"55D556DA004971C7038140012482550E021C7EB8028A821C7BC516DFF8000000",
INIT_27 => X"45E3DF471C70851400BA0071C5028FFD17FF6DAADB504001C71EDA82AAA09554",
INIT_28 => X"B555D516DA82410A3FFD7AAA4B8E824971F8E38E3DF45155EBF1D5492BED17FF",
INIT_29 => X"54AAAAA480082FF84000BAEBF1FFF7DEB8000092552ABFFEF08517DF6DB6FBE8",
INIT_2A => X"EFA8241516DB55A2FFEAB6DEB843DF551C20801C71C5157428FFDB420101C555",
INIT_2B => X"550428412A85082BEDF401D71C0A2DBC7EB80000280824ADBD7490E28BEF087F",
INIT_2C => X"51504005D71F8E004975D556DB68405092087FF8E00BE8A02082005F47145085",
INIT_2D => X"57BD75EFF78000000000000000000000000000000000000000000000E2AB7D00",
INIT_2E => X"55557DE00A2801554555557FE100055554BA5504000105D2A80145AA842AA005",
INIT_2F => X"5AAD557410F7D57DF55AAFBD55450055420BA0055574BAF7D17DFFFAAFFC2000",
INIT_30 => X"FF08517FFFFF7FBEAB455D517FE00082EBDF45AA8428A10085568ABAA2FBD754",
INIT_31 => X"4AAFFFFC00105D55554BAA28400000F784020BAAAD57FFEFA28402010552ABDF",
INIT_32 => X"FF55002AA8BEF007FFDE1000557DF45AAFBE8BEFA2803FF45550400155555155",
INIT_33 => X"80000087BD55450855400BA002A95400F7FBC01555D2EBFF55A284000AA08003",
INIT_34 => X"000000002EAABFF0051400105D5568A000051575FFF78415410087FEAA10F7AE",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000060000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(15),        -- Port A data input
DOA(0)   => data_read_a_hi(15),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(15),        -- Port B data input
DOB(0)   => data_read_b_hi(15),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_16_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"DA22C618B1000482B688B186588884862A400438255FC38381441205BA803003",
INIT_01 => X"264AC80028404C211203A952A90341080B173340412000E1005D628000820484",
INIT_02 => X"400034C206C405000001A48202084004003008255040826EE008B440200E2042",
INIT_03 => X"2916704900606AC82B49CC56DF8CC1E50E4800202115005760010010000C0400",
INIT_04 => X"052DCA856DC7504B82BF6614C86D2B7F85AAD17F4B100000B88148C4804A428A",
INIT_05 => X"373CB02A00C0502F301180141A42A5720E0F43C17A8479580001AC20000000E2",
INIT_06 => X"303E2094282B85242C85001038D5710E8410D5959BC4800015001219D0550077",
INIT_07 => X"880100000159954501280B0080146F7112D949A0015018220540000382805001",
INIT_08 => X"30015452880C8D90409A05B2CB2CA400200209E5601044A24000000462A60018",
INIT_09 => X"452D54000C0907000330000000000096480050000685400005FC014743E0DC92",
INIT_0A => X"00014808A02004200E540480212000A448C0080024AEA00C9688000000000005",
INIT_0B => X"000D58460018F6D3D84400044000440004400044000440004400042000220002",
INIT_0C => X"0001004010A8812831605DA0000A054052E40000817680220040025699200002",
INIT_0D => X"AAADA0C343F1AC1B01040A002024895514554485D00000012400240000000000",
INIT_0E => X"AAADA0CC421CA003B694B68018FAAA708E2CB5320018CAC99BA0A3B9320018CA",
INIT_0F => X"B1443A1891E4A928C29020E6A8524CE7A3EE59320018CAC99BA0ACB9320018CA",
INIT_10 => X"04B2A5A40B1E6644AF0F021EA003AC24352AB2449A3FF2FA04E5E09B128834AD",
INIT_11 => X"60ED838E890B703C6260D8E3A21275714C902375B801324301AB0067622E5E54",
INIT_12 => X"064F70DBDB1C74424E91E1C194C71D1216F50A8C241815FEB6A9158863F638FB",
INIT_13 => X"45FDF9D364DBD9435A6D45C9E81BED555E4C15F11133D171727A2550EE2F1BA0",
INIT_14 => X"08150013F162119014204373517700ACCC59432A2B2D001F803471A9A960E572",
INIT_15 => X"000000000000000000000000000000880002054000229088542210206B2AB015",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"2A898D21B4C98389ED146C080000000000000000000000000000000000000000",
INIT_19 => X"A29A29A29A29A29A29A29A29A29A28A28A28A28A28A53CBF0F0D3CF3CF0AB1A2",
INIT_1A => X"8F47A3D1E8F4FA7D3E9F4FA7D3E9F4FA7D3E8F4FA3D3E8F4FA3D3E9A29A29A29",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000FA7D3E9F4FA7D1E8F47A3D1E",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFF7FBE8B45AAD568BFFFFAA975FF00003FE0055000000000000000000000000",
INIT_1F => X"0005D2A95410FFFFC00000804154AA5D00001EFF78428AAA007BC2145F7843FF",
INIT_20 => X"7400007BEAAAAAAAE955555D5568A105D2E974BAF7FBEAB45FFFFC00BAF78002",
INIT_21 => X"C2000F78000010552E800AA002E821FFA2AAAAA00000417555FFD17DF45AAD15",
INIT_22 => X"43FEBA5D55575FFF7AABFE00557BD74AAAAD17DF45F7D1421EF0055400AA007F",
INIT_23 => X"D56AAAA5D043FFFFAAAABDEAA557BFDE00FFD140155F7AABDF55F7AE820AA080",
INIT_24 => X"8517DF55A2FBEAB555D04154BAA2FBE8B55FFFFD55FF557FC2000FF8015410FF",
INIT_25 => X"000000000000000000000000000000000000007FFDF45FF84000BA552ABDFEF0",
INIT_26 => X"21C7BC516DFF8438FC7E3F1EAB55B6DF6DBFFF7AA955C71C043FE10490000000",
INIT_27 => X"55FFF1C70BAF78A000005D2097438FFF1C7038140012482550E021C7EB8028A8",
INIT_28 => X"57DEBD17FF6DAADB504001C71EDA82AAA0955455D556DA00492490492F7FBE8B",
INIT_29 => X"71C70851400BA0071C5028FF84020285D2085092002A801FFB6AAA8A10080E17",
INIT_2A => X"BAF6DE3AA8709208043FEBA555B555FFE3AABFE005D71D5492BED17FF45E3DF4",
INIT_2B => X"BC0028E38412428EBD16DA82410A3FFD7AAA4B8E824971F8E38E3DF45155EBA4",
INIT_2C => X"8000092552ABFFEF08517DF6DB6FBE8B555D04124BAB6FBE8B45E3FBD55D7557",
INIT_2D => X"5003DE000000000000000000000000000000000000000000000000071FFF7DEB",
INIT_2E => X"5D2A80145AA842AA00557BD75EFF78428B55AAD168B55F7FFFDFEFFFAA955555",
INIT_2F => X"0000000010F7FBEAB45FFD1554AAFFAE820105500154AAF7D5554BA550400010",
INIT_30 => X"EFF7AEA8A10002E955FFA2D17DFFFAAFFC200055557DE00A2801554555557FE1",
INIT_31 => X"410F7D57DF55AAFBD55450055420BA0055574BAF784000BA5D0017410082E801",
INIT_32 => X"8ABAA2FBD7545AA802ABEFA2AA9541000003DEBA557BD75EFA2AEBDE105D5557",
INIT_33 => X"EAB45AAFFD55555D7FC20AAA280000AAAAD17FE00082EBDF45AA8428A1008556",
INIT_34 => X"00000000557FFEFA28402010552ABDFFF08517FFFFF7FBEAB455D04020AAFFFB",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000020000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(16),        -- Port A data input
DOA(0)   => data_read_a_hi(16),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(16),        -- Port B data input
DOB(0)   => data_read_b_hi(16),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_17_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"5284CE4FB7BD2C8994A13392DBD02E14006B82AC7E800D44D3DD2FD5F9B961C0",
INIT_01 => X"F9BA301F7E03FC6793F2199B39FC233C11D93AE6F3BB92B32091DBC339B24542",
INIT_02 => X"1D5FC0C08F040404446965C0607FB8A217C400C33A908078551BD04222186338",
INIT_03 => X"A14124C28DFD960832C90446DF8400A5055C25295B695FF97E1B5AC757F06D6B",
INIT_04 => X"04A106866DA3D02A01FB660C08A4AB7F840EDB6F48100DFC8081081D78AC7402",
INIT_05 => X"51E072F0C0C58D9C125EBFC00A46CF0388054100F680E0CE0107B8D040DAFCDA",
INIT_06 => X"019A4D00786B048112C58B16307F15DE8408B233661C10BBA5DAAFA9DDA1194D",
INIT_07 => X"8E00001660700CE170284A00891C7C03D29DE26814515835902AC089A2801540",
INIT_08 => X"C009F3A1B0120A1C51DFF881861CBE0305A12A0321810217C01D34EDC98FFA1C",
INIT_09 => X"747E6610052CDEE97FF1F9F63E3EF790380078002CE976AB6BF769769E4D437D",
INIT_0A => X"00185C44B91BC1740B7605040BE0018CFC7429F326B9D045FF8000E9AB415606",
INIT_0B => X"3A28FC1AAF5CF6F3D3EF3D3EF3D3EF3D3EF3D3EF3D3EF3D3EF3D3EF9E9F79E9E",
INIT_0C => X"0000020012E9E10A31EB5FF9296A67F5B4FFBD2FAD7FE653C3FBFF33E10C001B",
INIT_0D => X"333EA16031F2BD47BDA2CA5D8164FCCFE833C5C3D00018006C68170000000000",
INIT_0E => X"333EA160391BEFF2C32FB695F919110D5ECE542A6FEEB2533EA160782A6FEEB2",
INIT_0F => X"D18C0D06638A207CFDE1F7DDAD76D5282400F82A6FEEB2533EA160782A6FEEB2",
INIT_10 => X"E6E43E59AFE4A59B57679D19EFF2C7573FAD5A86840354D1706FFFA3EF6E24B6",
INIT_11 => X"F7D7A0ABD6DAAAB96529382B74E4E1FE4ACA4D77FAAB77CE3AF3EE78F58DB737",
INIT_12 => X"2D1281017F056E9C9C3FC95949C157ADB55572CA52606DFED6CA55334C04C04F",
INIT_13 => X"59FDEB974F486905001FDF5FA0D719F9956EAA1A184045D5D7A870D2F5A5D752",
INIT_14 => X"60158015177F916A039EF41FDB34A91F432EA58949D5B5C85F97871876F7D7E8",
INIT_15 => X"000000000000000000000000000004DC200005E705B7B3D9FC22F00BE419FB55",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"06013DB9880A5D22E229F3030018000000000000000000000000000000000000",
INIT_19 => X"D35D74D35D74D34D35D74D35D74D34D34D34D34D34D0D30D0D303AEBAE886E40",
INIT_1A => X"51A8D46A351A0D068341A0D068341A0D068341A8D468341A8D46834D35D74D34",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000008D46A351A8D46A351A8D46A3",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFF7FBFDF55A28402000F7D56ABFF55000000000000000000000000",
INIT_1F => X"A00F7843FEBA55043FFFFF7FBE8B45AAD568BFFFFAA975FF00003FE0055043FF",
INIT_20 => X"54AA5D00001EFF78428AAA007BC2145F7D568B45000002010552EBDF45A28028",
INIT_21 => X"95410FFAE800105D2A95410002A95410AAAEBFF55AAFFC00BAF7FFC000008041",
INIT_22 => X"57DE00F7AE800AAAAAABDFEF5D2E974BAF7FBEAB45FFFFC00BAF780020005D2A",
INIT_23 => X"517DF45AAD157400007BEAAAAAAAE955555D5568A105D7FFFFEFA2D568BFFFFD",
INIT_24 => X"2AAAAA00000417555FF8028B55082A974105D003FF55F7802AAAAAAD168AAA5D",
INIT_25 => X"000000000000000000000000000000000000000000010552E800AA002E821FFA",
INIT_26 => X"71C043FE10490A3FFFFFFFFFDFEFE3F5FAF45AA8000038F7DB6FBD7490000000",
INIT_27 => X"384124BFF7DB68A28A38F7803DE82490438FC7E3F1EAB55B6DF6DBFFF7AA955C",
INIT_28 => X"0BAFFF1C7038140012482550E021C7EB8028A821C7BC516DFFDF68B551C0E050",
INIT_29 => X"70BAF78A000005D2097438FFAA85000492495428082E95400AAA0BDF7DB6F5C7",
INIT_2A => X"FAFFFB6D56FBFFEBDB78E38F7AA800BAB6AEBDFD75D2490492F7FBE8B55FFF1C",
INIT_2B => X"028AAAB6D16FA8249517FF6DAADB504001C71EDA82AAA0955455D556DA00497F",
INIT_2C => X"2085092002A801FFB6AAA8A10080E1757DEB8A2DB5514249243841003FF6DEB8",
INIT_2D => X"7FFFDF550000000000000000000000000000000000000000000000004020285D",
INIT_2E => X"F7FFFDFEFFFAA9555555003DE00002ABFFEFF7FBFDFFFAAD168B55AA80000BAF",
INIT_2F => X"FF7FBEAB45552E954BA08003DFFFFFAAA8AAAF7843FE10000428B55AAD168B55",
INIT_30 => X"10AA843FFFFF7D5554BAF7D5554BA5504000105D2A80145AA842AA00557BD75E",
INIT_31 => X"010F7FBEAB45FFD1554AAFFAE820105500154AAF7AE974000800154AA002E954",
INIT_32 => X"554555557FE10007FEABEFFFD57FFEFAAFFE8ABAFFAA820BAF7AEBFF55550000",
INIT_33 => X"020AA08003DFFFA28028AAAF7D17DE0000517DFFFAAFFC200055557DE00A2801",
INIT_34 => X"0000000004000BA5D0017410082E801EFF7AEA8A10002E955FFA2AABFF455500",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000067FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(17),        -- Port A data input
DOA(0)   => data_read_a_hi(17),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(17),        -- Port B data input
DOB(0)   => data_read_b_hi(17),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_18_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"69844019080000A21A611406840014122A641074155FC28A2024001001801003",
INIT_01 => X"01067920034004180005E9E3C90360C0041C0181002001602025800008440084",
INIT_02 => X"40AC3CAA22D605200000856E2481902400344A20F802C22054001000021E2379",
INIT_03 => X"A95308ECD3207AC81D91C4002004C08A06008080BA868007E58040102B0E0100",
INIT_04 => X"044CC183800CA00780808004C8DB841405A80A100B586200FAC24AE4805242CA",
INIT_05 => X"771C10000000000B1135883C08A115320E0401C0200038394230070A19000020",
INIT_06 => X"3001499C602A8A003E800A042D8132A00098408F79E3901218050018024110D6",
INIT_07 => X"5029401000C983E60004010030400353C05806800104004E0000042E52800E20",
INIT_08 => X"0000117088080990419005B0C309402030060860E01004A828408800440405E3",
INIT_09 => X"6B8186185C42900693A002004040001E1950850C848601008708114A2030B480",
INIT_0A => X"100180A8062026000DC425C0301311324AA237108857220BA089420440000030",
INIT_0B => X"C44703657083080C2800C2000C2000C2000C2000C2000C2000C2000610006100",
INIT_0C => X"C1B0609C05013065CC042004040808084001E000108010230400800FD9B286C4",
INIT_0D => X"CCC15F9CBA45505640000A402019003F140FC2060014250B9080008306C18360",
INIT_0E => X"CCC15F9FB1962FCB69E08AAAEAEBCDDF7C728582081483ACC15F9C3982081483",
INIT_0F => X"EBF1CFFF7670ACC3811A28AB57523CDFEBFBF982081483ACC15F9F3982081483",
INIT_10 => X"C9002BF05800D875E63CC9962FCB52CAA02FE3F8E7F5E3AC3620805298B15A3F",
INIT_11 => X"F1B72A8A800B7546DB9F1CA320037F01BD67DC4041D4CF03138DD865103EFEEA",
INIT_12 => X"81CCFAFDBF9464006FD037AEFAE5150016EA8DB7BFE25208E8F46A228BF8A757",
INIT_13 => X"641256EC844B8AF92FD7CEDC24A9E181A8A29509EAAE7FD3B749471C48F8A459",
INIT_14 => X"0297D086E00036D2440E0880AAD62BEFF5778802A3AF8E8FB0440CE78773B709",
INIT_15 => X"8360D8360D8360D8360D8360D83609220D20D00000080C0601400B402307E480",
INIT_16 => X"360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D",
INIT_17 => X"60D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8",
INIT_18 => X"D9D701DC2E784601EFBE2C00000000000000000000000008360D8360D8360D83",
INIT_19 => X"5155555545145145155555545145145145145145145220B22A0B820820965177",
INIT_1A => X"44A25128944A25128944A25128944A25128944AA552A954A2512895554514514",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000025128944A25128944A251289",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFEFF7AE954BA5D04174AA00000000000000000000000000",
INIT_1F => X"145AA801741000043FFFFFFFFFFFFFF7FBFDF55A28402000F7D56ABFF55043FF",
INIT_20 => X"8B45AAD568BFFFFAA975FF00003FE0055043FFFFFFFFFDFEFA2D56AB45AA8400",
INIT_21 => X"3FEBA55557FFEFA2D168B55AAFBFFFFFFF80021EF0855421EF00043FFFFF7FBE",
INIT_22 => X"A82155F7AEBFEBAFFD56AA00A2D568B45000002010552EBDF45A28028A00F784",
INIT_23 => X"FFC00000804154AA5D00001EFF78428AAA007BC2145F7D5400000004020AA5D2",
INIT_24 => X"AAEBFF55AAFFC00BAF7AE80010082E954BA0004174AAAA8428B45082ABFEBAA2",
INIT_25 => X"000000000000000000000000000000000000002E800105D2A95410002A95410A",
INIT_26 => X"8F7DB6FBD7490E3FFFFFFFFFFFFFFFFBFDFEFFFAE954AA550415492140000000",
INIT_27 => X"D7AAD16FB6DBE8E00155BE8015410140A3FFFFFFFFFDFEFE3F5FAF45AA800003",
INIT_28 => X"1C7140438FC7E3F1EAB55B6DF6DBFFF7AA955C71C043FE1049043FFEFE3F1F8F",
INIT_29 => X"FF7DB68A28A38F7803DE82495B78FC7AAD56FB6DBEF1FAFD7E384001EF145B47",
INIT_2A => X"420381C0A02082492A85155E3A4BDE92FFD56FA28B6DF68B551C0E050384124B",
INIT_2B => X"E28B7D1420BDEAAA2F1C7038140012482550E021C7EB8028A821C7BC516DFFD1",
INIT_2C => X"2495428082E95400AAA0BDF7DB6F5C70BAFFAE870280024904BA1400174AABE8",
INIT_2D => X"50415410550000000000000000000000000000000000000000000002A8500049",
INIT_2E => X"AAD168B55AA80000BAF7FFFDF55002ABFFFFFFFFFFFEFF7FBFDFFFF7AA974BA5",
INIT_2F => X"000043DFEFA2D56AB45AAD57DFEFF7AA82155F78015400552ABFFEFF7FBFDFFF",
INIT_30 => X"55A280021EF557FD7555550428B55AAD168B55F7FFFDFEFFFAA9555555003DE0",
INIT_31 => X"B45552E954BA08003DFFFFFAAA8AAAF7843FE10007FEAB55A2D17FFEFFFD568B",
INIT_32 => X"AA00557BD75EFF7D1400AA5D2A82000002A95545A2843FE00F7D17FEAAF7FBEA",
INIT_33 => X"020AA5D04154BAF7AEA8BEF55003DEAAA2D5554BA5504000105D2A80145AA842",
INIT_34 => X"000000002E974000800154AA002E95410AA843FFFFF7D5554BAF7AE974BA0004",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000020000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(18),        -- Port A data input
DOA(0)   => data_read_a_hi(18),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(18),        -- Port B data input
DOB(0)   => data_read_b_hi(18),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_19_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"042200000000000041088001001AA00000000000000000000000500802000003",
INIT_01 => X"074018000024000000000404000000000A22000800000800004A200000000001",
INIT_02 => X"0000048002C405000000000006A84000000000200893C246A20000000020031A",
INIT_03 => X"020A9639044012C80001C4000004C08006000000001025000000000000000000",
INIT_04 => X"0400C0800000000380800004C8000000058800000B1000009880480480024200",
INIT_05 => X"420410000000000B10804004080001320E0401C0200038080000000000000000",
INIT_06 => X"2002409006F00A8428050A000280493104004500480090080A01120220140020",
INIT_07 => X"0000000000418026090240923240002190400000000000C0054A912054004021",
INIT_08 => X"0000115080000990000000B0C308000000000860200160000000000038380000",
INIT_09 => X"8000F80001012590001000000000001618000000020280008180810200000000",
INIT_0A => X"0000000000000000000000000000000100008000110000000000000000000017",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000840007600000000000000000800259000000",
INIT_0D => X"0008A0034078104B41A41000000000031400C002000000000000000000000000",
INIT_0E => X"0008A0004263C0343EDD414004042228DC0D385598035D0008A003B05598035D",
INIT_0F => X"040231068187C39F5A4F985C008902041124505598035D0008A000B05598035D",
INIT_10 => X"1BFBD406451B02000E033263C0343CB740500401180DE053A98F6ECC739D8140",
INIT_11 => X"420851546B2400000040D8549B5800000010227848D4303807FC8CC5508AEAED",
INIT_12 => X"52210402120A936B0000000004C2A8D6480000000018A700FCF980CC300318A2",
INIT_13 => X"B1427ED430B41402D025082359700181C21140E40511802208D6B30C48F8A8A4",
INIT_14 => X"9C000018440021011821B35254E99AF9E9410006362A2B6424287B08286208D6",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000023006000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"7747E18E0218CC18E88324000000000000000000000000000000000000000000",
INIT_19 => X"34C30C30C30C30D34C30C30C30C30C30C30C30C30C3504118982A69A6980E411",
INIT_1A => X"C26130984C26130984C26130984C261309A4D26130984C26130984C30C30C30D",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000130984C26130984C26130984",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAA954BA5500020BA5D000000000000000000000000",
INIT_1F => X"4BA5D517FFFF08043FFFFFFFFFFFFFFFFFFFFEFF7AE954BA5D04174AA007BFFF",
INIT_20 => X"FFFFF7FBFDF55A28402000F7D56ABFF557BFFFFFFFFFFFFFFFFFBFDFEFFFAA97",
INIT_21 => X"17410007BFFFFFFFFFFFFEFF7D16AB45AA8002000F7D5575455D043FFFFFFFFF",
INIT_22 => X"568B55F7AE955FFAA840201008043FFFFFFFFFDFEFA2D56AB45AA8400145AA80",
INIT_23 => X"043FFFFF7FBE8B45AAD568BFFFFAA975FF00003FE00557BFFFFFFFFBFDF45AAD",
INIT_24 => X"F80021EF0855421EF002ABFFEFF7D168B55AAD17FFEFF7AE975FF00557FFFF5D",
INIT_25 => X"00000000000000000000000000000000000000557FFEFA2D168B55AAFBFFFFFF",
INIT_26 => X"A5504154921471FFFFFFFFFFFFFFFFFFFFFFFF7AA954BA550000082550000000",
INIT_27 => X"EFF7FBFAFD7E3A4954BA555B7AFC7080E3FFFFFFFFFFFFFFFFBFDFEFFFAE954A",
INIT_28 => X"545550A3FFFFFFFFFDFEFE3F5FAF45AA8000038F7DB6FBD74975FFFFFFFFFFFF",
INIT_29 => X"FB6DBE8E00155BE8015410147FFFFFFF7FBF8FC7EBD568B55A28000000FFDF52",
INIT_2A => X"FDFC7E3F1FAF55A2DB6FB7DF7AE955C7BE800000008043FFEFE3F1F8FD7AAD16",
INIT_2B => X"0955FF145B7AFC7410438FC7E3F1EAB55B6DF6DBFFF7AA955C71C043FE10497B",
INIT_2C => X"D56FB6DBEF1FAFD7E384001EF145B471C71424B8FC7E3D56AB6DB6DF7AFC7EBA",
INIT_2D => X"50002000550000000000000000000000000000000000000000000005B78FC7AA",
INIT_2E => X"F7FBFDFFFF7AA974BA55041541055517FFFFFFFFFFFFFFFFFFFFEFF7AA974AA5",
INIT_2F => X"500517FFFFFFFBFDFEFFFFFEAB45AA80154AA557BEAB45002ABFFFFFFFFFFFEF",
INIT_30 => X"55A28002000F7FFC2155552ABFFEFF7FBFDFFFAAD168B55AA80000BAF7FFFDF5",
INIT_31 => X"FEFA2D56AB45AAD57DFEFF7AA82155F78015400557BFDFEFF7FBEAB55A2D56AB",
INIT_32 => X"555555003DE00007FFDF45AAD568B45AAFBFFFFFFFAA95545F7840201000043D",
INIT_33 => X"6ABFFFFFBEAB45A280155EF557FE8B55000428B55AAD168B55F7FFFDFEFFFAA9",
INIT_34 => X"000000007FEAB55A2D17FFEFFFD568B55A280021EF557FD755555042AB55AAD1",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000040000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(19),        -- Port A data input
DOA(0)   => data_read_a_hi(19),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(19),        -- Port B data input
DOB(0)   => data_read_b_hi(19),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_20_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000003",
INIT_01 => X"A65FF80000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000048002CC070000000000000000000000002FF86100200000000220002362",
INIT_03 => X"00000000000203D80025DC18004DC3D01E000000000000000000000000000000",
INIT_04 => X"07E5DF808071026F87C4191DD8005080679800000F300002998058068002C000",
INIT_05 => X"C205F23A2100557F70000004390021F61E1E87C3FD0CFBF80880072042000044",
INIT_06 => X"1209244C2000100006800000020010000008407FC800B0000000100600040000",
INIT_07 => X"8802000009FFBFE51886018002040020000800000554003E0000000002800000",
INIT_08 => X"30801F5780259FB0000000F7DF78020004011FEFE00000000020031502000083",
INIT_09 => X"00000000001000000000000000000056F8000001000000040000040141800802",
INIT_0A => X"0000000000000008000800000000000000000000000000000010010014800000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"00010240001721214E000004000000080000008000001000040080FFDB000000",
INIT_0D => X"0000000F3008001E00000000001803FF14FFC006000000008010200000000000",
INIT_0E => X"0000000F3040200000020000000026A70C0008020000200000000F3002000020",
INIT_0F => X"000030B86000400080000200000000004A58F0020000200000000F3002000020",
INIT_10 => X"0000000002183E61E6000040200001000000000019B140000800800000020000",
INIT_11 => X"C00010080000000000525801000000000014AC08000000508001030A0A400100",
INIT_12 => X"000002BC360020000000000292C0100000000000A56000090100000000001F86",
INIT_13 => X"8010000000000000574500001001060600000000001716800000803102020000",
INIT_14 => X"00000000000040040040002000080506049CDF70C08040100000706707600000",
INIT_15 => X"00000000000000000000000000802040200200604040000000000024FB7FE008",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"060070400020112240209A408004000000000000000000000000000000000000",
INIT_19 => X"65965965965965965965965965965861861861861860D30424343CF3CF340E00",
INIT_1A => X"90C86432190C86432190C86432190C86432190C86432190C8643219659659659",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000086432190C86432190C864321",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974AA55040201008000000000000000000000000",
INIT_1F => X"4AA550002000007BFFFFFFFFFFFFFFFFFFFFFFFFFAA954BA5500020BA5D7FFFF",
INIT_20 => X"FFFFFFFFFFFEFF7AE954BA5D04174AA00003FFFFFFFFFFFFFFFFFFFFFFF7AA97",
INIT_21 => X"7FFFF087FFFFFFFFFFFFFFFFFFFFDFEFFFAE974AA5D003FE005D043FFFFFFFFF",
INIT_22 => X"BFDFFFAA84000105D556AB55557BFFFFFFFFFFFFFFFFFBFDFEFFFAA974BA5D51",
INIT_23 => X"043FFFFFFFFFFFFFF7FBFDF55A28402000F7D56ABFF55003FFFFFFFFFFFFFF7F",
INIT_24 => X"A8002000F7D5575455D2EBFFFFFFFFFFFEFF7FBEAB55A28000010F7D16ABEF08",
INIT_25 => X"000000000000000000000000000000000000007BFFFFFFFFFFFFEFF7D16AB45A",
INIT_26 => X"A550000082557FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550400028000000000",
INIT_27 => X"FFFFFFFDFEFF7AE974BA5500050380071FFFFFFFFFFFFFFFFFFFFFFFF7AA954B",
INIT_28 => X"E285D0E3FFFFFFFFFFFFFFFFBFDFEFFFAE954AA55041549214043FFFFFFFFFFF",
INIT_29 => X"AFD7E3A4954BA555B7AFC70871FFFFFFFFFFFFFFF7FBFDFFFFFAA974BA550038",
INIT_2A => X"3FFFFFFFFFDFEFF7F1FAFC7A28002028555F6FB7D5D75FFFFFFFFFFFFEFF7FBF",
INIT_2B => X"402010FFDB6ABEF140A3FFFFFFFFFDFEFE3F5FAF45AA8000038F7DB6FBD7490E",
INIT_2C => X"FBF8FC7EBD568B55A28000000FFDF525455524BFFFFFFFBFDFC7E3F5E8B45A28",
INIT_2D => X"504000BA080000000000000000000000000000000000000000000007FFFFFFF7",
INIT_2E => X"FFFFFFFEFF7AA974AA550002000557FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5",
INIT_2F => X"055043FFFFFFFFFFFFFF7FBFDFEFFFAE954BA5500174AA08517FFFFFFFFFFFFF",
INIT_30 => X"EFF7AE974AA550028AAA5D2ABFFFFFFFFFFFEFF7FBFDFFFF7AA974BA55041541",
INIT_31 => X"FFFFFFBFDFEFFFFFEAB45AA80154AA557BEAB4500557FFFFFFFFFDFEFF7FFFFF",
INIT_32 => X"00BAF7FFFDF55002EBFFFFF7FBFDFEFFFD568B55A284020BA557FFFFFF5D517F",
INIT_33 => X"FFF55A2D16AB45AA8402000F7FBEABEF5D2ABFFEFF7FBFDFFFAAD168B55AA800",
INIT_34 => X"000000007BFDFEFF7FBEAB55A2D56AB55A28002000F7FFC215555043DFEFF7FB",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000007FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(20),        -- Port A data input
DOA(0)   => data_read_a_hi(20),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(20),        -- Port B data input
DOB(0)   => data_read_b_hi(20),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_21_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"4A302428B824900A128C090A5C1800261500213C005FE812D10420054085A202",
INIT_01 => X"081FFE3440B609703B0427F801A40B8115BC4F655300340288A40D30040E4DD8",
INIT_02 => X"04CA478082CC1740002019824E0203100640303FF8C0B31061096E21A1840814",
INIT_03 => X"230CA7A4810083F80095DE00102DC3823EA821094EC68248923200013290C800",
INIT_04 => X"07CFFFC04904AA7F8780409DF84A0202879800000F3000029980780EA2C3C002",
INIT_05 => X"DE87F0280000407FF900D914382091FE1E1C0FC3E01EFFF8000480200008D062",
INIT_06 => X"010E2182002BC107A03448808F0D7C002822987FC830F40134CC74D002016612",
INIT_07 => X"0401000011FBFFE00520000200422033025C4209104500000012004C004D8C0B",
INIT_08 => X"00EF1F5FA0041FF080AC70FFDF78220010841EFFE7116E144071268DFD3E4C24",
INIT_09 => X"FC8BFE18008083B4443151462A28C6DFF80010002605302248088950484550A3",
INIT_0A => X"10018C241102068006C620C03882019480E631A0855E924E2598038938404037",
INIT_0B => X"A641165448C80C103648A3648A3648A3648A3648A3648A3648A366451B2451B2",
INIT_0C => X"011100841200D001000624000100C002804A08221890004806A310FFDF000454",
INIT_0D => X"5004D8158809C86065941840B1014FFF56FFC0281280080180B2948004400220",
INIT_0E => X"5004D815810D42E04A08A80098C02450025360694101816002D41A4068C10181",
INIT_0F => X"134160C8125B0B271802242880A04482418A0068C101816002D41A4069410181",
INIT_10 => X"10080E05C0B06AA8B12CFD0D42E0441A300012682960828F05C96A001B029010",
INIT_11 => X"00010362A8A20826A88660D86B202049F115100920C54E8EA256ECF078BA081C",
INIT_12 => X"064802C0081B0D64040936443306C55144104F30A8801406D002900062803201",
INIT_13 => X"4581BA0038005A706680012280506A8010602011819E290048A2118EC8140C08",
INIT_14 => X"CC158092C044600466208CC5091011C322A4C40A0300600C0A80509F41800880",
INIT_15 => X"80200802008020080200802008020412002001000000381C02004000FBFFF80D",
INIT_16 => X"0200802008020080200802008020080200802008020080200802008020080200",
INIT_17 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_18 => X"FDDFEFFFBEFFE7C7BFBEFC000000000000000000000000080200802008020080",
INIT_19 => X"F7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7FFBFBFFF9E79E7FFFDF3",
INIT_1A => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFDFEFF7FBFDFEFF7FBFDF7DF7DF7D",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00001FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D000200008000000000000000000000000",
INIT_1F => X"4AA5D00020AA5D7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550402010087FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAA954BA5500020BA5D7FFFFFFFFFFFFFFFFFFFFFFFFFFAE95",
INIT_21 => X"0200000003FFFFFFFFFFFFFFFFFFFFFFF7AA974BA5D0402000557BFFFFFFFFFF",
INIT_22 => X"FFFFEFF7AE974BA5D00174BA00003FFFFFFFFFFFFFFFFFFFFFFF7AA974AA5500",
INIT_23 => X"043FFFFFFFFFFFFFFFFFFFFEFF7AE954BA5D04174AA00003FFFFFFFFFFFFFFFF",
INIT_24 => X"FAE974AA5D003FE005D2EBFFFFFFFFFFFFFFFFFFDFEFF7AE954AA5500174BA5D",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFDFEFF",
INIT_26 => X"A550400028007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0000010000000000",
INIT_27 => X"FFFFFFFFFFFFFAA954BA5D00000BA557FFFFFFFFFFFFFFFFFFFFFFFFFFAE974A",
INIT_28 => X"0005571FFFFFFFFFFFFFFFFFFFFFFFF7AA954BA550000082557BFFFFFFFFFFFF",
INIT_29 => X"DFEFF7AE974BA55000503800003FFFFFFFFFFFFFFFFFFFFEFF7AA974AA5D0405",
INIT_2A => X"3FFFFFFFFFFFFFFFFFFDFEFF7AE954BA5D00154AA00043FFFFFFFFFFFFFFFFFF",
INIT_2B => X"A974BA5D00104925D0E3FFFFFFFFFFFFFFFFBFDFEFFFAE954AA550415492140E",
INIT_2C => X"FFFFFFFF7FBFDFFFFFAA974BA550038E285D2ABFFFFFFFFFFFFFFFFBFDFEFFFA",
INIT_2D => X"D00000100000000000000000000000000000000000000000000000071FFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE954AA5504000BA087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0557BFFFFFFFFFFFFFFFFFFFFFFFF7AA954BA5D00000BA5D7FFFFFFFFFFFFFFF",
INIT_30 => X"EFF7AE954AA5D041740055517FFFFFFFFFFFFFFFFFFFFEFF7AA974AA55000200",
INIT_31 => X"FFFFFFFFFFFFF7FBFDFEFFFAE954BA5500174AA08043FFFFFFFFFFFFFFFFBFDF",
INIT_32 => X"74BA550415410552ABFFFFFFFFFFFFFF7FBFDFFFFFAA974AA5D00174BA08043F",
INIT_33 => X"FDFEFF7FBFFFFFF7AE954BA5D0000010552ABFFFFFFFFFFFEFF7FBFDFFFF7AA9",
INIT_34 => X"00000000557FFFFFFFFFDFEFF7FFFFFEFF7AE974AA550028AAA5D2EBFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(21),        -- Port A data input
DOA(0)   => data_read_a_hi(21),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(21),        -- Port B data input
DOB(0)   => data_read_b_hi(21),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_22_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"5290F4CDE914905A14A43D33F488243E17122300F55FEB189B343A1140548380",
INIT_01 => X"A94007B259F6A975386262000C344BA9573C6FF57B18A5FB0ABFCD3C2C5F4F0C",
INIT_02 => X"D56B4302AC01005111011BD506AA5205274056900596A539584E2E6DFE4B2418",
INIT_03 => X"9AC0FCBD854688207C90007A1000047A00E588632CA213C8903AD6B55AD0EB5A",
INIT_04 => X"30002047A6FCA110086C402022F2124A8022492580040440002021C922D9109B",
INIT_05 => X"14A206B6838151008D95DD1847811C08002380041F1104002205AC4140DAD060",
INIT_06 => X"1727FF2EB9EF113A10BD32F44289D1F840C1710010344DB9A808FDFF3DE03130",
INIT_07 => X"050700154A00401D00495A06A8D464C5F6B54AA8551040818F4C997AC80CBE05",
INIT_08 => X"0141008801018040E48D50080002B00A0C00801014541E9504703680017F6CB4",
INIT_09 => X"02680000010937986481514E2A29CE010708C0804C6A033F7FCFF9426A41F1AB",
INIT_0A => X"00500001840000C80B410014088040F4A944B1AA313C004554002381B8000500",
INIT_0B => X"A004D1594832824A070AA070AA070AA070AA070AA070AA070AA0725503855038",
INIT_0C => X"501428054278142151262CA50343854E506A2C6898B2950AA6A35B0004284058",
INIT_0D => X"90078E1F840A2B0114020104022460002200050F60E220A06880D2A14050A028",
INIT_0E => X"90078E1F891C239F8908003099C1ACF06273612B3482C0C0078E1F412B1582C0",
INIT_0F => X"1BA1B0FD16770236A4091621C08055C2C0DB012B1582C0C0078E1F412B3482C0",
INIT_10 => X"00101F09C030AB28B03C111C239F870828041BA859F213AFC14AA38043006018",
INIT_11 => X"10E8822A984B0025B0DE6089462660095337B08AA600CA88B143AB11880C2806",
INIT_12 => X"055412D4481128C4CC012A66F304553096004B61BD8068B92400D0004E303689",
INIT_13 => X"589C48082C006A9057CA4385809520F07830001AC2173B00E162563454C40804",
INIT_14 => X"00460848952220592745AC11A544B1BF006850840180A00E1C81900C4190E160",
INIT_15 => X"22088220882208822088220882208CD888088D940D2A3A9D5002001300800C8C",
INIT_16 => X"0080200882208822088220882208822088220882208822088220882208822088",
INIT_17 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_18 => X"FBDFD1FE3EFBD7BBEFBEFA0A245120000000007FFFFFFFF20080200802008020",
INIT_19 => X"F3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF7FFBFAFBBBEFBEFBEFBF7",
INIT_1A => X"CFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCF3CF3CF3C",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000007F3F9FCFE7F3F9FCFE7F3F9F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040000000000000000000000000000000",
INIT_1F => X"4BA550000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0002000087FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974AA550402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"020AA5D7FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5D00000AA007FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAA954BA5504000AA557FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5D00",
INIT_23 => X"7BFFFFFFFFFFFFFFFFFFFFFFFFFAA954BA5500020BA5D7FFFFFFFFFFFFFFFFFF",
INIT_24 => X"7AA974BA5D040200055517FFFFFFFFFFFFFFFFFFFFFFFFAA954BA5500000BA5D",
INIT_25 => X"00000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000080000000",
INIT_27 => X"FFFFFFFFFFFFFAE974AA550002010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"0BA087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550400028007FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAA954BA5D00000BA557FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5D0002",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAA954BA5504020AA5D7BFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"A974AA5D00070925D71FFFFFFFFFFFFFFFFFFFFFFFF7AA954BA5500000825571",
INIT_2C => X"FFFFFFFFFFFFFFEFF7AA974AA5D040500055517FFFFFFFFFFFFFFFFFFFFFFF7A",
INIT_2D => X"D040200008000000000000000000000000000000000000000000000003FFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"A087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550002000087FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAA954AA5D00020AA007FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5504000B",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFF7AA954BA5D00000BA5D7BFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"74AA55000200055517FFFFFFFFFFFFFFFFFFFFEFF7AA974BA5504020BA557BFF",
INIT_33 => X"FFFFFFFFFFDFEFF7AE974AA5D00154105D517FFFFFFFFFFFFFFFFFFFFEFF7AA9",
INIT_34 => X"00000000043FFFFFFFFFFFFFFFFBFDFEFF7AE954AA5D041740055557FFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000007FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(22),        -- Port A data input
DOA(0)   => data_read_a_hi(22),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(22),        -- Port B data input
DOB(0)   => data_read_b_hi(22),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_23_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"EF20906D902424807BC8241BC81801B97D38AD3C0800103362A6741C80A12A02",
INIT_01 => X"001FFF8409F089003B4422000D80C80106804A7951C5B9D1C828043EA28838F9",
INIT_02 => X"028406A002DC176444683862400003111001303FFC00F240D50146013B300500",
INIT_03 => X"0006C90C010203F80005DC00C52FC380BEAC25886C02034800200200A1008008",
INIT_04 => X"17DFFF8049000BFF878314BFF8488890979800002F702002BB807A068403C280",
INIT_05 => X"DA07F0000000007FF020C814380011FE5E1C2FC3E05FFFF90020000808900010",
INIT_06 => X"10004C9690A8CA008024685184097E81E872C8FFE900FC31348EFDF03BE15E22",
INIT_07 => X"402000001FFBFFFD00080200B8140011F0D8C108155542018D1A302193E94004",
INIT_08 => X"41BE1F5F80003FF0002023FFDF79000000000EFFE309606020008005FC000000",
INIT_09 => X"FC83FE1840C0902400300000000000DFFD4004040C4D32BF7C0EE860003CE680",
INIT_0A => X"10018C24110A860006C620C0312241C482B20420CC56924E2199000C00415037",
INIT_0B => X"4669070510C90C14304043040430404304043040430404304043040218202182",
INIT_0C => X"008000105400C00400100000A018000801000C024000004A940000FFDF820604",
INIT_0D => X"100152100801C17E61841950B1C10FFF57FFC02812F00429DC92C40002000100",
INIT_0E => X"10015210088528E00E02C8200A430A424202A1CAF13F214001521001CBF03F21",
INIT_0F => X"01C1C044006D0C94FB94320880603C420B8001CBF03F214001521001CAF13F21",
INIT_10 => X"30182800A018D9CA8000648528E00D12480202C86040902AC60BACDF0E02D020",
INIT_11 => X"0445C19960A00026880C006739000009B00300010AF5052419D1964419028014",
INIT_12 => X"01844068880CE72000013600600332C140004D101808458A5602E00089202911",
INIT_13 => X"41D0B9023402085020825132C8CB5B4040301009408021144CB042F880100C06",
INIT_14 => X"8E17C0D240406519400500840A9524EE38A1F80E02120018390320F050144CB2",
INIT_15 => X"01004010040100401004010040100100040040000000000001000900FBFFE000",
INIT_16 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_17 => X"0040100401004010040100401004010040100401004010040100401004010040",
INIT_18 => X"0000000000000000000000000000000000000000000000001004010040100401",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000000000000000000000000",
INIT_1F => X"4BA5D0400010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000007FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974BA5D0002000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"00010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA550002000007FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAE974AA550400000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5500",
INIT_23 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550402010087FFFFFFFFFFFFFFFFFF",
INIT_24 => X"FAE954AA5D00000AA007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA55040200008",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010000000000",
INIT_27 => X"FFFFFFFFFFFFFAE974BA5D0400010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0000010007FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAE974AA550002010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA550002",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550400010087FFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"E954AA5D0402038007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550400028007F",
INIT_2C => X"FFFFFFFFFFFFFFFFFFAE954AA5D00020BA087FFFFFFFFFFFFFFFFFFFFFFFFFFA",
INIT_2D => X"D0402010000000000000000000000000000000000000000000000007FFFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000087FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAE974BA550002010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D000001",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFFFAE974AA550002000087FFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"54AA5504000BA087FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA550400010007FFF",
INIT_33 => X"FFFFFFFFFFFFFFFFAA954AA5D04000AA087FFFFFFFFFFFFFFFFFFFFFFFFFFAE9",
INIT_34 => X"000000007BFFFFFFFFFFFFFFFFFFFFFFFFFAA954AA5D00020AA007BFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000007FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(23),        -- Port A data input
DOA(0)   => data_read_a_hi(23),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(23),        -- Port B data input
DOB(0)   => data_read_b_hi(23),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_24_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100600007FFF000080108004000800020000840041000080808",
INIT_02 => X"0000068002CC07400000090C080002000000103FF811F150231000520ABE4404",
INIT_03 => X"210A0600000203F80005DC00000DC3801EA000000745C4010220000000008000",
INIT_04 => X"07C5FF804900026F8780001DF8000000079800000F300002998078068003C080",
INIT_05 => X"C207F0000000007FF0000004380001FE1E1C07C3E00CFFF80000000000000000",
INIT_06 => X"0002648240F20035A0102000BD0000002802C87FC800FCAA035400001B918600",
INIT_07 => X"0000000001FBFFEC4D2B4AD0B8129063B2CC0000100042018408142F16C01848",
INIT_08 => X"008E1F5F80001FF0000000FFDF78000000000EFFE001600000000005FC000000",
INIT_09 => X"E883FE180000000000300000000000DFFD0000002A80D500000671000004A000",
INIT_0A => X"10018C0411020600048620C030020502000200000400920A2198000800404037",
INIT_0B => X"0641060400C00C00304003040030400304003040030400304003040018200182",
INIT_0C => X"000000001000C00000000000000240058000000000000000000000FFDF000404",
INIT_0D => X"E00880104809C1666594584031010FFF56FFC000104000000010440000000000",
INIT_0E => X"E0088010492064206100E81084200048C0804012500021B00880108012500021",
INIT_0F => X"04100144800803419043064900C0020501840012500021B00880108012500021",
INIT_10 => X"1018140F02C0000809408D206420530270040410004C840041A0D80054109038",
INIT_11 => X"110002C9E8010C00010480B35A0300400041020902F60002260D65B361BAA104",
INIT_12 => X"0228204300166B4060080008240593D0021800020818B06D9802F00030C02060",
INIT_13 => X"143B62023C00142800B04400095DFF90203020042108603100061516EE800C06",
INIT_14 => X"DC1180C7804400044029208301040214AE4C7C02000040206602C10B48110006",
INIT_15 => X"00000000000000000000000000000000000000000000000000000000FBFFE000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"DD5EDCF9822659B6888332000000000000000000000000000000000000000000",
INIT_19 => X"F3CF3CF3CF3CF3DF7DF7DF7DF7DF7DF3DF3DF3DF3DF4D30C2432AEBAEBFE5A15",
INIT_1A => X"C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783DF7DF7DF7C",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000F0783C1E0F0783C1E0F0783",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201008000000000000000000000000",
INIT_1F => X"4BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974BA5D0400000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"00010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000007FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAE974BA5D0000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_23 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0002000087FFFFFFFFFFFFFFFFFF",
INIT_24 => X"FAE974BA550002000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D000200000",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010080000000",
INIT_27 => X"FFFFFFFFFFFFFAE974BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000087FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAE974BA5D0400010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0000010007FFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"E974BA550002000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0000010007F",
INIT_2C => X"FFFFFFFFFFFFFFFFFFAE974BA550002000007FFFFFFFFFFFFFFFFFFFFFFFFFFA",
INIT_2D => X"D0402010080000000000000000000000000000000000000000000007FFFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAE974BA5D0400000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040200",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000087FFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"74BA5D0000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0000010087FFF",
INIT_33 => X"FFFFFFFFFFFFFFFFAE974BA550000010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE9",
INIT_34 => X"000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA550002010087FFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(24),        -- Port A data input
DOA(0)   => data_read_a_hi(24),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(24),        -- Port B data input
DOB(0)   => data_read_b_hi(24),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_25_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100200002000000080100004000000020000800041000080808",
INIT_02 => X"0000068002CC474000000800000002000000103FFCE302008000000880844A04",
INIT_03 => X"00000040700803FC0105DE00020DC3801EA00000040000000020000000008000",
INIT_04 => X"47C5FFC04904026F8780081DFC040000079C92484F30499299837C168003E400",
INIT_05 => X"C207F0382004407FF0000004382281FF1E1C07C3E00CFFFC090004B05000200A",
INIT_06 => X"1009015C4000000020000000390C10002802C87FC800F8000000000019810600",
INIT_07 => X"0501000001FBFFFD480A0280A816002010800001000054018408102000000002",
INIT_08 => X"0C8E1F5FA21C9FF8004000FFDF7C062031863EFFF75D78004001010DFC000020",
INIT_09 => X"E883FE180C00000000300000000000DFFF00180800000000000660100000A000",
INIT_0A => X"1001DCCC31222730A49620C030020100000200000400921A21D8000804404037",
INIT_0B => X"0641062400C00C00304003040030400304003040030400304003040018200182",
INIT_0C => X"C11160845004D04820000000000000000000000000000000940000FFDF000404",
INIT_0D => X"000800000801C0786184185031810FFF56FFC02812E0182000F2C48304418220",
INIT_0E => X"0008000000002020000008000000000800800002400001000800000002400001",
INIT_0F => X"0000010000000000900000080000000400000002400001000800000002400001",
INIT_10 => X"1000000002002000004000002020000200000000000404000000880000001000",
INIT_11 => X"010000082000000001000001080000000040000100C600800001040000040009",
INIT_12 => X"0000000100002100000000080000104000000002000000081001000000000040",
INIT_13 => X"0010200000000000001004000001080000400080000040010000001080001008",
INIT_14 => X"8C11808200400000400000C20000000420000000030280000000010000010000",
INIT_15 => X"82208822088220882208822088A20C52082081A30080000002005008FBFFF001",
INIT_16 => X"2208822088220882208822088220882208822088220882208822088220882208",
INIT_17 => X"2088220882208822088220882208822088220882208822088220882208822088",
INIT_18 => X"29432D518B45265D82BB4101000005FFFFFFFFFFFFFFFFF82208822088220882",
INIT_19 => X"24924924924924820820820820820820924820924824000A6242B4D34D7F7451",
INIT_1A => X"AC562B158AC562B158AC562B158AC562B1188C46231188C46231189249249249",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000162B158AC562B158AC562B158",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000000000000000000000000",
INIT_1F => X"4BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"02000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAE974BA5D0402000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_23 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000007FFFFFFFFFFFFFFFFFF",
INIT_24 => X"FAE974BA5D0400000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040000008",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010000000000",
INIT_27 => X"FFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAE974BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000007FFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"E974BA5D0400000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000087F",
INIT_2C => X"FFFFFFFFFFFFFFFFFFAE974BA5D0400000007FFFFFFFFFFFFFFFFFFFFFFFFFFA",
INIT_2D => X"D0402010000000000000000000000000000000000000000000000007FFFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"74BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000007FFF",
INIT_33 => X"FFFFFFFFFFFFFFFFAE974BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE9",
INIT_34 => X"000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000007FFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000007FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(25),        -- Port A data input
DOA(0)   => data_read_a_hi(25),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(25),        -- Port B data input
DOB(0)   => data_read_b_hi(25),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_26_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"E9264EAB20190CA3BA4997AA9002AE9C001006B0778015CFA17E0811039879C7",
INIT_01 => X"F1FFF9BB1F773C7F9BB07DFFFDD863FC5FFF3FEFFBBF9FFB22FFFBC7B9F30686",
INIT_02 => X"9B3184F8AFDEAF300029E4E300FC78A6258548EFFA71C00172082400003A2161",
INIT_03 => X"0084F0FF7FFF1FDD3FEFDCDE981DC3FF5F0D294A7B2B18A0001B9CE6CC606E73",
INIT_04 => X"0FC5DFD7EDFFD66F87FE605DDDBFF3690F9EDB7F5F7AFF639BD7DE37C2FEF591",
INIT_05 => X"F205F0F8E9D199FF76DFEE1C3FCC3FF7BE1FD7C3FFACFBFFDFF7B4FEFFDAA10E",
INIT_06 => X"042648C40179912406C1830639AFBEC14489737FDC00B13BB79DFDB83BF4112A",
INIT_07 => X"763A844769FFBFE4398E4390BB9C28B1D0F049080414583F9468D1AEFC000060",
INIT_08 => X"02C05FD7BC471FBD13D981F7DF7D7E6171AF3FEFE8A3E679FAC1FD1FFFBEB000",
INIT_09 => X"F8CFFE38FF7F6BD928F1ABB47476B5FEF9F59F5FCEEDE73FEE0EFC53B079F5CC",
INIT_0A => X"315BDDCC3B336F7C548667D47B7737AF3FD62601EDC2B66A67B9D60FE4C4427F",
INIT_0B => X"06E19F4DA0E80E903DE3035E3035E3035E3035E3035E3035E3035E981AF181AE",
INIT_0C => X"EBFBF7FEBD66DBFCA3F87501AE7B080607307DCFE1D4077B4D026FFFFBFFAFCD",
INIT_0D => X"0007E010084BCD7FF1B61B5C33813FFFFCFFC7D7D51D6F5FDCB935D7AFEBD7F5",
INIT_0E => X"0007E01001BD8020500008001F010040520201F45EC0010007E01001F45EC001",
INIT_0F => X"1DC0004600400F781429C0080000770001A001F45EC0010007E01001F45EC001",
INIT_10 => X"10003C064000E408010081BD8020600200001EC00040B02007EC09A0E0001000",
INIT_11 => X"360403E434588007200D00F88C84C081C203404B3BFD0402346235408402C080",
INIT_12 => X"07B00040091F1190982038406807C868B1000E401A08FE0012040000FC002001",
INIT_13 => X"7D00212000007C400082D81009FC08281D00001F010021560406758091454000",
INIT_14 => X"FFBFF5FA1040076065F730FC08043A903A80008320C0403C3400008860160406",
INIT_15 => X"D7F5FD7F5FD7F5FD7F5FD7F5FDFF7F7F7F77F9F761FFBFDFFDE5BFFFFF7FF005",
INIT_16 => X"7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5F",
INIT_17 => X"F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD",
INIT_18 => X"B79E923C2CD990AA7F0DDB6B910C8DFFFFFFFFFFFFFFFFFD7F5FD7F5FD7F5FD7",
INIT_19 => X"30C30C30C30C30C30C30C30C30C30C30D34D34C30C35F7AA9ABF0E38E3A8EB62",
INIT_1A => X"C26130984C26130984C26130984C26130984C26130984C26130984C30C30C30C",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000130984C26130984C26130984",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000000000000000000000000",
INIT_1F => X"4BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"02010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_23 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFF",
INIT_24 => X"FAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010000000000",
INIT_27 => X"FFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"E974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007F",
INIT_2C => X"FFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFA",
INIT_2D => X"D0402010000000000000000000000000000000000000000000000007FFFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"74BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFF",
INIT_33 => X"FFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE9",
INIT_34 => X"000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(26),        -- Port A data input
DOA(0)   => data_read_a_hi(26),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(26),        -- Port B data input
DOB(0)   => data_read_b_hi(26),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_27_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"00080A40000A41248002029000050A088000008242A0004404480002000A1155",
INIT_01 => X"F1FFF1C11F781C129C107DFFFE0860941E81258CA2B71C2220EC1B86E1A00002",
INIT_02 => X"183080988B2EAE00002BE001117C78C6848140CFFA0000800042008000011081",
INIT_03 => X"000000FF7CF91F1D3DEF3CDA881D23FB5C0C21085B0B0820001318C60C204C63",
INIT_04 => X"8FC51FD7EDFDD66E47EE205D1DB7F1490E5EDB7D5CBADB2385D79C3643D4E580",
INIT_05 => X"E001F0C0C991BBFC76DFEA1A3F8C3BC7391F9723FF2CE3FCD6D13096B79C8106",
INIT_06 => X"40000001000000084041830600A40C415004637FC4003021259CFDB01BF80028",
INIT_07 => X"3158954761FA3FE402088220AC1108001080400A400041018468D1A060000050",
INIT_08 => X"02005F0784411E390A4881C7BEFC5F6171CE2F8FE823E778DAC16C1FFBBC9000",
INIT_09 => X"F0C7FEBABF3F6BD108F40E04C0C084F0F8B58B5B8849673F6C0E7A01B00914C4",
INIT_0A => X"B51BFDCC39732F3554866AD57C37BEAF1C152201A4C0B6EA63AAD60B60D4427F",
INIT_0B => X"06F18FC5A0E00F0038D1030D1030D1030D1030D1030D1030D1030F0818688186",
INIT_0C => X"AB6AD7EAB962CBD8A3A83101F47E08040510768EA0C406630D0226FFE375ADE5",
INIT_0D => X"000760000843C561E5C55C42B9011FFF48FFCC57550D63564D1D2556ADAB56D5",
INIT_0E => X"0007600004BD8020100008001F010000130201E44A40010007600005E44A4001",
INIT_0F => X"1DC0000208400D781020C00800007700002005E44A40010007600005E44A4001",
INIT_10 => X"10003C064000C400018080BD8020200200001EC00000382006EC0820A0001000",
INIT_11 => X"3E0403A424108007200102E888808081C20040431BC504021462354004004080",
INIT_12 => X"07B00000015D1110102038400817484821000E400204FE0010040000FC000000",
INIT_13 => X"7D00202000007C400000F81001FC08080500001F0100005E0404758081014000",
INIT_14 => X"8DBBB5FA10400360649310FC08003A903A8000012040403C34000080201E0404",
INIT_15 => X"56D5B56D5B56D5B56D5B56D5B56D7E3D7B57B1C4E17F0944B8D596EEFC7FF001",
INIT_16 => X"6D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B",
INIT_17 => X"D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B5",
INIT_18 => X"2D0200903950C080420948E2D10E8FFFFFFFFFFFFFFFFFF56D5B56D5B56D5B56",
INIT_19 => X"00000000000000000000000000000104000000000004000E5E420000002921C4",
INIT_1A => X"28140A05028140A05028140A05028140A0100804020100804020100000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000140A05028140A05028140A050",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000000000000000000000000",
INIT_1F => X"4BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_23 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFF",
INIT_24 => X"FAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201008",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010000000000",
INIT_27 => X"FFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"E974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087F",
INIT_2C => X"FFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFA",
INIT_2D => X"D0402010000000000000000000000000000000000000000000000007FFFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"74BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFF",
INIT_33 => X"FFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE9",
INIT_34 => X"000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000007FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(27),        -- Port A data input
DOA(0)   => data_read_a_hi(27),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(27),        -- Port B data input
DOB(0)   => data_read_b_hi(27),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_28_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"02200AA400180030808802A900002A08001280A08A801044104A1000001818C3",
INIT_01 => X"50A00011460214428114180000882214413D0A71592A01D92213D28005210202",
INIT_02 => X"8A54800A210200111100C2110054289220810440030404010844000444410001",
INIT_03 => X"1080010208B51400007800000A000001000108C21008092000018C6295200631",
INIT_04 => X"0008000000017000000028000001610300000010000802202040012040040011",
INIT_05 => X"2000044440048880026A22000026A20000000000000000004994140203000064",
INIT_06 => X"1400922401041008004891224228810080010200040001020800000004000008",
INIT_07 => X"150B001328000001404010040084088404200020455514000224489028492201",
INIT_08 => X"00414000201800004080A0000002480B04008100011000088800081002C19020",
INIT_09 => X"000400001036584108415B4A6A694A0000100101C08200000001000190200044",
INIT_0A => X"004800210C19808400500010009110091500020B408820000200400040811600",
INIT_0B => X"40000800B00100040D8140581405814058140581405814058140580A02C0A02C",
INIT_0C => X"00200248010201008298150006210802043058C46054032981002D00201C8081",
INIT_0D => X"0000A00000400600841041108280300008000140000401028008330000800040",
INIT_0E => X"0000A000000080001000000000000000500000040A40000000A00000040A4000",
INIT_0F => X"00000006000000080020C00000000000012000040A40000000A00000040A4000",
INIT_10 => X"00000000000024000000000080002000000000000000A00000040020A0000000",
INIT_11 => X"2200000404108000000900008080808000024040152000000020000004004080",
INIT_12 => X"0000000009001010102000004800080821000000120002000004000000000001",
INIT_13 => X"2000002000000000000288000020000805000000000001420000200001014000",
INIT_14 => X"408010000000022000D610280000080000000001204000000000000820020000",
INIT_15 => X"00401004010040100401004010042024210218734CD52150A840827504000000",
INIT_16 => X"0401004010040100401004010040100401004010040100401004010040100401",
INIT_17 => X"4010040100401004010040100401004010040100401004010040100401004010",
INIT_18 => X"05822140048D2E57B1348141845C200000000000000000000401004010040100",
INIT_19 => X"04104104104104104104104104104104104104104101A6A0A0EB1861863BC422",
INIT_1A => X"2C160B0582C160B0582C160B0582C160B0180C06030180C06030181041041041",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000160B0582C160B0582C160B058",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000000000000000000000000",
INIT_1F => X"4BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_23 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFF",
INIT_24 => X"FAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010000000000",
INIT_27 => X"FFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"E974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007F",
INIT_2C => X"FFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFA",
INIT_2D => X"D0402010000000000000000000000000000000000000000000000007FFFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"74BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFF",
INIT_33 => X"FFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE9",
INIT_34 => X"000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000007FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(28),        -- Port A data input
DOA(0)   => data_read_a_hi(28),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(28),        -- Port B data input
DOB(0)   => data_read_b_hi(28),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_29_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"79964E4BA01DACAB9E659792D00AAE160002829C7FDFEFCEE97C2815039D70C3",
INIT_01 => X"50BFF9AB0775343F9AB01DF80D5821FC0FFF3FEFD1AF9FF1207FFBC7B9720586",
INIT_02 => X"0D15846807D207200021C4E200D428A2018408600271C000720A0000003A2161",
INIT_03 => X"0000B0027BBF17C43E6DC05E1A0DC07D1F0000803B2819A00019084345606421",
INIT_04 => X"07CDC047A4FB526F807C681DC4B97369078249370F482E62BA414627C2FE3000",
INIT_05 => X"F204007861C088FF0EFF260407C427F19E03C7C01F8CF80749B390EA4BCA202C",
INIT_06 => X"000248C00079800406C081023B233E804488527FDC008019968D74982C94110A",
INIT_07 => X"5229000221FF8000398641903B082831D05000200000083F942850AEB4000221",
INIT_08 => X"00805FD0180E1F8C1111A0F041056A0100A11FE000916249A800B915FE82B020",
INIT_09 => X"F80C000055FF7C492840AAB45456B55E015015058665A31DA603A4539058F54C",
INIT_0A => X"000850400A11414C005005000B51158936D20601A98A204006114005C4800217",
INIT_0B => X"40201948B029029409A3401A3401A3401A3401A3401A3401A3401A9A00D1A00C",
INIT_0C => X"40B1225C1506512C83E85500AC3A080406305587A154023141006DFFF89E82C9",
INIT_0D => X"0000A01008480D3EB4A24A0C910037FFFC0007C7C0140D0B50A8218102C08160",
INIT_0E => X"0000A010010080005000000000000040520000141EC0000000A01000141EC000",
INIT_0F => X"00000046000002080429C0000000000001A000141EC0000000A01000141EC000",
INIT_10 => X"00000000000024080100010080006000000000000040B000010401A0E0000000",
INIT_11 => X"3600004414588000000D00108484C080000340483B590000202000008402C080",
INIT_12 => X"00000040090210909820000068008828B10000001A0802000204000000002001",
INIT_13 => X"20000120000000000082D800082000281D000000000021560002200011454000",
INIT_14 => X"B29450580000066021F6303C000408000000008320C000000000000860160002",
INIT_15 => X"816058160581605816058160589625662522506344FF9FCFFF62EB6DFF001004",
INIT_16 => X"1605816058160581605816058160581605816058160581605816058160581605",
INIT_17 => X"6058160581605816058160581605816058160581605816058160581605816058",
INIT_18 => X"F2DDCFFFBEFFCF07FFBFFD41800C05FFFFFFFFFFFFFFFFF81605816058160581",
INIT_19 => X"7DF7DF7DF7DF7DF7DF7DF7DF7DF7DD75D75D75D75D77FFBF3F7DFFFFFFD779F3",
INIT_1A => X"FEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDF7DF7DF7DF",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00001F7FBFDFEFF7FBFDFEFF7FBFD",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000000000000000000000000",
INIT_1F => X"4BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_23 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFF",
INIT_24 => X"FAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010000000000",
INIT_27 => X"FFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"E974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007F",
INIT_2C => X"FFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFA",
INIT_2D => X"D0402010000000000000000000000000000000000000000000000007FFFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"74BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFF",
INIT_33 => X"FFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE9",
INIT_34 => X"000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(29),        -- Port A data input
DOA(0)   => data_read_a_hi(29),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(29),        -- Port B data input
DOB(0)   => data_read_b_hi(29),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_30_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"FFDFF3FC3EFFF7FFFFBFFA000000000000000000000000000000000000000000",
INIT_19 => X"F3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF5F7AEBEBFBEFBEFFEFFF7",
INIT_1A => X"CFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCF3CF3CF3C",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000007F3F9FCFE7F3F9FCFE7F3F9F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000000000000000000000000",
INIT_1F => X"4BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_23 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFF",
INIT_24 => X"FAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010000000000",
INIT_27 => X"FFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"E974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007F",
INIT_2C => X"FFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFA",
INIT_2D => X"D0402010000000000000000000000000000000000000000000000007FFFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"74BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFF",
INIT_33 => X"FFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE9",
INIT_34 => X"000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(30),        -- Port A data input
DOA(0)   => data_read_a_hi(30),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(30),        -- Port B data input
DOB(0)   => data_read_b_hi(30),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_31_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"129000008004A00804A40000400800020000000C005FEA005800200400050100",
INIT_01 => X"A15FF18019700810180065FFFC0040801E80258CA2951C2200EC0906A0804140",
INIT_02 => X"146000808A0C060444692000402850040400408FF80000000010000000004000",
INIT_03 => X"000000FD74480B1C3D951C5A800D03FA1C0C21084B0300000012108518004842",
INIT_04 => X"07C51FC7EDFCA26E07EE001D1CB6904A061EDB6D4C30490281831C1602D0E480",
INIT_05 => X"C001F0808181117C7C95C8183FA099C7181F8703FF0CE3FC0201209010988002",
INIT_06 => X"00000000000000010001020400840C41C000617FC0003021259CFDB01BF00020",
INIT_07 => X"0000000441FA3FE400080200A810000010804008100040018448912040000040",
INIT_08 => X"00011F0780011E38004801C79E7C162231862E8FE00166704041240DF93D0000",
INIT_09 => X"F0C3FE180D89279000B00000000000D0F80088080849673F6C0E780020091480",
INIT_0A => X"1011DCCC31222730048620C4382204A608142002A440924A6188020920404437",
INIT_0B => X"0661874500E00E00304003040030400304003040030400304003060018200182",
INIT_0C => X"810040801060C04821202001A05A00040100240A80800442040202FFC3200444",
INIT_0D => X"000740000803C0616184184031010FFF40FFC407500020004C10060204010200",
INIT_0E => X"0007400000BD0020000008001F010000020201E04000010007400001E0400001",
INIT_0F => X"1DC0000000400D701000000800007700000001E04000010007400001E0400001",
INIT_10 => X"10003C064000C000010080BD0020000200001EC00000102006E8080000001000",
INIT_11 => X"140403A020000007200000E808000001C200000308C504021442354000000000",
INIT_12 => X"07B00000001D0100000038400007404000000E400000FC0010000000FC000000",
INIT_13 => X"5D00200000007C400000501001DC08000000001F010000140404558080000000",
INIT_14 => X"8C1380DA10400140640100D4080032903A8000000000403C3400008000140404",
INIT_15 => X"02008020080200802008020080200C1808008184012A08041202500AF87FF001",
INIT_16 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_17 => X"0080200802008020080200802008020080200802008020080200802008020080",
INIT_18 => X"000000000000000000000002001005FFFFFFFFFFFFFFFFF02008020080200802",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000000000000000000000000",
INIT_1F => X"4BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_23 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFF",
INIT_24 => X"FAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010000000000",
INIT_27 => X"FFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"E974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007F",
INIT_2C => X"FFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFA",
INIT_2D => X"D0402010000000000000000000000000000000000000000000000007FFFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"74BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFF",
INIT_33 => X"FFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE9",
INIT_34 => X"000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(31),        -- Port A data input
DOA(0)   => data_read_a_hi(31),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(31),        -- Port B data input
DOB(0)   => data_read_b_hi(31),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_0_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"ED39BA795990D275FB4A6E96ACC4731DEA4598B0AFB54867F6EE4618C3749807",
INIT_01 => X"58A0047D8607944AC7DA180001ECA2444042106208408208C20022E9173734B3",
INIT_02 => X"8B1E49562021F8051500147A0E162923024F28000415F5787B09FBF999BB1EFC",
INIT_03 => X"1013BF028A959403C06A23A147723C01E140088280C4CF6996088862C7922221",
INIT_04 => X"781A003802015D9078011DE20340699198600000B08694916434804825241311",
INIT_05 => X"2CA000587E10C880036A3103C00F2000E1E0383C00730002B4409845E4425171",
INIT_06 => X"179B48CFF95DCF9EF730E1C3BB731138AF7B888025340C0888430047040FEE18",
INIT_07 => X"AF155113160400185F87C1F05707D415E664A6E7C5551EBE783060CEB164833F",
INIT_08 => X"4D7E40002B7AE005FDB47600208229010C6101001EFE198C96B0528202C0DCB4",
INIT_09 => X"062400608234D864444081048A80CC00062D42D30222108091C107A1DA040267",
INIT_0A => X"204A21008E514844EB5145000255DA599581D3A9583C24351240B58298011308",
INIT_0B => X"E08C4830F81380CE0F89E07A9E0789E07A9E0789E07A9E0789E070CF0184F038",
INIT_0C => X"3A4E9D63EA180EB150CA1CA45C254D4AF4AA414568729139F2A12C0000016110",
INIT_0D => X"F0009E0FC048211E9C11C31F82E4A000890022B827EB52F52347F174E93A749D",
INIT_0E => X"F0009E0FCC42EFDFBF0AE03080E2AEB2E0F1F80FA97FE0F0009E0FC40FA97FE0",
INIT_0F => X"0231F0BD9E3FC08FEBD6F661C0E008C3CB5F040FAB3FE0F0009E0FC40FAB3FE0",
INIT_10 => X"20180309A0F83BE2B87C7C42EFDFBF187806013879BA878FE807F65FBF12E038",
INIT_11 => X"0BE9F01FC8B38C2098DAE007F323A0C83136B248831ACBFC8BBDCAB779BC699F",
INIT_12 => X"004C72BEC800FE7464290626D7003F9947184131B59003FFEC07F00003F01FB9",
INIT_13 => X"A0FFDA2A3C0202B8776A2FA7F023F7D065703080E29F1B2BE9F8A27E6E915C0E",
INIT_14 => X"016C2D25E52630BB1AE49C2BA7F98D6F846DFC0C2352A0024B83F07F198BE9F8",
INIT_15 => X"749D2749D2749D2749D2749D2749F285F25D2C500815A5522CB5A4B400000CD4",
INIT_16 => X"49D2749D2749D2749D2749D2749D2749D2749D2749D2749D2749D2749D2749D2",
INIT_17 => X"9D2749D2749D2749D2749D2749D2749D2749D2749D2749D2749D2749D2749D27",
INIT_18 => X"31C136AD8E9B562BA39E2600654BA800000000000000000749D2749D2749D274",
INIT_19 => X"4104104104104104104104104104104104104104104104109C83B8E38E2ABE71",
INIT_1A => X"0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0410410410",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000007C3E1F0F87C3E1F0F87C3E1F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000187FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"BAF7FFD55EF007FD75EFFFAE97555557BD75EF5D000000000000000000000000",
INIT_1F => X"000AA843FE00AAFBE8B45AA803DFEFA28428B455D0017410A28428AAAA2FBD54",
INIT_20 => X"FEBAA2D5401450051401555D7FC0145F7AEBFFFF08002AA10A2AABFEAAA2FFC0",
INIT_21 => X"D755555517FFEFA280021FF082E974AA5D7BFFE000804000BAAAAAAAB45557FF",
INIT_22 => X"EA8B45005168A10AA8028A10087FD7410557FC21555D51574AAA2FFE8B455D7B",
INIT_23 => X"AE95410AA80000005D003FEAAFFAEBFE00A2803FEBA002A820AA0800174BA5D2",
INIT_24 => X"2AEA8A10000417410A2FFE8BEFF7FFE8B45FFFBC00005D003FF45557FC01FFFF",
INIT_25 => X"00000000000000000000000000000000000000557DF5500003DFEFFF84175EFA",
INIT_26 => X"5F524AFE38B780154BAFFF1D54AF0075D75EFEBAE9554540754717F1F8000000",
INIT_27 => X"50B6AABDE12BEA0AF010B7D1F8F47E00A2DB45AA8A3AFD7B68E2AB78550E1255",
INIT_28 => X"E9257F1E816D557095EAAA2D1401D500002A150038038E285D7F78FD7000B6AB",
INIT_29 => X"5A87AAD178A8002D1D21C5E8257D5C7AA854008700249243A412EBFF5542A43F",
INIT_2A => X"52A82000E3A5D2150AB8F401471EDBC0B680900AAF52B474385D75C502D15754",
INIT_2B => X"FD7E9541242FE920AD082E10A28F6A150012A2F02AFFDF40E85F475451D502D1",
INIT_2C => X"0550E87B7A405B52AAD152BD00151EAFEDB52E3F1EFFFF485A2DA3D5D24BD417",
INIT_2D => X"57F40545850000000000000000000000000000000000000000000005AAF55508",
INIT_2E => X"F7AEAABFF5D2A81151FB8635A02FA69574BAF7D5555AF0D79D55FFA2AC974450",
INIT_2F => X"8D46F6ABE7082AAAAF2FAC77FE00FF16565B2FA9075F4F7B3EBDF50FEAEAAB55",
INIT_30 => X"56803CE3AEB038662E5D81406014D5D51F5E08A394003A908B8410E707EF34A0",
INIT_31 => X"4AF0151555AF58794040077D774FAE8C798A11A0EAEF75F7AA84001A7052C952",
INIT_32 => X"4E1870108B11020AD4AA05542A0A05051023F9A9D57B63BFBF906CB45FABC095",
INIT_33 => X"F5F0DA6BC9525688C1A2A0C06E9FEE5555BE48AB2A2AE0A0F20C43EAC562245B",
INIT_34 => X"000000FF80F55E25C00A0BA7FBED407A97F6F35F498B96BEB12DAAB77558ABD5",
INIT_35 => X"8000000FF8000000FF8000000FF8000000FF8000000FF8000000FF8000000FF8",
INIT_36 => X"00000000000000000000000000FF8000000FF8000000FF8000000FF8000000FF",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000008000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(0),        -- Port A data input
DOA(0)   => data_read_a_lo_256(0),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(0),        -- Port B data input
DOB(0)   => data_read_b_lo_256(0),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_1_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"212C001411984004084D000508C53810A03D1450E839B003342114428A000803",
INIT_01 => X"08000010400A0008010600000084005000400002000000000000000000140000",
INIT_02 => X"C084484000002014400205851002007030450E0000A606C8C44CB4C6666C00E0",
INIT_03 => X"CCF7CE0002058001000000800240200001018CA1800001091408463061120118",
INIT_04 => X"082800100000000040000900010000100040000000008411600401C02100000C",
INIT_05 => X"10800202080422000020012200000000810000200000000004020C00200011A0",
INIT_06 => X"56BDBFBC48C315A8660C18305750C008940D8000011000820001000104050004",
INIT_07 => X"8B4344400004000150248912154404C6060A2FE24555013E13060C158AC97F01",
INIT_08 => X"00082080087A000559102400200281000469000008B000000090108000400430",
INIT_09 => X"0000000000001004140545402820020000010010208000008041060008200001",
INIT_0A => X"2102210182004840007845004044020000200080080844200000048088000000",
INIT_0B => X"48800000190191064620646A06468064680646A0646A06468064690321503234",
INIT_0C => X"02008100200800A1100707040101E20BE0B002605C1C110848200C0000000800",
INIT_0D => X"F000A000C0000012187087010AE4B00000000810010040108104100408020401",
INIT_0E => X"F000A000CC4200002F08E03080000010F18058000003C0F000A000C4000003C0",
INIT_0F => X"000000078808C00000023461C0E00000012704000003C0F000A000C4000003C0",
INIT_10 => X"201803000000240218C0044200001E1878060000000AAC00680000001F10E038",
INIT_11 => X"2100B00048230C200009A0001303204800025200040A00D000000202090C281F",
INIT_12 => X"00000002C9000260640900004D0000904618400012900001EC03F00000000039",
INIT_13 => X"80025A0A3C020000002A8400B00007806070308000000961002880204A901C0E",
INIT_14 => X"000801046004308A185000020128000904285C0C0312A0020000000838810028",
INIT_15 => X"0401004010040100401004010040100010410C002000040280100000000008D0",
INIT_16 => X"4010040100401004010040100401004010040100401004010040100401004010",
INIT_17 => X"0100401004010040100401004010040100401004010040100401004010040100",
INIT_18 => X"48D757DF8A9410218E8A56085142020000000000000000004010040100401004",
INIT_19 => X"555555555555555555555555555554514514514514550431A581924924B02651",
INIT_1A => X"4BA5D2E974BA5D2E974BA5D2E974BA5D2EB75BADD6EB75BADD6EB75555555555",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800005D2E974BA5D2E974BA5D2E97",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000607FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"10AAAABFFFFFF803FE10F7D17FEBA55556AAAAAA800000000000000000000000",
INIT_1F => X"EBAFFD555400557BD54BA5D7FFDF45A2FBD75EFA2AE97555F7FBFFF45FFAE800",
INIT_20 => X"ABEFA2D568A005D5157400AA8028AAAF7FBD54AA002A955555D7FE8ABA082EBF",
INIT_21 => X"FDF55AAFBC0010555540010550417555AA8028BEFAAAE97555082A80000AA802",
INIT_22 => X"BD7410550428ABA5D5168ABA552EBDFEF5D7FEAA00AAAABFEAA007BC0145FFFF",
INIT_23 => X"FFEAB55557FFFEBAAAD568B45A2D5575555D7FC2155F7AEA8BEFAAAA954BA557",
INIT_24 => X"D7BD74000804154BA082ABFF55FFD57DF45F7D568ABAF7AABFFFF082ABFFFFFF",
INIT_25 => X"000000000000000000000000000000000000002EBFFEFA280021FF082E974AA5",
INIT_26 => X"5E175EFF57BF8FC2000BEA4BAE97F78A3FE28E3D17DEAA485FE8E02B50000000",
INIT_27 => X"455571E8A2A087BF8EAAEB8E0016D5D75D54BA5D7BFFF7DA2FFD55EFAAA49554",
INIT_28 => X"157428145A00AA8A2FBD7B6DF6AA28550E10405F7A4AFE38EAA0924921C2FD55",
INIT_29 => X"8E971471C7010B7D168F47400A07A28415A001684104155C5B6DF6DBEFBFAA07",
INIT_2A => X"BFBD7B6A0BF492415FC20105D24AAABF1FFBC7010FF8A38FEF557FEAB78B6AAB",
INIT_2B => X"017EBA4A8EB8F6FFD5FE8B7D557495EAAA2D16D1FDBED56A55557A43DE385FD4",
INIT_2C => X"854008700249243A417FFF41542F5D717FE2AAAA56DEBD17FE3DF7FB7FEBFE38",
INIT_2D => X"07DFCA127B8000000000000000000000000000000000000000000002A3D5C7AA",
INIT_2E => X"AAFBD55FFAA8416545A6FB60F47AF2A00010F78028B15F7823FEAAA2D57DFBA0",
INIT_2F => X"22A38C20B2552E975F758516AAAA0869AAAB8A7C19C55550E8574BA557BFFFEF",
INIT_30 => X"55FFEFBCEE5FBAACB10085EE5DE10A2AEBFF55F7BAAA8565DBAC1112FFAC21A0",
INIT_31 => X"BEA097BEAAFAF2863FA00DD574201E7AD1FFF5575841DE08007FC20480028957",
INIT_32 => X"54FF57EFBFA18D4FBFFF40FF809D4000D7FC00FC5D062BBA05ED5034472A02EA",
INIT_33 => X"7DFBFF6963FCAAA2283CF14050062B0A2F7AE8B5D5D51F5E18ABD5EAFFF2AF95",
INIT_34 => X"000000002CB75F7AA84001A7052C95256807DC31AA8114DE55F5BED201FFFED1",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000008000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(1),        -- Port A data input
DOA(0)   => data_read_a_lo_256(1),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(1),        -- Port B data input
DOB(0)   => data_read_b_lo_256(1),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_2_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10E44660018259B2843913100062C98004802322D3E030235201006009B2813",
INIT_01 => X"000AC188084900481C8024A542400340404000720885800802000906E4910204",
INIT_02 => X"82040072AC248C31010204880000007401044C0550200000480E0080001300E0",
INIT_03 => X"0080812C130D0A0D1193088802182142494D218220021100001A8020C1004A00",
INIT_04 => X"090D0AD62824A44A428408540D1610020C6E510818923441A4908B0503404201",
INIT_05 => X"5000A004081122242420480A14A99C428908122144244150906124248C002168",
INIT_06 => X"1400088400450000460000001308890094082015800011012D41D518044C1100",
INIT_07 => X"26731111491C1541324C1114BD880004002040204050413F1400100480000201",
INIT_08 => X"02410582881E0C1511D02082AAAB016A2463288549B044605201D10AE11B0020",
INIT_09 => X"E80394280E40158020B591000800481051241A4A404B5035C60904502054E000",
INIT_0A => X"0102C9E12202EA6014D027C418428E220A5500024808922801A0900A84454458",
INIT_0B => X"4600070110C10D04340043400434A043420434A04342043480434102184021A0",
INIT_0C => X"E9CA34328E44CA1401306100A246000402100C088104010AC8005C5681812B04",
INIT_0D => X"0000A0000801487334E34C1A980001550055481204090A4C01351253A728D194",
INIT_0E => X"0000A000013800004000080000000000500000B01480010000A0000150148001",
INIT_0F => X"0000000608000A500409000800000000012001501480010000A00000B0148001",
INIT_10 => X"1000000000002400000001A100004002000000000000A0000360018040001000",
INIT_11 => X"380001C01048000000090298040440000002400008C400022042004080028000",
INIT_12 => X"0000000009530080880000004813802090000000120C94000200000000000001",
INIT_13 => X"4C000100000000000002E0000950002018000000000001580002508010440000",
INIT_14 => X"7120642000000400015020500004221018000082008000000000000820180002",
INIT_15 => X"5094A5294A5294A52942509425094209461468000822241A03835D88482AB001",
INIT_16 => X"09465094A5294A5294A5294250942509425094A5294A5294A529425094250942",
INIT_17 => X"94650946509465294E5294E5294E5094650946509465294E5294E5294E509465",
INIT_18 => X"080271AE180616A38A18FA204452A7F03F03F07E07E07E05294E5294E5294E50",
INIT_19 => X"20820820820820820820820820820820820820820820490C04102CB2CB2EB2C0",
INIT_1A => X"8944A25128944A25128944A25128944A25128944A25128944A25128208208208",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF1F804A25128944A25128944A2512",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000787FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"AAAA843DFFFAAD1554005D7FD74AA00040015500000000000000000000000000",
INIT_1F => X"F45AAAAA8A10A2AE80010A2AA975FF5D003FE10F7D17FEBAF7D5420AA0855420",
INIT_20 => X"FF45A2AA975EFA2FFD7555FFFBFFF45AAFBC20AAF7D1575EF55517DF555D2EBF",
INIT_21 => X"95555552E974105D517DF55AAAAAABEFAAD1575EFAAAE974AA5D51554BA5D7FF",
INIT_22 => X"E82010F7AABFE10FFD542145FFD5554AA555555555557FE8ABA082EBFFFFAAAE",
INIT_23 => X"FBC0010AA802ABEFAAD540000FFD540000AA802AABAF7FFC2010AAAE821EF552",
INIT_24 => X"A8028BEFAAAE821550851420AA002E800AA08042AB45007FC00BAFFD168BEFF7",
INIT_25 => X"000000000000000000000000000000000000002E80010555540010550417555A",
INIT_26 => X"AE95F40002157F470AABE803AE97A2DF55400557FD54AA1D04001C5150000000",
INIT_27 => X"EF55517DFC5552ABDF45B6AEAFFD5F7A482000BEAE905C755003FE28E3D17DEA",
INIT_28 => X"0BA5FD0154BA5D7BFAF7DA2AE955EFAAA495545E3F5EFF57F7FE80082FFDE105",
INIT_29 => X"8AAF082AB8EAAEB8E0016D5D2A924105D5B7FF7DB6AAAABC7BEDB505EFBEA407",
INIT_2A => X"95038AAAEAF1D7410E80000FF8438E00B6DF68FEF4871D24BA495B5556D5571E",
INIT_2B => X"1ED1EFEAF1EFFFDEAD1C5010AA8E2FBD7B6DF47A00EBDB50000A380AAE28E804",
INIT_2C => X"5A001684104155C5B68E2DBEFBFFBC703AE2DF42AAA002A851C214003FF68007",
INIT_2D => X"50002155510000000000000000000000000000000000000000000002087A2841",
INIT_2E => X"55003FEAAAAD57DEBAA2FDDC01051FBD74BAF7802AB05AAFBD5400557BD54AA5",
INIT_2F => X"7AF7FC20B2F7FBC015D58517FF555D2ABDF55F782BEB47AFAD00010F7AA82155",
INIT_30 => X"55FFFFC20FFF3AE544108410174BA557BEABEFAAEBD55FFAA1456547A2D360F4",
INIT_31 => X"0BA547FD75FF58516AAAA0828AAAB4A78016545540400010557BFDFFFF7822A9",
INIT_32 => X"550AAFACAAA122AA8954BAA2AE9D545002A800A8FF862BA00F2F9E8F0050D442",
INIT_33 => X"954505C417FFFF08555555BAAD335B57AB5155400A2AEBFF45FFFB404007FFBD",
INIT_34 => X"00000000061DE08007FC2048002895755FFAEBCFE57BBA57002DF3C4AAAA002E",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000010000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(2),        -- Port A data input
DOA(0)   => data_read_a_lo_256(2),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(2),        -- Port B data input
DOB(0)   => data_read_b_lo_256(2),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_3_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"210C44A20020248B08431120001604B8156023104C40771B3430400A02380206",
INIT_01 => X"015A2A4050B009683C0422C992000B61404040028804A0080A000C16A8990A0C",
INIT_02 => X"C0A406500CE0A95011000D1501005274B5041AB330860281CC08008222170060",
INIT_03 => X"AB488054270F08E1289084C8020420E005A48DA16C021100003A46B06900C91A",
INIT_04 => X"848966150DA0A02941A4080C612A104201C689044382FD403C17E491829B259B",
INIT_05 => X"D006620608843116942508120A208D18A5050160C600D4C894600094B49CA068",
INIT_06 => X"12002D9401C70008060408141788E2C094887033080071913209CC8004640100",
INIT_07 => X"221111454874CCC4122C0932155400C2023940284000003E15020525CE805E11",
INIT_08 => X"020103C9984A0AC511102029869D974214EDBA132891000052C1750B48290020",
INIT_09 => X"60808C8A2E41351020004148A289428730A51E5E644C8233A0090E1020208100",
INIT_0A => X"A4000041A600417914506F955D6422000934000A090A94A020229603A414144D",
INIT_0B => X"469100841001000406D04065040650406D0406D04065040670406C8201782032",
INIT_0C => X"6A4AF532A8040AF821042D01F14084030070262810340402C0000CCE4CC12520",
INIT_0D => X"000800000401C333494594532980733302CCC81300094E5C91200257AD2AD795",
INIT_0E => X"00080000051C0000400000000000000800000190148000000800000450148000",
INIT_0F => X"0000010000000B100409000000000004000005101480000008000004F0148000",
INIT_10 => X"0000000002000000000001B00000400000000000000400000168018040000000",
INIT_11 => X"1000034010480000010002D804044000004000812E4400002440014080028000",
INIT_12 => X"0000000100570080880000080015C02090000002000CCC000200000000000040",
INIT_13 => X"1C0001000000000000104000094C002018000000000040100006418010440000",
INIT_14 => X"4128652000004404010E20500004208018800082008000000000010000100006",
INIT_15 => X"5795A5595A5595A5595A5595A5595E1152556D008028341B13924D80C2E67009",
INIT_16 => X"69565795A5595A5595A5595A5595A5595A559525795257952579525795257952",
INIT_17 => X"95256956579525495E5595A5495E5595A5495E5595A569565795256956579525",
INIT_18 => X"7818F18E0C8514298B0C52A0115009AA9556AAD552AAD5556956579525695657",
INIT_19 => X"24924924924924924924924924924820820820820825042C0000249249202A60",
INIT_1A => X"8D46A351A8D46A351A8D46A351A8D46A353A9D4EA753A9D4EA753A9249249249",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF248086A351A8D46A351A8D46A351A",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"EFAAFFD54AAF7D168B45AAAABDF5500002AA1000000000000000000000000000",
INIT_1F => X"F45FFD168AAA0855420AAAA843DFFFAAD1554005D7FD74AAA284001550055421",
INIT_20 => X"55FF5D003FE10F7803FEBAFFD5420AA080400155AAD5554AAF7802AB4500043D",
INIT_21 => X"28B45A2AE82155A2FBFFEBA0800021550855555FFAA84001FFAAAE80010A2AA9",
INIT_22 => X"168ABAFFFBD54BAAAAE97400A2FBC20AAA284175EF55517DF555D2EBFE00AA80",
INIT_23 => X"AA954AA5D7FFFF45AAAA975EF007BD7555FFFBFDF55AAFBD55EF5D2EBFE10085",
INIT_24 => X"AD1575EFAAAE974AA5D00175555D0015410F7AAAAAAA55043DE00FFFFD5555AA",
INIT_25 => X"0000000000000000000000000000000000000004174105D517DF55AAAAAABEFA",
INIT_26 => X"ABC04001C51551471D7AAF1D05D2EBD56DB7DBEAEBFF551C042AA101D0000000",
INIT_27 => X"92EB842FB5508043FF55EBD56ABD75D5B470AABE8A3AFD7A2DF55400557FD54A",
INIT_28 => X"557FD2082000BEAE905C755003FE28E3D17DEAAEBDF40002550F47155AADB504",
INIT_29 => X"DF40552ABDF45B6AEAFFD5F7A48017DAAFFFAE821C0A0717D1C5B575FFB68E82",
INIT_2A => X"C55D7492E90E3808756DA92EBFFD74BAE3AE85480FFFFC00AABE8E105C755517",
INIT_2B => X"43AE10EAF5C5547FF80954AA5D7FFAF7DA2AE905EF0075D5545E3F5EFF57F7D5",
INIT_2C => X"5B7FF7DB6AAAABC7BEDB505EFBEF5C7092FF801756D490A10438EBA4B8E92410",
INIT_2D => X"D0028A00510000000000000000000000000000000000000000000000E124105D",
INIT_2E => X"AAFBD54005D7BD54AAF78002155515157555AAD142040A2D57FFFFFFAEBFF555",
INIT_2F => X"051AE955F7AAFBC0000AF843FF5500003FF55AAFD6AB455157D74BAF7AAA8B45",
INIT_30 => X"FF557BD74EFFBACD41577B8400010F7AA8215555003FEAAAAC53DEB8A2FDDC01",
INIT_31 => X"0BAF7AA8015558517FF555D2ABDF51F782BCB47ABAE801FFAAFBEAA105D2E955",
INIT_32 => X"214FA2D3EAF57AFFDD7555082AA0AAA00557FEA8A2FDD64BAAF8282012AFFEC2",
INIT_33 => X"820AAAB842AA00000028AB0AAFF48547AE04174BA557BEABEFA2AA951FF88554",
INIT_34 => X"000000002A80010557BFDFFFF7822A955FFFFC21FFF3BE40412DE02955FF082A",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000008000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(3),        -- Port A data input
DOA(0)   => data_read_a_lo_256(3),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(3),        -- Port B data input
DOB(0)   => data_read_b_lo_256(3),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_4_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"A108400020612C80284210081034849800A000303100048B3432C82904204006",
INIT_01 => X"210668000008004C1C20250E12100368403008418984014902030906A8910200",
INIT_02 => X"120404C0024C0600000206100008402404040C00F104008040080080001310E0",
INIT_03 => X"7728805052470B5C1B873C04121D03845D0020CA0822018000080084C1000002",
INIT_04 => X"0B899E43891686690790485D5C3E02000E9892201D306D03A9835C16029AC186",
INIT_05 => X"C001E080005030767434C0003C8A01D6B81C5703C82CDBC000072400089C8120",
INIT_06 => X"1000088100410000460002041300004084080070D00030032009700024641102",
INIT_07 => X"4261950408CCBC2012048310951000000003402A4000143E1008912480000211",
INIT_08 => X"00811007AC0A1EB5131120C79E7D176251E53E80E8B361604041340838452020",
INIT_09 => X"C08360820C0912800035F1801630A8260900180C00C8021C800FEE522020A108",
INIT_0A => X"8400F88C166262E940D00D410D62AD02091704024D0A02882192020DA0544043",
INIT_0B => X"4011078510C90D143142430C243042430C24304243042430C24305121A612186",
INIT_0C => X"C08060101000C00401008800F004140009400E4002A0010240000DC3C080002C",
INIT_0D => X"000800100001C07261C51C42390240F050C3C000950008088130040100018000",
INIT_0E => X"00080010003510004000000000000048010002E0100000000800100220100000",
INIT_0F => X"0000014008001550000800000000000400800280100000000800100360100000",
INIT_10 => X"00000000020000080080009410004000000000000044080000D8008000000000",
INIT_11 => X"000005800008000001040168000040000041000100EC00004002214000008000",
INIT_12 => X"00000041003C000008000008200D00001000000208050C000200000000002040",
INIT_13 => X"17000100000000000090000002C8000008000000000060000004480000400000",
INIT_14 => X"8400C00208004844C00800000000528008000000008000000000010040000000",
INIT_15 => X"0100800004030080000C010000A00D1804404912802A261B53104810DB1E0028",
INIT_16 => X"000C030000200C01000020040300800004030000000C03000000040100802004",
INIT_17 => X"008020040100C010000200800004010040300800000020040100C03000020000",
INIT_18 => X"40C700FC0A000280C68A08A950520E964C3269B2C9864D30000C030040100800",
INIT_19 => X"555555555555555555555555555554514514514514526991A199A28A28981451",
INIT_1A => X"41A0D068341A0D068341A0D068341A0D06A351A8D46A351A8D46A35555555555",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF771F60D068341A0D068341A0D0683",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FF087FFDF5508003FEBA087FD54BAAA841540055000000000000000000000000",
INIT_1F => X"F5500003DF455555421EFAAFFD54AAF7D168B45AAAABDF55A2802AA1000002AB",
INIT_20 => X"DFFFAAD1554005D7FD74AAAA840015500002AABA082E954005500021FF5D2EBF",
INIT_21 => X"68BEF080028BFF0855555455500174BAA2AABDE0055517FF555555420AAAA843",
INIT_22 => X"168ABA0055574BA5555554BA5D0400155AAD1554AAF7802AB4500043DF45FFD1",
INIT_23 => X"0400010A2AA955FF55003FE10F7803FEBAFFD5420BA085168A00007BFDE10085",
INIT_24 => X"855555FFAA84001FFAAFBEAB45002A97545F7D1555EF55043DF5555517DEAA5D",
INIT_25 => X"000000000000000000000000000000000000002A82155A2FBFFEBA0800021550",
INIT_26 => X"5BC042AA101D0A28BC7007FFDF45080A3AEAA007BD2482BE84124285C0000000",
INIT_27 => X"004100021FF492AB8F7D1C0438E381451471D7AAFBD0492EBD56DB7DBEAEBFF5",
INIT_28 => X"FED1C5F470AABE8A3AFD7A2DF55400557FD54AABE84001C5550A28ABA1424974",
INIT_29 => X"FB5508043FF55EBD56ABD75D0428BEF005557545490012482B6A0BAE2849557A",
INIT_2A => X"6DA101475FDE10145F68A921C55504924955524AA140E0717DAADB50492EB842",
INIT_2B => X"43AF6D405F78E3A1C2002000BEAA905C755003FE28E3803DEAAEBDF40002557F",
INIT_2C => X"FFFAE821C0A0717D1C5B575FFB6DF425575D7BEFB55002097555FFD5401EF5D0",
INIT_2D => X"784000AA59000000000000000000000000000000000000000000000208017DAA",
INIT_2E => X"A2D57FFFFF7AEBFF55FF8028A00512EAAB45007FFFF55082EA8AAA087FC2010F",
INIT_2F => X"5512AAAA085D04174100800021FF002EA8BEF5D0428ABA595557555AAFBC2000",
INIT_30 => X"00FF802ABAA04552ABFF597FD74BAF7AAA8B45AAFBD54005D7BD54AAF7800215",
INIT_31 => X"5FFAAFBC0000AF843FF5500003FF55AAFD6AB4551002ABEF0055555550004020",
INIT_32 => X"DEB0A2FD5600051537DE005D557DE005D7BE8AA85555400100879560AA592F95",
INIT_33 => X"17545FFD5421FF5D0428BEF0079FCABA598400010F7AA8215555003FEAAAA843",
INIT_34 => X"0000000004001FFAAFBEAA105D2E955FF557BD75EFFBBCD415521FBFDF450004",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000010000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(4),        -- Port A data input
DOA(0)   => data_read_a_lo_256(4),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(4),        -- Port B data input
DOB(0)   => data_read_b_lo_256(4),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_5_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50DB0A0791B1B41694368283C81F9996A091A32152007AB36B20E03C040C002",
INIT_01 => X"880015C49830884C446A40000C34C24841280A00084000C8C212892EEA953231",
INIT_02 => X"408F417400B1D9100002171C1FA20171124E6AA00D8633F8CD09DBFBBB972F7C",
INIT_03 => X"88538F0182058082D800C3314722DC08A34084A100C4D7C99208521063D00148",
INIT_04 => X"F45E41AFAF420996B8411CA282F80A9091224800A2C61490363080C8A4000308",
INIT_05 => X"0EA416069640420901A01505C4410020C6E228DC30532839B043289D9C005031",
INIT_06 => X"13992D9AF8C74E92B7B568D19708C038AFFA89F0B9348C9204C389672407EF12",
INIT_07 => X"6255000016053C18162589725146F442222CE6AF844012BE795224458BA4DE0F",
INIT_08 => X"4F3F00503B4AE104B5347230418190420821006016FC18843630D285FC416CB4",
INIT_09 => X"EEA33E700340902C4424C442B0344724066C56C2248130A2D9C185B24A24832B",
INIT_0A => X"315325008348CC40AB570500204462508135D5AA593E043731E9B18A98440137",
INIT_0B => X"E0CD463C5813804E0258E0358E02D8E03D8E0258E03D8E02D8E03447012C701E",
INIT_0C => X"F8DE3C27CA181E5D710664A5F140C14BD32A2E281992940AFAA15C3FC0836310",
INIT_0D => X"F000BE0FC80020130841840308653FF0313FE92C23FB1EECB367C0F3E378F0BC",
INIT_0E => X"F000BE0FCD806FFFAF0AE83080E2AEB2F0F1E01BE53FE1F000BE0FC41BE53FE1",
INIT_0F => X"0231F0BF9E3F02A7FFD63669C0E008C3CB7F041BE1BFE1F000BE0FC41BE1BFE1",
INIT_10 => X"30180309A0F83FE2B87C7D006FFF9F1A7806013879BAA78FC103FF5F1F12F038",
INIT_11 => X"39E9C1DBF8A30C2098DBE2FF7F2320483136F200A822CBACAB9DDEB7F9BC291F",
INIT_12 => X"004C72BEC95FEF64E4090626DF15B7D1C6184131B7980DFFFC03F00003F01FB9",
INIT_13 => X"1DFFFA0A3C0202B8776AE7A7C9CBFFF060703080E29F1B79E9F6427EFE901C0E",
INIT_14 => X"2B716CA5C56620590350ACD3A7D5B7EFAC6DFC8C0312A0024B83F07F3999E9F2",
INIT_15 => X"F0BCAF3BC2F3BC6F0BCEF2BC2F3BC6DBC67C251104A2261253904580207E1C81",
INIT_16 => X"1BCEF0BC2F3BC2F1BCEF0BC6F2BC2F1BCAF1BC6F2BC6F2BCAF1BC2F3BC6F2BCE",
INIT_17 => X"BCEF0BC2F3BC2F1BCAF1BCAF3BC6F0BCEF0BCEF2BC6F2BCAF1BCAF1BC2F3BCAF",
INIT_18 => X"69CFEF73B6FFE7436DB6FD0831518424965B4D2492CB69AF1BCEF0BC6F2BC6F0",
INIT_19 => X"F7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF3EF9FBFBB9E79E7BEBCB7",
INIT_1A => X"DEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDF7DF7DF7D",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF29FDAF77BBDDEEF77BBDDEEF77BBD",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"AAA2802AA10FFFFFDE0008556AABA5D2ABFFEFFF800000000000000000000000",
INIT_1F => X"ABAF7AAA8BFFAA802ABFF087FFDF5508003FEBA087FD54BA0804154005555574",
INIT_20 => X"54AAF7D168B45AAAABDF55AA802AA1000003FEBA00002AABA5D2EBFEBAAAD16A",
INIT_21 => X"3DE005555575EFA2D142145A2FFE8B45FF80001555D2E955FFFFD5421EFAAFFD",
INIT_22 => X"FC00BA5D5568AAAF7AAAAAAAAA802AABA082E954005500021FF5D2EBFF550000",
INIT_23 => X"D5420AAAA843DFFFAAD1554005D7FD74AAAA840014500517FFEF007BEABFF5D7",
INIT_24 => X"2AABDE0055517FF555504154BAA2FBEAA105D2E97410FFD16AAAA5D2ABDEBAFF",
INIT_25 => X"000000000000000000000000000000000000000028BFF0855555455500174BAA",
INIT_26 => X"21E84124285C51574BAB68A2DA00FFFFFFE38085F6FA92552AB8FEFF78000000",
INIT_27 => X"925D2AB8EBABEDB6AA92F7AAA8BC7B68A28BC70075FDF45080A3AEAA007BD248",
INIT_28 => X"5FFFFD1471D7AAFBD0492EBD56DB7DBEAEBFF55BE842AA105D0A38EBA1C0428A",
INIT_29 => X"21FF492AB8F7D1C0438E38145B575EFA2DB45145B6F5EFB6DF78E05145552A92",
INIT_2A => X"7DFC70875EABC7557FC20AA415F68AAAF7AAAAA82BE8A28A9214249740041000",
INIT_2B => X"B6FABA542ABAE2AF7DF470AABE8A3AFD7A2DF55400557FD54AABE84001C55551",
INIT_2C => X"5557545490012482B6A0BAE2849043AFED1C0E10492B6FFEFA105D2A95410FFD",
INIT_2D => X"D2AAABEFFB8000000000000000000000000000000000000000000000428BEF00",
INIT_2E => X"082EA8AAA087FC20105504000AA5955554BAFFAEBDE10F7FBFDEBA007BFDE005",
INIT_2F => X"0512AA8AAA5D0028A005D2AA8ABAF7FBE8A00FFAEAAB45F3AAAAB4500557FF55",
INIT_30 => X"EFFFAA97545552A821EFFBD557555AAFBC2000A2D57FFFFF7AEBFF55FF8028A0",
INIT_31 => X"A005D04174100800021FF002EA8BEF5D0428ABA597FD55FFA2FFD5555FFD57FF",
INIT_32 => X"54AAF7800015551517DF45005168B55557FC0012087FEAABAF7AAAAA10F3AAAA",
INIT_33 => X"FFE005D2A95410F7FFFFEBA5D2EA8ABAFBFFD74BAF7AAA8B45AAFBD54005D7BD",
INIT_34 => X"00000000002ABEF005555555000402000FF802AAAA04452ABFF592E80010FFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000060000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(5),        -- Port A data input
DOA(0)   => data_read_a_lo_256(5),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(5),        -- Port B data input
DOB(0)   => data_read_b_lo_256(5),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_6_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10800B0061A01002840002C030028180004003220200403312301C4389B2082",
INIT_01 => X"060009C838394848188160000C42426041000000090800090210090000510200",
INIT_02 => X"00043040009001100000061000018070002408000000000648080000001210E0",
INIT_03 => X"0000800002054081020080801200A0000300008000201184681A0000410C4800",
INIT_04 => X"0808801040000001401048008100022401400002024024053200020089000100",
INIT_05 => X"0240040408402202002000C200400020A50000A0000010010001260808000520",
INIT_06 => X"44000881064500004600000013088002840C240F5048011200010000440C0146",
INIT_07 => X"0241914041FE83E010040110110003040020402A0000003E1000000488000201",
INIT_08 => X"8001BF002C4A01041B112020200110024029006FE09081002004902000012068",
INIT_09 => X"0083FE38A040100281353150ACB645AEF8C01404448000008011061204200108",
INIT_0A => X"3103AD0413424E4014D627C470462200011504420C0A962A2189002881404060",
INIT_0B => X"46C1060C16C96D15B0425B0425B1425B1425B0C25B0C25B1C25B1512D8212D82",
INIT_0C => X"009000140401100601016600A040220203A004480598010248000D0010420C0C",
INIT_0D => X"0000A01033A00013000000000018800F2400091081100C0090A5008200410020",
INIT_0E => X"0000A0103142000000000000000000455D0018100000000000A0103410000000",
INIT_0F => X"000000466800C200000000000000000001A0F4100000000000A0103410000000",
INIT_10 => X"00000000000024094680014200000000000000000041E8002900000000000000",
INIT_11 => X"F000322000000000000D1A000000000000034D240C2000502000000000000000",
INIT_12 => X"000000403F4000000000000068D24000000000001A60F0000000000000002007",
INIT_13 => X"C0000000000000000087C0003014000000000000000025D00008958000000000",
INIT_14 => X"02000000000814C219500150002800101280000000000000000000086670000C",
INIT_15 => X"8120C82208812048120882208892055A0060011280222413130449010301F051",
INIT_16 => X"3200802008320C82200802048320C82200812048320880200812048220880204",
INIT_17 => X"20C83208812048020883204802048120882204812008220C8220081204822088",
INIT_18 => X"79CFF1FE1E9F52ABEF9EFE8150120EC718638E38E30C71C812088220C8120080",
INIT_19 => X"71C71C71C71C71C71C71C71C71C71C71C71C71C71C736D9DBD9BBEFBEFBEBEF1",
INIT_1A => X"CFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FC71C71C71C",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCF29A7F3F9FCFE7F3F9FCFE7F3F9F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000607FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"EFA2FBD54BA5555554BAAAFBC20BA5D7BEAAAAFF800000000000000000000000",
INIT_1F => X"EBA0855421455555574AAA2802AA10FFFFFDE0008556AABA5D2ABFFEFFF843DF",
INIT_20 => X"DF5508003FEBA087FD54BA000415400550428AAAAA84021FF007BD54BAAAD17D",
INIT_21 => X"A8BFFAAD1554BA002A95555A28417400AAFBE8ABAF7FFD54AAAA802ABFF087FF",
INIT_22 => X"BD5545080417555A2D17FE1000003FEBA00002AABA5D2EBFEBAAAD16AABAF7AA",
INIT_23 => X"D5421EFAAFFD54AAF7D168B45AAAABDF55AA802AA100000001EF087FEAA00FFF",
INIT_24 => X"F80001555D2E955FFFF843DEAAA2803DFEF0855401FF082EA8B555D7FC21FFFF",
INIT_25 => X"0000000000000000000000000000000000000055575EFA2D142145A2FFE8B45F",
INIT_26 => X"2552AB8FEFF78E3DFFFAAFFD04AA415B52492B6F5C20825D7FE8A92FF8000000",
INIT_27 => X"EF147BD2482BED57AE921451421555551574BAB68A2DA00FFFFFFE38085F6FA9",
INIT_28 => X"4BAB68A28BC70075FDF45080A3AEAA007BD24821C04124281C0E2DA82BE8E001",
INIT_29 => X"8EBABEDB6AA92F7AAA8BC7B6D5524AA14209557DA28E15400BEF1EFA92FFFFD2",
INIT_2A => X"071FF0071EDA38F7F1D5555000417545B6D178E281C0A38EBA1C0428A925D2AB",
INIT_2B => X"4A8B555C7FC2147F7D1471D7AAFBD0492EBD56DB7DBEAEBFF55BE842AA105D0E",
INIT_2C => X"DB45145B6F5EFB6DF78E05145552A925FFFF8E3DE82BE8E38FFF0851401C7082",
INIT_2D => X"57FE8A00F38000000000000000000000000000000000000000000005B575EFA2",
INIT_2E => X"F7FBFDEBA007BFDE005D2AAABEFFBAABDFEFAAFBC00BA007BC0000FFD5420005",
INIT_2F => X"A592ABFE00F7AA821FF557FC0010F7D168A105D55421455155554BAFFAEBDE10",
INIT_30 => X"10F7D57DE00FFFBC00AAFBAAAAB4500557FF55082EA8AAA087FC20105504000A",
INIT_31 => X"AAA5D0028A005D2AA8ABAF7FBE8A00FFAEAAB45F3D5400BA5504155EFAAAE954",
INIT_32 => X"FF55FF8028A00512E975FF08557FEAAF7D157545080417545F7D56AAAA592AA8",
INIT_33 => X"AABEF005542155000028B555D7FC2145F3D557555AAFBC2000A2D57FFFFF7AEB",
INIT_34 => X"000000007FD55FFA2FFD5555FFD57FFEFFFAA97545552A821EFFBAABDE00F7AA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000048000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(6),        -- Port A data input
DOA(0)   => data_read_a_lo_256(6),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(6),        -- Port B data input
DOB(0)   => data_read_b_lo_256(6),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_7_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10844B00482258A2842112C02450418800002300500030B313300C418992002",
INIT_01 => X"020009C23838684D1C20E0000E11424840000000080000080200000000110204",
INIT_02 => X"000520700CA08910000206101180803081144880010400044808000000122160",
INIT_03 => X"000080040305208000008000328080040304008020303194289A000041484800",
INIT_04 => X"08088000000000010000CA008008060441000000028234493410820191000000",
INIT_05 => X"03500404000022020020044000000C208400408000001000984005949C002928",
INIT_06 => X"54000881044500004680000013008002940C24001A4A010200018920646410C7",
INIT_07 => X"22510040400500011204813015012204002040280000013E1000000488000201",
INIT_08 => X"9001A0602C4A01051B132820208001024069004008908002120851420001226A",
INIT_09 => X"01100020A2401008A20404E08200A05000A4264640800022C8198C4E05200018",
INIT_0A => X"20002000024040400050450440C48A0041140C420B0904208800904286000008",
INIT_0B => X"50822002120D2134800648006480064800648106481064810648193240432404",
INIT_0C => X"284A142288042A5C24202451505E00A621A5220A8091444040188C001B41210A",
INIT_0D => X"00F001F021141A12004104020810B000100000000109064C80010050A3285194",
INIT_0E => X"00F001F027420000400004C3201C514408081C1014800000F001F02810148000",
INIT_0F => X"E00E0E404100E200040900000B0380383480C81014800000F001F02810148000",
INIT_10 => X"4160C0301D07001D0402034200004000019860078641004039000180400002C0",
INIT_11 => X"08103BA0104810C8462416E8040446120C890814600010512000000080028400",
INIT_12 => X"98038D4030DD008088C2419120B740209021908C4846FC000200030F000FE006",
INIT_13 => X"DD000100411C81078884204035DC00201804C3201C60A408100DD58010440130",
INIT_14 => X"412024202211148019064200402A32901A8000B2048902C0807C0E00C448100D",
INIT_15 => X"50942509425194651946519465894619421421102000269243854D8002000250",
INIT_16 => X"19465194E50942509425094E51946519465094A50942509425194E5194651942",
INIT_17 => X"9425094251946539465094250946539465194250942509465194650942509425",
INIT_18 => X"0000000000000000000000080150890820800041041000052942509465194653",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF21E6C000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"AAF7D5575455D557DFEF002AAAB55002E820AAAA800000000000000000000000",
INIT_1F => X"B55007FD74AAAA843DFEFA2FBD54BA5555554BAAAFBC20BA5D7BEAAAAFFFBC00",
INIT_20 => X"AA10FFFFFDE0008556AABA5D2ABFFEFFFAAAAAAAF7D57FFEFF7D555555A2AEAA",
INIT_21 => X"42145552ABDFEFFFAA801EFFFFBFDF550000175555504175450055574AAA2802",
INIT_22 => X"A975EF00003DF55555168A00000428AAAAA84021FF007BD54BAAAD17DEBA0855",
INIT_23 => X"802ABFF087FFDF5508003FEBA087FD54BA000415400557BD74BAFFD140000082",
INIT_24 => X"AFBE8ABAF7FFD54AAAAAEA8ABA55557FEAAA2843FF55A2AEA8B55AAAABDEAAFF",
INIT_25 => X"0000000000000000000000000000000000000051554BA002A95555A28417400A",
INIT_26 => X"25D7FE8A92FFFFC70BAE3D155555415178FD7082EAAB550820870BAAA8000000",
INIT_27 => X"FFEBD55557DBEA4AFB550871D7482AA8E3DFFFAAFFD04AA415B52492B6F5C208",
INIT_28 => X"5550051574BAB68A2DA00FFFFFFE38085F6FA92552AB8FEFF7A0ADABAEBD578F",
INIT_29 => X"2482BED57AE921451421555524BDFD7FFA4801D7F7F5FDF55000E17545410E17",
INIT_2A => X"D2482E3D1450381C20905EF08003AF55415F6DA38080E2DA82BE8E001EF147BD",
INIT_2B => X"AAFB55ABA0BDE02EB8A28BC70075FDF45080A3AEAA007BD24821C04124281C7B",
INIT_2C => X"209557DA28E15400BEF1EFA92FFFFD24BAB6A4A8A82495F78E92AA843DF45BEA",
INIT_2D => X"800174BAA680000000000000000000000000000000000000000000055524AA14",
INIT_2E => X"007BC0000FFD542000557FE8A00F3FFD54BAAAD15754508556AB45002AA8B450",
INIT_2F => X"FFB803DEAAAAD56ABEFAAD5575EFF7803DF45085557410AEAABDFEFAAFBC00BA",
INIT_30 => X"55082E97555002E955550C55554BAFFAEBDE10F7FBFDEBA007BFDE005D2AAABE",
INIT_31 => X"E00F7AA821FF557FC0010F7D168A105D554214551003FF45FF8400145FFD57FF",
INIT_32 => X"20105504000AA597FC2010A2D1554AA5500021EF000028B55087BFDEBA042ABF",
INIT_33 => X"E8A00A2803FF45F7AABDF55AA843FE10AEAAAAB4500557FF55082EA8AAA087FC",
INIT_34 => X"0000000055400BA5504155EFAAAE95410F7D57DE00FFFBC00AAFB8028A00007F",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000007FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(7),        -- Port A data input
DOA(0)   => data_read_a_lo_256(7),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(7),        -- Port B data input
DOB(0)   => data_read_b_lo_256(7),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_8_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000B0000040042840002C0000001800000070000000033022000000000086",
INIT_01 => X"000009C21838284D1C2160000E12426840000000180800080200080040510200",
INIT_02 => X"0001004000900110000006100080003000240800014400004808000000122160",
INIT_03 => X"00008000020440810002A0801010A0044300000000200086011A000040404800",
INIT_04 => X"8000801000020401400040408108022029400000124004041200000089000100",
INIT_05 => X"02080424085022020000040200480020850010A0002010010120060800040400",
INIT_06 => X"50000880006500000680000011008006840C200018C1010200018920E0640102",
INIT_07 => X"426000404005000112048130150120240020400A0000013E1000000488000010",
INIT_08 => X"220100402C42010413110020200100024029004000A200002004902200012141",
INIT_09 => X"0000000080400008010410A2940A45240040140440800022C8388E1200A00008",
INIT_0A => X"00420100020048405000070440C0000001140412090000000021002081000048",
INIT_0B => X"0000000800000100011000010000100001000010000100001000010000880008",
INIT_0C => X"001000040001100008012008004020102180800804802000C0080D00100A0008",
INIT_0D => X"0FF0000002200A1200410402080080003000091085100C008124008000400020",
INIT_0E => X"0FF000000140000040F517CF600000000104081010001E0FF00000001010001E",
INIT_0F => X"E000000000804200000809963F1F80000000001010001E0FF00000001010001E",
INIT_10 => X"CFE7C0F00000000000810140000040E587F9E000000008100900008000ED0FC7",
INIT_11 => X"00021040030C73D80000021000585F3600000020240020102000000802419660",
INIT_12 => X"F80000000042000B0BD6C0000010800618E7B000000C000003F80FFF00000000",
INIT_13 => X"800005D5C3FD800000000008180000078A8FCF600000000002028001006AA3F1",
INIT_14 => X"020000000008808219002100100C000041120370DCAD1FC18000000000000202",
INIT_15 => X"8020080200812048120481204812055A04604930A02026934215410102000110",
INIT_16 => X"0200802008020080200802048120481204812048120481204802008020080200",
INIT_17 => X"2008020081204812048120481200802008020080200802048120481204812048",
INIT_18 => X"414A87D78AF42143CEBAC88151120A0000000000000000081204812008020080",
INIT_19 => X"F3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF7E799B1BEB65B65948051",
INIT_1A => X"C3E9F0FA7C3E9F0FA7C3E9F0FA7C3E9F0F87C3E1F0F87C3E1F0F87CF3CF3CF3C",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF1B5DA9F0FA7C3E9F0FA7C3E9F0FA7",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"0000043DF55087BC01EF007FD75FFFF84000AAFF800000000000000000000000",
INIT_1F => X"E10A28028AAAAAFBC00AAF7D5575455D557DFEF002AAAB55002E820AAAA84000",
INIT_20 => X"54BA5555554BAAAFBC20BA5D7BEAAAAFFAA95545552ABFE00087BC00AA082EBF",
INIT_21 => X"D74AAAAD57FF45002A975FF007BE8BFFA2FBFFFFFAAD5400AAFF843DFEFA2FBD",
INIT_22 => X"BE8A00082A97410F7D5555EFAAAAAAAAAF7D57FFEFF7D555555A2AEAAB55007F",
INIT_23 => X"55574AAA2802AA10FFFFFDE0008556AABA5D2ABFFEFFFAA82000555555545AAF",
INIT_24 => X"00017555550417545000015545087BC2010AAD54014500516ABFFA2AABDF4500",
INIT_25 => X"000000000000000000000000000000000000002ABDFEFFFAA801EFFFFBFDF550",
INIT_26 => X"50820870BAAA8407000140038F450075C71FF087BD75D7FF84050BAEB8000000",
INIT_27 => X"10007FC50BA002ABFE00AA8A2AABABEFFC70BAE3D155555415178FD7082EAAB5",
INIT_28 => X"082EB8E3DFFFAAFFD04AA415B52492B6F5C20825D7FE8A92FFA497545552AB8E",
INIT_29 => X"557DBEA4AFB550871D7482AAD17DF451C24955EF0875EFBD7B6F1FFFC7BEDB45",
INIT_2A => X"87000415B5057DAAFBE8A10082092410EBD5505EFB6A0ADABAEBD578FFFEBD55",
INIT_2B => X"B6ABC7B6AABFFED0051574BAB68A2DA00FFFFFFE38085F6FA92552AB8FEFF7AA",
INIT_2C => X"A4801D7F7F5FDF55000E17545410E17555000E17545007BC0000BED14217D005",
INIT_2D => X"784174AAA280000000000000000000000000000000000000000000024BDFD7FF",
INIT_2E => X"08556AB45002AA8B450800174BAA684174105D042AB550055555FF007BD7555F",
INIT_2F => X"0F384175555D2EA8A00087BD74BA082EBDE10AAAEA8ABAF7FFD54BAAAD157545",
INIT_30 => X"55FFD57DF55FFFBD5400A2AABDFEFAAFBC00BA007BC0000FFD542000557FE8A0",
INIT_31 => X"EAAAAD56ABEFAAD5575EFF7803DF45085557410AED17FF455D04155FF00557DF",
INIT_32 => X"DE005D2AAABEFFBAE97410087BC21EFA2FFEAA00000002010A2D5421FFFF803D",
INIT_33 => X"C0010FFD1401EF087FE8B55FFAEBDFEF0855554BAFFAEBDE10F7FBFDEBA007BF",
INIT_34 => X"00000000003FF45FF8400145FFD57FF55082E97555002E955550C2E95555087B",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000020000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(8),        -- Port A data input
DOA(0)   => data_read_a_lo_256(8),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(8),        -- Port B data input
DOB(0)   => data_read_b_lo_256(8),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_9_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00018248A2840112C00002C18000002300500030B3132000400812002",
INIT_01 => X"A140098218302849180060000C004240413C0A61590001D90213C90008510204",
INIT_02 => X"102008700CB089100002061031285074810448800104008048080080001210E2",
INIT_03 => X"00008015074608840390A0040040800203140000A00010800408108448020042",
INIT_04 => X"082080400004A00100000100840602020100000002C2344156108201811801C0",
INIT_05 => X"0200048480011502049500280020CC2084000080008010019161249C9C002188",
INIT_06 => X"70000881004500004E01020411D08000940C00001800010200018B20206C0102",
INIT_07 => X"EA70C0040005000312048130150100040020404A0000017E10408104C8000110",
INIT_08 => X"000000402C220104131004202081120050A5104000A204617201D10801002000",
INIT_09 => X"000800002F4924003085E51420A0100400641E4E40800022C8088C1220200908",
INIT_0A => X"20102000024040484028450001648C2229150400080244000401900284000440",
INIT_0B => X"0880110901081110411204112040120411204012041120401204111020090208",
INIT_0C => X"685B34A688841A5C21200101A01A0004009024028004044248404D00104B2100",
INIT_0D => X"0000A01000000213000000000000B0001000010000190E44802002D1A168D0B4",
INIT_0E => X"0000A010014000000000000000000040500008100400000000A0100410040000",
INIT_0F => X"0000004608004200040000000000000001A004100080000000A0100410008000",
INIT_10 => X"00000000000024080000014000000000000000000040A0000900010000000000",
INIT_11 => X"300013E010000000000D00F804000000000340000C0000102000000080000000",
INIT_12 => X"00000040091F0000800000006807C000800000001A0CFC000000000000002001",
INIT_13 => X"DD000000000000000082C00019DC002000000000000021500006D58010000000",
INIT_14 => X"03206420000000C019502050000C32901A800080000000000000000860100006",
INIT_15 => X"D1B46D1B46D0B42D0B42D0B42D8B424342342832002A24921082158802001011",
INIT_16 => X"0B42D0B42D0B42D0B42D0B46D1B46D1B46D1B46D1B46D1B46D1B46D1B46D1B46",
INIT_17 => X"B42D0B42D1B46D1B46D1B46D1B46D1B46D1B46D1B46D1B42D0B42D0B42D0B42D",
INIT_18 => X"89999E91BCD1512B871C4A0100000000000000000000000D0B42D0B42D0B42D0",
INIT_19 => X"A28A28A28A28A28A28A28A28A28A29A69A69A69A69A51C200807249041202AE6",
INIT_1A => X"8349A4D068341A0D269341A0D269341A0D068341A0D068341A0D068A28A28A28",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF2DA921A0D269341A0D068349A4D06",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"45A280154BA5555401EFFFD5421EFA2FFFFF555D000000000000000000000000",
INIT_1F => X"5EF00557DF555D040000000043DF55087BC01EF007FD75FFFF84000AAFFD57DF",
INIT_20 => X"75455D557DFEF002AAAB55002E820AAAA843DFEF00517DEBA007BFDFEFFFD157",
INIT_21 => X"28AAAAAAABDF45F7803FFEF555568AAAF7802AA00FFFBD7555087BC00AAF7D55",
INIT_22 => X"BD54BA550417400085155555082A95545552ABFE00087BC00AA082EBFE10A280",
INIT_23 => X"043DFEFA2FBD54BA5555554BAAAFBC20BA5D7BEAAAAFFFBC00AA552E95545087",
INIT_24 => X"2FBFFFFFAAD5400AAFF8402000A2FFFDF555D7BE8BFF5D51575EFA280175555D",
INIT_25 => X"00000000000000000000000000000000000000557FF45002A975FF007BE8BFFA",
INIT_26 => X"7FF84050BAEBDF78F45B68010482415B471C7E3DF451EFBEFBFAF45490000000",
INIT_27 => X"82007FFAFEFE3DB505EF1C5B7AF45490407000140038F450075C71FF087BD75D",
INIT_28 => X"5451C7FC70BAE3D155555415178FD7082EAAB550820870BAAA8438FFF00517DE",
INIT_29 => X"50BA002ABFE00AA8A2AABABEAEB8F45F78A3DFD741516DAAAE38E2DA28EBFFD5",
INIT_2A => X"C20BA5D2E905550071D54825D0A1543808515756D1C2497545552AB8E10007FC",
INIT_2B => X"5505FFBE801256D490E3DFFFAAFFD04AA415B52492B6F5C20825D7FE8A92FFFF",
INIT_2C => X"24955EF0875EFBD7B6F1FFFC7BEDB45082EB8002000AAFFFDF6D417FEABEF5D5",
INIT_2D => X"7FBE8B5500000000000000000000000000000000000000000000000517DF451C",
INIT_2E => X"0055555FF007BD7555F784174AAA2FBEAB45F78402010007BD5545AAFFD55EFF",
INIT_2F => X"AA68028BEF00517FE10007BE8BFFAAFFC01FF557FE8B550004174105D042AB55",
INIT_30 => X"AAAAAEBFEAAAAFFD5545557FD54BAAAD15754508556AB45002AA8B450800174B",
INIT_31 => X"5555D2EA8A00087BD74BA082EBDE10AAAEA8ABAF7AAAAB45F7AEBFF4508557FE",
INIT_32 => X"2000557FE8A00F3FFC00BA552E80145005557400552A954BA0051575EF550417",
INIT_33 => X"FDFFF007FE8BFF5551401EFF784021FF002ABDFEFAAFBC00BA007BC0000FFD54",
INIT_34 => X"00000000517FF455D04155FF00557DF55FFD57DF55FFFBD5400A28400010A2FB",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000040000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(9),        -- Port A data input
DOA(0)   => data_read_a_lo_256(9),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(9),        -- Port B data input
DOB(0)   => data_read_b_lo_256(9),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_10_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00018248A2840112C00002C18000202300500030B3132000400992006",
INIT_01 => X"A140098218302849180060000C00424040000000080000080200090008510204",
INIT_02 => X"102100400C8001100000061000A8503401044880010400004808000000122160",
INIT_03 => X"000080150746088401908000100080020304000020201080001A108448404842",
INIT_04 => X"800080400004A001000040008406020201000000020004401000000180180080",
INIT_05 => X"02000484800133020495040800208C20A4000080000010000001249010042008",
INIT_06 => X"50000881004500004681020411808000940C20001800010200018920206C0102",
INIT_07 => X"024084044005000112048130150120040020400A0000013E10408104C8000010",
INIT_08 => X"000100402C020105131100200000124250A51040088084614001110801012000",
INIT_09 => X"00080082CD09240820800000000000040000180840800022C8088C1220200108",
INIT_0A => X"841201000200484910000F050560262229140402080200A00402000484140400",
INIT_0B => X"0010118900080010000200102001020000200002001020010200001000010008",
INIT_0C => X"408120900404004821202001F05E00040180260A8080044240004C0010800228",
INIT_0D => X"0000A01000000813004104020800800030000800010008088124020102008100",
INIT_0E => X"0000A010014000004000000000000040500008101480000000A0100410148000",
INIT_0F => X"0000004608004200040900000000000001A004101480000000A0100410148000",
INIT_10 => X"00000000000024080000014000004000000000000040A0000900018040000000",
INIT_11 => X"3800100010480000000D00000404400000034000282000102000000080028000",
INIT_12 => X"00000040090000808800000068000020900000001A0000000200000000002001",
INIT_13 => X"80000100000000000082E0001000002018000000000021580000800010440000",
INIT_14 => X"00004000000004C0195000500008000000000082008000000000000860180000",
INIT_15 => X"0100401004010040100401004090055804404110802A24921317580802001011",
INIT_16 => X"0000000000000000000000040100401004010040100401004010040100401004",
INIT_17 => X"0040100400000000000000000000000000000000000000000000000000000000",
INIT_18 => X"215281FC1A72E2486AAA40A85052020000000000000000001004010040100401",
INIT_19 => X"51451451451451451451451451451451451451451452AA83330A8A28A29EA8D1",
INIT_1A => X"5CA6532994CA6532B95CAE572994CA6532994CA6532994CA6532994514514514",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF31CE2E572994CA6532994CAE572B9",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"10AAFBE8AAAA2D540000F7D57DF55A2AABFFEF08000000000000000000000000",
INIT_1F => X"F45FFFBC2010AAD57DF45A280154BA5555401EFFFD5421EFA2FFFFF555D003FE",
INIT_20 => X"DF55087BC01EF007FD75FFFF84000AAFF8002155AAFFE8B45AAD540000087FFD",
INIT_21 => X"7DF555D517FEBA082A801EFF7FBD5400FFD568B555D00155EF08040000000043",
INIT_22 => X"BFDE00A2FBC0145005168A10AA843DFEF00517DEBA007BFDFEFFFD1575EF0055",
INIT_23 => X"7BC00AAF7D5575455D557DFEF002AAAB55002E820AAAA803FEBA082AAAAAAF7F",
INIT_24 => X"7802AA00FFFBD7555082E82155FFAEAAB55AAD568B455D00154BAFFFBD75EF5D",
INIT_25 => X"000000000000000000000000000000000000002ABDF45F7803FFEF555568AAAF",
INIT_26 => X"FBEFBFAF4549003DE10BEF5EDAAAAAD547038EBD57DF7DA2AEB8FC7000000000",
INIT_27 => X"6DAADF470280075FFF45E3F1C7038A2DF78F45B68010482415B471C7E3DF451E",
INIT_28 => X"5C7000407000140038F450075C71FF087BD75D7FF84050BAEB8002155BEF5EDB",
INIT_29 => X"AFEFE3DB505EF1C5B7AF45495B7DEAA0824851EFEBFBD2410EBD168B7D410A17",
INIT_2A => X"38EAA0824A8AAAEBF5FAE28AAF1C2155005F68A10A28438FFF00517DE82007FF",
INIT_2B => X"4104AAF7F1D75EF557FC70BAE3D155555415178FD7082EAAB550820870BAAA80",
INIT_2C => X"8A3DFD741516DAAAE38E2DA28EBFFD55451C2087155EBA4A8B7DAADF68B7D410",
INIT_2D => X"2AEAAB55000000000000000000000000000000000000000000000002EB8F45F7",
INIT_2E => X"007BD5545AAFFD55EFF7FBE8B5500043FE00F7D17FEBAA2D5574BAAAD17DFEFA",
INIT_2F => X"AA28002155FFD17FFFFA2FBD74BA00557FF45A2D5554AAA2FBEAB45F78402010",
INIT_30 => X"00AAD16ABFF002A975450004174105D042AB550055555FF007BD7555F784174A",
INIT_31 => X"BEF00517FE10007BE8BFFAAFFC01FF557FE8B55007FFDEAA0004175FFA2FBC20",
INIT_32 => X"8B450800174BAA68428AAA08042AABAAAD56AABAAAD140155087FEAA10A28028",
INIT_33 => X"2ABEFAAFBE8BFF0004020AAFFD5555EF557FD54BAAAD15754508556AB45002AA",
INIT_34 => X"000000002AAAB45F7AEBFF4508557FEAAAAAEBFEAAAAFFD5545550015555A284",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000047FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(10),        -- Port A data input
DOA(0)   => data_read_a_lo_256(10),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(10),        -- Port B data input
DOB(0)   => data_read_b_lo_256(10),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_11_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10180B05A0010402840602C2D001019000000300000000330A20080EC180002",
INIT_01 => X"AB400984B830084C1820E0000C36424840000000080000088200000802112220",
INIT_02 => X"102A68440080011000000618062AD03502640800010410424908136019920868",
INIT_03 => X"001282118644C88481908001106088022300000080F4925CDC9A10844A9A4842",
INIT_04 => X"401280480004A1011000418084460002E12000000200040010000040A8000000",
INIT_05 => X"0FC8048484011502059511488020802084400888001110000000050000005400",
INIT_06 => X"1011088AE24500001631024511C08004A70AA40008B90D0200018B60A0650D45",
INIT_07 => X"020011005405000910040150110041040024400D800002BE18408104C9205908",
INIT_08 => X"89390040280241041D175820000001020061004004800567403512A801014C46",
INIT_09 => X"050800E20D09A424C5840400808000040680180840800022D8288E946CA00833",
INIT_0A => X"85002000024040410A000D0504408C32E915D9C208050084840201A099100400",
INIT_0B => X"B01011934A005101431CA821CA831CA821CA831CA831CA821CA83165410E5410",
INIT_0C => X"00010080028000010402214850444091019B02080885200042A9CC001000003A",
INIT_0D => X"5A5018C5A0A00812004104020808B00030000808024008008325820000000000",
INIT_0E => X"5A5018C5AB0062C38A4DB680A0D8241500D5761B011986695014A96E1A811986",
INIT_0F => X"42056A289A1BB2078A922DA2A8B180A2600AAE1A811986695014A96E1B011986",
INIT_10 => X"05AA429189B60AC43C6C7F0272C3841DB528802CAB18468F4101621B1BAC8455",
INIT_11 => X"C003104289A668B8CAB270106338317A3D94392020224ACDE215883078681B5C",
INIT_12 => X"804B020A06020C67061BC785938085134CD551BCA1C90006C0C2958502861120",
INIT_13 => X"80819A5539D503336D61056ABA006282806CA64090B89E015AAA880E48382EB8",
INIT_14 => X"40000000E808989003066E03513E41470126C6284B2D20410AB4503089C00A82",
INIT_15 => X"0000000000000000000000000000041800400110200026124202500802000800",
INIT_16 => X"1004010040100401004010000000000000000000000000000000000000000000",
INIT_17 => X"0040100401004010040100401004010040100401004010040100401004010040",
INIT_18 => X"C110083018162148420840280050800000000000000000001004010040100401",
INIT_19 => X"000000000000000000000000000001041041041041003882928E0000000AA0C4",
INIT_1A => X"0000000000008040000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3E0FC000000000000020100000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"EFAA842ABEFA280155EFFFFBC01EF08554000055000000000000000000000000",
INIT_1F => X"F4508514000000003FE10AAFBE8AAAA2D540000F7D57DF55A2AABFFEF0804155",
INIT_20 => X"54BA5555401EFFFD5421EFA2FFFFF555D51575FFA2FFD75FF550015400FFFBFF",
INIT_21 => X"C2010AAD568AAAAAD142145FF80155EF0051555FF0804155FFF7D57DF45A2801",
INIT_22 => X"01540008514215555003DFFFA28002155AAFFE8B45AAD540000087FFDF45FFFB",
INIT_23 => X"040000000043DF55087BC01EF007FD75FFFF84000AAFF802ABFFA2AABFE10080",
INIT_24 => X"FD568B555D00155EF085168B45085142010FFAE800AA5D7BFDF45F7FFEAA0000",
INIT_25 => X"00000000000000000000000000000000000000517FEBA082A801EFF7FBD5400F",
INIT_26 => X"DA2AEB8FC70000175EFB6802DBC7BE8A155EFE3FBC71FF145B42038550000000",
INIT_27 => X"EF550E15400E3F1FFF7D085B420381C003DE10BEF5EDAAAAAD547038EBD57DF7",
INIT_28 => X"5C7F7DF78F45B68010482415B471C7E3DF451EFBEFBFAF45495F575FFBEF5D05",
INIT_29 => X"70280075FFF45E3F1C7038A2DB68ABAB6D145145FF84155D7085B555C7140410",
INIT_2A => X"28BEFBEA4BDE28140A1543800514515549003FFC7BE8002155BEF5EDB6DAADF4",
INIT_2B => X"FFFF7DE3F1EFA10140407000140038F450075C71FF087BD75D7FF84050BAEB84",
INIT_2C => X"24851EFEBFBD2410EBD168B7D410A175C7005B6DB55145140000FFAE85082417",
INIT_2D => X"57BC20AA5D0000000000000000000000000000000000000000000005B7DEAA08",
INIT_2E => X"A2D5574BAAAD17DFEFA2AEAAB550004175FFF7803DF45FFAE955EFAAFBD55EF5",
INIT_2F => X"5007FD75FFF7D5401EF5D2E97410AAD17DFEF007FC20AA5D043FE00F7D17FEBA",
INIT_30 => X"55007FD5545550400145FFFBEAB45F78402010007BD5545AAFFD55EFF7FBE8B5",
INIT_31 => X"155FFD17FFFFA2FBD74BA00557FF45A2D5554AAA2FBEAAAAFFD555545FF80155",
INIT_32 => X"7555F784174AAA2842ABEFFF803DEAA5D2E974AA00515754500003FF55FF8002",
INIT_33 => X"40000FFAE97410007BFFFFFA2D57FE105D04174105D042AB550055555FF007BD",
INIT_34 => X"000000007FFDEAA0004175FFA2FBC2000AAD16ABFF002A97545007FFFF455555",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000040000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(11),        -- Port A data input
DOA(0)   => data_read_a_lo_256(11),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(11),        -- Port B data input
DOB(0)   => data_read_b_lo_256(11),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_12_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50080B01BC002006940202C0DE041196A83183000000023322287E0FC000006",
INIT_01 => X"0E000C068000E04D40238000001702484000000008000008820009280A553231",
INIT_02 => X"400B71440C8001100000171C0283813013766A800586235ECC09C8423B962966",
INIT_03 => X"CC618E048306E082000081000040900003548421A080025EDF08421042DC0108",
INIT_04 => X"00028020000000812000012080080000E100001002000448100000C1BC18008C",
INIT_05 => X"0FF8060610000402010015E100004C2084800090000310000000079010007C19",
INIT_06 => X"33992D98DEC74A003EA468D01510C03E8F580C800A3F018200418927E0668645",
INIT_07 => X"0204000406050013142409121142F746222EE2498000007E111204058B84C50C",
INIT_08 => X"E826A0602902A10491165C200000820018A5104010C01086003C13E000004EDF",
INIT_09 => X"023000000000000867000000000000040000600060801022C9F88D244FA40133",
INIT_0A => X"00100000820040482B28050001600010C13499F01B334015980001E09F000000",
INIT_0B => X"B80460124F16F06BC20CBC30CBC20CBC20CBC30CBC20CBC20CBC3065E1865E10",
INIT_0C => X"00000000029D204B7C0382FD0100F3F9F80FA0200E0BF40063F99C0010000012",
INIT_0D => X"93900F6EE230301208008001007A80001100002002801000A042000000000000",
INIT_0E => X"93900F6EEC421392C96B1237E0D8BD9629F97E0B348EDAC3900F6EFA0B158EDA",
INIT_0F => X"622DBC31D73F6006A5891533EF9500EAE64BCA0B158EDAC3900F6EFA0B348EDA",
INIT_10 => X"C2B083798D341B10DEFE14400392C74CAEAD412EDD2B4FCFF812A383430C669E",
INIT_11 => X"49FAB442994B3238D4E2FB104636652E19B8BA30C022DAD8C100CA39E8CEBE66",
INIT_12 => X"30469392526208C6CC95C33717D88532966471A9C5DD00B12728D5360234D62A",
INIT_13 => X"828C4999AF580395542D27CDBA0020F0FABAC800DA550C29F36A8A2554E48A64",
INIT_14 => X"40000000873FB80B8A00EF03F56CC12B416A51B60585A5C28895962502E9F36A",
INIT_15 => X"0000000000000000000000000000008000000410802A26924010000002000EE0",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"28C1111026C152A121960A884042020000000000000000000000000000000000",
INIT_19 => X"2082082082082082082082082082092492492492492400200005A8A28A200A37",
INIT_1A => X"964B2592C964B2592C964B2592C964B2590C86432190C86432190C8208208208",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF400FEB2592C964B2592C964B2592C",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FF00042ABEFFF8400010082EAABFF55002ABEF08000000000000000000000000",
INIT_1F => X"BEFFFFBD54000004155EFAA842ABEFA280155EFFFFBC01EF0855400005555421",
INIT_20 => X"8AAAA2D540000F7D57DF55A2AABFFEF08556AA10000028AAAFFD15541000002A",
INIT_21 => X"40000005168AAA087BFFFFF5D04001FF00041554555557FE005D003FE10AAFBE",
INIT_22 => X"1555FF082AA8B55F7AEA8BEF5551575FFA2FFD75FF550015400FFFBFFF450851",
INIT_23 => X"D57DF45A280154BA5555401EFFFD5421EFA2FFFFF555D0000145082E955FF085",
INIT_24 => X"051555FF0804155FFF7842AA100000020BAAA801541055042ABEFFFFBD5410AA",
INIT_25 => X"000000000000000000000000000000000000005568AAAAAD142145FF80155EF0",
INIT_26 => X"F145B42038555F401D71C0A2DBC7EB80000280824ADBD7490E28BEF080000000",
INIT_27 => X"82FFDB5243800002FBD7EBFBD24101C00175EFB6802DBC7BE8A155EFE3FBC71F",
INIT_28 => X"E1041003DE10BEF5EDAAAAAD547038EBD57DF7DA2AEB8FC7005F6AA381C0A2DA",
INIT_29 => X"5400E3F1FFF7D085B420381C5B6AA82147FF8FEF410E001FF000E17555555B7A",
INIT_2A => X"0017D142E905EF1451525C7082AADB45F7AEA8BEF555F575FFBEF5D05EF550E1",
INIT_2B => X"02FBEFEBFBD2410AADF78F45B68010482415B471C7E3DF451EFBEFBFAF454900",
INIT_2C => X"D145145FF84155D7085B555C71404105C7F7842FA381C0A00082AA8A10410410",
INIT_2D => X"02AA8BEF000000000000000000000000000000000000000000000005B68ABAB6",
INIT_2E => X"FFAE955EFAAFBD55EF557BC20AA5D7BC01555D2EBFF55A284000AA08003FF550",
INIT_2F => X"5007BE8AAA5D2EBDE00FFFFC00AA08003FF55A2FBC00105D04175FFF7803DF45",
INIT_30 => X"FF082A97555557FE8A0000043FE00F7D17FEBAA2D5574BAAAD17DFEFA2AEAAB5",
INIT_31 => X"5FFF7D5401EF5D2E97410AAD17DFEF007FC20AA5D7BE8A005D7FEABFF002E821",
INIT_32 => X"55EFF7FBE8B550004001FF5D2A801EF5D5142145082EBFF55F7AAAABEF5D7FD7",
INIT_33 => X"82010A2AA8000008043FFFFA2FBC2010A2FBEAB45F78402010007BD5545AAFFD",
INIT_34 => X"000000007BEAAAAFFD555545FF8015555007FD5545550400145FF843DEAA552A",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000007FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(12),        -- Port A data input
DOA(0)   => data_read_a_lo_256(12),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(12),        -- Port B data input
DOB(0)   => data_read_b_lo_256(12),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_13_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10110A0441812402840402822007818000E00700000000330A3000000008042",
INIT_01 => X"A1400986B830E84D182260000C1042484001000008220008A20019080A510200",
INIT_02 => X"10A108600C9141100000C6180CA85035010E4880010431004908135980122D60",
INIT_03 => X"0013881507460886C190832175809C02030400002020124C441A108468424842",
INIT_04 => X"203080680204A0113801D600864E0C96C12000008244244052200201801802C0",
INIT_05 => X"030004849601110204950409C0208C2084E0009C0000100120A00C9918002098",
INIT_06 => X"10000882804544921681428591908000AF28A8002BC00D020003896020658FC4",
INIT_07 => X"CA20400450050009100501501102E0042020448D0000023E10408144C800D800",
INIT_08 => X"1D2B00402B220104B53100200001020218A5104016CC1C616401910801010100",
INIT_09 => X"050800404D49A42EB08000000000000406481C8C408000A2D8088D1820200B00",
INIT_0A => X"0010000002004048AA08050401604462E9144002090740148441200484000500",
INIT_0B => X"000A112100000000010000000001000000000000001000000000000000800000",
INIT_0C => X"509528954404144C200425010040000001B020081094040072005C0030864208",
INIT_0D => X"1C10B3831034081200000000000430003000206822F20CA8826AC2A14250A128",
INIT_0E => X"1C10B383110218CB0E54C2EA404A4F03D404A41AA5B7344C10B383081BA4B734",
INIT_0F => X"8001CE3E20A5B284ED1132909C72885A2B2C381BA4B7344C10B383081AA5B734",
INIT_10 => X"AC3CC0C0B8182597A801610218CB0C3548B3A008E730A01AB113A5524E6ACA67",
INIT_11 => X"A151EC5952E44128CA194517354C180A3C066430202021252991C22C99731014",
INIT_12 => X"1804C8A0ADA2E6A983014780CA28B2A5C8825194332B018A444AEA2701288A15",
INIT_13 => X"02D09852745F80112C428562EE0353635232D50048A411C158BB0A7910142C77",
INIT_14 => X"4240480068001C9B9150A0000297046E4023F8BE8E3E1E0109472C3EB50158BB",
INIT_15 => X"A1284A1284A1284A1284A1284A12851A84284110406A26924302590806000110",
INIT_16 => X"1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284",
INIT_17 => X"284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A",
INIT_18 => X"7DDFE7EFBEFFE7D3EFBEFC48A0550000000000000000000A1284A1284A1284A1",
INIT_19 => X"D75D75D75D75D75D75D75D75D75D75D75D75D75D75D7EFBFBFBBAAAAAABEFDF7",
INIT_1A => X"5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5D75D75D75",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000FEFD7EBF5FAFD7EBF5FAFD7EBF",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"AA5D043FFFFAAAABDEAA557BFDE00FFD140155F7800000000000000000000000",
INIT_1F => X"400AAD540155A2D5421FF00042ABEFFF8400010082EAABFF55002ABEF08556AA",
INIT_20 => X"ABEFA280155EFFFFBC01EF08554000055043DEBAF7843FFFFF7AABDF55A2AA97",
INIT_21 => X"D5400005568A1055043DEBAAAFFE8B45557FD7410552EAAABAAA84155EFAA842",
INIT_22 => X"FE8ABAAA8428A00087BD7555FFD56AA10000028AAAFFD15541000002ABEFFFFB",
INIT_23 => X"803FE10AAFBE8AAAA2D540000F7D57DF55A2AABFFEF085557545FFD17DEBAA2F",
INIT_24 => X"0041554555557FE005D0000155557BEAABA5D2ABDF450851420AA5D7FD5555A2",
INIT_25 => X"000000000000000000000000000000000000005168AAA087BFFFFF5D04001FF0",
INIT_26 => X"7490E28BEF08516DA82410A3FFD7AAA4B8E824971F8E38E3DF45155EB8000000",
INIT_27 => X"D7EBA4BDF45AAAA90410BEDF45155A2DF401D71C0A2DBC7EB80000280824ADBD",
INIT_28 => X"A82B680175EFB6802DBC7BE8A155EFE3FBC71FF145B42038550E38E92EB803FF",
INIT_29 => X"243800002FBD7EBFBD24101C556FA38490A3FE92BEFFEAB45417FD24385D2AAF",
INIT_2A => X"5056DE3D17FE92BEF1EFA92AA8428A10007FD557DFFDF6AA381C0A2DA82FFDB5",
INIT_2B => X"B400925D7FD557DA2803DE10BEF5EDAAAAAD547038EBD57DF7DA2AEB8FC70051",
INIT_2C => X"7FF8FEF410E001FF000E17555555B7AE10410E00155497FEFABA4120B8F55085",
INIT_2D => X"2FBD7545AA8000000000000000000000000000000000000000000005B6AA8214",
INIT_2E => X"A284000AA08003FF55002AA8BEF00517FE00082EBDF45AA8428A10085568ABAA",
INIT_2F => X"A5D2EA8A00A2803DF45AA843DF55AAAE82000F7FBD5545AAFBC01555D2EBFF55",
INIT_30 => X"55087FC00BA552ABFE10F784175FFF7803DF45FFAE955EFAAFBD55EF557BC20A",
INIT_31 => X"AAA5D2EBDE00FFFFC00AA08003FF55A2FBC00105D517FEAA082EBFE10F7FFE8B",
INIT_32 => X"DFEFA2AEAAB550051401FFA2D57FE10F7D57DE00AA842AA00007FD75FFF7FBE8",
INIT_33 => X"FDEAA08042AB45087FC0010557FD55FFAA843FE00F7D17FEBAA2D5574BAAAD17",
INIT_34 => X"000000007BE8A005D7FEABFF002E821FF082A97555557FE8A00002E82155007B",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000067FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(13),        -- Port A data input
DOA(0)   => data_read_a_lo_256(13),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(13),        -- Port B data input
DOB(0)   => data_read_b_lo_256(13),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_14_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10020A000180000284008280000281800000030000000033022000000580002",
INIT_01 => X"A14009821830284D186860000C30C24840000000084000084200090008510200",
INIT_02 => X"102100600C9001100000061020A8503401044880010400204908012018122F64",
INIT_03 => X"00008015074608840190800010008002030400002074F401209A108448404842",
INIT_04 => X"000080400004A00100004000840E000201000000024024401200020180180080",
INIT_05 => X"0A000484800111020495040800208C2084000080000010010020049818002008",
INIT_06 => X"1000088020450402B6A1420511C080008468A80008000D0200018B202067AF10",
INIT_07 => X"422000044005000910040110510260040024400C800000BE3850A144C924080E",
INIT_08 => X"000B004028020104111100200001020210A51040008004616001910801010000",
INIT_09 => X"000800004D492408208000000000000406401C0C40800022C8088DB420200900",
INIT_0A => X"0010000002004048000005040160042229140002090200000401000484000400",
INIT_0B => X"0000110100000000010000100000000000000100000000000000100000000000",
INIT_0C => X"409120940404104C2000210100400000011020080084040040005C0010820208",
INIT_0D => X"E0E0A0000190081200000000000000003000000000100C088020028102408120",
INIT_0E => X"E0E0A0000B02740421A0E5D1A024002050805210040000B0E0A0000210040000",
INIT_0F => X"E01200860008920106460D4501CB000111300210008000B0E0A0000210008000",
INIT_10 => X"0ABBC00905C33C6000400F02740412C0715C40110080A4006110510C14D18178",
INIT_11 => X"20000041DB011CC000090012565306500002411420220080220C0093C3892324",
INIT_12 => X"5809240C09024A4AE0CA00004800839682398000120800658992F3C700C30181",
INIT_13 => X"002B46867DBC002A830280000800F7B7A0B1E240240A8340000200067EAA8CB6",
INIT_14 => X"42004005800004801150A00341244000845C7DB0D0200900422ACA4B28000002",
INIT_15 => X"8120481204812048120481204812051A04204110002A26924302590802000000",
INIT_16 => X"1204812048120481204812048120481204812048120481204812048120481204",
INIT_17 => X"2048120481204812048120481204812048120481204812048120481204812048",
INIT_18 => X"69CB91FE1EF7D3ABEFBECA080050000000000000000000081204812048120481",
INIT_19 => X"F3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF7EFBBBBBF9E79E7BEAAF3",
INIT_1A => X"CFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCF3CF3CF3C",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FF007F3F9FCFE7F3F9FCFE7F3F9F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"45AAD157400007BEAAAAAAAE955555D5568A105D000000000000000000000000",
INIT_1F => X"0AAF784020AAF7D56AAAA5D043FFFFAAAABDEAA557BFDE00FFD140155F7D17DF",
INIT_20 => X"ABEFFF8400010082EAABFF55002ABEF085155400FFD1420100055574AAA2AA80",
INIT_21 => X"40155A28028B550051574005D7FFFE105D7BD7545A284020BA0055421FF00042",
INIT_22 => X"1421FF5D7FFDEBA085168B45FF843DEBAF7843FFFFF7AABDF55A2AA97400AAD5",
INIT_23 => X"04155EFAA842ABEFA280155EFFFFBC01EF08554000055002AB455D5142010085",
INIT_24 => X"57FD7410552EAAABAAA8017400AAD140000002EBFFEFA2AAA8BEFF780021FF55",
INIT_25 => X"000000000000000000000000000000000000005568A1055043DEBAAAFFE8B455",
INIT_26 => X"8E3DF45155EBD17FF6DAADB504001C71EDA82AAA0955455D556DA00490000000",
INIT_27 => X"101C55554AAAAA480082FF84000BAEBD16DA82410A3FFD7AAA4B8E824971F8E3",
INIT_28 => X"092085F401D71C0A2DBC7EB80000280824ADBD7490E28BEF085157428FFDB420",
INIT_29 => X"DF45AAAA90410BEDF45155A28E2AB7D0051504005D71F8E004975D556DB68405",
INIT_2A => X"28B6D5D51420101C5B401EF417BFAEAA08516AB45E38E38E92EB803FFD7EBA4B",
INIT_2B => X"EAFBC7EB80071FF5500175EFB6802DBC7BE8A155EFE3FBC71FF145B420385500",
INIT_2C => X"0A3FE92BEFFEAB45417FD24385D2AAFA82B68015400AADB40000082EBFFC7A2A",
INIT_2D => X"5557FE1000000000000000000000000000000000000000000000000556FA3849",
INIT_2E => X"AA8428A10085568ABAA2FBD7545AAD17DFFFAAFFC200055557DE00A280155455",
INIT_2F => X"F0051554AAFFFFC00105D55554BAA28400000F784020BAAAD17FE00082EBDF45",
INIT_30 => X"000051575FFF78415410087BC01555D2EBFF55A284000AA08003FF55002AA8BE",
INIT_31 => X"A00A2803DF45AA843DF55AAAE82000F7FBD5545AAAEAABFF0051400105D5568A",
INIT_32 => X"55EF557BC20AA5D042ABFF555142000557FC01EF007FEAABA00556AB55A2AEA8",
INIT_33 => X"C0010082EBDF55A2AABDF45A284175FF5D04175FFF7803DF45FFAE955EFAAFBD",
INIT_34 => X"00000000517FEAA082EBFE10F7FFE8B55087FC00BA552ABFE10F78415400A2FB",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000007FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(14),        -- Port A data input
DOA(0)   => data_read_a_lo_256(14),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(14),        -- Port B data input
DOB(0)   => data_read_b_lo_256(14),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_15_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000A000000000284000280000001800020030000000033022000000180002",
INIT_01 => X"A140098018300848180060000C00426040000000080000080200000000110200",
INIT_02 => X"1020004000801110000006100028503400040800010430004808000180120278",
INIT_03 => X"00008011064408840190800000228002A3000000000010000008108448000042",
INIT_04 => X"701280400004A991000000A28406000211000000220004941000000880000000",
INIT_05 => X"02000484800155020495000800218020C4002880005310000000040000000001",
INIT_06 => X"10000880004540000711224491C08000850A880008000D020001892020656300",
INIT_07 => X"8A04000016050009140501505100000420204008000000BE70408104C8000000",
INIT_08 => X"001F004028026104111002200000000200210040008004614001100801010000",
INIT_09 => X"000800000D09240000800000000000040600180840800022C8088C1020200000",
INIT_0A => X"0000000002004040000105000040042229140002080000000400000080000400",
INIT_0B => X"0000110100000000010000100001000010000000000000000000100000800008",
INIT_0C => X"0001008000000000000025000040000001300008009400006200580010000000",
INIT_0D => X"0000000002300012000000000004200030000000000008008020020000000000",
INIT_0E => X"0000000001000000400000000000000000000010108000000000000010108000",
INIT_0F => X"0000000000000200000900000000000000000010140000000000000010140000",
INIT_10 => X"0140000000000000000001000000400000000000000000000100008040000000",
INIT_11 => X"0000004000480000000000100004400000000030002000406000000000068409",
INIT_12 => X"8000000000020080080000000000802010000000000800000201000800000000",
INIT_13 => X"00000100000000000000000008000000184400A0000000000002000000441108",
INIT_14 => X"4000000000000000010620000004000000000242038B82800000000000000002",
INIT_15 => X"0000000000000000000000000000041800000110000024130202500802000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000080050000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"000804154AA5D00001EFF78428AAA007BC2145F7800000000000000000000000",
INIT_1F => X"0AA007FC2000F7D17DF45AAD157400007BEAAAAAAAE955555D5568A105D7FC00",
INIT_20 => X"FFFFAAAABDEAA557BFDE00FFD140155F7FBD74AAAAD17DF45F7D1421EF005540",
INIT_21 => X"020AAF7FFFDF45FF84000BA552ABDFEF08517DF55A2FBEAB555D556AAAA5D043",
INIT_22 => X"FEAB45F7843FF45082A801FF005155400FFD1420100055574AAA2AA800AAF784",
INIT_23 => X"D5421FF00042ABEFFF8400010082EAABFF55002ABEF087BE8ABA555168B55AAF",
INIT_24 => X"D7BD7545A284020BA007FFFE10A284000AA0055401550055574005D2E800AAA2",
INIT_25 => X"000000000000000000000000000000000000000028B550051574005D7FFFE105",
INIT_26 => X"55D556DA004971C7038140012482550E021C7EB8028A821C7BC516DFF8000000",
INIT_27 => X"45E3DF471C70851400BA0071C5028FFD17FF6DAADB504001C71EDA82AAA09554",
INIT_28 => X"B555D516DA82410A3FFD7AAA4B8E824971F8E38E3DF45155EBF1D5492BED17FF",
INIT_29 => X"54AAAAA480082FF84000BAEBF1FFF7DEB8000092552ABFFEF08517DF6DB6FBE8",
INIT_2A => X"EFA8241516DB55A2FFEAB6DEB843DF551C20801C71C5157428FFDB420101C555",
INIT_2B => X"550428412A85082BEDF401D71C0A2DBC7EB80000280824ADBD7490E28BEF087F",
INIT_2C => X"51504005D71F8E004975D556DB68405092087FF8E00BE8A02082005F47145085",
INIT_2D => X"57BD75EFF78000000000000000000000000000000000000000000000E2AB7D00",
INIT_2E => X"55557DE00A2801554555557FE100055554BA5504000105D2A80145AA842AA005",
INIT_2F => X"5AAD557410F7D57DF55AAFBD55450055420BA0055574BAF7D17DFFFAAFFC2000",
INIT_30 => X"FF08517FFFFF7FBEAB455D517FE00082EBDF45AA8428A10085568ABAA2FBD754",
INIT_31 => X"4AAFFFFC00105D55554BAA28400000F784020BAAAD57FFEFA28402010552ABDF",
INIT_32 => X"FF55002AA8BEF007FFDE1000557DF45AAFBE8BEFA2803FF45550400155555155",
INIT_33 => X"80000087BD55450855400BA002A95400F7FBC01555D2EBFF55A284000AA08003",
INIT_34 => X"000000002EAABFF0051400105D5568A000051575FFF78415410087FEAA10F7AE",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000060000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(15),        -- Port A data input
DOA(0)   => data_read_a_lo_256(15),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(15),        -- Port B data input
DOB(0)   => data_read_b_lo_256(15),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_16_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"DA22C618B1000482B688B186588884862A400438255FC38381441205BA803003",
INIT_01 => X"264AC80028404C211203A952A90341080B173340412000E1005D628000820484",
INIT_02 => X"400034C206C405000001A48202084004003008255040826EE008B440200E2042",
INIT_03 => X"2916704900606AC82B49CC56DF8CC1E50E4800202115005760010010000C0400",
INIT_04 => X"052DCA856DC7504B82BF6614C86D2B7F85AAD17F4B100000B88148C4804A428A",
INIT_05 => X"373CB02A00C0502F301180141A42A5720E0F43C17A8479580001AC20000000E2",
INIT_06 => X"303E2094282B85242C85001038D5710E8410D5959BC4800015001219D0550077",
INIT_07 => X"880100000159954501280B0080146F7112D949A0015018220540000382805001",
INIT_08 => X"30015452880C8D90409A05B2CB2CA400200209E5601044A24000000462A60018",
INIT_09 => X"452D54000C0907000330000000000096480050000685400005FC014743E0DC92",
INIT_0A => X"00014808A02004200E540480212000A448C0080024AEA00C9688000000000005",
INIT_0B => X"000D58460018F6D3D84400044000440004400044000440004400042000220002",
INIT_0C => X"0001004010A8812831605DA0000A054052E40000817680220040025699200002",
INIT_0D => X"AAADA0C343F1AC1B01040A002024895514554485D00000012400240000000000",
INIT_0E => X"AAADA0CC421CA003B694B68018FAAA708E2CB5320018CAC99BA0A3B9320018CA",
INIT_0F => X"B1443A1891E4A928C29020E6A8524CE7A3EE59320018CAC99BA0ACB9320018CA",
INIT_10 => X"04B2A5A40B1E6644AF0F021EA003AC24352AB2449A3FF2FA04E5E09B128834AD",
INIT_11 => X"60ED838E890B703C6260D8E3A21275714C902375B801324301AB0067622E5E54",
INIT_12 => X"064F70DBDB1C74424E91E1C194C71D1216F50A8C241815FEB6A9158863F638FB",
INIT_13 => X"45FDF9D364DBD9435A6D45C9E81BED555E4C15F11133D171727A2550EE2F1BA0",
INIT_14 => X"08150013F162119014204373517700ACCC59432A2B2D001F803471A9A960E572",
INIT_15 => X"000000000000000000000000000000880002054000229088542210206B2AB015",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"2A898D21B4C98389ED146C080000000000000000000000000000000000000000",
INIT_19 => X"A29A29A29A29A29A29A29A29A29A28A28A28A28A28A53CBF0F0D3CF3CF0AB1A2",
INIT_1A => X"8F47A3D1E8F4FA7D3E9F4FA7D3E9F4FA7D3E8F4FA3D3E8F4FA3D3E9A29A29A29",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000FA7D3E9F4FA7D1E8F47A3D1E",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFF7FBE8B45AAD568BFFFFAA975FF00003FE0055000000000000000000000000",
INIT_1F => X"0005D2A95410FFFFC00000804154AA5D00001EFF78428AAA007BC2145F7843FF",
INIT_20 => X"7400007BEAAAAAAAE955555D5568A105D2E974BAF7FBEAB45FFFFC00BAF78002",
INIT_21 => X"C2000F78000010552E800AA002E821FFA2AAAAA00000417555FFD17DF45AAD15",
INIT_22 => X"43FEBA5D55575FFF7AABFE00557BD74AAAAD17DF45F7D1421EF0055400AA007F",
INIT_23 => X"D56AAAA5D043FFFFAAAABDEAA557BFDE00FFD140155F7AABDF55F7AE820AA080",
INIT_24 => X"8517DF55A2FBEAB555D04154BAA2FBE8B55FFFFD55FF557FC2000FF8015410FF",
INIT_25 => X"000000000000000000000000000000000000007FFDF45FF84000BA552ABDFEF0",
INIT_26 => X"21C7BC516DFF8438FC7E3F1EAB55B6DF6DBFFF7AA955C71C043FE10490000000",
INIT_27 => X"55FFF1C70BAF78A000005D2097438FFF1C7038140012482550E021C7EB8028A8",
INIT_28 => X"57DEBD17FF6DAADB504001C71EDA82AAA0955455D556DA00492490492F7FBE8B",
INIT_29 => X"71C70851400BA0071C5028FF84020285D2085092002A801FFB6AAA8A10080E17",
INIT_2A => X"BAF6DE3AA8709208043FEBA555B555FFE3AABFE005D71D5492BED17FF45E3DF4",
INIT_2B => X"BC0028E38412428EBD16DA82410A3FFD7AAA4B8E824971F8E38E3DF45155EBA4",
INIT_2C => X"8000092552ABFFEF08517DF6DB6FBE8B555D04124BAB6FBE8B45E3FBD55D7557",
INIT_2D => X"5003DE000000000000000000000000000000000000000000000000071FFF7DEB",
INIT_2E => X"5D2A80145AA842AA00557BD75EFF78428B55AAD168B55F7FFFDFEFFFAA955555",
INIT_2F => X"0000000010F7FBEAB45FFD1554AAFFAE820105500154AAF7D5554BA550400010",
INIT_30 => X"EFF7AEA8A10002E955FFA2D17DFFFAAFFC200055557DE00A2801554555557FE1",
INIT_31 => X"410F7D57DF55AAFBD55450055420BA0055574BAF784000BA5D0017410082E801",
INIT_32 => X"8ABAA2FBD7545AA802ABEFA2AA9541000003DEBA557BD75EFA2AEBDE105D5557",
INIT_33 => X"EAB45AAFFD55555D7FC20AAA280000AAAAD17FE00082EBDF45AA8428A1008556",
INIT_34 => X"00000000557FFEFA28402010552ABDFFF08517FFFFF7FBEAB455D04020AAFFFB",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000020000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(16),        -- Port A data input
DOA(0)   => data_read_a_lo_256(16),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(16),        -- Port B data input
DOB(0)   => data_read_b_lo_256(16),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_17_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"5284CE4FB7BD2C8994A13392DBD02E14006B82AC7E800D44D3DD2FD5F9B961C0",
INIT_01 => X"F9BA301F7E03FC6793F2199B39FC233C11D93AE6F3BB92B32091DBC339B24542",
INIT_02 => X"1D5FC0C08F040404446965C0607FB8A217C400C33A908078551BD04222186338",
INIT_03 => X"A14124C28DFD960832C90446DF8400A5055C25295B695FF97E1B5AC757F06D6B",
INIT_04 => X"04A106866DA3D02A01FB660C08A4AB7F840EDB6F48100DFC8081081D78AC7402",
INIT_05 => X"51E072F0C0C58D9C125EBFC00A46CF0388054100F680E0CE0107B8D040DAFCDA",
INIT_06 => X"019A4D00786B048112C58B16307F15DE8408B233661C10BBA5DAAFA9DDA1194D",
INIT_07 => X"8E00001660700CE170284A00891C7C03D29DE26814515835902AC089A2801540",
INIT_08 => X"C009F3A1B0120A1C51DFF881861CBE0305A12A0321810217C01D34EDC98FFA1C",
INIT_09 => X"747E6610052CDEE97FF1F9F63E3EF790380078002CE976AB6BF769769E4D437D",
INIT_0A => X"00185C44B91BC1740B7605040BE0018CFC7429F326B9D045FF8000E9AB415606",
INIT_0B => X"3A28FC1AAF5CF6F3D3EF3D3EF3D3EF3D3EF3D3EF3D3EF3D3EF3D3EF9E9F79E9E",
INIT_0C => X"0000020012E9E10A31EB5FF9296A67F5B4FFBD2FAD7FE653C3FBFF33E10C001B",
INIT_0D => X"333EA16031F2BD47BDA2CA5D8164FCCFE833C5C3D00018006C68170000000000",
INIT_0E => X"333EA160391BEFF2C32FB695F919110D5ECE542A6FEEB2533EA160782A6FEEB2",
INIT_0F => X"D18C0D06638A207CFDE1F7DDAD76D5282400F82A6FEEB2533EA160782A6FEEB2",
INIT_10 => X"E6E43E59AFE4A59B57679D19EFF2C7573FAD5A86840354D1706FFFA3EF6E24B6",
INIT_11 => X"F7D7A0ABD6DAAAB96529382B74E4E1FE4ACA4D77FAAB77CE3AF3EE78F58DB737",
INIT_12 => X"2D1281017F056E9C9C3FC95949C157ADB55572CA52606DFED6CA55334C04C04F",
INIT_13 => X"59FDEB974F486905001FDF5FA0D719F9956EAA1A184045D5D7A870D2F5A5D752",
INIT_14 => X"60158015177F916A039EF41FDB34A91F432EA58949D5B5C85F97871876F7D7E8",
INIT_15 => X"000000000000000000000000000004DC200005E705B7B3D9FC22F00BE419FB55",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"06013DB9880A5D22E229F3030018000000000000000000000000000000000000",
INIT_19 => X"D35D74D35D74D34D35D74D35D74D34D34D34D34D34D0D30D0D303AEBAE886E40",
INIT_1A => X"51A8D46A351A0D068341A0D068341A0D068341A8D468341A8D46834D35D74D34",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000008D46A351A8D46A351A8D46A3",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFF7FBFDF55A28402000F7D56ABFF55000000000000000000000000",
INIT_1F => X"A00F7843FEBA55043FFFFF7FBE8B45AAD568BFFFFAA975FF00003FE0055043FF",
INIT_20 => X"54AA5D00001EFF78428AAA007BC2145F7D568B45000002010552EBDF45A28028",
INIT_21 => X"95410FFAE800105D2A95410002A95410AAAEBFF55AAFFC00BAF7FFC000008041",
INIT_22 => X"57DE00F7AE800AAAAAABDFEF5D2E974BAF7FBEAB45FFFFC00BAF780020005D2A",
INIT_23 => X"517DF45AAD157400007BEAAAAAAAE955555D5568A105D7FFFFEFA2D568BFFFFD",
INIT_24 => X"2AAAAA00000417555FF8028B55082A974105D003FF55F7802AAAAAAD168AAA5D",
INIT_25 => X"000000000000000000000000000000000000000000010552E800AA002E821FFA",
INIT_26 => X"71C043FE10490A3FFFFFFFFFDFEFE3F5FAF45AA8000038F7DB6FBD7490000000",
INIT_27 => X"384124BFF7DB68A28A38F7803DE82490438FC7E3F1EAB55B6DF6DBFFF7AA955C",
INIT_28 => X"0BAFFF1C7038140012482550E021C7EB8028A821C7BC516DFFDF68B551C0E050",
INIT_29 => X"70BAF78A000005D2097438FFAA85000492495428082E95400AAA0BDF7DB6F5C7",
INIT_2A => X"FAFFFB6D56FBFFEBDB78E38F7AA800BAB6AEBDFD75D2490492F7FBE8B55FFF1C",
INIT_2B => X"028AAAB6D16FA8249517FF6DAADB504001C71EDA82AAA0955455D556DA00497F",
INIT_2C => X"2085092002A801FFB6AAA8A10080E1757DEB8A2DB5514249243841003FF6DEB8",
INIT_2D => X"7FFFDF550000000000000000000000000000000000000000000000004020285D",
INIT_2E => X"F7FFFDFEFFFAA9555555003DE00002ABFFEFF7FBFDFFFAAD168B55AA80000BAF",
INIT_2F => X"FF7FBEAB45552E954BA08003DFFFFFAAA8AAAF7843FE10000428B55AAD168B55",
INIT_30 => X"10AA843FFFFF7D5554BAF7D5554BA5504000105D2A80145AA842AA00557BD75E",
INIT_31 => X"010F7FBEAB45FFD1554AAFFAE820105500154AAF7AE974000800154AA002E954",
INIT_32 => X"554555557FE10007FEABEFFFD57FFEFAAFFE8ABAFFAA820BAF7AEBFF55550000",
INIT_33 => X"020AA08003DFFFA28028AAAF7D17DE0000517DFFFAAFFC200055557DE00A2801",
INIT_34 => X"0000000004000BA5D0017410082E801EFF7AEA8A10002E955FFA2AABFF455500",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000067FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(17),        -- Port A data input
DOA(0)   => data_read_a_lo_256(17),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(17),        -- Port B data input
DOB(0)   => data_read_b_lo_256(17),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_18_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"69844019080000A21A611406840014122A641074155FC28A2024001001801003",
INIT_01 => X"01067920034004180005E9E3C90360C0041C0181002001602025800008440084",
INIT_02 => X"40AC3CAA22D605200000856E2481902400344A20F802C22054001000021E2379",
INIT_03 => X"A95308ECD3207AC81D91C4002004C08A06008080BA868007E58040102B0E0100",
INIT_04 => X"044CC183800CA00780808004C8DB841405A80A100B586200FAC24AE4805242CA",
INIT_05 => X"771C10000000000B1135883C08A115320E0401C0200038394230070A19000020",
INIT_06 => X"3001499C602A8A003E800A042D8132A00098408F79E3901218050018024110D6",
INIT_07 => X"5029401000C983E60004010030400353C05806800104004E0000042E52800E20",
INIT_08 => X"0000117088080990419005B0C309402030060860E01004A828408800440405E3",
INIT_09 => X"6B8186185C42900693A002004040001E1950850C848601008708114A2030B480",
INIT_0A => X"100180A8062026000DC425C0301311324AA237108857220BA089420440000030",
INIT_0B => X"C44703657083080C2800C2000C2000C2000C2000C2000C2000C2000610006100",
INIT_0C => X"C1B0609C05013065CC042004040808084001E000108010230400800FD9B286C4",
INIT_0D => X"CCC15F9CBA45505640000A402019003F140FC2060014250B9080008306C18360",
INIT_0E => X"CCC15F9FB1962FCB69E08AAAEAEBCDDF7C728582081483ACC15F9C3982081483",
INIT_0F => X"EBF1CFFF7670ACC3811A28AB57523CDFEBFBF982081483ACC15F9F3982081483",
INIT_10 => X"C9002BF05800D875E63CC9962FCB52CAA02FE3F8E7F5E3AC3620805298B15A3F",
INIT_11 => X"F1B72A8A800B7546DB9F1CA320037F01BD67DC4041D4CF03138DD865103EFEEA",
INIT_12 => X"81CCFAFDBF9464006FD037AEFAE5150016EA8DB7BFE25208E8F46A228BF8A757",
INIT_13 => X"641256EC844B8AF92FD7CEDC24A9E181A8A29509EAAE7FD3B749471C48F8A459",
INIT_14 => X"0297D086E00036D2440E0880AAD62BEFF5778802A3AF8E8FB0440CE78773B709",
INIT_15 => X"8360D8360D8360D8360D8360D83609220D20D00000080C0601400B402307E480",
INIT_16 => X"360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D",
INIT_17 => X"60D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8",
INIT_18 => X"D9D701DC2E784601EFBE2C00000000000000000000000008360D8360D8360D83",
INIT_19 => X"5155555545145145155555545145145145145145145220B22A0B820820965177",
INIT_1A => X"44A25128944A25128944A25128944A25128944AA552A954A2512895554514514",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000025128944A25128944A251289",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFEFF7AE954BA5D04174AA00000000000000000000000000",
INIT_1F => X"145AA801741000043FFFFFFFFFFFFFF7FBFDF55A28402000F7D56ABFF55043FF",
INIT_20 => X"8B45AAD568BFFFFAA975FF00003FE0055043FFFFFFFFFDFEFA2D56AB45AA8400",
INIT_21 => X"3FEBA55557FFEFA2D168B55AAFBFFFFFFF80021EF0855421EF00043FFFFF7FBE",
INIT_22 => X"A82155F7AEBFEBAFFD56AA00A2D568B45000002010552EBDF45A28028A00F784",
INIT_23 => X"FFC00000804154AA5D00001EFF78428AAA007BC2145F7D5400000004020AA5D2",
INIT_24 => X"AAEBFF55AAFFC00BAF7AE80010082E954BA0004174AAAA8428B45082ABFEBAA2",
INIT_25 => X"000000000000000000000000000000000000002E800105D2A95410002A95410A",
INIT_26 => X"8F7DB6FBD7490E3FFFFFFFFFFFFFFFFBFDFEFFFAE954AA550415492140000000",
INIT_27 => X"D7AAD16FB6DBE8E00155BE8015410140A3FFFFFFFFFDFEFE3F5FAF45AA800003",
INIT_28 => X"1C7140438FC7E3F1EAB55B6DF6DBFFF7AA955C71C043FE1049043FFEFE3F1F8F",
INIT_29 => X"FF7DB68A28A38F7803DE82495B78FC7AAD56FB6DBEF1FAFD7E384001EF145B47",
INIT_2A => X"420381C0A02082492A85155E3A4BDE92FFD56FA28B6DF68B551C0E050384124B",
INIT_2B => X"E28B7D1420BDEAAA2F1C7038140012482550E021C7EB8028A821C7BC516DFFD1",
INIT_2C => X"2495428082E95400AAA0BDF7DB6F5C70BAFFAE870280024904BA1400174AABE8",
INIT_2D => X"50415410550000000000000000000000000000000000000000000002A8500049",
INIT_2E => X"AAD168B55AA80000BAF7FFFDF55002ABFFFFFFFFFFFEFF7FBFDFFFF7AA974BA5",
INIT_2F => X"000043DFEFA2D56AB45AAD57DFEFF7AA82155F78015400552ABFFEFF7FBFDFFF",
INIT_30 => X"55A280021EF557FD7555550428B55AAD168B55F7FFFDFEFFFAA9555555003DE0",
INIT_31 => X"B45552E954BA08003DFFFFFAAA8AAAF7843FE10007FEAB55A2D17FFEFFFD568B",
INIT_32 => X"AA00557BD75EFF7D1400AA5D2A82000002A95545A2843FE00F7D17FEAAF7FBEA",
INIT_33 => X"020AA5D04154BAF7AEA8BEF55003DEAAA2D5554BA5504000105D2A80145AA842",
INIT_34 => X"000000002E974000800154AA002E95410AA843FFFFF7D5554BAF7AE974BA0004",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000020000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(18),        -- Port A data input
DOA(0)   => data_read_a_lo_256(18),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(18),        -- Port B data input
DOB(0)   => data_read_b_lo_256(18),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_19_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"042200000000000041088001001AA00000000000000000000000500802000003",
INIT_01 => X"074018000024000000000404000000000A22000800000800004A200000000001",
INIT_02 => X"0000048002C405000000000006A84000000000200893C246A20000000020031A",
INIT_03 => X"020A9639044012C80001C4000004C08006000000001025000000000000000000",
INIT_04 => X"0400C0800000000380800004C8000000058800000B1000009880480480024200",
INIT_05 => X"420410000000000B10804004080001320E0401C0200038080000000000000000",
INIT_06 => X"2002409006F00A8428050A000280493104004500480090080A01120220140020",
INIT_07 => X"0000000000418026090240923240002190400000000000C0054A912054004021",
INIT_08 => X"0000115080000990000000B0C308000000000860200160000000000038380000",
INIT_09 => X"8000F80001012590001000000000001618000000020280008180810200000000",
INIT_0A => X"0000000000000000000000000000000100008000110000000000000000000017",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000840007600000000000000000800259000000",
INIT_0D => X"0008A0034078104B41A41000000000031400C002000000000000000000000000",
INIT_0E => X"0008A0004263C0343EDD414004042228DC0D385598035D0008A003B05598035D",
INIT_0F => X"040231068187C39F5A4F985C008902041124505598035D0008A000B05598035D",
INIT_10 => X"1BFBD406451B02000E033263C0343CB740500401180DE053A98F6ECC739D8140",
INIT_11 => X"420851546B2400000040D8549B5800000010227848D4303807FC8CC5508AEAED",
INIT_12 => X"52210402120A936B0000000004C2A8D6480000000018A700FCF980CC300318A2",
INIT_13 => X"B1427ED430B41402D025082359700181C21140E40511802208D6B30C48F8A8A4",
INIT_14 => X"9C000018440021011821B35254E99AF9E9410006362A2B6424287B08286208D6",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000023006000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"7747E18E0218CC18E88324000000000000000000000000000000000000000000",
INIT_19 => X"34C30C30C30C30D34C30C30C30C30C30C30C30C30C3504118982A69A6980E411",
INIT_1A => X"C26130984C26130984C26130984C261309A4D26130984C26130984C30C30C30D",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000130984C26130984C26130984",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAA954BA5500020BA5D000000000000000000000000",
INIT_1F => X"4BA5D517FFFF08043FFFFFFFFFFFFFFFFFFFFEFF7AE954BA5D04174AA007BFFF",
INIT_20 => X"FFFFF7FBFDF55A28402000F7D56ABFF557BFFFFFFFFFFFFFFFFFBFDFEFFFAA97",
INIT_21 => X"17410007BFFFFFFFFFFFFEFF7D16AB45AA8002000F7D5575455D043FFFFFFFFF",
INIT_22 => X"568B55F7AE955FFAA840201008043FFFFFFFFFDFEFA2D56AB45AA8400145AA80",
INIT_23 => X"043FFFFF7FBE8B45AAD568BFFFFAA975FF00003FE00557BFFFFFFFFBFDF45AAD",
INIT_24 => X"F80021EF0855421EF002ABFFEFF7D168B55AAD17FFEFF7AE975FF00557FFFF5D",
INIT_25 => X"00000000000000000000000000000000000000557FFEFA2D168B55AAFBFFFFFF",
INIT_26 => X"A5504154921471FFFFFFFFFFFFFFFFFFFFFFFF7AA954BA550000082550000000",
INIT_27 => X"EFF7FBFAFD7E3A4954BA555B7AFC7080E3FFFFFFFFFFFFFFFFBFDFEFFFAE954A",
INIT_28 => X"545550A3FFFFFFFFFDFEFE3F5FAF45AA8000038F7DB6FBD74975FFFFFFFFFFFF",
INIT_29 => X"FB6DBE8E00155BE8015410147FFFFFFF7FBF8FC7EBD568B55A28000000FFDF52",
INIT_2A => X"FDFC7E3F1FAF55A2DB6FB7DF7AE955C7BE800000008043FFEFE3F1F8FD7AAD16",
INIT_2B => X"0955FF145B7AFC7410438FC7E3F1EAB55B6DF6DBFFF7AA955C71C043FE10497B",
INIT_2C => X"D56FB6DBEF1FAFD7E384001EF145B471C71424B8FC7E3D56AB6DB6DF7AFC7EBA",
INIT_2D => X"50002000550000000000000000000000000000000000000000000005B78FC7AA",
INIT_2E => X"F7FBFDFFFF7AA974BA55041541055517FFFFFFFFFFFFFFFFFFFFEFF7AA974AA5",
INIT_2F => X"500517FFFFFFFBFDFEFFFFFEAB45AA80154AA557BEAB45002ABFFFFFFFFFFFEF",
INIT_30 => X"55A28002000F7FFC2155552ABFFEFF7FBFDFFFAAD168B55AA80000BAF7FFFDF5",
INIT_31 => X"FEFA2D56AB45AAD57DFEFF7AA82155F78015400557BFDFEFF7FBEAB55A2D56AB",
INIT_32 => X"555555003DE00007FFDF45AAD568B45AAFBFFFFFFFAA95545F7840201000043D",
INIT_33 => X"6ABFFFFFBEAB45A280155EF557FE8B55000428B55AAD168B55F7FFFDFEFFFAA9",
INIT_34 => X"000000007FEAB55A2D17FFEFFFD568B55A280021EF557FD755555042AB55AAD1",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000040000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(19),        -- Port A data input
DOA(0)   => data_read_a_lo_256(19),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(19),        -- Port B data input
DOB(0)   => data_read_b_lo_256(19),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_20_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000003",
INIT_01 => X"A65FF80000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000048002CC070000000000000000000000002FF86100200000000220002362",
INIT_03 => X"00000000000203D80025DC18004DC3D01E000000000000000000000000000000",
INIT_04 => X"07E5DF808071026F87C4191DD8005080679800000F300002998058068002C000",
INIT_05 => X"C205F23A2100557F70000004390021F61E1E87C3FD0CFBF80880072042000044",
INIT_06 => X"1209244C2000100006800000020010000008407FC800B0000000100600040000",
INIT_07 => X"8802000009FFBFE51886018002040020000800000554003E0000000002800000",
INIT_08 => X"30801F5780259FB0000000F7DF78020004011FEFE00000000020031502000083",
INIT_09 => X"00000000001000000000000000000056F8000001000000040000040141800802",
INIT_0A => X"0000000000000008000800000000000000000000000000000010010014800000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"00010240001721214E000004000000080000008000001000040080FFDB000000",
INIT_0D => X"0000000F3008001E00000000001803FF14FFC006000000008010200000000000",
INIT_0E => X"0000000F3040200000020000000026A70C0008020000200000000F3002000020",
INIT_0F => X"000030B86000400080000200000000004A58F0020000200000000F3002000020",
INIT_10 => X"0000000002183E61E6000040200001000000000019B140000800800000020000",
INIT_11 => X"C00010080000000000525801000000000014AC08000000508001030A0A400100",
INIT_12 => X"000002BC360020000000000292C0100000000000A56000090100000000001F86",
INIT_13 => X"8010000000000000574500001001060600000000001716800000803102020000",
INIT_14 => X"00000000000040040040002000080506049CDF70C08040100000706707600000",
INIT_15 => X"00000000000000000000000000802040200200604040000000000024FB7FE008",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"060070400020112240209A408004000000000000000000000000000000000000",
INIT_19 => X"65965965965965965965965965965861861861861860D30424343CF3CF340E00",
INIT_1A => X"90C86432190C86432190C86432190C86432190C86432190C8643219659659659",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000086432190C86432190C864321",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974AA55040201008000000000000000000000000",
INIT_1F => X"4AA550002000007BFFFFFFFFFFFFFFFFFFFFFFFFFAA954BA5500020BA5D7FFFF",
INIT_20 => X"FFFFFFFFFFFEFF7AE954BA5D04174AA00003FFFFFFFFFFFFFFFFFFFFFFF7AA97",
INIT_21 => X"7FFFF087FFFFFFFFFFFFFFFFFFFFDFEFFFAE974AA5D003FE005D043FFFFFFFFF",
INIT_22 => X"BFDFFFAA84000105D556AB55557BFFFFFFFFFFFFFFFFFBFDFEFFFAA974BA5D51",
INIT_23 => X"043FFFFFFFFFFFFFF7FBFDF55A28402000F7D56ABFF55003FFFFFFFFFFFFFF7F",
INIT_24 => X"A8002000F7D5575455D2EBFFFFFFFFFFFEFF7FBEAB55A28000010F7D16ABEF08",
INIT_25 => X"000000000000000000000000000000000000007BFFFFFFFFFFFFEFF7D16AB45A",
INIT_26 => X"A550000082557FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550400028000000000",
INIT_27 => X"FFFFFFFDFEFF7AE974BA5500050380071FFFFFFFFFFFFFFFFFFFFFFFF7AA954B",
INIT_28 => X"E285D0E3FFFFFFFFFFFFFFFFBFDFEFFFAE954AA55041549214043FFFFFFFFFFF",
INIT_29 => X"AFD7E3A4954BA555B7AFC70871FFFFFFFFFFFFFFF7FBFDFFFFFAA974BA550038",
INIT_2A => X"3FFFFFFFFFDFEFF7F1FAFC7A28002028555F6FB7D5D75FFFFFFFFFFFFEFF7FBF",
INIT_2B => X"402010FFDB6ABEF140A3FFFFFFFFFDFEFE3F5FAF45AA8000038F7DB6FBD7490E",
INIT_2C => X"FBF8FC7EBD568B55A28000000FFDF525455524BFFFFFFFBFDFC7E3F5E8B45A28",
INIT_2D => X"504000BA080000000000000000000000000000000000000000000007FFFFFFF7",
INIT_2E => X"FFFFFFFEFF7AA974AA550002000557FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5",
INIT_2F => X"055043FFFFFFFFFFFFFF7FBFDFEFFFAE954BA5500174AA08517FFFFFFFFFFFFF",
INIT_30 => X"EFF7AE974AA550028AAA5D2ABFFFFFFFFFFFEFF7FBFDFFFF7AA974BA55041541",
INIT_31 => X"FFFFFFBFDFEFFFFFEAB45AA80154AA557BEAB4500557FFFFFFFFFDFEFF7FFFFF",
INIT_32 => X"00BAF7FFFDF55002EBFFFFF7FBFDFEFFFD568B55A284020BA557FFFFFF5D517F",
INIT_33 => X"FFF55A2D16AB45AA8402000F7FBEABEF5D2ABFFEFF7FBFDFFFAAD168B55AA800",
INIT_34 => X"000000007BFDFEFF7FBEAB55A2D56AB55A28002000F7FFC215555043DFEFF7FB",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000007FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(20),        -- Port A data input
DOA(0)   => data_read_a_lo_256(20),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(20),        -- Port B data input
DOB(0)   => data_read_b_lo_256(20),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_21_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"4A302428B824900A128C090A5C1800261500213C005FE812D10420054085A202",
INIT_01 => X"081FFE3440B609703B0427F801A40B8115BC4F655300340288A40D30040E4DD8",
INIT_02 => X"04CA478082CC1740002019824E0203100640303FF8C0B31061096E21A1840814",
INIT_03 => X"230CA7A4810083F80095DE00102DC3823EA821094EC68248923200013290C800",
INIT_04 => X"07CFFFC04904AA7F8780409DF84A0202879800000F3000029980780EA2C3C002",
INIT_05 => X"DE87F0280000407FF900D914382091FE1E1C0FC3E01EFFF8000480200008D062",
INIT_06 => X"010E2182002BC107A03448808F0D7C002822987FC830F40134CC74D002016612",
INIT_07 => X"0401000011FBFFE00520000200422033025C4209104500000012004C004D8C0B",
INIT_08 => X"00EF1F5FA0041FF080AC70FFDF78220010841EFFE7116E144071268DFD3E4C24",
INIT_09 => X"FC8BFE18008083B4443151462A28C6DFF80010002605302248088950484550A3",
INIT_0A => X"10018C241102068006C620C03882019480E631A0855E924E2598038938404037",
INIT_0B => X"A641165448C80C103648A3648A3648A3648A3648A3648A3648A366451B2451B2",
INIT_0C => X"011100841200D001000624000100C002804A08221890004806A310FFDF000454",
INIT_0D => X"5004D8158809C86065941840B1014FFF56FFC0281280080180B2948004400220",
INIT_0E => X"5004D815810D42E04A08A80098C02450025360694101816002D41A4068C10181",
INIT_0F => X"134160C8125B0B271802242880A04482418A0068C101816002D41A4069410181",
INIT_10 => X"10080E05C0B06AA8B12CFD0D42E0441A300012682960828F05C96A001B029010",
INIT_11 => X"00010362A8A20826A88660D86B202049F115100920C54E8EA256ECF078BA081C",
INIT_12 => X"064802C0081B0D64040936443306C55144104F30A8801406D002900062803201",
INIT_13 => X"4581BA0038005A706680012280506A8010602011819E290048A2118EC8140C08",
INIT_14 => X"CC158092C044600466208CC5091011C322A4C40A0300600C0A80509F41800880",
INIT_15 => X"80200802008020080200802008020412002001000000381C02004000FBFFF80D",
INIT_16 => X"0200802008020080200802008020080200802008020080200802008020080200",
INIT_17 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_18 => X"FDDFEFFFBEFFE7C7BFBEFC000000000000000000000000080200802008020080",
INIT_19 => X"F7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7FFBFBFFF9E79E7FFFDF3",
INIT_1A => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFDFEFF7FBFDFEFF7FBFDF7DF7DF7D",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00001FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D000200008000000000000000000000000",
INIT_1F => X"4AA5D00020AA5D7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550402010087FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAA954BA5500020BA5D7FFFFFFFFFFFFFFFFFFFFFFFFFFAE95",
INIT_21 => X"0200000003FFFFFFFFFFFFFFFFFFFFFFF7AA974BA5D0402000557BFFFFFFFFFF",
INIT_22 => X"FFFFEFF7AE974BA5D00174BA00003FFFFFFFFFFFFFFFFFFFFFFF7AA974AA5500",
INIT_23 => X"043FFFFFFFFFFFFFFFFFFFFEFF7AE954BA5D04174AA00003FFFFFFFFFFFFFFFF",
INIT_24 => X"FAE974AA5D003FE005D2EBFFFFFFFFFFFFFFFFFFDFEFF7AE954AA5500174BA5D",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFDFEFF",
INIT_26 => X"A550400028007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0000010000000000",
INIT_27 => X"FFFFFFFFFFFFFAA954BA5D00000BA557FFFFFFFFFFFFFFFFFFFFFFFFFFAE974A",
INIT_28 => X"0005571FFFFFFFFFFFFFFFFFFFFFFFF7AA954BA550000082557BFFFFFFFFFFFF",
INIT_29 => X"DFEFF7AE974BA55000503800003FFFFFFFFFFFFFFFFFFFFEFF7AA974AA5D0405",
INIT_2A => X"3FFFFFFFFFFFFFFFFFFDFEFF7AE954BA5D00154AA00043FFFFFFFFFFFFFFFFFF",
INIT_2B => X"A974BA5D00104925D0E3FFFFFFFFFFFFFFFFBFDFEFFFAE954AA550415492140E",
INIT_2C => X"FFFFFFFF7FBFDFFFFFAA974BA550038E285D2ABFFFFFFFFFFFFFFFFBFDFEFFFA",
INIT_2D => X"D00000100000000000000000000000000000000000000000000000071FFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE954AA5504000BA087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0557BFFFFFFFFFFFFFFFFFFFFFFFF7AA954BA5D00000BA5D7FFFFFFFFFFFFFFF",
INIT_30 => X"EFF7AE954AA5D041740055517FFFFFFFFFFFFFFFFFFFFEFF7AA974AA55000200",
INIT_31 => X"FFFFFFFFFFFFF7FBFDFEFFFAE954BA5500174AA08043FFFFFFFFFFFFFFFFBFDF",
INIT_32 => X"74BA550415410552ABFFFFFFFFFFFFFF7FBFDFFFFFAA974AA5D00174BA08043F",
INIT_33 => X"FDFEFF7FBFFFFFF7AE954BA5D0000010552ABFFFFFFFFFFFEFF7FBFDFFFF7AA9",
INIT_34 => X"00000000557FFFFFFFFFDFEFF7FFFFFEFF7AE974AA550028AAA5D2EBFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(21),        -- Port A data input
DOA(0)   => data_read_a_lo_256(21),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(21),        -- Port B data input
DOB(0)   => data_read_b_lo_256(21),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_22_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"5290F4CDE914905A14A43D33F488243E17122300F55FEB189B343A1140548380",
INIT_01 => X"A94007B259F6A975386262000C344BA9573C6FF57B18A5FB0ABFCD3C2C5F4F0C",
INIT_02 => X"D56B4302AC01005111011BD506AA5205274056900596A539584E2E6DFE4B2418",
INIT_03 => X"9AC0FCBD854688207C90007A1000047A00E588632CA213C8903AD6B55AD0EB5A",
INIT_04 => X"30002047A6FCA110086C402022F2124A8022492580040440002021C922D9109B",
INIT_05 => X"14A206B6838151008D95DD1847811C08002380041F1104002205AC4140DAD060",
INIT_06 => X"1727FF2EB9EF113A10BD32F44289D1F840C1710010344DB9A808FDFF3DE03130",
INIT_07 => X"050700154A00401D00495A06A8D464C5F6B54AA8551040818F4C997AC80CBE05",
INIT_08 => X"0141008801018040E48D50080002B00A0C00801014541E9504703680017F6CB4",
INIT_09 => X"02680000010937986481514E2A29CE010708C0804C6A033F7FCFF9426A41F1AB",
INIT_0A => X"00500001840000C80B410014088040F4A944B1AA313C004554002381B8000500",
INIT_0B => X"A004D1594832824A070AA070AA070AA070AA070AA070AA070AA0725503855038",
INIT_0C => X"501428054278142151262CA50343854E506A2C6898B2950AA6A35B0004284058",
INIT_0D => X"90078E1F840A2B0114020104022460002200050F60E220A06880D2A14050A028",
INIT_0E => X"90078E1F891C239F8908003099C1ACF06273612B3482C0C0078E1F412B1582C0",
INIT_0F => X"1BA1B0FD16770236A4091621C08055C2C0DB012B1582C0C0078E1F412B3482C0",
INIT_10 => X"00101F09C030AB28B03C111C239F870828041BA859F213AFC14AA38043006018",
INIT_11 => X"10E8822A984B0025B0DE6089462660095337B08AA600CA88B143AB11880C2806",
INIT_12 => X"055412D4481128C4CC012A66F304553096004B61BD8068B92400D0004E303689",
INIT_13 => X"589C48082C006A9057CA4385809520F07830001AC2173B00E162563454C40804",
INIT_14 => X"00460848952220592745AC11A544B1BF006850840180A00E1C81900C4190E160",
INIT_15 => X"22088220882208822088220882208CD888088D940D2A3A9D5002001300800C8C",
INIT_16 => X"0080200882208822088220882208822088220882208822088220882208822088",
INIT_17 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_18 => X"FBDFD1FE3EFBD7BBEFBEFA0A245120000000007FFFFFFFF20080200802008020",
INIT_19 => X"F3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF7FFBFAFBBBEFBEFBEFBF7",
INIT_1A => X"CFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCF3CF3CF3C",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000007F3F9FCFE7F3F9FCFE7F3F9F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040000000000000000000000000000000",
INIT_1F => X"4BA550000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0002000087FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974AA550402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"020AA5D7FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5D00000AA007FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAA954BA5504000AA557FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5D00",
INIT_23 => X"7BFFFFFFFFFFFFFFFFFFFFFFFFFAA954BA5500020BA5D7FFFFFFFFFFFFFFFFFF",
INIT_24 => X"7AA974BA5D040200055517FFFFFFFFFFFFFFFFFFFFFFFFAA954BA5500000BA5D",
INIT_25 => X"00000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000080000000",
INIT_27 => X"FFFFFFFFFFFFFAE974AA550002010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"0BA087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550400028007FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAA954BA5D00000BA557FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5D0002",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAA954BA5504020AA5D7BFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"A974AA5D00070925D71FFFFFFFFFFFFFFFFFFFFFFFF7AA954BA5500000825571",
INIT_2C => X"FFFFFFFFFFFFFFEFF7AA974AA5D040500055517FFFFFFFFFFFFFFFFFFFFFFF7A",
INIT_2D => X"D040200008000000000000000000000000000000000000000000000003FFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"A087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550002000087FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAA954AA5D00020AA007FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5504000B",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFF7AA954BA5D00000BA5D7BFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"74AA55000200055517FFFFFFFFFFFFFFFFFFFFEFF7AA974BA5504020BA557BFF",
INIT_33 => X"FFFFFFFFFFDFEFF7AE974AA5D00154105D517FFFFFFFFFFFFFFFFFFFFEFF7AA9",
INIT_34 => X"00000000043FFFFFFFFFFFFFFFFBFDFEFF7AE954AA5D041740055557FFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000007FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(22),        -- Port A data input
DOA(0)   => data_read_a_lo_256(22),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(22),        -- Port B data input
DOB(0)   => data_read_b_lo_256(22),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_23_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"EF20906D902424807BC8241BC81801B97D38AD3C0800103362A6741C80A12A02",
INIT_01 => X"001FFF8409F089003B4422000D80C80106804A7951C5B9D1C828043EA28838F9",
INIT_02 => X"028406A002DC176444683862400003111001303FFC00F240D50146013B300500",
INIT_03 => X"0006C90C010203F80005DC00C52FC380BEAC25886C02034800200200A1008008",
INIT_04 => X"17DFFF8049000BFF878314BFF8488890979800002F702002BB807A068403C280",
INIT_05 => X"DA07F0000000007FF020C814380011FE5E1C2FC3E05FFFF90020000808900010",
INIT_06 => X"10004C9690A8CA008024685184097E81E872C8FFE900FC31348EFDF03BE15E22",
INIT_07 => X"402000001FFBFFFD00080200B8140011F0D8C108155542018D1A302193E94004",
INIT_08 => X"41BE1F5F80003FF0002023FFDF79000000000EFFE309606020008005FC000000",
INIT_09 => X"FC83FE1840C0902400300000000000DFFD4004040C4D32BF7C0EE860003CE680",
INIT_0A => X"10018C24110A860006C620C0312241C482B20420CC56924E2199000C00415037",
INIT_0B => X"4669070510C90C14304043040430404304043040430404304043040218202182",
INIT_0C => X"008000105400C00400100000A018000801000C024000004A940000FFDF820604",
INIT_0D => X"100152100801C17E61841950B1C10FFF57FFC02812F00429DC92C40002000100",
INIT_0E => X"10015210088528E00E02C8200A430A424202A1CAF13F214001521001CBF03F21",
INIT_0F => X"01C1C044006D0C94FB94320880603C420B8001CBF03F214001521001CAF13F21",
INIT_10 => X"30182800A018D9CA8000648528E00D12480202C86040902AC60BACDF0E02D020",
INIT_11 => X"0445C19960A00026880C006739000009B00300010AF5052419D1964419028014",
INIT_12 => X"01844068880CE72000013600600332C140004D101808458A5602E00089202911",
INIT_13 => X"41D0B9023402085020825132C8CB5B4040301009408021144CB042F880100C06",
INIT_14 => X"8E17C0D240406519400500840A9524EE38A1F80E02120018390320F050144CB2",
INIT_15 => X"01004010040100401004010040100100040040000000000001000900FBFFE000",
INIT_16 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_17 => X"0040100401004010040100401004010040100401004010040100401004010040",
INIT_18 => X"0000000000000000000000000000000000000000000000001004010040100401",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000000000000000000000000",
INIT_1F => X"4BA5D0400010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000007FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974BA5D0002000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"00010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA550002000007FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAE974AA550400000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5500",
INIT_23 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550402010087FFFFFFFFFFFFFFFFFF",
INIT_24 => X"FAE954AA5D00000AA007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA55040200008",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010000000000",
INIT_27 => X"FFFFFFFFFFFFFAE974BA5D0400010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0000010007FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAE974AA550002010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA550002",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550400010087FFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"E954AA5D0402038007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550400028007F",
INIT_2C => X"FFFFFFFFFFFFFFFFFFAE954AA5D00020BA087FFFFFFFFFFFFFFFFFFFFFFFFFFA",
INIT_2D => X"D0402010000000000000000000000000000000000000000000000007FFFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000087FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAE974BA550002010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D000001",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFFFAE974AA550002000087FFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"54AA5504000BA087FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA550400010007FFF",
INIT_33 => X"FFFFFFFFFFFFFFFFAA954AA5D04000AA087FFFFFFFFFFFFFFFFFFFFFFFFFFAE9",
INIT_34 => X"000000007BFFFFFFFFFFFFFFFFFFFFFFFFFAA954AA5D00020AA007BFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000007FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(23),        -- Port A data input
DOA(0)   => data_read_a_lo_256(23),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(23),        -- Port B data input
DOB(0)   => data_read_b_lo_256(23),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_24_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100600007FFF000080108004000800020000840041000080808",
INIT_02 => X"0000068002CC07400000090C080002000000103FF811F150231000520ABE4404",
INIT_03 => X"210A0600000203F80005DC00000DC3801EA000000745C4010220000000008000",
INIT_04 => X"07C5FF804900026F8780001DF8000000079800000F300002998078068003C080",
INIT_05 => X"C207F0000000007FF0000004380001FE1E1C07C3E00CFFF80000000000000000",
INIT_06 => X"0002648240F20035A0102000BD0000002802C87FC800FCAA035400001B918600",
INIT_07 => X"0000000001FBFFEC4D2B4AD0B8129063B2CC0000100042018408142F16C01848",
INIT_08 => X"008E1F5F80001FF0000000FFDF78000000000EFFE001600000000005FC000000",
INIT_09 => X"E883FE180000000000300000000000DFFD0000002A80D500000671000004A000",
INIT_0A => X"10018C0411020600048620C030020502000200000400920A2198000800404037",
INIT_0B => X"0641060400C00C00304003040030400304003040030400304003040018200182",
INIT_0C => X"000000001000C00000000000000240058000000000000000000000FFDF000404",
INIT_0D => X"E00880104809C1666594584031010FFF56FFC000104000000010440000000000",
INIT_0E => X"E0088010492064206100E81084200048C0804012500021B00880108012500021",
INIT_0F => X"04100144800803419043064900C0020501840012500021B00880108012500021",
INIT_10 => X"1018140F02C0000809408D206420530270040410004C840041A0D80054109038",
INIT_11 => X"110002C9E8010C00010480B35A0300400041020902F60002260D65B361BAA104",
INIT_12 => X"0228204300166B4060080008240593D0021800020818B06D9802F00030C02060",
INIT_13 => X"143B62023C00142800B04400095DFF90203020042108603100061516EE800C06",
INIT_14 => X"DC1180C7804400044029208301040214AE4C7C02000040206602C10B48110006",
INIT_15 => X"00000000000000000000000000000000000000000000000000000000FBFFE000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"DD5EDCF9822659B6888332000000000000000000000000000000000000000000",
INIT_19 => X"F3CF3CF3CF3CF3DF7DF7DF7DF7DF7DF3DF3DF3DF3DF4D30C2432AEBAEBFE5A15",
INIT_1A => X"C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783DF7DF7DF7C",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000F0783C1E0F0783C1E0F0783",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201008000000000000000000000000",
INIT_1F => X"4BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974BA5D0400000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"00010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000007FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAE974BA5D0000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_23 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0002000087FFFFFFFFFFFFFFFFFF",
INIT_24 => X"FAE974BA550002000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D000200000",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010080000000",
INIT_27 => X"FFFFFFFFFFFFFAE974BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000087FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAE974BA5D0400010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0000010007FFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"E974BA550002000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0000010007F",
INIT_2C => X"FFFFFFFFFFFFFFFFFFAE974BA550002000007FFFFFFFFFFFFFFFFFFFFFFFFFFA",
INIT_2D => X"D0402010080000000000000000000000000000000000000000000007FFFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAE974BA5D0400000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040200",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000087FFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"74BA5D0000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0000010087FFF",
INIT_33 => X"FFFFFFFFFFFFFFFFAE974BA550000010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE9",
INIT_34 => X"000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA550002010087FFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(24),        -- Port A data input
DOA(0)   => data_read_a_lo_256(24),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(24),        -- Port B data input
DOB(0)   => data_read_b_lo_256(24),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_25_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100200002000000080100004000000020000800041000080808",
INIT_02 => X"0000068002CC474000000800000002000000103FFCE302008000000880844A04",
INIT_03 => X"00000040700803FC0105DE00020DC3801EA00000040000000020000000008000",
INIT_04 => X"47C5FFC04904026F8780081DFC040000079C92484F30499299837C168003E400",
INIT_05 => X"C207F0382004407FF0000004382281FF1E1C07C3E00CFFFC090004B05000200A",
INIT_06 => X"1009015C4000000020000000390C10002802C87FC800F8000000000019810600",
INIT_07 => X"0501000001FBFFFD480A0280A816002010800001000054018408102000000002",
INIT_08 => X"0C8E1F5FA21C9FF8004000FFDF7C062031863EFFF75D78004001010DFC000020",
INIT_09 => X"E883FE180C00000000300000000000DFFF00180800000000000660100000A000",
INIT_0A => X"1001DCCC31222730A49620C030020100000200000400921A21D8000804404037",
INIT_0B => X"0641062400C00C00304003040030400304003040030400304003040018200182",
INIT_0C => X"C11160845004D04820000000000000000000000000000000940000FFDF000404",
INIT_0D => X"000800000801C0786184185031810FFF56FFC02812E0182000F2C48304418220",
INIT_0E => X"0008000000002020000008000000000800800002400001000800000002400001",
INIT_0F => X"0000010000000000900000080000000400000002400001000800000002400001",
INIT_10 => X"1000000002002000004000002020000200000000000404000000880000001000",
INIT_11 => X"010000082000000001000001080000000040000100C600800001040000040009",
INIT_12 => X"0000000100002100000000080000104000000002000000081001000000000040",
INIT_13 => X"0010200000000000001004000001080000400080000040010000001080001008",
INIT_14 => X"8C11808200400000400000C20000000420000000030280000000010000010000",
INIT_15 => X"82208822088220882208822088A20C52082081A30080000002005008FBFFF001",
INIT_16 => X"2208822088220882208822088220882208822088220882208822088220882208",
INIT_17 => X"2088220882208822088220882208822088220882208822088220882208822088",
INIT_18 => X"29432D518B45265D82BB4101000005FFFFFFFFFFFFFFFFF82208822088220882",
INIT_19 => X"24924924924924820820820820820820924820924824000A6242B4D34D7F7451",
INIT_1A => X"AC562B158AC562B158AC562B158AC562B1188C46231188C46231189249249249",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000162B158AC562B158AC562B158",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000000000000000000000000",
INIT_1F => X"4BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"02000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAE974BA5D0402000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_23 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000007FFFFFFFFFFFFFFFFFF",
INIT_24 => X"FAE974BA5D0400000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040000008",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010000000000",
INIT_27 => X"FFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAE974BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000007FFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"E974BA5D0400000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000087F",
INIT_2C => X"FFFFFFFFFFFFFFFFFFAE974BA5D0400000007FFFFFFFFFFFFFFFFFFFFFFFFFFA",
INIT_2D => X"D0402010000000000000000000000000000000000000000000000007FFFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"74BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000007FFF",
INIT_33 => X"FFFFFFFFFFFFFFFFAE974BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE9",
INIT_34 => X"000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000007FFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000007FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(25),        -- Port A data input
DOA(0)   => data_read_a_lo_256(25),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(25),        -- Port B data input
DOB(0)   => data_read_b_lo_256(25),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_26_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"E9264EAB20190CA3BA4997AA9002AE9C001006B0778015CFA17E0811039879C7",
INIT_01 => X"F1FFF9BB1F773C7F9BB07DFFFDD863FC5FFF3FEFFBBF9FFB22FFFBC7B9F30686",
INIT_02 => X"9B3184F8AFDEAF300029E4E300FC78A6258548EFFA71C00172082400003A2161",
INIT_03 => X"0084F0FF7FFF1FDD3FEFDCDE981DC3FF5F0D294A7B2B18A0001B9CE6CC606E73",
INIT_04 => X"0FC5DFD7EDFFD66F87FE605DDDBFF3690F9EDB7F5F7AFF639BD7DE37C2FEF591",
INIT_05 => X"F205F0F8E9D199FF76DFEE1C3FCC3FF7BE1FD7C3FFACFBFFDFF7B4FEFFDAA10E",
INIT_06 => X"042648C40179912406C1830639AFBEC14489737FDC00B13BB79DFDB83BF4112A",
INIT_07 => X"763A844769FFBFE4398E4390BB9C28B1D0F049080414583F9468D1AEFC000060",
INIT_08 => X"02C05FD7BC471FBD13D981F7DF7D7E6171AF3FEFE8A3E679FAC1FD1FFFBEB000",
INIT_09 => X"F8CFFE38FF7F6BD928F1ABB47476B5FEF9F59F5FCEEDE73FEE0EFC53B079F5CC",
INIT_0A => X"315BDDCC3B336F7C548667D47B7737AF3FD62601EDC2B66A67B9D60FE4C4427F",
INIT_0B => X"06E19F4DA0E80E903DE3035E3035E3035E3035E3035E3035E3035E981AF181AE",
INIT_0C => X"EBFBF7FEBD66DBFCA3F87501AE7B080607307DCFE1D4077B4D026FFFFBFFAFCD",
INIT_0D => X"0007E010084BCD7FF1B61B5C33813FFFFCFFC7D7D51D6F5FDCB935D7AFEBD7F5",
INIT_0E => X"0007E01001BD8020500008001F010040520201F45EC0010007E01001F45EC001",
INIT_0F => X"1DC0004600400F781429C0080000770001A001F45EC0010007E01001F45EC001",
INIT_10 => X"10003C064000E408010081BD8020600200001EC00040B02007EC09A0E0001000",
INIT_11 => X"360403E434588007200D00F88C84C081C203404B3BFD0402346235408402C080",
INIT_12 => X"07B00040091F1190982038406807C868B1000E401A08FE0012040000FC002001",
INIT_13 => X"7D00212000007C400082D81009FC08281D00001F010021560406758091454000",
INIT_14 => X"FFBFF5FA1040076065F730FC08043A903A80008320C0403C3400008860160406",
INIT_15 => X"D7F5FD7F5FD7F5FD7F5FD7F5FDFF7F7F7F77F9F761FFBFDFFDE5BFFFFF7FF005",
INIT_16 => X"7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5F",
INIT_17 => X"F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD",
INIT_18 => X"B79E923C2CD990AA7F0DDB6B910C8DFFFFFFFFFFFFFFFFFD7F5FD7F5FD7F5FD7",
INIT_19 => X"30C30C30C30C30C30C30C30C30C30C30D34D34C30C35F7AA9ABF0E38E3A8EB62",
INIT_1A => X"C26130984C26130984C26130984C26130984C26130984C26130984C30C30C30C",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000130984C26130984C26130984",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000000000000000000000000",
INIT_1F => X"4BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"02010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_23 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFF",
INIT_24 => X"FAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010000000000",
INIT_27 => X"FFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"E974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007F",
INIT_2C => X"FFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFA",
INIT_2D => X"D0402010000000000000000000000000000000000000000000000007FFFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"74BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFF",
INIT_33 => X"FFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE9",
INIT_34 => X"000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(26),        -- Port A data input
DOA(0)   => data_read_a_lo_256(26),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(26),        -- Port B data input
DOB(0)   => data_read_b_lo_256(26),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_27_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"00080A40000A41248002029000050A088000008242A0004404480002000A1155",
INIT_01 => X"F1FFF1C11F781C129C107DFFFE0860941E81258CA2B71C2220EC1B86E1A00002",
INIT_02 => X"183080988B2EAE00002BE001117C78C6848140CFFA0000800042008000011081",
INIT_03 => X"000000FF7CF91F1D3DEF3CDA881D23FB5C0C21085B0B0820001318C60C204C63",
INIT_04 => X"8FC51FD7EDFDD66E47EE205D1DB7F1490E5EDB7D5CBADB2385D79C3643D4E580",
INIT_05 => X"E001F0C0C991BBFC76DFEA1A3F8C3BC7391F9723FF2CE3FCD6D13096B79C8106",
INIT_06 => X"40000001000000084041830600A40C415004637FC4003021259CFDB01BF80028",
INIT_07 => X"3158954761FA3FE402088220AC1108001080400A400041018468D1A060000050",
INIT_08 => X"02005F0784411E390A4881C7BEFC5F6171CE2F8FE823E778DAC16C1FFBBC9000",
INIT_09 => X"F0C7FEBABF3F6BD108F40E04C0C084F0F8B58B5B8849673F6C0E7A01B00914C4",
INIT_0A => X"B51BFDCC39732F3554866AD57C37BEAF1C152201A4C0B6EA63AAD60B60D4427F",
INIT_0B => X"06F18FC5A0E00F0038D1030D1030D1030D1030D1030D1030D1030F0818688186",
INIT_0C => X"AB6AD7EAB962CBD8A3A83101F47E08040510768EA0C406630D0226FFE375ADE5",
INIT_0D => X"000760000843C561E5C55C42B9011FFF48FFCC57550D63564D1D2556ADAB56D5",
INIT_0E => X"0007600004BD8020100008001F010000130201E44A40010007600005E44A4001",
INIT_0F => X"1DC0000208400D781020C00800007700002005E44A40010007600005E44A4001",
INIT_10 => X"10003C064000C400018080BD8020200200001EC00000382006EC0820A0001000",
INIT_11 => X"3E0403A424108007200102E888808081C20040431BC504021462354004004080",
INIT_12 => X"07B00000015D1110102038400817484821000E400204FE0010040000FC000000",
INIT_13 => X"7D00202000007C400000F81001FC08080500001F0100005E0404758081014000",
INIT_14 => X"8DBBB5FA10400360649310FC08003A903A8000012040403C34000080201E0404",
INIT_15 => X"56D5B56D5B56D5B56D5B56D5B56D7E3D7B57B1C4E17F0944B8D596EEFC7FF001",
INIT_16 => X"6D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B",
INIT_17 => X"D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B5",
INIT_18 => X"2D0200903950C080420948E2D10E8FFFFFFFFFFFFFFFFFF56D5B56D5B56D5B56",
INIT_19 => X"00000000000000000000000000000104000000000004000E5E420000002921C4",
INIT_1A => X"28140A05028140A05028140A05028140A0100804020100804020100000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000140A05028140A05028140A050",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000000000000000000000000",
INIT_1F => X"4BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_23 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFF",
INIT_24 => X"FAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201008",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010000000000",
INIT_27 => X"FFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"E974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087F",
INIT_2C => X"FFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFA",
INIT_2D => X"D0402010000000000000000000000000000000000000000000000007FFFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"74BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFF",
INIT_33 => X"FFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE9",
INIT_34 => X"000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000007FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(27),        -- Port A data input
DOA(0)   => data_read_a_lo_256(27),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(27),        -- Port B data input
DOB(0)   => data_read_b_lo_256(27),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_28_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"02200AA400180030808802A900002A08001280A08A801044104A1000001818C3",
INIT_01 => X"50A00011460214428114180000882214413D0A71592A01D92213D28005210202",
INIT_02 => X"8A54800A210200111100C2110054289220810440030404010844000444410001",
INIT_03 => X"1080010208B51400007800000A000001000108C21008092000018C6295200631",
INIT_04 => X"0008000000017000000028000001610300000010000802202040012040040011",
INIT_05 => X"2000044440048880026A22000026A20000000000000000004994140203000064",
INIT_06 => X"1400922401041008004891224228810080010200040001020800000004000008",
INIT_07 => X"150B001328000001404010040084088404200020455514000224489028492201",
INIT_08 => X"00414000201800004080A0000002480B04008100011000088800081002C19020",
INIT_09 => X"000400001036584108415B4A6A694A0000100101C08200000001000190200044",
INIT_0A => X"004800210C19808400500010009110091500020B408820000200400040811600",
INIT_0B => X"40000800B00100040D8140581405814058140581405814058140580A02C0A02C",
INIT_0C => X"00200248010201008298150006210802043058C46054032981002D00201C8081",
INIT_0D => X"0000A00000400600841041108280300008000140000401028008330000800040",
INIT_0E => X"0000A000000080001000000000000000500000040A40000000A00000040A4000",
INIT_0F => X"00000006000000080020C00000000000012000040A40000000A00000040A4000",
INIT_10 => X"00000000000024000000000080002000000000000000A00000040020A0000000",
INIT_11 => X"2200000404108000000900008080808000024040152000000020000004004080",
INIT_12 => X"0000000009001010102000004800080821000000120002000004000000000001",
INIT_13 => X"2000002000000000000288000020000805000000000001420000200001014000",
INIT_14 => X"408010000000022000D610280000080000000001204000000000000820020000",
INIT_15 => X"00401004010040100401004010042024210218734CD52150A840827504000000",
INIT_16 => X"0401004010040100401004010040100401004010040100401004010040100401",
INIT_17 => X"4010040100401004010040100401004010040100401004010040100401004010",
INIT_18 => X"05822140048D2E57B1348141845C200000000000000000000401004010040100",
INIT_19 => X"04104104104104104104104104104104104104104101A6A0A0EB1861863BC422",
INIT_1A => X"2C160B0582C160B0582C160B0582C160B0180C06030180C06030181041041041",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000160B0582C160B0582C160B058",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000000000000000000000000",
INIT_1F => X"4BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_23 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFF",
INIT_24 => X"FAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010000000000",
INIT_27 => X"FFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"E974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007F",
INIT_2C => X"FFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFA",
INIT_2D => X"D0402010000000000000000000000000000000000000000000000007FFFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"74BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFF",
INIT_33 => X"FFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE9",
INIT_34 => X"000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000007FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(28),        -- Port A data input
DOA(0)   => data_read_a_lo_256(28),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(28),        -- Port B data input
DOB(0)   => data_read_b_lo_256(28),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_29_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"79964E4BA01DACAB9E659792D00AAE160002829C7FDFEFCEE97C2815039D70C3",
INIT_01 => X"50BFF9AB0775343F9AB01DF80D5821FC0FFF3FEFD1AF9FF1207FFBC7B9720586",
INIT_02 => X"0D15846807D207200021C4E200D428A2018408600271C000720A0000003A2161",
INIT_03 => X"0000B0027BBF17C43E6DC05E1A0DC07D1F0000803B2819A00019084345606421",
INIT_04 => X"07CDC047A4FB526F807C681DC4B97369078249370F482E62BA414627C2FE3000",
INIT_05 => X"F204007861C088FF0EFF260407C427F19E03C7C01F8CF80749B390EA4BCA202C",
INIT_06 => X"000248C00079800406C081023B233E804488527FDC008019968D74982C94110A",
INIT_07 => X"5229000221FF8000398641903B082831D05000200000083F942850AEB4000221",
INIT_08 => X"00805FD0180E1F8C1111A0F041056A0100A11FE000916249A800B915FE82B020",
INIT_09 => X"F80C000055FF7C492840AAB45456B55E015015058665A31DA603A4539058F54C",
INIT_0A => X"000850400A11414C005005000B51158936D20601A98A204006114005C4800217",
INIT_0B => X"40201948B029029409A3401A3401A3401A3401A3401A3401A3401A9A00D1A00C",
INIT_0C => X"40B1225C1506512C83E85500AC3A080406305587A154023141006DFFF89E82C9",
INIT_0D => X"0000A01008480D3EB4A24A0C910037FFFC0007C7C0140D0B50A8218102C08160",
INIT_0E => X"0000A010010080005000000000000040520000141EC0000000A01000141EC000",
INIT_0F => X"00000046000002080429C0000000000001A000141EC0000000A01000141EC000",
INIT_10 => X"00000000000024080100010080006000000000000040B000010401A0E0000000",
INIT_11 => X"3600004414588000000D00108484C080000340483B590000202000008402C080",
INIT_12 => X"00000040090210909820000068008828B10000001A0802000204000000002001",
INIT_13 => X"20000120000000000082D800082000281D000000000021560002200011454000",
INIT_14 => X"B29450580000066021F6303C000408000000008320C000000000000860160002",
INIT_15 => X"816058160581605816058160589625662522506344FF9FCFFF62EB6DFF001004",
INIT_16 => X"1605816058160581605816058160581605816058160581605816058160581605",
INIT_17 => X"6058160581605816058160581605816058160581605816058160581605816058",
INIT_18 => X"F2DDCFFFBEFFCF07FFBFFD41800C05FFFFFFFFFFFFFFFFF81605816058160581",
INIT_19 => X"7DF7DF7DF7DF7DF7DF7DF7DF7DF7DD75D75D75D75D77FFBF3F7DFFFFFFD779F3",
INIT_1A => X"FEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDF7DF7DF7DF",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00001F7FBFDFEFF7FBFDFEFF7FBFD",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000000000000000000000000",
INIT_1F => X"4BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_23 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFF",
INIT_24 => X"FAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010000000000",
INIT_27 => X"FFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"E974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007F",
INIT_2C => X"FFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFA",
INIT_2D => X"D0402010000000000000000000000000000000000000000000000007FFFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"74BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFF",
INIT_33 => X"FFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE9",
INIT_34 => X"000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(29),        -- Port A data input
DOA(0)   => data_read_a_lo_256(29),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(29),        -- Port B data input
DOB(0)   => data_read_b_lo_256(29),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_30_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"FFDFF3FC3EFFF7FFFFBFFA000000000000000000000000000000000000000000",
INIT_19 => X"F3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF5F7AEBEBFBEFBEFFEFFF7",
INIT_1A => X"CFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCF3CF3CF3C",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000007F3F9FCFE7F3F9FCFE7F3F9F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000000000000000000000000",
INIT_1F => X"4BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_23 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFF",
INIT_24 => X"FAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010000000000",
INIT_27 => X"FFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"E974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007F",
INIT_2C => X"FFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFA",
INIT_2D => X"D0402010000000000000000000000000000000000000000000000007FFFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"74BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFF",
INIT_33 => X"FFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE9",
INIT_34 => X"000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(30),        -- Port A data input
DOA(0)   => data_read_a_lo_256(30),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(30),        -- Port B data input
DOB(0)   => data_read_b_lo_256(30),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_31_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"129000008004A00804A40000400800020000000C005FEA005800200400050100",
INIT_01 => X"A15FF18019700810180065FFFC0040801E80258CA2951C2200EC0906A0804140",
INIT_02 => X"146000808A0C060444692000402850040400408FF80000000010000000004000",
INIT_03 => X"000000FD74480B1C3D951C5A800D03FA1C0C21084B0300000012108518004842",
INIT_04 => X"07C51FC7EDFCA26E07EE001D1CB6904A061EDB6D4C30490281831C1602D0E480",
INIT_05 => X"C001F0808181117C7C95C8183FA099C7181F8703FF0CE3FC0201209010988002",
INIT_06 => X"00000000000000010001020400840C41C000617FC0003021259CFDB01BF00020",
INIT_07 => X"0000000441FA3FE400080200A810000010804008100040018448912040000040",
INIT_08 => X"00011F0780011E38004801C79E7C162231862E8FE00166704041240DF93D0000",
INIT_09 => X"F0C3FE180D89279000B00000000000D0F80088080849673F6C0E780020091480",
INIT_0A => X"1011DCCC31222730048620C4382204A608142002A440924A6188020920404437",
INIT_0B => X"0661874500E00E00304003040030400304003040030400304003060018200182",
INIT_0C => X"810040801060C04821202001A05A00040100240A80800442040202FFC3200444",
INIT_0D => X"000740000803C0616184184031010FFF40FFC407500020004C10060204010200",
INIT_0E => X"0007400000BD0020000008001F010000020201E04000010007400001E0400001",
INIT_0F => X"1DC0000000400D701000000800007700000001E04000010007400001E0400001",
INIT_10 => X"10003C064000C000010080BD0020000200001EC00000102006E8080000001000",
INIT_11 => X"140403A020000007200000E808000001C200000308C504021442354000000000",
INIT_12 => X"07B00000001D0100000038400007404000000E400000FC0010000000FC000000",
INIT_13 => X"5D00200000007C400000501001DC08000000001F010000140404558080000000",
INIT_14 => X"8C1380DA10400140640100D4080032903A8000000000403C3400008000140404",
INIT_15 => X"02008020080200802008020080200C1808008184012A08041202500AF87FF001",
INIT_16 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_17 => X"0080200802008020080200802008020080200802008020080200802008020080",
INIT_18 => X"000000000000000000000002001005FFFFFFFFFFFFFFFFF02008020080200802",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000000000000000000000000",
INIT_1F => X"4BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_23 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFF",
INIT_24 => X"FAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010000000000",
INIT_27 => X"FFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"E974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007F",
INIT_2C => X"FFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFA",
INIT_2D => X"D0402010000000000000000000000000000000000000000000000007FFFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"74BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFF",
INIT_33 => X"FFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE9",
INIT_34 => X"000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(31),        -- Port A data input
DOA(0)   => data_read_a_lo_256(31),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(31),        -- Port B data input
DOB(0)   => data_read_b_lo_256(31),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_0_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"ED39BA795990D275FB4A6E96ACC4731DEA4598B0AFB54867F6EE4618C3749807",
INIT_01 => X"58A0047D8607944AC7DA180001ECA2444042106208408208C20022E9173734B3",
INIT_02 => X"8B1E49562021F8051500147A0E162923024F28000415F5787B09FBF999BB1EFC",
INIT_03 => X"1013BF028A959403C06A23A147723C01E140088280C4CF6996088862C7922221",
INIT_04 => X"781A003802015D9078011DE20340699198600000B08694916434804825241311",
INIT_05 => X"2CA000587E10C880036A3103C00F2000E1E0383C00730002B4409845E4425171",
INIT_06 => X"179B48CFF95DCF9EF730E1C3BB731138AF7B888025340C0888430047040FEE18",
INIT_07 => X"AF155113160400185F87C1F05707D415E664A6E7C5551EBE783060CEB164833F",
INIT_08 => X"4D7E40002B7AE005FDB47600208229010C6101001EFE198C96B0528202C0DCB4",
INIT_09 => X"062400608234D864444081048A80CC00062D42D30222108091C107A1DA040267",
INIT_0A => X"204A21008E514844EB5145000255DA599581D3A9583C24351240B58298011308",
INIT_0B => X"E08C4830F81380CE0F89E07A9E0789E07A9E0789E07A9E0789E070CF0184F038",
INIT_0C => X"3A4E9D63EA180EB150CA1CA45C254D4AF4AA414568729139F2A12C0000016110",
INIT_0D => X"F0009E0FC048211E9C11C31F82E4A000890022B827EB52F52347F174E93A749D",
INIT_0E => X"F0009E0FCC42EFDFBF0AE03080E2AEB2E0F1F80FA97FE0F0009E0FC40FA97FE0",
INIT_0F => X"0231F0BD9E3FC08FEBD6F661C0E008C3CB5F040FAB3FE0F0009E0FC40FAB3FE0",
INIT_10 => X"20180309A0F83BE2B87C7C42EFDFBF187806013879BA878FE807F65FBF12E038",
INIT_11 => X"0BE9F01FC8B38C2098DAE007F323A0C83136B248831ACBFC8BBDCAB779BC699F",
INIT_12 => X"004C72BEC800FE7464290626D7003F9947184131B59003FFEC07F00003F01FB9",
INIT_13 => X"A0FFDA2A3C0202B8776A2FA7F023F7D065703080E29F1B2BE9F8A27E6E915C0E",
INIT_14 => X"016C2D25E52630BB1AE49C2BA7F98D6F846DFC0C2352A0024B83F07F198BE9F8",
INIT_15 => X"749D2749D2749D2749D2749D2749F285F25D2C500815A5522CB5A4B400000CD4",
INIT_16 => X"49D2749D2749D2749D2749D2749D2749D2749D2749D2749D2749D2749D2749D2",
INIT_17 => X"9D2749D2749D2749D2749D2749D2749D2749D2749D2749D2749D2749D2749D27",
INIT_18 => X"31C136AD8E9B562BA39E2600654BA800000000000000000749D2749D2749D274",
INIT_19 => X"4104104104104104104104104104104104104104104104109C83B8E38E2ABE71",
INIT_1A => X"0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0410410410",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000007C3E1F0F87C3E1F0F87C3E1F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000187FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"BAF7FFD55EF007FD75EFFFAE97555557BD75EF5D000000000000000000000000",
INIT_1F => X"000AA843FE00AAFBE8B45AA803DFEFA28428B455D0017410A28428AAAA2FBD54",
INIT_20 => X"FEBAA2D5401450051401555D7FC0145F7AEBFFFF08002AA10A2AABFEAAA2FFC0",
INIT_21 => X"D755555517FFEFA280021FF082E974AA5D7BFFE000804000BAAAAAAAB45557FF",
INIT_22 => X"EA8B45005168A10AA8028A10087FD7410557FC21555D51574AAA2FFE8B455D7B",
INIT_23 => X"AE95410AA80000005D003FEAAFFAEBFE00A2803FEBA002A820AA0800174BA5D2",
INIT_24 => X"2AEA8A10000417410A2FFE8BEFF7FFE8B45FFFBC00005D003FF45557FC01FFFF",
INIT_25 => X"00000000000000000000000000000000000000557DF5500003DFEFFF84175EFA",
INIT_26 => X"5F524AFE38B780154BAFFF1D54AF0075D75EFEBAE9554540754717F1F8000000",
INIT_27 => X"50B6AABDE12BEA0AF010B7D1F8F47E00A2DB45AA8A3AFD7B68E2AB78550E1255",
INIT_28 => X"E9257F1E816D557095EAAA2D1401D500002A150038038E285D7F78FD7000B6AB",
INIT_29 => X"5A87AAD178A8002D1D21C5E8257D5C7AA854008700249243A412EBFF5542A43F",
INIT_2A => X"52A82000E3A5D2150AB8F401471EDBC0B680900AAF52B474385D75C502D15754",
INIT_2B => X"FD7E9541242FE920AD082E10A28F6A150012A2F02AFFDF40E85F475451D502D1",
INIT_2C => X"0550E87B7A405B52AAD152BD00151EAFEDB52E3F1EFFFF485A2DA3D5D24BD417",
INIT_2D => X"57F40545850000000000000000000000000000000000000000000005AAF55508",
INIT_2E => X"F7AEAABFF5D2A81151FB8635A02FA69574BAF7D5555AF0D79D55FFA2AC974450",
INIT_2F => X"8D46F6ABE7082AAAAF2FAC77FE00FF16565B2FA9075F4F7B3EBDF50FEAEAAB55",
INIT_30 => X"56803CE3AEB038662E5D81406014D5D51F5E08A394003A908B8410E707EF34A0",
INIT_31 => X"4AF0151555AF58794040077D774FAE8C798A11A0EAEF75F7AA84001A7052C952",
INIT_32 => X"4E1870108B11020AD4AA05542A0A05051023F9A9D57B63BFBF906CB45FABC095",
INIT_33 => X"F5F0DA6BC9525688C1A2A0C06E9FEE5555BE48AB2A2AE0A0F20C43EAC562245B",
INIT_34 => X"000000FF80F55E25C00A0BA7FBED407A97F6F35F498B96BEB12DAAB77558ABD5",
INIT_35 => X"8000000FF8000000FF8000000FF8000000FF8000000FF8000000FF8000000FF8",
INIT_36 => X"00000000000000000000000000FF8000000FF8000000FF8000000FF8000000FF",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000008000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(0),        -- Port A data input
DOA(0)   => data_read_a_hi_256(0),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(0),        -- Port B data input
DOB(0)   => data_read_b_hi_256(0),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_1_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"212C001411984004084D000508C53810A03D1450E839B003342114428A000803",
INIT_01 => X"08000010400A0008010600000084005000400002000000000000000000140000",
INIT_02 => X"C084484000002014400205851002007030450E0000A606C8C44CB4C6666C00E0",
INIT_03 => X"CCF7CE0002058001000000800240200001018CA1800001091408463061120118",
INIT_04 => X"082800100000000040000900010000100040000000008411600401C02100000C",
INIT_05 => X"10800202080422000020012200000000810000200000000004020C00200011A0",
INIT_06 => X"56BDBFBC48C315A8660C18305750C008940D8000011000820001000104050004",
INIT_07 => X"8B4344400004000150248912154404C6060A2FE24555013E13060C158AC97F01",
INIT_08 => X"00082080087A000559102400200281000469000008B000000090108000400430",
INIT_09 => X"0000000000001004140545402820020000010010208000008041060008200001",
INIT_0A => X"2102210182004840007845004044020000200080080844200000048088000000",
INIT_0B => X"48800000190191064620646A06468064680646A0646A06468064690321503234",
INIT_0C => X"02008100200800A1100707040101E20BE0B002605C1C110848200C0000000800",
INIT_0D => X"F000A000C0000012187087010AE4B00000000810010040108104100408020401",
INIT_0E => X"F000A000CC4200002F08E03080000010F18058000003C0F000A000C4000003C0",
INIT_0F => X"000000078808C00000023461C0E00000012704000003C0F000A000C4000003C0",
INIT_10 => X"201803000000240218C0044200001E1878060000000AAC00680000001F10E038",
INIT_11 => X"2100B00048230C200009A0001303204800025200040A00D000000202090C281F",
INIT_12 => X"00000002C9000260640900004D0000904618400012900001EC03F00000000039",
INIT_13 => X"80025A0A3C020000002A8400B00007806070308000000961002880204A901C0E",
INIT_14 => X"000801046004308A185000020128000904285C0C0312A0020000000838810028",
INIT_15 => X"0401004010040100401004010040100010410C002000040280100000000008D0",
INIT_16 => X"4010040100401004010040100401004010040100401004010040100401004010",
INIT_17 => X"0100401004010040100401004010040100401004010040100401004010040100",
INIT_18 => X"48D757DF8A9410218E8A56085142020000000000000000004010040100401004",
INIT_19 => X"555555555555555555555555555554514514514514550431A581924924B02651",
INIT_1A => X"4BA5D2E974BA5D2E974BA5D2E974BA5D2EB75BADD6EB75BADD6EB75555555555",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800005D2E974BA5D2E974BA5D2E97",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000607FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"10AAAABFFFFFF803FE10F7D17FEBA55556AAAAAA800000000000000000000000",
INIT_1F => X"EBAFFD555400557BD54BA5D7FFDF45A2FBD75EFA2AE97555F7FBFFF45FFAE800",
INIT_20 => X"ABEFA2D568A005D5157400AA8028AAAF7FBD54AA002A955555D7FE8ABA082EBF",
INIT_21 => X"FDF55AAFBC0010555540010550417555AA8028BEFAAAE97555082A80000AA802",
INIT_22 => X"BD7410550428ABA5D5168ABA552EBDFEF5D7FEAA00AAAABFEAA007BC0145FFFF",
INIT_23 => X"FFEAB55557FFFEBAAAD568B45A2D5575555D7FC2155F7AEA8BEFAAAA954BA557",
INIT_24 => X"D7BD74000804154BA082ABFF55FFD57DF45F7D568ABAF7AABFFFF082ABFFFFFF",
INIT_25 => X"000000000000000000000000000000000000002EBFFEFA280021FF082E974AA5",
INIT_26 => X"5E175EFF57BF8FC2000BEA4BAE97F78A3FE28E3D17DEAA485FE8E02B50000000",
INIT_27 => X"455571E8A2A087BF8EAAEB8E0016D5D75D54BA5D7BFFF7DA2FFD55EFAAA49554",
INIT_28 => X"157428145A00AA8A2FBD7B6DF6AA28550E10405F7A4AFE38EAA0924921C2FD55",
INIT_29 => X"8E971471C7010B7D168F47400A07A28415A001684104155C5B6DF6DBEFBFAA07",
INIT_2A => X"BFBD7B6A0BF492415FC20105D24AAABF1FFBC7010FF8A38FEF557FEAB78B6AAB",
INIT_2B => X"017EBA4A8EB8F6FFD5FE8B7D557495EAAA2D16D1FDBED56A55557A43DE385FD4",
INIT_2C => X"854008700249243A417FFF41542F5D717FE2AAAA56DEBD17FE3DF7FB7FEBFE38",
INIT_2D => X"07DFCA127B8000000000000000000000000000000000000000000002A3D5C7AA",
INIT_2E => X"AAFBD55FFAA8416545A6FB60F47AF2A00010F78028B15F7823FEAAA2D57DFBA0",
INIT_2F => X"22A38C20B2552E975F758516AAAA0869AAAB8A7C19C55550E8574BA557BFFFEF",
INIT_30 => X"55FFEFBCEE5FBAACB10085EE5DE10A2AEBFF55F7BAAA8565DBAC1112FFAC21A0",
INIT_31 => X"BEA097BEAAFAF2863FA00DD574201E7AD1FFF5575841DE08007FC20480028957",
INIT_32 => X"54FF57EFBFA18D4FBFFF40FF809D4000D7FC00FC5D062BBA05ED5034472A02EA",
INIT_33 => X"7DFBFF6963FCAAA2283CF14050062B0A2F7AE8B5D5D51F5E18ABD5EAFFF2AF95",
INIT_34 => X"000000002CB75F7AA84001A7052C95256807DC31AA8114DE55F5BED201FFFED1",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000008000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(1),        -- Port A data input
DOA(0)   => data_read_a_hi_256(1),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(1),        -- Port B data input
DOB(0)   => data_read_b_hi_256(1),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_2_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10E44660018259B2843913100062C98004802322D3E030235201006009B2813",
INIT_01 => X"000AC188084900481C8024A542400340404000720885800802000906E4910204",
INIT_02 => X"82040072AC248C31010204880000007401044C0550200000480E0080001300E0",
INIT_03 => X"0080812C130D0A0D1193088802182142494D218220021100001A8020C1004A00",
INIT_04 => X"090D0AD62824A44A428408540D1610020C6E510818923441A4908B0503404201",
INIT_05 => X"5000A004081122242420480A14A99C428908122144244150906124248C002168",
INIT_06 => X"1400088400450000460000001308890094082015800011012D41D518044C1100",
INIT_07 => X"26731111491C1541324C1114BD880004002040204050413F1400100480000201",
INIT_08 => X"02410582881E0C1511D02082AAAB016A2463288549B044605201D10AE11B0020",
INIT_09 => X"E80394280E40158020B591000800481051241A4A404B5035C60904502054E000",
INIT_0A => X"0102C9E12202EA6014D027C418428E220A5500024808922801A0900A84454458",
INIT_0B => X"4600070110C10D04340043400434A043420434A04342043480434102184021A0",
INIT_0C => X"E9CA34328E44CA1401306100A246000402100C088104010AC8005C5681812B04",
INIT_0D => X"0000A0000801487334E34C1A980001550055481204090A4C01351253A728D194",
INIT_0E => X"0000A000013800004000080000000000500000B01480010000A0000150148001",
INIT_0F => X"0000000608000A500409000800000000012001501480010000A00000B0148001",
INIT_10 => X"1000000000002400000001A100004002000000000000A0000360018040001000",
INIT_11 => X"380001C01048000000090298040440000002400008C400022042004080028000",
INIT_12 => X"0000000009530080880000004813802090000000120C94000200000000000001",
INIT_13 => X"4C000100000000000002E0000950002018000000000001580002508010440000",
INIT_14 => X"7120642000000400015020500004221018000082008000000000000820180002",
INIT_15 => X"5094A5294A5294A52942509425094209461468000822241A03835D88482AB001",
INIT_16 => X"09465094A5294A5294A5294250942509425094A5294A5294A529425094250942",
INIT_17 => X"94650946509465294E5294E5294E5094650946509465294E5294E5294E509465",
INIT_18 => X"080271AE180616A38A18FA204452A7F03F03F07E07E07E05294E5294E5294E50",
INIT_19 => X"20820820820820820820820820820820820820820820490C04102CB2CB2EB2C0",
INIT_1A => X"8944A25128944A25128944A25128944A25128944A25128944A25128208208208",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF1F804A25128944A25128944A2512",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000787FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"AAAA843DFFFAAD1554005D7FD74AA00040015500000000000000000000000000",
INIT_1F => X"F45AAAAA8A10A2AE80010A2AA975FF5D003FE10F7D17FEBAF7D5420AA0855420",
INIT_20 => X"FF45A2AA975EFA2FFD7555FFFBFFF45AAFBC20AAF7D1575EF55517DF555D2EBF",
INIT_21 => X"95555552E974105D517DF55AAAAAABEFAAD1575EFAAAE974AA5D51554BA5D7FF",
INIT_22 => X"E82010F7AABFE10FFD542145FFD5554AA555555555557FE8ABA082EBFFFFAAAE",
INIT_23 => X"FBC0010AA802ABEFAAD540000FFD540000AA802AABAF7FFC2010AAAE821EF552",
INIT_24 => X"A8028BEFAAAE821550851420AA002E800AA08042AB45007FC00BAFFD168BEFF7",
INIT_25 => X"000000000000000000000000000000000000002E80010555540010550417555A",
INIT_26 => X"AE95F40002157F470AABE803AE97A2DF55400557FD54AA1D04001C5150000000",
INIT_27 => X"EF55517DFC5552ABDF45B6AEAFFD5F7A482000BEAE905C755003FE28E3D17DEA",
INIT_28 => X"0BA5FD0154BA5D7BFAF7DA2AE955EFAAA495545E3F5EFF57F7FE80082FFDE105",
INIT_29 => X"8AAF082AB8EAAEB8E0016D5D2A924105D5B7FF7DB6AAAABC7BEDB505EFBEA407",
INIT_2A => X"95038AAAEAF1D7410E80000FF8438E00B6DF68FEF4871D24BA495B5556D5571E",
INIT_2B => X"1ED1EFEAF1EFFFDEAD1C5010AA8E2FBD7B6DF47A00EBDB50000A380AAE28E804",
INIT_2C => X"5A001684104155C5B68E2DBEFBFFBC703AE2DF42AAA002A851C214003FF68007",
INIT_2D => X"50002155510000000000000000000000000000000000000000000002087A2841",
INIT_2E => X"55003FEAAAAD57DEBAA2FDDC01051FBD74BAF7802AB05AAFBD5400557BD54AA5",
INIT_2F => X"7AF7FC20B2F7FBC015D58517FF555D2ABDF55F782BEB47AFAD00010F7AA82155",
INIT_30 => X"55FFFFC20FFF3AE544108410174BA557BEABEFAAEBD55FFAA1456547A2D360F4",
INIT_31 => X"0BA547FD75FF58516AAAA0828AAAB4A78016545540400010557BFDFFFF7822A9",
INIT_32 => X"550AAFACAAA122AA8954BAA2AE9D545002A800A8FF862BA00F2F9E8F0050D442",
INIT_33 => X"954505C417FFFF08555555BAAD335B57AB5155400A2AEBFF45FFFB404007FFBD",
INIT_34 => X"00000000061DE08007FC2048002895755FFAEBCFE57BBA57002DF3C4AAAA002E",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000010000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(2),        -- Port A data input
DOA(0)   => data_read_a_hi_256(2),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(2),        -- Port B data input
DOB(0)   => data_read_b_hi_256(2),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_3_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"210C44A20020248B08431120001604B8156023104C40771B3430400A02380206",
INIT_01 => X"015A2A4050B009683C0422C992000B61404040028804A0080A000C16A8990A0C",
INIT_02 => X"C0A406500CE0A95011000D1501005274B5041AB330860281CC08008222170060",
INIT_03 => X"AB488054270F08E1289084C8020420E005A48DA16C021100003A46B06900C91A",
INIT_04 => X"848966150DA0A02941A4080C612A104201C689044382FD403C17E491829B259B",
INIT_05 => X"D006620608843116942508120A208D18A5050160C600D4C894600094B49CA068",
INIT_06 => X"12002D9401C70008060408141788E2C094887033080071913209CC8004640100",
INIT_07 => X"221111454874CCC4122C0932155400C2023940284000003E15020525CE805E11",
INIT_08 => X"020103C9984A0AC511102029869D974214EDBA132891000052C1750B48290020",
INIT_09 => X"60808C8A2E41351020004148A289428730A51E5E644C8233A0090E1020208100",
INIT_0A => X"A4000041A600417914506F955D6422000934000A090A94A020229603A414144D",
INIT_0B => X"469100841001000406D04065040650406D0406D04065040670406C8201782032",
INIT_0C => X"6A4AF532A8040AF821042D01F14084030070262810340402C0000CCE4CC12520",
INIT_0D => X"000800000401C333494594532980733302CCC81300094E5C91200257AD2AD795",
INIT_0E => X"00080000051C0000400000000000000800000190148000000800000450148000",
INIT_0F => X"0000010000000B100409000000000004000005101480000008000004F0148000",
INIT_10 => X"0000000002000000000001B00000400000000000000400000168018040000000",
INIT_11 => X"1000034010480000010002D804044000004000812E4400002440014080028000",
INIT_12 => X"0000000100570080880000080015C02090000002000CCC000200000000000040",
INIT_13 => X"1C0001000000000000104000094C002018000000000040100006418010440000",
INIT_14 => X"4128652000004404010E20500004208018800082008000000000010000100006",
INIT_15 => X"5795A5595A5595A5595A5595A5595E1152556D008028341B13924D80C2E67009",
INIT_16 => X"69565795A5595A5595A5595A5595A5595A559525795257952579525795257952",
INIT_17 => X"95256956579525495E5595A5495E5595A5495E5595A569565795256956579525",
INIT_18 => X"7818F18E0C8514298B0C52A0115009AA9556AAD552AAD5556956579525695657",
INIT_19 => X"24924924924924924924924924924820820820820825042C0000249249202A60",
INIT_1A => X"8D46A351A8D46A351A8D46A351A8D46A353A9D4EA753A9D4EA753A9249249249",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF248086A351A8D46A351A8D46A351A",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"EFAAFFD54AAF7D168B45AAAABDF5500002AA1000000000000000000000000000",
INIT_1F => X"F45FFD168AAA0855420AAAA843DFFFAAD1554005D7FD74AAA284001550055421",
INIT_20 => X"55FF5D003FE10F7803FEBAFFD5420AA080400155AAD5554AAF7802AB4500043D",
INIT_21 => X"28B45A2AE82155A2FBFFEBA0800021550855555FFAA84001FFAAAE80010A2AA9",
INIT_22 => X"168ABAFFFBD54BAAAAE97400A2FBC20AAA284175EF55517DF555D2EBFE00AA80",
INIT_23 => X"AA954AA5D7FFFF45AAAA975EF007BD7555FFFBFDF55AAFBD55EF5D2EBFE10085",
INIT_24 => X"AD1575EFAAAE974AA5D00175555D0015410F7AAAAAAA55043DE00FFFFD5555AA",
INIT_25 => X"0000000000000000000000000000000000000004174105D517DF55AAAAAABEFA",
INIT_26 => X"ABC04001C51551471D7AAF1D05D2EBD56DB7DBEAEBFF551C042AA101D0000000",
INIT_27 => X"92EB842FB5508043FF55EBD56ABD75D5B470AABE8A3AFD7A2DF55400557FD54A",
INIT_28 => X"557FD2082000BEAE905C755003FE28E3D17DEAAEBDF40002550F47155AADB504",
INIT_29 => X"DF40552ABDF45B6AEAFFD5F7A48017DAAFFFAE821C0A0717D1C5B575FFB68E82",
INIT_2A => X"C55D7492E90E3808756DA92EBFFD74BAE3AE85480FFFFC00AABE8E105C755517",
INIT_2B => X"43AE10EAF5C5547FF80954AA5D7FFAF7DA2AE905EF0075D5545E3F5EFF57F7D5",
INIT_2C => X"5B7FF7DB6AAAABC7BEDB505EFBEF5C7092FF801756D490A10438EBA4B8E92410",
INIT_2D => X"D0028A00510000000000000000000000000000000000000000000000E124105D",
INIT_2E => X"AAFBD54005D7BD54AAF78002155515157555AAD142040A2D57FFFFFFAEBFF555",
INIT_2F => X"051AE955F7AAFBC0000AF843FF5500003FF55AAFD6AB455157D74BAF7AAA8B45",
INIT_30 => X"FF557BD74EFFBACD41577B8400010F7AA8215555003FEAAAAC53DEB8A2FDDC01",
INIT_31 => X"0BAF7AA8015558517FF555D2ABDF51F782BCB47ABAE801FFAAFBEAA105D2E955",
INIT_32 => X"214FA2D3EAF57AFFDD7555082AA0AAA00557FEA8A2FDD64BAAF8282012AFFEC2",
INIT_33 => X"820AAAB842AA00000028AB0AAFF48547AE04174BA557BEABEFA2AA951FF88554",
INIT_34 => X"000000002A80010557BFDFFFF7822A955FFFFC21FFF3BE40412DE02955FF082A",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000008000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(3),        -- Port A data input
DOA(0)   => data_read_a_hi_256(3),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(3),        -- Port B data input
DOB(0)   => data_read_b_hi_256(3),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_4_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"A108400020612C80284210081034849800A000303100048B3432C82904204006",
INIT_01 => X"210668000008004C1C20250E12100368403008418984014902030906A8910200",
INIT_02 => X"120404C0024C0600000206100008402404040C00F104008040080080001310E0",
INIT_03 => X"7728805052470B5C1B873C04121D03845D0020CA0822018000080084C1000002",
INIT_04 => X"0B899E43891686690790485D5C3E02000E9892201D306D03A9835C16029AC186",
INIT_05 => X"C001E080005030767434C0003C8A01D6B81C5703C82CDBC000072400089C8120",
INIT_06 => X"1000088100410000460002041300004084080070D00030032009700024641102",
INIT_07 => X"4261950408CCBC2012048310951000000003402A4000143E1008912480000211",
INIT_08 => X"00811007AC0A1EB5131120C79E7D176251E53E80E8B361604041340838452020",
INIT_09 => X"C08360820C0912800035F1801630A8260900180C00C8021C800FEE522020A108",
INIT_0A => X"8400F88C166262E940D00D410D62AD02091704024D0A02882192020DA0544043",
INIT_0B => X"4011078510C90D143142430C243042430C24304243042430C24305121A612186",
INIT_0C => X"C08060101000C00401008800F004140009400E4002A0010240000DC3C080002C",
INIT_0D => X"000800100001C07261C51C42390240F050C3C000950008088130040100018000",
INIT_0E => X"00080010003510004000000000000048010002E0100000000800100220100000",
INIT_0F => X"0000014008001550000800000000000400800280100000000800100360100000",
INIT_10 => X"00000000020000080080009410004000000000000044080000D8008000000000",
INIT_11 => X"000005800008000001040168000040000041000100EC00004002214000008000",
INIT_12 => X"00000041003C000008000008200D00001000000208050C000200000000002040",
INIT_13 => X"17000100000000000090000002C8000008000000000060000004480000400000",
INIT_14 => X"8400C00208004844C00800000000528008000000008000000000010040000000",
INIT_15 => X"0100800004030080000C010000A00D1804404912802A261B53104810DB1E0028",
INIT_16 => X"000C030000200C01000020040300800004030000000C03000000040100802004",
INIT_17 => X"008020040100C010000200800004010040300800000020040100C03000020000",
INIT_18 => X"40C700FC0A000280C68A08A950520E964C3269B2C9864D30000C030040100800",
INIT_19 => X"555555555555555555555555555554514514514514526991A199A28A28981451",
INIT_1A => X"41A0D068341A0D068341A0D068341A0D06A351A8D46A351A8D46A35555555555",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF771F60D068341A0D068341A0D0683",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FF087FFDF5508003FEBA087FD54BAAA841540055000000000000000000000000",
INIT_1F => X"F5500003DF455555421EFAAFFD54AAF7D168B45AAAABDF55A2802AA1000002AB",
INIT_20 => X"DFFFAAD1554005D7FD74AAAA840015500002AABA082E954005500021FF5D2EBF",
INIT_21 => X"68BEF080028BFF0855555455500174BAA2AABDE0055517FF555555420AAAA843",
INIT_22 => X"168ABA0055574BA5555554BA5D0400155AAD1554AAF7802AB4500043DF45FFD1",
INIT_23 => X"0400010A2AA955FF55003FE10F7803FEBAFFD5420BA085168A00007BFDE10085",
INIT_24 => X"855555FFAA84001FFAAFBEAB45002A97545F7D1555EF55043DF5555517DEAA5D",
INIT_25 => X"000000000000000000000000000000000000002A82155A2FBFFEBA0800021550",
INIT_26 => X"5BC042AA101D0A28BC7007FFDF45080A3AEAA007BD2482BE84124285C0000000",
INIT_27 => X"004100021FF492AB8F7D1C0438E381451471D7AAFBD0492EBD56DB7DBEAEBFF5",
INIT_28 => X"FED1C5F470AABE8A3AFD7A2DF55400557FD54AABE84001C5550A28ABA1424974",
INIT_29 => X"FB5508043FF55EBD56ABD75D0428BEF005557545490012482B6A0BAE2849557A",
INIT_2A => X"6DA101475FDE10145F68A921C55504924955524AA140E0717DAADB50492EB842",
INIT_2B => X"43AF6D405F78E3A1C2002000BEAA905C755003FE28E3803DEAAEBDF40002557F",
INIT_2C => X"FFFAE821C0A0717D1C5B575FFB6DF425575D7BEFB55002097555FFD5401EF5D0",
INIT_2D => X"784000AA59000000000000000000000000000000000000000000000208017DAA",
INIT_2E => X"A2D57FFFFF7AEBFF55FF8028A00512EAAB45007FFFF55082EA8AAA087FC2010F",
INIT_2F => X"5512AAAA085D04174100800021FF002EA8BEF5D0428ABA595557555AAFBC2000",
INIT_30 => X"00FF802ABAA04552ABFF597FD74BAF7AAA8B45AAFBD54005D7BD54AAF7800215",
INIT_31 => X"5FFAAFBC0000AF843FF5500003FF55AAFD6AB4551002ABEF0055555550004020",
INIT_32 => X"DEB0A2FD5600051537DE005D557DE005D7BE8AA85555400100879560AA592F95",
INIT_33 => X"17545FFD5421FF5D0428BEF0079FCABA598400010F7AA8215555003FEAAAA843",
INIT_34 => X"0000000004001FFAAFBEAA105D2E955FF557BD75EFFBBCD415521FBFDF450004",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000010000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(4),        -- Port A data input
DOA(0)   => data_read_a_hi_256(4),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(4),        -- Port B data input
DOB(0)   => data_read_b_hi_256(4),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_5_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50DB0A0791B1B41694368283C81F9996A091A32152007AB36B20E03C040C002",
INIT_01 => X"880015C49830884C446A40000C34C24841280A00084000C8C212892EEA953231",
INIT_02 => X"408F417400B1D9100002171C1FA20171124E6AA00D8633F8CD09DBFBBB972F7C",
INIT_03 => X"88538F0182058082D800C3314722DC08A34084A100C4D7C99208521063D00148",
INIT_04 => X"F45E41AFAF420996B8411CA282F80A9091224800A2C61490363080C8A4000308",
INIT_05 => X"0EA416069640420901A01505C4410020C6E228DC30532839B043289D9C005031",
INIT_06 => X"13992D9AF8C74E92B7B568D19708C038AFFA89F0B9348C9204C389672407EF12",
INIT_07 => X"6255000016053C18162589725146F442222CE6AF844012BE795224458BA4DE0F",
INIT_08 => X"4F3F00503B4AE104B5347230418190420821006016FC18843630D285FC416CB4",
INIT_09 => X"EEA33E700340902C4424C442B0344724066C56C2248130A2D9C185B24A24832B",
INIT_0A => X"315325008348CC40AB570500204462508135D5AA593E043731E9B18A98440137",
INIT_0B => X"E0CD463C5813804E0258E0358E02D8E03D8E0258E03D8E02D8E03447012C701E",
INIT_0C => X"F8DE3C27CA181E5D710664A5F140C14BD32A2E281992940AFAA15C3FC0836310",
INIT_0D => X"F000BE0FC80020130841840308653FF0313FE92C23FB1EECB367C0F3E378F0BC",
INIT_0E => X"F000BE0FCD806FFFAF0AE83080E2AEB2F0F1E01BE53FE1F000BE0FC41BE53FE1",
INIT_0F => X"0231F0BF9E3F02A7FFD63669C0E008C3CB7F041BE1BFE1F000BE0FC41BE1BFE1",
INIT_10 => X"30180309A0F83FE2B87C7D006FFF9F1A7806013879BAA78FC103FF5F1F12F038",
INIT_11 => X"39E9C1DBF8A30C2098DBE2FF7F2320483136F200A822CBACAB9DDEB7F9BC291F",
INIT_12 => X"004C72BEC95FEF64E4090626DF15B7D1C6184131B7980DFFFC03F00003F01FB9",
INIT_13 => X"1DFFFA0A3C0202B8776AE7A7C9CBFFF060703080E29F1B79E9F6427EFE901C0E",
INIT_14 => X"2B716CA5C56620590350ACD3A7D5B7EFAC6DFC8C0312A0024B83F07F3999E9F2",
INIT_15 => X"F0BCAF3BC2F3BC6F0BCEF2BC2F3BC6DBC67C251104A2261253904580207E1C81",
INIT_16 => X"1BCEF0BC2F3BC2F1BCEF0BC6F2BC2F1BCAF1BC6F2BC6F2BCAF1BC2F3BC6F2BCE",
INIT_17 => X"BCEF0BC2F3BC2F1BCAF1BCAF3BC6F0BCEF0BCEF2BC6F2BCAF1BCAF1BC2F3BCAF",
INIT_18 => X"69CFEF73B6FFE7436DB6FD0831518424965B4D2492CB69AF1BCEF0BC6F2BC6F0",
INIT_19 => X"F7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF3EF9FBFBB9E79E7BEBCB7",
INIT_1A => X"DEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDF7DF7DF7D",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF29FDAF77BBDDEEF77BBDDEEF77BBD",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"AAA2802AA10FFFFFDE0008556AABA5D2ABFFEFFF800000000000000000000000",
INIT_1F => X"ABAF7AAA8BFFAA802ABFF087FFDF5508003FEBA087FD54BA0804154005555574",
INIT_20 => X"54AAF7D168B45AAAABDF55AA802AA1000003FEBA00002AABA5D2EBFEBAAAD16A",
INIT_21 => X"3DE005555575EFA2D142145A2FFE8B45FF80001555D2E955FFFFD5421EFAAFFD",
INIT_22 => X"FC00BA5D5568AAAF7AAAAAAAAA802AABA082E954005500021FF5D2EBFF550000",
INIT_23 => X"D5420AAAA843DFFFAAD1554005D7FD74AAAA840014500517FFEF007BEABFF5D7",
INIT_24 => X"2AABDE0055517FF555504154BAA2FBEAA105D2E97410FFD16AAAA5D2ABDEBAFF",
INIT_25 => X"000000000000000000000000000000000000000028BFF0855555455500174BAA",
INIT_26 => X"21E84124285C51574BAB68A2DA00FFFFFFE38085F6FA92552AB8FEFF78000000",
INIT_27 => X"925D2AB8EBABEDB6AA92F7AAA8BC7B68A28BC70075FDF45080A3AEAA007BD248",
INIT_28 => X"5FFFFD1471D7AAFBD0492EBD56DB7DBEAEBFF55BE842AA105D0A38EBA1C0428A",
INIT_29 => X"21FF492AB8F7D1C0438E38145B575EFA2DB45145B6F5EFB6DF78E05145552A92",
INIT_2A => X"7DFC70875EABC7557FC20AA415F68AAAF7AAAAA82BE8A28A9214249740041000",
INIT_2B => X"B6FABA542ABAE2AF7DF470AABE8A3AFD7A2DF55400557FD54AABE84001C55551",
INIT_2C => X"5557545490012482B6A0BAE2849043AFED1C0E10492B6FFEFA105D2A95410FFD",
INIT_2D => X"D2AAABEFFB8000000000000000000000000000000000000000000000428BEF00",
INIT_2E => X"082EA8AAA087FC20105504000AA5955554BAFFAEBDE10F7FBFDEBA007BFDE005",
INIT_2F => X"0512AA8AAA5D0028A005D2AA8ABAF7FBE8A00FFAEAAB45F3AAAAB4500557FF55",
INIT_30 => X"EFFFAA97545552A821EFFBD557555AAFBC2000A2D57FFFFF7AEBFF55FF8028A0",
INIT_31 => X"A005D04174100800021FF002EA8BEF5D0428ABA597FD55FFA2FFD5555FFD57FF",
INIT_32 => X"54AAF7800015551517DF45005168B55557FC0012087FEAABAF7AAAAA10F3AAAA",
INIT_33 => X"FFE005D2A95410F7FFFFEBA5D2EA8ABAFBFFD74BAF7AAA8B45AAFBD54005D7BD",
INIT_34 => X"00000000002ABEF005555555000402000FF802AAAA04452ABFF592E80010FFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000060000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(5),        -- Port A data input
DOA(0)   => data_read_a_hi_256(5),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(5),        -- Port B data input
DOB(0)   => data_read_b_hi_256(5),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_6_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10800B0061A01002840002C030028180004003220200403312301C4389B2082",
INIT_01 => X"060009C838394848188160000C42426041000000090800090210090000510200",
INIT_02 => X"00043040009001100000061000018070002408000000000648080000001210E0",
INIT_03 => X"0000800002054081020080801200A0000300008000201184681A0000410C4800",
INIT_04 => X"0808801040000001401048008100022401400002024024053200020089000100",
INIT_05 => X"0240040408402202002000C200400020A50000A0000010010001260808000520",
INIT_06 => X"44000881064500004600000013088002840C240F5048011200010000440C0146",
INIT_07 => X"0241914041FE83E010040110110003040020402A0000003E1000000488000201",
INIT_08 => X"8001BF002C4A01041B112020200110024029006FE09081002004902000012068",
INIT_09 => X"0083FE38A040100281353150ACB645AEF8C01404448000008011061204200108",
INIT_0A => X"3103AD0413424E4014D627C470462200011504420C0A962A2189002881404060",
INIT_0B => X"46C1060C16C96D15B0425B0425B1425B1425B0C25B0C25B1C25B1512D8212D82",
INIT_0C => X"009000140401100601016600A040220203A004480598010248000D0010420C0C",
INIT_0D => X"0000A01033A00013000000000018800F2400091081100C0090A5008200410020",
INIT_0E => X"0000A0103142000000000000000000455D0018100000000000A0103410000000",
INIT_0F => X"000000466800C200000000000000000001A0F4100000000000A0103410000000",
INIT_10 => X"00000000000024094680014200000000000000000041E8002900000000000000",
INIT_11 => X"F000322000000000000D1A000000000000034D240C2000502000000000000000",
INIT_12 => X"000000403F4000000000000068D24000000000001A60F0000000000000002007",
INIT_13 => X"C0000000000000000087C0003014000000000000000025D00008958000000000",
INIT_14 => X"02000000000814C219500150002800101280000000000000000000086670000C",
INIT_15 => X"8120C82208812048120882208892055A0060011280222413130449010301F051",
INIT_16 => X"3200802008320C82200802048320C82200812048320880200812048220880204",
INIT_17 => X"20C83208812048020883204802048120882204812008220C8220081204822088",
INIT_18 => X"79CFF1FE1E9F52ABEF9EFE8150120EC718638E38E30C71C812088220C8120080",
INIT_19 => X"71C71C71C71C71C71C71C71C71C71C71C71C71C71C736D9DBD9BBEFBEFBEBEF1",
INIT_1A => X"CFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FC71C71C71C",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCF29A7F3F9FCFE7F3F9FCFE7F3F9F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000607FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"EFA2FBD54BA5555554BAAAFBC20BA5D7BEAAAAFF800000000000000000000000",
INIT_1F => X"EBA0855421455555574AAA2802AA10FFFFFDE0008556AABA5D2ABFFEFFF843DF",
INIT_20 => X"DF5508003FEBA087FD54BA000415400550428AAAAA84021FF007BD54BAAAD17D",
INIT_21 => X"A8BFFAAD1554BA002A95555A28417400AAFBE8ABAF7FFD54AAAA802ABFF087FF",
INIT_22 => X"BD5545080417555A2D17FE1000003FEBA00002AABA5D2EBFEBAAAD16AABAF7AA",
INIT_23 => X"D5421EFAAFFD54AAF7D168B45AAAABDF55AA802AA100000001EF087FEAA00FFF",
INIT_24 => X"F80001555D2E955FFFF843DEAAA2803DFEF0855401FF082EA8B555D7FC21FFFF",
INIT_25 => X"0000000000000000000000000000000000000055575EFA2D142145A2FFE8B45F",
INIT_26 => X"2552AB8FEFF78E3DFFFAAFFD04AA415B52492B6F5C20825D7FE8A92FF8000000",
INIT_27 => X"EF147BD2482BED57AE921451421555551574BAB68A2DA00FFFFFFE38085F6FA9",
INIT_28 => X"4BAB68A28BC70075FDF45080A3AEAA007BD24821C04124281C0E2DA82BE8E001",
INIT_29 => X"8EBABEDB6AA92F7AAA8BC7B6D5524AA14209557DA28E15400BEF1EFA92FFFFD2",
INIT_2A => X"071FF0071EDA38F7F1D5555000417545B6D178E281C0A38EBA1C0428A925D2AB",
INIT_2B => X"4A8B555C7FC2147F7D1471D7AAFBD0492EBD56DB7DBEAEBFF55BE842AA105D0E",
INIT_2C => X"DB45145B6F5EFB6DF78E05145552A925FFFF8E3DE82BE8E38FFF0851401C7082",
INIT_2D => X"57FE8A00F38000000000000000000000000000000000000000000005B575EFA2",
INIT_2E => X"F7FBFDEBA007BFDE005D2AAABEFFBAABDFEFAAFBC00BA007BC0000FFD5420005",
INIT_2F => X"A592ABFE00F7AA821FF557FC0010F7D168A105D55421455155554BAFFAEBDE10",
INIT_30 => X"10F7D57DE00FFFBC00AAFBAAAAB4500557FF55082EA8AAA087FC20105504000A",
INIT_31 => X"AAA5D0028A005D2AA8ABAF7FBE8A00FFAEAAB45F3D5400BA5504155EFAAAE954",
INIT_32 => X"FF55FF8028A00512E975FF08557FEAAF7D157545080417545F7D56AAAA592AA8",
INIT_33 => X"AABEF005542155000028B555D7FC2145F3D557555AAFBC2000A2D57FFFFF7AEB",
INIT_34 => X"000000007FD55FFA2FFD5555FFD57FFEFFFAA97545552A821EFFBAABDE00F7AA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000048000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(6),        -- Port A data input
DOA(0)   => data_read_a_hi_256(6),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(6),        -- Port B data input
DOB(0)   => data_read_b_hi_256(6),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_7_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10844B00482258A2842112C02450418800002300500030B313300C418992002",
INIT_01 => X"020009C23838684D1C20E0000E11424840000000080000080200000000110204",
INIT_02 => X"000520700CA08910000206101180803081144880010400044808000000122160",
INIT_03 => X"000080040305208000008000328080040304008020303194289A000041484800",
INIT_04 => X"08088000000000010000CA008008060441000000028234493410820191000000",
INIT_05 => X"03500404000022020020044000000C208400408000001000984005949C002928",
INIT_06 => X"54000881044500004680000013008002940C24001A4A010200018920646410C7",
INIT_07 => X"22510040400500011204813015012204002040280000013E1000000488000201",
INIT_08 => X"9001A0602C4A01051B132820208001024069004008908002120851420001226A",
INIT_09 => X"01100020A2401008A20404E08200A05000A4264640800022C8198C4E05200018",
INIT_0A => X"20002000024040400050450440C48A0041140C420B0904208800904286000008",
INIT_0B => X"50822002120D2134800648006480064800648106481064810648193240432404",
INIT_0C => X"284A142288042A5C24202451505E00A621A5220A8091444040188C001B41210A",
INIT_0D => X"00F001F021141A12004104020810B000100000000109064C80010050A3285194",
INIT_0E => X"00F001F027420000400004C3201C514408081C1014800000F001F02810148000",
INIT_0F => X"E00E0E404100E200040900000B0380383480C81014800000F001F02810148000",
INIT_10 => X"4160C0301D07001D0402034200004000019860078641004039000180400002C0",
INIT_11 => X"08103BA0104810C8462416E8040446120C890814600010512000000080028400",
INIT_12 => X"98038D4030DD008088C2419120B740209021908C4846FC000200030F000FE006",
INIT_13 => X"DD000100411C81078884204035DC00201804C3201C60A408100DD58010440130",
INIT_14 => X"412024202211148019064200402A32901A8000B2048902C0807C0E00C448100D",
INIT_15 => X"50942509425194651946519465894619421421102000269243854D8002000250",
INIT_16 => X"19465194E50942509425094E51946519465094A50942509425194E5194651942",
INIT_17 => X"9425094251946539465094250946539465194250942509465194650942509425",
INIT_18 => X"0000000000000000000000080150890820800041041000052942509465194653",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF21E6C000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"AAF7D5575455D557DFEF002AAAB55002E820AAAA800000000000000000000000",
INIT_1F => X"B55007FD74AAAA843DFEFA2FBD54BA5555554BAAAFBC20BA5D7BEAAAAFFFBC00",
INIT_20 => X"AA10FFFFFDE0008556AABA5D2ABFFEFFFAAAAAAAF7D57FFEFF7D555555A2AEAA",
INIT_21 => X"42145552ABDFEFFFAA801EFFFFBFDF550000175555504175450055574AAA2802",
INIT_22 => X"A975EF00003DF55555168A00000428AAAAA84021FF007BD54BAAAD17DEBA0855",
INIT_23 => X"802ABFF087FFDF5508003FEBA087FD54BA000415400557BD74BAFFD140000082",
INIT_24 => X"AFBE8ABAF7FFD54AAAAAEA8ABA55557FEAAA2843FF55A2AEA8B55AAAABDEAAFF",
INIT_25 => X"0000000000000000000000000000000000000051554BA002A95555A28417400A",
INIT_26 => X"25D7FE8A92FFFFC70BAE3D155555415178FD7082EAAB550820870BAAA8000000",
INIT_27 => X"FFEBD55557DBEA4AFB550871D7482AA8E3DFFFAAFFD04AA415B52492B6F5C208",
INIT_28 => X"5550051574BAB68A2DA00FFFFFFE38085F6FA92552AB8FEFF7A0ADABAEBD578F",
INIT_29 => X"2482BED57AE921451421555524BDFD7FFA4801D7F7F5FDF55000E17545410E17",
INIT_2A => X"D2482E3D1450381C20905EF08003AF55415F6DA38080E2DA82BE8E001EF147BD",
INIT_2B => X"AAFB55ABA0BDE02EB8A28BC70075FDF45080A3AEAA007BD24821C04124281C7B",
INIT_2C => X"209557DA28E15400BEF1EFA92FFFFD24BAB6A4A8A82495F78E92AA843DF45BEA",
INIT_2D => X"800174BAA680000000000000000000000000000000000000000000055524AA14",
INIT_2E => X"007BC0000FFD542000557FE8A00F3FFD54BAAAD15754508556AB45002AA8B450",
INIT_2F => X"FFB803DEAAAAD56ABEFAAD5575EFF7803DF45085557410AEAABDFEFAAFBC00BA",
INIT_30 => X"55082E97555002E955550C55554BAFFAEBDE10F7FBFDEBA007BFDE005D2AAABE",
INIT_31 => X"E00F7AA821FF557FC0010F7D168A105D554214551003FF45FF8400145FFD57FF",
INIT_32 => X"20105504000AA597FC2010A2D1554AA5500021EF000028B55087BFDEBA042ABF",
INIT_33 => X"E8A00A2803FF45F7AABDF55AA843FE10AEAAAAB4500557FF55082EA8AAA087FC",
INIT_34 => X"0000000055400BA5504155EFAAAE95410F7D57DE00FFFBC00AAFB8028A00007F",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000007FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(7),        -- Port A data input
DOA(0)   => data_read_a_hi_256(7),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(7),        -- Port B data input
DOB(0)   => data_read_b_hi_256(7),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_8_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000B0000040042840002C0000001800000070000000033022000000000086",
INIT_01 => X"000009C21838284D1C2160000E12426840000000180800080200080040510200",
INIT_02 => X"0001004000900110000006100080003000240800014400004808000000122160",
INIT_03 => X"00008000020440810002A0801010A0044300000000200086011A000040404800",
INIT_04 => X"8000801000020401400040408108022029400000124004041200000089000100",
INIT_05 => X"02080424085022020000040200480020850010A0002010010120060800040400",
INIT_06 => X"50000880006500000680000011008006840C200018C1010200018920E0640102",
INIT_07 => X"426000404005000112048130150120240020400A0000013E1000000488000010",
INIT_08 => X"220100402C42010413110020200100024029004000A200002004902200012141",
INIT_09 => X"0000000080400008010410A2940A45240040140440800022C8388E1200A00008",
INIT_0A => X"00420100020048405000070440C0000001140412090000000021002081000048",
INIT_0B => X"0000000800000100011000010000100001000010000100001000010000880008",
INIT_0C => X"001000040001100008012008004020102180800804802000C0080D00100A0008",
INIT_0D => X"0FF0000002200A1200410402080080003000091085100C008124008000400020",
INIT_0E => X"0FF000000140000040F517CF600000000104081010001E0FF00000001010001E",
INIT_0F => X"E000000000804200000809963F1F80000000001010001E0FF00000001010001E",
INIT_10 => X"CFE7C0F00000000000810140000040E587F9E000000008100900008000ED0FC7",
INIT_11 => X"00021040030C73D80000021000585F3600000020240020102000000802419660",
INIT_12 => X"F80000000042000B0BD6C0000010800618E7B000000C000003F80FFF00000000",
INIT_13 => X"800005D5C3FD800000000008180000078A8FCF600000000002028001006AA3F1",
INIT_14 => X"020000000008808219002100100C000041120370DCAD1FC18000000000000202",
INIT_15 => X"8020080200812048120481204812055A04604930A02026934215410102000110",
INIT_16 => X"0200802008020080200802048120481204812048120481204802008020080200",
INIT_17 => X"2008020081204812048120481200802008020080200802048120481204812048",
INIT_18 => X"414A87D78AF42143CEBAC88151120A0000000000000000081204812008020080",
INIT_19 => X"F3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF7E799B1BEB65B65948051",
INIT_1A => X"C3E9F0FA7C3E9F0FA7C3E9F0FA7C3E9F0F87C3E1F0F87C3E1F0F87CF3CF3CF3C",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF1B5DA9F0FA7C3E9F0FA7C3E9F0FA7",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"0000043DF55087BC01EF007FD75FFFF84000AAFF800000000000000000000000",
INIT_1F => X"E10A28028AAAAAFBC00AAF7D5575455D557DFEF002AAAB55002E820AAAA84000",
INIT_20 => X"54BA5555554BAAAFBC20BA5D7BEAAAAFFAA95545552ABFE00087BC00AA082EBF",
INIT_21 => X"D74AAAAD57FF45002A975FF007BE8BFFA2FBFFFFFAAD5400AAFF843DFEFA2FBD",
INIT_22 => X"BE8A00082A97410F7D5555EFAAAAAAAAAF7D57FFEFF7D555555A2AEAAB55007F",
INIT_23 => X"55574AAA2802AA10FFFFFDE0008556AABA5D2ABFFEFFFAA82000555555545AAF",
INIT_24 => X"00017555550417545000015545087BC2010AAD54014500516ABFFA2AABDF4500",
INIT_25 => X"000000000000000000000000000000000000002ABDFEFFFAA801EFFFFBFDF550",
INIT_26 => X"50820870BAAA8407000140038F450075C71FF087BD75D7FF84050BAEB8000000",
INIT_27 => X"10007FC50BA002ABFE00AA8A2AABABEFFC70BAE3D155555415178FD7082EAAB5",
INIT_28 => X"082EB8E3DFFFAAFFD04AA415B52492B6F5C20825D7FE8A92FFA497545552AB8E",
INIT_29 => X"557DBEA4AFB550871D7482AAD17DF451C24955EF0875EFBD7B6F1FFFC7BEDB45",
INIT_2A => X"87000415B5057DAAFBE8A10082092410EBD5505EFB6A0ADABAEBD578FFFEBD55",
INIT_2B => X"B6ABC7B6AABFFED0051574BAB68A2DA00FFFFFFE38085F6FA92552AB8FEFF7AA",
INIT_2C => X"A4801D7F7F5FDF55000E17545410E17555000E17545007BC0000BED14217D005",
INIT_2D => X"784174AAA280000000000000000000000000000000000000000000024BDFD7FF",
INIT_2E => X"08556AB45002AA8B450800174BAA684174105D042AB550055555FF007BD7555F",
INIT_2F => X"0F384175555D2EA8A00087BD74BA082EBDE10AAAEA8ABAF7FFD54BAAAD157545",
INIT_30 => X"55FFD57DF55FFFBD5400A2AABDFEFAAFBC00BA007BC0000FFD542000557FE8A0",
INIT_31 => X"EAAAAD56ABEFAAD5575EFF7803DF45085557410AED17FF455D04155FF00557DF",
INIT_32 => X"DE005D2AAABEFFBAE97410087BC21EFA2FFEAA00000002010A2D5421FFFF803D",
INIT_33 => X"C0010FFD1401EF087FE8B55FFAEBDFEF0855554BAFFAEBDE10F7FBFDEBA007BF",
INIT_34 => X"00000000003FF45FF8400145FFD57FF55082E97555002E955550C2E95555087B",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000020000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(8),        -- Port A data input
DOA(0)   => data_read_a_hi_256(8),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(8),        -- Port B data input
DOB(0)   => data_read_b_hi_256(8),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_9_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00018248A2840112C00002C18000002300500030B3132000400812002",
INIT_01 => X"A140098218302849180060000C004240413C0A61590001D90213C90008510204",
INIT_02 => X"102008700CB089100002061031285074810448800104008048080080001210E2",
INIT_03 => X"00008015074608840390A0040040800203140000A00010800408108448020042",
INIT_04 => X"082080400004A00100000100840602020100000002C2344156108201811801C0",
INIT_05 => X"0200048480011502049500280020CC2084000080008010019161249C9C002188",
INIT_06 => X"70000881004500004E01020411D08000940C00001800010200018B20206C0102",
INIT_07 => X"EA70C0040005000312048130150100040020404A0000017E10408104C8000110",
INIT_08 => X"000000402C220104131004202081120050A5104000A204617201D10801002000",
INIT_09 => X"000800002F4924003085E51420A0100400641E4E40800022C8088C1220200908",
INIT_0A => X"20102000024040484028450001648C2229150400080244000401900284000440",
INIT_0B => X"0880110901081110411204112040120411204012041120401204111020090208",
INIT_0C => X"685B34A688841A5C21200101A01A0004009024028004044248404D00104B2100",
INIT_0D => X"0000A01000000213000000000000B0001000010000190E44802002D1A168D0B4",
INIT_0E => X"0000A010014000000000000000000040500008100400000000A0100410040000",
INIT_0F => X"0000004608004200040000000000000001A004100080000000A0100410008000",
INIT_10 => X"00000000000024080000014000000000000000000040A0000900010000000000",
INIT_11 => X"300013E010000000000D00F804000000000340000C0000102000000080000000",
INIT_12 => X"00000040091F0000800000006807C000800000001A0CFC000000000000002001",
INIT_13 => X"DD000000000000000082C00019DC002000000000000021500006D58010000000",
INIT_14 => X"03206420000000C019502050000C32901A800080000000000000000860100006",
INIT_15 => X"D1B46D1B46D0B42D0B42D0B42D8B424342342832002A24921082158802001011",
INIT_16 => X"0B42D0B42D0B42D0B42D0B46D1B46D1B46D1B46D1B46D1B46D1B46D1B46D1B46",
INIT_17 => X"B42D0B42D1B46D1B46D1B46D1B46D1B46D1B46D1B46D1B42D0B42D0B42D0B42D",
INIT_18 => X"89999E91BCD1512B871C4A0100000000000000000000000D0B42D0B42D0B42D0",
INIT_19 => X"A28A28A28A28A28A28A28A28A28A29A69A69A69A69A51C200807249041202AE6",
INIT_1A => X"8349A4D068341A0D269341A0D269341A0D068341A0D068341A0D068A28A28A28",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF2DA921A0D269341A0D068349A4D06",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"45A280154BA5555401EFFFD5421EFA2FFFFF555D000000000000000000000000",
INIT_1F => X"5EF00557DF555D040000000043DF55087BC01EF007FD75FFFF84000AAFFD57DF",
INIT_20 => X"75455D557DFEF002AAAB55002E820AAAA843DFEF00517DEBA007BFDFEFFFD157",
INIT_21 => X"28AAAAAAABDF45F7803FFEF555568AAAF7802AA00FFFBD7555087BC00AAF7D55",
INIT_22 => X"BD54BA550417400085155555082A95545552ABFE00087BC00AA082EBFE10A280",
INIT_23 => X"043DFEFA2FBD54BA5555554BAAAFBC20BA5D7BEAAAAFFFBC00AA552E95545087",
INIT_24 => X"2FBFFFFFAAD5400AAFF8402000A2FFFDF555D7BE8BFF5D51575EFA280175555D",
INIT_25 => X"00000000000000000000000000000000000000557FF45002A975FF007BE8BFFA",
INIT_26 => X"7FF84050BAEBDF78F45B68010482415B471C7E3DF451EFBEFBFAF45490000000",
INIT_27 => X"82007FFAFEFE3DB505EF1C5B7AF45490407000140038F450075C71FF087BD75D",
INIT_28 => X"5451C7FC70BAE3D155555415178FD7082EAAB550820870BAAA8438FFF00517DE",
INIT_29 => X"50BA002ABFE00AA8A2AABABEAEB8F45F78A3DFD741516DAAAE38E2DA28EBFFD5",
INIT_2A => X"C20BA5D2E905550071D54825D0A1543808515756D1C2497545552AB8E10007FC",
INIT_2B => X"5505FFBE801256D490E3DFFFAAFFD04AA415B52492B6F5C20825D7FE8A92FFFF",
INIT_2C => X"24955EF0875EFBD7B6F1FFFC7BEDB45082EB8002000AAFFFDF6D417FEABEF5D5",
INIT_2D => X"7FBE8B5500000000000000000000000000000000000000000000000517DF451C",
INIT_2E => X"0055555FF007BD7555F784174AAA2FBEAB45F78402010007BD5545AAFFD55EFF",
INIT_2F => X"AA68028BEF00517FE10007BE8BFFAAFFC01FF557FE8B550004174105D042AB55",
INIT_30 => X"AAAAAEBFEAAAAFFD5545557FD54BAAAD15754508556AB45002AA8B450800174B",
INIT_31 => X"5555D2EA8A00087BD74BA082EBDE10AAAEA8ABAF7AAAAB45F7AEBFF4508557FE",
INIT_32 => X"2000557FE8A00F3FFC00BA552E80145005557400552A954BA0051575EF550417",
INIT_33 => X"FDFFF007FE8BFF5551401EFF784021FF002ABDFEFAAFBC00BA007BC0000FFD54",
INIT_34 => X"00000000517FF455D04155FF00557DF55FFD57DF55FFFBD5400A28400010A2FB",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000040000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(9),        -- Port A data input
DOA(0)   => data_read_a_hi_256(9),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(9),        -- Port B data input
DOB(0)   => data_read_b_hi_256(9),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_10_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00018248A2840112C00002C18000202300500030B3132000400992006",
INIT_01 => X"A140098218302849180060000C00424040000000080000080200090008510204",
INIT_02 => X"102100400C8001100000061000A8503401044880010400004808000000122160",
INIT_03 => X"000080150746088401908000100080020304000020201080001A108448404842",
INIT_04 => X"800080400004A001000040008406020201000000020004401000000180180080",
INIT_05 => X"02000484800133020495040800208C20A4000080000010000001249010042008",
INIT_06 => X"50000881004500004681020411808000940C20001800010200018920206C0102",
INIT_07 => X"024084044005000112048130150120040020400A0000013E10408104C8000010",
INIT_08 => X"000100402C020105131100200000124250A51040088084614001110801012000",
INIT_09 => X"00080082CD09240820800000000000040000180840800022C8088C1220200108",
INIT_0A => X"841201000200484910000F050560262229140402080200A00402000484140400",
INIT_0B => X"0010118900080010000200102001020000200002001020010200001000010008",
INIT_0C => X"408120900404004821202001F05E00040180260A8080044240004C0010800228",
INIT_0D => X"0000A01000000813004104020800800030000800010008088124020102008100",
INIT_0E => X"0000A010014000004000000000000040500008101480000000A0100410148000",
INIT_0F => X"0000004608004200040900000000000001A004101480000000A0100410148000",
INIT_10 => X"00000000000024080000014000004000000000000040A0000900018040000000",
INIT_11 => X"3800100010480000000D00000404400000034000282000102000000080028000",
INIT_12 => X"00000040090000808800000068000020900000001A0000000200000000002001",
INIT_13 => X"80000100000000000082E0001000002018000000000021580000800010440000",
INIT_14 => X"00004000000004C0195000500008000000000082008000000000000860180000",
INIT_15 => X"0100401004010040100401004090055804404110802A24921317580802001011",
INIT_16 => X"0000000000000000000000040100401004010040100401004010040100401004",
INIT_17 => X"0040100400000000000000000000000000000000000000000000000000000000",
INIT_18 => X"215281FC1A72E2486AAA40A85052020000000000000000001004010040100401",
INIT_19 => X"51451451451451451451451451451451451451451452AA83330A8A28A29EA8D1",
INIT_1A => X"5CA6532994CA6532B95CAE572994CA6532994CA6532994CA6532994514514514",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF31CE2E572994CA6532994CAE572B9",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"10AAFBE8AAAA2D540000F7D57DF55A2AABFFEF08000000000000000000000000",
INIT_1F => X"F45FFFBC2010AAD57DF45A280154BA5555401EFFFD5421EFA2FFFFF555D003FE",
INIT_20 => X"DF55087BC01EF007FD75FFFF84000AAFF8002155AAFFE8B45AAD540000087FFD",
INIT_21 => X"7DF555D517FEBA082A801EFF7FBD5400FFD568B555D00155EF08040000000043",
INIT_22 => X"BFDE00A2FBC0145005168A10AA843DFEF00517DEBA007BFDFEFFFD1575EF0055",
INIT_23 => X"7BC00AAF7D5575455D557DFEF002AAAB55002E820AAAA803FEBA082AAAAAAF7F",
INIT_24 => X"7802AA00FFFBD7555082E82155FFAEAAB55AAD568B455D00154BAFFFBD75EF5D",
INIT_25 => X"000000000000000000000000000000000000002ABDF45F7803FFEF555568AAAF",
INIT_26 => X"FBEFBFAF4549003DE10BEF5EDAAAAAD547038EBD57DF7DA2AEB8FC7000000000",
INIT_27 => X"6DAADF470280075FFF45E3F1C7038A2DF78F45B68010482415B471C7E3DF451E",
INIT_28 => X"5C7000407000140038F450075C71FF087BD75D7FF84050BAEB8002155BEF5EDB",
INIT_29 => X"AFEFE3DB505EF1C5B7AF45495B7DEAA0824851EFEBFBD2410EBD168B7D410A17",
INIT_2A => X"38EAA0824A8AAAEBF5FAE28AAF1C2155005F68A10A28438FFF00517DE82007FF",
INIT_2B => X"4104AAF7F1D75EF557FC70BAE3D155555415178FD7082EAAB550820870BAAA80",
INIT_2C => X"8A3DFD741516DAAAE38E2DA28EBFFD55451C2087155EBA4A8B7DAADF68B7D410",
INIT_2D => X"2AEAAB55000000000000000000000000000000000000000000000002EB8F45F7",
INIT_2E => X"007BD5545AAFFD55EFF7FBE8B5500043FE00F7D17FEBAA2D5574BAAAD17DFEFA",
INIT_2F => X"AA28002155FFD17FFFFA2FBD74BA00557FF45A2D5554AAA2FBEAB45F78402010",
INIT_30 => X"00AAD16ABFF002A975450004174105D042AB550055555FF007BD7555F784174A",
INIT_31 => X"BEF00517FE10007BE8BFFAAFFC01FF557FE8B55007FFDEAA0004175FFA2FBC20",
INIT_32 => X"8B450800174BAA68428AAA08042AABAAAD56AABAAAD140155087FEAA10A28028",
INIT_33 => X"2ABEFAAFBE8BFF0004020AAFFD5555EF557FD54BAAAD15754508556AB45002AA",
INIT_34 => X"000000002AAAB45F7AEBFF4508557FEAAAAAEBFEAAAAFFD5545550015555A284",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000047FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(10),        -- Port A data input
DOA(0)   => data_read_a_hi_256(10),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(10),        -- Port B data input
DOB(0)   => data_read_b_hi_256(10),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_11_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10180B05A0010402840602C2D001019000000300000000330A20080EC180002",
INIT_01 => X"AB400984B830084C1820E0000C36424840000000080000088200000802112220",
INIT_02 => X"102A68440080011000000618062AD03502640800010410424908136019920868",
INIT_03 => X"001282118644C88481908001106088022300000080F4925CDC9A10844A9A4842",
INIT_04 => X"401280480004A1011000418084460002E12000000200040010000040A8000000",
INIT_05 => X"0FC8048484011502059511488020802084400888001110000000050000005400",
INIT_06 => X"1011088AE24500001631024511C08004A70AA40008B90D0200018B60A0650D45",
INIT_07 => X"020011005405000910040150110041040024400D800002BE18408104C9205908",
INIT_08 => X"89390040280241041D175820000001020061004004800567403512A801014C46",
INIT_09 => X"050800E20D09A424C5840400808000040680180840800022D8288E946CA00833",
INIT_0A => X"85002000024040410A000D0504408C32E915D9C208050084840201A099100400",
INIT_0B => X"B01011934A005101431CA821CA831CA821CA831CA831CA821CA83165410E5410",
INIT_0C => X"00010080028000010402214850444091019B02080885200042A9CC001000003A",
INIT_0D => X"5A5018C5A0A00812004104020808B00030000808024008008325820000000000",
INIT_0E => X"5A5018C5AB0062C38A4DB680A0D8241500D5761B011986695014A96E1A811986",
INIT_0F => X"42056A289A1BB2078A922DA2A8B180A2600AAE1A811986695014A96E1B011986",
INIT_10 => X"05AA429189B60AC43C6C7F0272C3841DB528802CAB18468F4101621B1BAC8455",
INIT_11 => X"C003104289A668B8CAB270106338317A3D94392020224ACDE215883078681B5C",
INIT_12 => X"804B020A06020C67061BC785938085134CD551BCA1C90006C0C2958502861120",
INIT_13 => X"80819A5539D503336D61056ABA006282806CA64090B89E015AAA880E48382EB8",
INIT_14 => X"40000000E808989003066E03513E41470126C6284B2D20410AB4503089C00A82",
INIT_15 => X"0000000000000000000000000000041800400110200026124202500802000800",
INIT_16 => X"1004010040100401004010000000000000000000000000000000000000000000",
INIT_17 => X"0040100401004010040100401004010040100401004010040100401004010040",
INIT_18 => X"C110083018162148420840280050800000000000000000001004010040100401",
INIT_19 => X"000000000000000000000000000001041041041041003882928E0000000AA0C4",
INIT_1A => X"0000000000008040000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3E0FC000000000000020100000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"EFAA842ABEFA280155EFFFFBC01EF08554000055000000000000000000000000",
INIT_1F => X"F4508514000000003FE10AAFBE8AAAA2D540000F7D57DF55A2AABFFEF0804155",
INIT_20 => X"54BA5555401EFFFD5421EFA2FFFFF555D51575FFA2FFD75FF550015400FFFBFF",
INIT_21 => X"C2010AAD568AAAAAD142145FF80155EF0051555FF0804155FFF7D57DF45A2801",
INIT_22 => X"01540008514215555003DFFFA28002155AAFFE8B45AAD540000087FFDF45FFFB",
INIT_23 => X"040000000043DF55087BC01EF007FD75FFFF84000AAFF802ABFFA2AABFE10080",
INIT_24 => X"FD568B555D00155EF085168B45085142010FFAE800AA5D7BFDF45F7FFEAA0000",
INIT_25 => X"00000000000000000000000000000000000000517FEBA082A801EFF7FBD5400F",
INIT_26 => X"DA2AEB8FC70000175EFB6802DBC7BE8A155EFE3FBC71FF145B42038550000000",
INIT_27 => X"EF550E15400E3F1FFF7D085B420381C003DE10BEF5EDAAAAAD547038EBD57DF7",
INIT_28 => X"5C7F7DF78F45B68010482415B471C7E3DF451EFBEFBFAF45495F575FFBEF5D05",
INIT_29 => X"70280075FFF45E3F1C7038A2DB68ABAB6D145145FF84155D7085B555C7140410",
INIT_2A => X"28BEFBEA4BDE28140A1543800514515549003FFC7BE8002155BEF5EDB6DAADF4",
INIT_2B => X"FFFF7DE3F1EFA10140407000140038F450075C71FF087BD75D7FF84050BAEB84",
INIT_2C => X"24851EFEBFBD2410EBD168B7D410A175C7005B6DB55145140000FFAE85082417",
INIT_2D => X"57BC20AA5D0000000000000000000000000000000000000000000005B7DEAA08",
INIT_2E => X"A2D5574BAAAD17DFEFA2AEAAB550004175FFF7803DF45FFAE955EFAAFBD55EF5",
INIT_2F => X"5007FD75FFF7D5401EF5D2E97410AAD17DFEF007FC20AA5D043FE00F7D17FEBA",
INIT_30 => X"55007FD5545550400145FFFBEAB45F78402010007BD5545AAFFD55EFF7FBE8B5",
INIT_31 => X"155FFD17FFFFA2FBD74BA00557FF45A2D5554AAA2FBEAAAAFFD555545FF80155",
INIT_32 => X"7555F784174AAA2842ABEFFF803DEAA5D2E974AA00515754500003FF55FF8002",
INIT_33 => X"40000FFAE97410007BFFFFFA2D57FE105D04174105D042AB550055555FF007BD",
INIT_34 => X"000000007FFDEAA0004175FFA2FBC2000AAD16ABFF002A97545007FFFF455555",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000040000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(11),        -- Port A data input
DOA(0)   => data_read_a_hi_256(11),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(11),        -- Port B data input
DOB(0)   => data_read_b_hi_256(11),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_12_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50080B01BC002006940202C0DE041196A83183000000023322287E0FC000006",
INIT_01 => X"0E000C068000E04D40238000001702484000000008000008820009280A553231",
INIT_02 => X"400B71440C8001100000171C0283813013766A800586235ECC09C8423B962966",
INIT_03 => X"CC618E048306E082000081000040900003548421A080025EDF08421042DC0108",
INIT_04 => X"00028020000000812000012080080000E100001002000448100000C1BC18008C",
INIT_05 => X"0FF8060610000402010015E100004C2084800090000310000000079010007C19",
INIT_06 => X"33992D98DEC74A003EA468D01510C03E8F580C800A3F018200418927E0668645",
INIT_07 => X"0204000406050013142409121142F746222EE2498000007E111204058B84C50C",
INIT_08 => X"E826A0602902A10491165C200000820018A5104010C01086003C13E000004EDF",
INIT_09 => X"023000000000000867000000000000040000600060801022C9F88D244FA40133",
INIT_0A => X"00100000820040482B28050001600010C13499F01B334015980001E09F000000",
INIT_0B => X"B80460124F16F06BC20CBC30CBC20CBC20CBC30CBC20CBC20CBC3065E1865E10",
INIT_0C => X"00000000029D204B7C0382FD0100F3F9F80FA0200E0BF40063F99C0010000012",
INIT_0D => X"93900F6EE230301208008001007A80001100002002801000A042000000000000",
INIT_0E => X"93900F6EEC421392C96B1237E0D8BD9629F97E0B348EDAC3900F6EFA0B158EDA",
INIT_0F => X"622DBC31D73F6006A5891533EF9500EAE64BCA0B158EDAC3900F6EFA0B348EDA",
INIT_10 => X"C2B083798D341B10DEFE14400392C74CAEAD412EDD2B4FCFF812A383430C669E",
INIT_11 => X"49FAB442994B3238D4E2FB104636652E19B8BA30C022DAD8C100CA39E8CEBE66",
INIT_12 => X"30469392526208C6CC95C33717D88532966471A9C5DD00B12728D5360234D62A",
INIT_13 => X"828C4999AF580395542D27CDBA0020F0FABAC800DA550C29F36A8A2554E48A64",
INIT_14 => X"40000000873FB80B8A00EF03F56CC12B416A51B60585A5C28895962502E9F36A",
INIT_15 => X"0000000000000000000000000000008000000410802A26924010000002000EE0",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"28C1111026C152A121960A884042020000000000000000000000000000000000",
INIT_19 => X"2082082082082082082082082082092492492492492400200005A8A28A200A37",
INIT_1A => X"964B2592C964B2592C964B2592C964B2590C86432190C86432190C8208208208",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF400FEB2592C964B2592C964B2592C",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FF00042ABEFFF8400010082EAABFF55002ABEF08000000000000000000000000",
INIT_1F => X"BEFFFFBD54000004155EFAA842ABEFA280155EFFFFBC01EF0855400005555421",
INIT_20 => X"8AAAA2D540000F7D57DF55A2AABFFEF08556AA10000028AAAFFD15541000002A",
INIT_21 => X"40000005168AAA087BFFFFF5D04001FF00041554555557FE005D003FE10AAFBE",
INIT_22 => X"1555FF082AA8B55F7AEA8BEF5551575FFA2FFD75FF550015400FFFBFFF450851",
INIT_23 => X"D57DF45A280154BA5555401EFFFD5421EFA2FFFFF555D0000145082E955FF085",
INIT_24 => X"051555FF0804155FFF7842AA100000020BAAA801541055042ABEFFFFBD5410AA",
INIT_25 => X"000000000000000000000000000000000000005568AAAAAD142145FF80155EF0",
INIT_26 => X"F145B42038555F401D71C0A2DBC7EB80000280824ADBD7490E28BEF080000000",
INIT_27 => X"82FFDB5243800002FBD7EBFBD24101C00175EFB6802DBC7BE8A155EFE3FBC71F",
INIT_28 => X"E1041003DE10BEF5EDAAAAAD547038EBD57DF7DA2AEB8FC7005F6AA381C0A2DA",
INIT_29 => X"5400E3F1FFF7D085B420381C5B6AA82147FF8FEF410E001FF000E17555555B7A",
INIT_2A => X"0017D142E905EF1451525C7082AADB45F7AEA8BEF555F575FFBEF5D05EF550E1",
INIT_2B => X"02FBEFEBFBD2410AADF78F45B68010482415B471C7E3DF451EFBEFBFAF454900",
INIT_2C => X"D145145FF84155D7085B555C71404105C7F7842FA381C0A00082AA8A10410410",
INIT_2D => X"02AA8BEF000000000000000000000000000000000000000000000005B68ABAB6",
INIT_2E => X"FFAE955EFAAFBD55EF557BC20AA5D7BC01555D2EBFF55A284000AA08003FF550",
INIT_2F => X"5007BE8AAA5D2EBDE00FFFFC00AA08003FF55A2FBC00105D04175FFF7803DF45",
INIT_30 => X"FF082A97555557FE8A0000043FE00F7D17FEBAA2D5574BAAAD17DFEFA2AEAAB5",
INIT_31 => X"5FFF7D5401EF5D2E97410AAD17DFEF007FC20AA5D7BE8A005D7FEABFF002E821",
INIT_32 => X"55EFF7FBE8B550004001FF5D2A801EF5D5142145082EBFF55F7AAAABEF5D7FD7",
INIT_33 => X"82010A2AA8000008043FFFFA2FBC2010A2FBEAB45F78402010007BD5545AAFFD",
INIT_34 => X"000000007BEAAAAFFD555545FF8015555007FD5545550400145FF843DEAA552A",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000007FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(12),        -- Port A data input
DOA(0)   => data_read_a_hi_256(12),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(12),        -- Port B data input
DOB(0)   => data_read_b_hi_256(12),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_13_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10110A0441812402840402822007818000E00700000000330A3000000008042",
INIT_01 => X"A1400986B830E84D182260000C1042484001000008220008A20019080A510200",
INIT_02 => X"10A108600C9141100000C6180CA85035010E4880010431004908135980122D60",
INIT_03 => X"0013881507460886C190832175809C02030400002020124C441A108468424842",
INIT_04 => X"203080680204A0113801D600864E0C96C12000008244244052200201801802C0",
INIT_05 => X"030004849601110204950409C0208C2084E0009C0000100120A00C9918002098",
INIT_06 => X"10000882804544921681428591908000AF28A8002BC00D020003896020658FC4",
INIT_07 => X"CA20400450050009100501501102E0042020448D0000023E10408144C800D800",
INIT_08 => X"1D2B00402B220104B53100200001020218A5104016CC1C616401910801010100",
INIT_09 => X"050800404D49A42EB08000000000000406481C8C408000A2D8088D1820200B00",
INIT_0A => X"0010000002004048AA08050401604462E9144002090740148441200484000500",
INIT_0B => X"000A112100000000010000000001000000000000001000000000000000800000",
INIT_0C => X"509528954404144C200425010040000001B020081094040072005C0030864208",
INIT_0D => X"1C10B3831034081200000000000430003000206822F20CA8826AC2A14250A128",
INIT_0E => X"1C10B383110218CB0E54C2EA404A4F03D404A41AA5B7344C10B383081BA4B734",
INIT_0F => X"8001CE3E20A5B284ED1132909C72885A2B2C381BA4B7344C10B383081AA5B734",
INIT_10 => X"AC3CC0C0B8182597A801610218CB0C3548B3A008E730A01AB113A5524E6ACA67",
INIT_11 => X"A151EC5952E44128CA194517354C180A3C066430202021252991C22C99731014",
INIT_12 => X"1804C8A0ADA2E6A983014780CA28B2A5C8825194332B018A444AEA2701288A15",
INIT_13 => X"02D09852745F80112C428562EE0353635232D50048A411C158BB0A7910142C77",
INIT_14 => X"4240480068001C9B9150A0000297046E4023F8BE8E3E1E0109472C3EB50158BB",
INIT_15 => X"A1284A1284A1284A1284A1284A12851A84284110406A26924302590806000110",
INIT_16 => X"1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284",
INIT_17 => X"284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A",
INIT_18 => X"7DDFE7EFBEFFE7D3EFBEFC48A0550000000000000000000A1284A1284A1284A1",
INIT_19 => X"D75D75D75D75D75D75D75D75D75D75D75D75D75D75D7EFBFBFBBAAAAAABEFDF7",
INIT_1A => X"5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5D75D75D75",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000FEFD7EBF5FAFD7EBF5FAFD7EBF",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"AA5D043FFFFAAAABDEAA557BFDE00FFD140155F7800000000000000000000000",
INIT_1F => X"400AAD540155A2D5421FF00042ABEFFF8400010082EAABFF55002ABEF08556AA",
INIT_20 => X"ABEFA280155EFFFFBC01EF08554000055043DEBAF7843FFFFF7AABDF55A2AA97",
INIT_21 => X"D5400005568A1055043DEBAAAFFE8B45557FD7410552EAAABAAA84155EFAA842",
INIT_22 => X"FE8ABAAA8428A00087BD7555FFD56AA10000028AAAFFD15541000002ABEFFFFB",
INIT_23 => X"803FE10AAFBE8AAAA2D540000F7D57DF55A2AABFFEF085557545FFD17DEBAA2F",
INIT_24 => X"0041554555557FE005D0000155557BEAABA5D2ABDF450851420AA5D7FD5555A2",
INIT_25 => X"000000000000000000000000000000000000005168AAA087BFFFFF5D04001FF0",
INIT_26 => X"7490E28BEF08516DA82410A3FFD7AAA4B8E824971F8E38E3DF45155EB8000000",
INIT_27 => X"D7EBA4BDF45AAAA90410BEDF45155A2DF401D71C0A2DBC7EB80000280824ADBD",
INIT_28 => X"A82B680175EFB6802DBC7BE8A155EFE3FBC71FF145B42038550E38E92EB803FF",
INIT_29 => X"243800002FBD7EBFBD24101C556FA38490A3FE92BEFFEAB45417FD24385D2AAF",
INIT_2A => X"5056DE3D17FE92BEF1EFA92AA8428A10007FD557DFFDF6AA381C0A2DA82FFDB5",
INIT_2B => X"B400925D7FD557DA2803DE10BEF5EDAAAAAD547038EBD57DF7DA2AEB8FC70051",
INIT_2C => X"7FF8FEF410E001FF000E17555555B7AE10410E00155497FEFABA4120B8F55085",
INIT_2D => X"2FBD7545AA8000000000000000000000000000000000000000000005B6AA8214",
INIT_2E => X"A284000AA08003FF55002AA8BEF00517FE00082EBDF45AA8428A10085568ABAA",
INIT_2F => X"A5D2EA8A00A2803DF45AA843DF55AAAE82000F7FBD5545AAFBC01555D2EBFF55",
INIT_30 => X"55087FC00BA552ABFE10F784175FFF7803DF45FFAE955EFAAFBD55EF557BC20A",
INIT_31 => X"AAA5D2EBDE00FFFFC00AA08003FF55A2FBC00105D517FEAA082EBFE10F7FFE8B",
INIT_32 => X"DFEFA2AEAAB550051401FFA2D57FE10F7D57DE00AA842AA00007FD75FFF7FBE8",
INIT_33 => X"FDEAA08042AB45087FC0010557FD55FFAA843FE00F7D17FEBAA2D5574BAAAD17",
INIT_34 => X"000000007BE8A005D7FEABFF002E821FF082A97555557FE8A00002E82155007B",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000067FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(13),        -- Port A data input
DOA(0)   => data_read_a_hi_256(13),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(13),        -- Port B data input
DOB(0)   => data_read_b_hi_256(13),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_14_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10020A000180000284008280000281800000030000000033022000000580002",
INIT_01 => X"A14009821830284D186860000C30C24840000000084000084200090008510200",
INIT_02 => X"102100600C9001100000061020A8503401044880010400204908012018122F64",
INIT_03 => X"00008015074608840190800010008002030400002074F401209A108448404842",
INIT_04 => X"000080400004A00100004000840E000201000000024024401200020180180080",
INIT_05 => X"0A000484800111020495040800208C2084000080000010010020049818002008",
INIT_06 => X"1000088020450402B6A1420511C080008468A80008000D0200018B202067AF10",
INIT_07 => X"422000044005000910040110510260040024400C800000BE3850A144C924080E",
INIT_08 => X"000B004028020104111100200001020210A51040008004616001910801010000",
INIT_09 => X"000800004D492408208000000000000406401C0C40800022C8088DB420200900",
INIT_0A => X"0010000002004048000005040160042229140002090200000401000484000400",
INIT_0B => X"0000110100000000010000100000000000000100000000000000100000000000",
INIT_0C => X"409120940404104C2000210100400000011020080084040040005C0010820208",
INIT_0D => X"E0E0A0000190081200000000000000003000000000100C088020028102408120",
INIT_0E => X"E0E0A0000B02740421A0E5D1A024002050805210040000B0E0A0000210040000",
INIT_0F => X"E01200860008920106460D4501CB000111300210008000B0E0A0000210008000",
INIT_10 => X"0ABBC00905C33C6000400F02740412C0715C40110080A4006110510C14D18178",
INIT_11 => X"20000041DB011CC000090012565306500002411420220080220C0093C3892324",
INIT_12 => X"5809240C09024A4AE0CA00004800839682398000120800658992F3C700C30181",
INIT_13 => X"002B46867DBC002A830280000800F7B7A0B1E240240A8340000200067EAA8CB6",
INIT_14 => X"42004005800004801150A00341244000845C7DB0D0200900422ACA4B28000002",
INIT_15 => X"8120481204812048120481204812051A04204110002A26924302590802000000",
INIT_16 => X"1204812048120481204812048120481204812048120481204812048120481204",
INIT_17 => X"2048120481204812048120481204812048120481204812048120481204812048",
INIT_18 => X"69CB91FE1EF7D3ABEFBECA080050000000000000000000081204812048120481",
INIT_19 => X"F3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF7EFBBBBBF9E79E7BEAAF3",
INIT_1A => X"CFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCF3CF3CF3C",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FF007F3F9FCFE7F3F9FCFE7F3F9F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"45AAD157400007BEAAAAAAAE955555D5568A105D000000000000000000000000",
INIT_1F => X"0AAF784020AAF7D56AAAA5D043FFFFAAAABDEAA557BFDE00FFD140155F7D17DF",
INIT_20 => X"ABEFFF8400010082EAABFF55002ABEF085155400FFD1420100055574AAA2AA80",
INIT_21 => X"40155A28028B550051574005D7FFFE105D7BD7545A284020BA0055421FF00042",
INIT_22 => X"1421FF5D7FFDEBA085168B45FF843DEBAF7843FFFFF7AABDF55A2AA97400AAD5",
INIT_23 => X"04155EFAA842ABEFA280155EFFFFBC01EF08554000055002AB455D5142010085",
INIT_24 => X"57FD7410552EAAABAAA8017400AAD140000002EBFFEFA2AAA8BEFF780021FF55",
INIT_25 => X"000000000000000000000000000000000000005568A1055043DEBAAAFFE8B455",
INIT_26 => X"8E3DF45155EBD17FF6DAADB504001C71EDA82AAA0955455D556DA00490000000",
INIT_27 => X"101C55554AAAAA480082FF84000BAEBD16DA82410A3FFD7AAA4B8E824971F8E3",
INIT_28 => X"092085F401D71C0A2DBC7EB80000280824ADBD7490E28BEF085157428FFDB420",
INIT_29 => X"DF45AAAA90410BEDF45155A28E2AB7D0051504005D71F8E004975D556DB68405",
INIT_2A => X"28B6D5D51420101C5B401EF417BFAEAA08516AB45E38E38E92EB803FFD7EBA4B",
INIT_2B => X"EAFBC7EB80071FF5500175EFB6802DBC7BE8A155EFE3FBC71FF145B420385500",
INIT_2C => X"0A3FE92BEFFEAB45417FD24385D2AAFA82B68015400AADB40000082EBFFC7A2A",
INIT_2D => X"5557FE1000000000000000000000000000000000000000000000000556FA3849",
INIT_2E => X"AA8428A10085568ABAA2FBD7545AAD17DFFFAAFFC200055557DE00A280155455",
INIT_2F => X"F0051554AAFFFFC00105D55554BAA28400000F784020BAAAD17FE00082EBDF45",
INIT_30 => X"000051575FFF78415410087BC01555D2EBFF55A284000AA08003FF55002AA8BE",
INIT_31 => X"A00A2803DF45AA843DF55AAAE82000F7FBD5545AAAEAABFF0051400105D5568A",
INIT_32 => X"55EF557BC20AA5D042ABFF555142000557FC01EF007FEAABA00556AB55A2AEA8",
INIT_33 => X"C0010082EBDF55A2AABDF45A284175FF5D04175FFF7803DF45FFAE955EFAAFBD",
INIT_34 => X"00000000517FEAA082EBFE10F7FFE8B55087FC00BA552ABFE10F78415400A2FB",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000007FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(14),        -- Port A data input
DOA(0)   => data_read_a_hi_256(14),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(14),        -- Port B data input
DOB(0)   => data_read_b_hi_256(14),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_15_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000A000000000284000280000001800020030000000033022000000180002",
INIT_01 => X"A140098018300848180060000C00426040000000080000080200000000110200",
INIT_02 => X"1020004000801110000006100028503400040800010430004808000180120278",
INIT_03 => X"00008011064408840190800000228002A3000000000010000008108448000042",
INIT_04 => X"701280400004A991000000A28406000211000000220004941000000880000000",
INIT_05 => X"02000484800155020495000800218020C4002880005310000000040000000001",
INIT_06 => X"10000880004540000711224491C08000850A880008000D020001892020656300",
INIT_07 => X"8A04000016050009140501505100000420204008000000BE70408104C8000000",
INIT_08 => X"001F004028026104111002200000000200210040008004614001100801010000",
INIT_09 => X"000800000D09240000800000000000040600180840800022C8088C1020200000",
INIT_0A => X"0000000002004040000105000040042229140002080000000400000080000400",
INIT_0B => X"0000110100000000010000100001000010000000000000000000100000800008",
INIT_0C => X"0001008000000000000025000040000001300008009400006200580010000000",
INIT_0D => X"0000000002300012000000000004200030000000000008008020020000000000",
INIT_0E => X"0000000001000000400000000000000000000010108000000000000010108000",
INIT_0F => X"0000000000000200000900000000000000000010140000000000000010140000",
INIT_10 => X"0140000000000000000001000000400000000000000000000100008040000000",
INIT_11 => X"0000004000480000000000100004400000000030002000406000000000068409",
INIT_12 => X"8000000000020080080000000000802010000000000800000201000800000000",
INIT_13 => X"00000100000000000000000008000000184400A0000000000002000000441108",
INIT_14 => X"4000000000000000010620000004000000000242038B82800000000000000002",
INIT_15 => X"0000000000000000000000000000041800000110000024130202500802000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000080050000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"000804154AA5D00001EFF78428AAA007BC2145F7800000000000000000000000",
INIT_1F => X"0AA007FC2000F7D17DF45AAD157400007BEAAAAAAAE955555D5568A105D7FC00",
INIT_20 => X"FFFFAAAABDEAA557BFDE00FFD140155F7FBD74AAAAD17DF45F7D1421EF005540",
INIT_21 => X"020AAF7FFFDF45FF84000BA552ABDFEF08517DF55A2FBEAB555D556AAAA5D043",
INIT_22 => X"FEAB45F7843FF45082A801FF005155400FFD1420100055574AAA2AA800AAF784",
INIT_23 => X"D5421FF00042ABEFFF8400010082EAABFF55002ABEF087BE8ABA555168B55AAF",
INIT_24 => X"D7BD7545A284020BA007FFFE10A284000AA0055401550055574005D2E800AAA2",
INIT_25 => X"000000000000000000000000000000000000000028B550051574005D7FFFE105",
INIT_26 => X"55D556DA004971C7038140012482550E021C7EB8028A821C7BC516DFF8000000",
INIT_27 => X"45E3DF471C70851400BA0071C5028FFD17FF6DAADB504001C71EDA82AAA09554",
INIT_28 => X"B555D516DA82410A3FFD7AAA4B8E824971F8E38E3DF45155EBF1D5492BED17FF",
INIT_29 => X"54AAAAA480082FF84000BAEBF1FFF7DEB8000092552ABFFEF08517DF6DB6FBE8",
INIT_2A => X"EFA8241516DB55A2FFEAB6DEB843DF551C20801C71C5157428FFDB420101C555",
INIT_2B => X"550428412A85082BEDF401D71C0A2DBC7EB80000280824ADBD7490E28BEF087F",
INIT_2C => X"51504005D71F8E004975D556DB68405092087FF8E00BE8A02082005F47145085",
INIT_2D => X"57BD75EFF78000000000000000000000000000000000000000000000E2AB7D00",
INIT_2E => X"55557DE00A2801554555557FE100055554BA5504000105D2A80145AA842AA005",
INIT_2F => X"5AAD557410F7D57DF55AAFBD55450055420BA0055574BAF7D17DFFFAAFFC2000",
INIT_30 => X"FF08517FFFFF7FBEAB455D517FE00082EBDF45AA8428A10085568ABAA2FBD754",
INIT_31 => X"4AAFFFFC00105D55554BAA28400000F784020BAAAD57FFEFA28402010552ABDF",
INIT_32 => X"FF55002AA8BEF007FFDE1000557DF45AAFBE8BEFA2803FF45550400155555155",
INIT_33 => X"80000087BD55450855400BA002A95400F7FBC01555D2EBFF55A284000AA08003",
INIT_34 => X"000000002EAABFF0051400105D5568A000051575FFF78415410087FEAA10F7AE",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000060000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(15),        -- Port A data input
DOA(0)   => data_read_a_hi_256(15),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(15),        -- Port B data input
DOB(0)   => data_read_b_hi_256(15),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_16_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"DA22C618B1000482B688B186588884862A400438255FC38381441205BA803003",
INIT_01 => X"264AC80028404C211203A952A90341080B173340412000E1005D628000820484",
INIT_02 => X"400034C206C405000001A48202084004003008255040826EE008B440200E2042",
INIT_03 => X"2916704900606AC82B49CC56DF8CC1E50E4800202115005760010010000C0400",
INIT_04 => X"052DCA856DC7504B82BF6614C86D2B7F85AAD17F4B100000B88148C4804A428A",
INIT_05 => X"373CB02A00C0502F301180141A42A5720E0F43C17A8479580001AC20000000E2",
INIT_06 => X"303E2094282B85242C85001038D5710E8410D5959BC4800015001219D0550077",
INIT_07 => X"880100000159954501280B0080146F7112D949A0015018220540000382805001",
INIT_08 => X"30015452880C8D90409A05B2CB2CA400200209E5601044A24000000462A60018",
INIT_09 => X"452D54000C0907000330000000000096480050000685400005FC014743E0DC92",
INIT_0A => X"00014808A02004200E540480212000A448C0080024AEA00C9688000000000005",
INIT_0B => X"000D58460018F6D3D84400044000440004400044000440004400042000220002",
INIT_0C => X"0001004010A8812831605DA0000A054052E40000817680220040025699200002",
INIT_0D => X"AAADA0C343F1AC1B01040A002024895514554485D00000012400240000000000",
INIT_0E => X"AAADA0CC421CA003B694B68018FAAA708E2CB5320018CAC99BA0A3B9320018CA",
INIT_0F => X"B1443A1891E4A928C29020E6A8524CE7A3EE59320018CAC99BA0ACB9320018CA",
INIT_10 => X"04B2A5A40B1E6644AF0F021EA003AC24352AB2449A3FF2FA04E5E09B128834AD",
INIT_11 => X"60ED838E890B703C6260D8E3A21275714C902375B801324301AB0067622E5E54",
INIT_12 => X"064F70DBDB1C74424E91E1C194C71D1216F50A8C241815FEB6A9158863F638FB",
INIT_13 => X"45FDF9D364DBD9435A6D45C9E81BED555E4C15F11133D171727A2550EE2F1BA0",
INIT_14 => X"08150013F162119014204373517700ACCC59432A2B2D001F803471A9A960E572",
INIT_15 => X"000000000000000000000000000000880002054000229088542210206B2AB015",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"2A898D21B4C98389ED146C080000000000000000000000000000000000000000",
INIT_19 => X"A29A29A29A29A29A29A29A29A29A28A28A28A28A28A53CBF0F0D3CF3CF0AB1A2",
INIT_1A => X"8F47A3D1E8F4FA7D3E9F4FA7D3E9F4FA7D3E8F4FA3D3E8F4FA3D3E9A29A29A29",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000FA7D3E9F4FA7D1E8F47A3D1E",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFF7FBE8B45AAD568BFFFFAA975FF00003FE0055000000000000000000000000",
INIT_1F => X"0005D2A95410FFFFC00000804154AA5D00001EFF78428AAA007BC2145F7843FF",
INIT_20 => X"7400007BEAAAAAAAE955555D5568A105D2E974BAF7FBEAB45FFFFC00BAF78002",
INIT_21 => X"C2000F78000010552E800AA002E821FFA2AAAAA00000417555FFD17DF45AAD15",
INIT_22 => X"43FEBA5D55575FFF7AABFE00557BD74AAAAD17DF45F7D1421EF0055400AA007F",
INIT_23 => X"D56AAAA5D043FFFFAAAABDEAA557BFDE00FFD140155F7AABDF55F7AE820AA080",
INIT_24 => X"8517DF55A2FBEAB555D04154BAA2FBE8B55FFFFD55FF557FC2000FF8015410FF",
INIT_25 => X"000000000000000000000000000000000000007FFDF45FF84000BA552ABDFEF0",
INIT_26 => X"21C7BC516DFF8438FC7E3F1EAB55B6DF6DBFFF7AA955C71C043FE10490000000",
INIT_27 => X"55FFF1C70BAF78A000005D2097438FFF1C7038140012482550E021C7EB8028A8",
INIT_28 => X"57DEBD17FF6DAADB504001C71EDA82AAA0955455D556DA00492490492F7FBE8B",
INIT_29 => X"71C70851400BA0071C5028FF84020285D2085092002A801FFB6AAA8A10080E17",
INIT_2A => X"BAF6DE3AA8709208043FEBA555B555FFE3AABFE005D71D5492BED17FF45E3DF4",
INIT_2B => X"BC0028E38412428EBD16DA82410A3FFD7AAA4B8E824971F8E38E3DF45155EBA4",
INIT_2C => X"8000092552ABFFEF08517DF6DB6FBE8B555D04124BAB6FBE8B45E3FBD55D7557",
INIT_2D => X"5003DE000000000000000000000000000000000000000000000000071FFF7DEB",
INIT_2E => X"5D2A80145AA842AA00557BD75EFF78428B55AAD168B55F7FFFDFEFFFAA955555",
INIT_2F => X"0000000010F7FBEAB45FFD1554AAFFAE820105500154AAF7D5554BA550400010",
INIT_30 => X"EFF7AEA8A10002E955FFA2D17DFFFAAFFC200055557DE00A2801554555557FE1",
INIT_31 => X"410F7D57DF55AAFBD55450055420BA0055574BAF784000BA5D0017410082E801",
INIT_32 => X"8ABAA2FBD7545AA802ABEFA2AA9541000003DEBA557BD75EFA2AEBDE105D5557",
INIT_33 => X"EAB45AAFFD55555D7FC20AAA280000AAAAD17FE00082EBDF45AA8428A1008556",
INIT_34 => X"00000000557FFEFA28402010552ABDFFF08517FFFFF7FBEAB455D04020AAFFFB",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000020000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(16),        -- Port A data input
DOA(0)   => data_read_a_hi_256(16),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(16),        -- Port B data input
DOB(0)   => data_read_b_hi_256(16),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_17_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"5284CE4FB7BD2C8994A13392DBD02E14006B82AC7E800D44D3DD2FD5F9B961C0",
INIT_01 => X"F9BA301F7E03FC6793F2199B39FC233C11D93AE6F3BB92B32091DBC339B24542",
INIT_02 => X"1D5FC0C08F040404446965C0607FB8A217C400C33A908078551BD04222186338",
INIT_03 => X"A14124C28DFD960832C90446DF8400A5055C25295B695FF97E1B5AC757F06D6B",
INIT_04 => X"04A106866DA3D02A01FB660C08A4AB7F840EDB6F48100DFC8081081D78AC7402",
INIT_05 => X"51E072F0C0C58D9C125EBFC00A46CF0388054100F680E0CE0107B8D040DAFCDA",
INIT_06 => X"019A4D00786B048112C58B16307F15DE8408B233661C10BBA5DAAFA9DDA1194D",
INIT_07 => X"8E00001660700CE170284A00891C7C03D29DE26814515835902AC089A2801540",
INIT_08 => X"C009F3A1B0120A1C51DFF881861CBE0305A12A0321810217C01D34EDC98FFA1C",
INIT_09 => X"747E6610052CDEE97FF1F9F63E3EF790380078002CE976AB6BF769769E4D437D",
INIT_0A => X"00185C44B91BC1740B7605040BE0018CFC7429F326B9D045FF8000E9AB415606",
INIT_0B => X"3A28FC1AAF5CF6F3D3EF3D3EF3D3EF3D3EF3D3EF3D3EF3D3EF3D3EF9E9F79E9E",
INIT_0C => X"0000020012E9E10A31EB5FF9296A67F5B4FFBD2FAD7FE653C3FBFF33E10C001B",
INIT_0D => X"333EA16031F2BD47BDA2CA5D8164FCCFE833C5C3D00018006C68170000000000",
INIT_0E => X"333EA160391BEFF2C32FB695F919110D5ECE542A6FEEB2533EA160782A6FEEB2",
INIT_0F => X"D18C0D06638A207CFDE1F7DDAD76D5282400F82A6FEEB2533EA160782A6FEEB2",
INIT_10 => X"E6E43E59AFE4A59B57679D19EFF2C7573FAD5A86840354D1706FFFA3EF6E24B6",
INIT_11 => X"F7D7A0ABD6DAAAB96529382B74E4E1FE4ACA4D77FAAB77CE3AF3EE78F58DB737",
INIT_12 => X"2D1281017F056E9C9C3FC95949C157ADB55572CA52606DFED6CA55334C04C04F",
INIT_13 => X"59FDEB974F486905001FDF5FA0D719F9956EAA1A184045D5D7A870D2F5A5D752",
INIT_14 => X"60158015177F916A039EF41FDB34A91F432EA58949D5B5C85F97871876F7D7E8",
INIT_15 => X"000000000000000000000000000004DC200005E705B7B3D9FC22F00BE419FB55",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"06013DB9880A5D22E229F3030018000000000000000000000000000000000000",
INIT_19 => X"D35D74D35D74D34D35D74D35D74D34D34D34D34D34D0D30D0D303AEBAE886E40",
INIT_1A => X"51A8D46A351A0D068341A0D068341A0D068341A8D468341A8D46834D35D74D34",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000008D46A351A8D46A351A8D46A3",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFF7FBFDF55A28402000F7D56ABFF55000000000000000000000000",
INIT_1F => X"A00F7843FEBA55043FFFFF7FBE8B45AAD568BFFFFAA975FF00003FE0055043FF",
INIT_20 => X"54AA5D00001EFF78428AAA007BC2145F7D568B45000002010552EBDF45A28028",
INIT_21 => X"95410FFAE800105D2A95410002A95410AAAEBFF55AAFFC00BAF7FFC000008041",
INIT_22 => X"57DE00F7AE800AAAAAABDFEF5D2E974BAF7FBEAB45FFFFC00BAF780020005D2A",
INIT_23 => X"517DF45AAD157400007BEAAAAAAAE955555D5568A105D7FFFFEFA2D568BFFFFD",
INIT_24 => X"2AAAAA00000417555FF8028B55082A974105D003FF55F7802AAAAAAD168AAA5D",
INIT_25 => X"000000000000000000000000000000000000000000010552E800AA002E821FFA",
INIT_26 => X"71C043FE10490A3FFFFFFFFFDFEFE3F5FAF45AA8000038F7DB6FBD7490000000",
INIT_27 => X"384124BFF7DB68A28A38F7803DE82490438FC7E3F1EAB55B6DF6DBFFF7AA955C",
INIT_28 => X"0BAFFF1C7038140012482550E021C7EB8028A821C7BC516DFFDF68B551C0E050",
INIT_29 => X"70BAF78A000005D2097438FFAA85000492495428082E95400AAA0BDF7DB6F5C7",
INIT_2A => X"FAFFFB6D56FBFFEBDB78E38F7AA800BAB6AEBDFD75D2490492F7FBE8B55FFF1C",
INIT_2B => X"028AAAB6D16FA8249517FF6DAADB504001C71EDA82AAA0955455D556DA00497F",
INIT_2C => X"2085092002A801FFB6AAA8A10080E1757DEB8A2DB5514249243841003FF6DEB8",
INIT_2D => X"7FFFDF550000000000000000000000000000000000000000000000004020285D",
INIT_2E => X"F7FFFDFEFFFAA9555555003DE00002ABFFEFF7FBFDFFFAAD168B55AA80000BAF",
INIT_2F => X"FF7FBEAB45552E954BA08003DFFFFFAAA8AAAF7843FE10000428B55AAD168B55",
INIT_30 => X"10AA843FFFFF7D5554BAF7D5554BA5504000105D2A80145AA842AA00557BD75E",
INIT_31 => X"010F7FBEAB45FFD1554AAFFAE820105500154AAF7AE974000800154AA002E954",
INIT_32 => X"554555557FE10007FEABEFFFD57FFEFAAFFE8ABAFFAA820BAF7AEBFF55550000",
INIT_33 => X"020AA08003DFFFA28028AAAF7D17DE0000517DFFFAAFFC200055557DE00A2801",
INIT_34 => X"0000000004000BA5D0017410082E801EFF7AEA8A10002E955FFA2AABFF455500",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000067FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(17),        -- Port A data input
DOA(0)   => data_read_a_hi_256(17),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(17),        -- Port B data input
DOB(0)   => data_read_b_hi_256(17),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_18_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"69844019080000A21A611406840014122A641074155FC28A2024001001801003",
INIT_01 => X"01067920034004180005E9E3C90360C0041C0181002001602025800008440084",
INIT_02 => X"40AC3CAA22D605200000856E2481902400344A20F802C22054001000021E2379",
INIT_03 => X"A95308ECD3207AC81D91C4002004C08A06008080BA868007E58040102B0E0100",
INIT_04 => X"044CC183800CA00780808004C8DB841405A80A100B586200FAC24AE4805242CA",
INIT_05 => X"771C10000000000B1135883C08A115320E0401C0200038394230070A19000020",
INIT_06 => X"3001499C602A8A003E800A042D8132A00098408F79E3901218050018024110D6",
INIT_07 => X"5029401000C983E60004010030400353C05806800104004E0000042E52800E20",
INIT_08 => X"0000117088080990419005B0C309402030060860E01004A828408800440405E3",
INIT_09 => X"6B8186185C42900693A002004040001E1950850C848601008708114A2030B480",
INIT_0A => X"100180A8062026000DC425C0301311324AA237108857220BA089420440000030",
INIT_0B => X"C44703657083080C2800C2000C2000C2000C2000C2000C2000C2000610006100",
INIT_0C => X"C1B0609C05013065CC042004040808084001E000108010230400800FD9B286C4",
INIT_0D => X"CCC15F9CBA45505640000A402019003F140FC2060014250B9080008306C18360",
INIT_0E => X"CCC15F9FB1962FCB69E08AAAEAEBCDDF7C728582081483ACC15F9C3982081483",
INIT_0F => X"EBF1CFFF7670ACC3811A28AB57523CDFEBFBF982081483ACC15F9F3982081483",
INIT_10 => X"C9002BF05800D875E63CC9962FCB52CAA02FE3F8E7F5E3AC3620805298B15A3F",
INIT_11 => X"F1B72A8A800B7546DB9F1CA320037F01BD67DC4041D4CF03138DD865103EFEEA",
INIT_12 => X"81CCFAFDBF9464006FD037AEFAE5150016EA8DB7BFE25208E8F46A228BF8A757",
INIT_13 => X"641256EC844B8AF92FD7CEDC24A9E181A8A29509EAAE7FD3B749471C48F8A459",
INIT_14 => X"0297D086E00036D2440E0880AAD62BEFF5778802A3AF8E8FB0440CE78773B709",
INIT_15 => X"8360D8360D8360D8360D8360D83609220D20D00000080C0601400B402307E480",
INIT_16 => X"360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D",
INIT_17 => X"60D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8",
INIT_18 => X"D9D701DC2E784601EFBE2C00000000000000000000000008360D8360D8360D83",
INIT_19 => X"5155555545145145155555545145145145145145145220B22A0B820820965177",
INIT_1A => X"44A25128944A25128944A25128944A25128944AA552A954A2512895554514514",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000025128944A25128944A251289",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFEFF7AE954BA5D04174AA00000000000000000000000000",
INIT_1F => X"145AA801741000043FFFFFFFFFFFFFF7FBFDF55A28402000F7D56ABFF55043FF",
INIT_20 => X"8B45AAD568BFFFFAA975FF00003FE0055043FFFFFFFFFDFEFA2D56AB45AA8400",
INIT_21 => X"3FEBA55557FFEFA2D168B55AAFBFFFFFFF80021EF0855421EF00043FFFFF7FBE",
INIT_22 => X"A82155F7AEBFEBAFFD56AA00A2D568B45000002010552EBDF45A28028A00F784",
INIT_23 => X"FFC00000804154AA5D00001EFF78428AAA007BC2145F7D5400000004020AA5D2",
INIT_24 => X"AAEBFF55AAFFC00BAF7AE80010082E954BA0004174AAAA8428B45082ABFEBAA2",
INIT_25 => X"000000000000000000000000000000000000002E800105D2A95410002A95410A",
INIT_26 => X"8F7DB6FBD7490E3FFFFFFFFFFFFFFFFBFDFEFFFAE954AA550415492140000000",
INIT_27 => X"D7AAD16FB6DBE8E00155BE8015410140A3FFFFFFFFFDFEFE3F5FAF45AA800003",
INIT_28 => X"1C7140438FC7E3F1EAB55B6DF6DBFFF7AA955C71C043FE1049043FFEFE3F1F8F",
INIT_29 => X"FF7DB68A28A38F7803DE82495B78FC7AAD56FB6DBEF1FAFD7E384001EF145B47",
INIT_2A => X"420381C0A02082492A85155E3A4BDE92FFD56FA28B6DF68B551C0E050384124B",
INIT_2B => X"E28B7D1420BDEAAA2F1C7038140012482550E021C7EB8028A821C7BC516DFFD1",
INIT_2C => X"2495428082E95400AAA0BDF7DB6F5C70BAFFAE870280024904BA1400174AABE8",
INIT_2D => X"50415410550000000000000000000000000000000000000000000002A8500049",
INIT_2E => X"AAD168B55AA80000BAF7FFFDF55002ABFFFFFFFFFFFEFF7FBFDFFFF7AA974BA5",
INIT_2F => X"000043DFEFA2D56AB45AAD57DFEFF7AA82155F78015400552ABFFEFF7FBFDFFF",
INIT_30 => X"55A280021EF557FD7555550428B55AAD168B55F7FFFDFEFFFAA9555555003DE0",
INIT_31 => X"B45552E954BA08003DFFFFFAAA8AAAF7843FE10007FEAB55A2D17FFEFFFD568B",
INIT_32 => X"AA00557BD75EFF7D1400AA5D2A82000002A95545A2843FE00F7D17FEAAF7FBEA",
INIT_33 => X"020AA5D04154BAF7AEA8BEF55003DEAAA2D5554BA5504000105D2A80145AA842",
INIT_34 => X"000000002E974000800154AA002E95410AA843FFFFF7D5554BAF7AE974BA0004",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000020000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(18),        -- Port A data input
DOA(0)   => data_read_a_hi_256(18),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(18),        -- Port B data input
DOB(0)   => data_read_b_hi_256(18),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_19_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"042200000000000041088001001AA00000000000000000000000500802000003",
INIT_01 => X"074018000024000000000404000000000A22000800000800004A200000000001",
INIT_02 => X"0000048002C405000000000006A84000000000200893C246A20000000020031A",
INIT_03 => X"020A9639044012C80001C4000004C08006000000001025000000000000000000",
INIT_04 => X"0400C0800000000380800004C8000000058800000B1000009880480480024200",
INIT_05 => X"420410000000000B10804004080001320E0401C0200038080000000000000000",
INIT_06 => X"2002409006F00A8428050A000280493104004500480090080A01120220140020",
INIT_07 => X"0000000000418026090240923240002190400000000000C0054A912054004021",
INIT_08 => X"0000115080000990000000B0C308000000000860200160000000000038380000",
INIT_09 => X"8000F80001012590001000000000001618000000020280008180810200000000",
INIT_0A => X"0000000000000000000000000000000100008000110000000000000000000017",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000840007600000000000000000800259000000",
INIT_0D => X"0008A0034078104B41A41000000000031400C002000000000000000000000000",
INIT_0E => X"0008A0004263C0343EDD414004042228DC0D385598035D0008A003B05598035D",
INIT_0F => X"040231068187C39F5A4F985C008902041124505598035D0008A000B05598035D",
INIT_10 => X"1BFBD406451B02000E033263C0343CB740500401180DE053A98F6ECC739D8140",
INIT_11 => X"420851546B2400000040D8549B5800000010227848D4303807FC8CC5508AEAED",
INIT_12 => X"52210402120A936B0000000004C2A8D6480000000018A700FCF980CC300318A2",
INIT_13 => X"B1427ED430B41402D025082359700181C21140E40511802208D6B30C48F8A8A4",
INIT_14 => X"9C000018440021011821B35254E99AF9E9410006362A2B6424287B08286208D6",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000023006000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"7747E18E0218CC18E88324000000000000000000000000000000000000000000",
INIT_19 => X"34C30C30C30C30D34C30C30C30C30C30C30C30C30C3504118982A69A6980E411",
INIT_1A => X"C26130984C26130984C26130984C261309A4D26130984C26130984C30C30C30D",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000130984C26130984C26130984",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAA954BA5500020BA5D000000000000000000000000",
INIT_1F => X"4BA5D517FFFF08043FFFFFFFFFFFFFFFFFFFFEFF7AE954BA5D04174AA007BFFF",
INIT_20 => X"FFFFF7FBFDF55A28402000F7D56ABFF557BFFFFFFFFFFFFFFFFFBFDFEFFFAA97",
INIT_21 => X"17410007BFFFFFFFFFFFFEFF7D16AB45AA8002000F7D5575455D043FFFFFFFFF",
INIT_22 => X"568B55F7AE955FFAA840201008043FFFFFFFFFDFEFA2D56AB45AA8400145AA80",
INIT_23 => X"043FFFFF7FBE8B45AAD568BFFFFAA975FF00003FE00557BFFFFFFFFBFDF45AAD",
INIT_24 => X"F80021EF0855421EF002ABFFEFF7D168B55AAD17FFEFF7AE975FF00557FFFF5D",
INIT_25 => X"00000000000000000000000000000000000000557FFEFA2D168B55AAFBFFFFFF",
INIT_26 => X"A5504154921471FFFFFFFFFFFFFFFFFFFFFFFF7AA954BA550000082550000000",
INIT_27 => X"EFF7FBFAFD7E3A4954BA555B7AFC7080E3FFFFFFFFFFFFFFFFBFDFEFFFAE954A",
INIT_28 => X"545550A3FFFFFFFFFDFEFE3F5FAF45AA8000038F7DB6FBD74975FFFFFFFFFFFF",
INIT_29 => X"FB6DBE8E00155BE8015410147FFFFFFF7FBF8FC7EBD568B55A28000000FFDF52",
INIT_2A => X"FDFC7E3F1FAF55A2DB6FB7DF7AE955C7BE800000008043FFEFE3F1F8FD7AAD16",
INIT_2B => X"0955FF145B7AFC7410438FC7E3F1EAB55B6DF6DBFFF7AA955C71C043FE10497B",
INIT_2C => X"D56FB6DBEF1FAFD7E384001EF145B471C71424B8FC7E3D56AB6DB6DF7AFC7EBA",
INIT_2D => X"50002000550000000000000000000000000000000000000000000005B78FC7AA",
INIT_2E => X"F7FBFDFFFF7AA974BA55041541055517FFFFFFFFFFFFFFFFFFFFEFF7AA974AA5",
INIT_2F => X"500517FFFFFFFBFDFEFFFFFEAB45AA80154AA557BEAB45002ABFFFFFFFFFFFEF",
INIT_30 => X"55A28002000F7FFC2155552ABFFEFF7FBFDFFFAAD168B55AA80000BAF7FFFDF5",
INIT_31 => X"FEFA2D56AB45AAD57DFEFF7AA82155F78015400557BFDFEFF7FBEAB55A2D56AB",
INIT_32 => X"555555003DE00007FFDF45AAD568B45AAFBFFFFFFFAA95545F7840201000043D",
INIT_33 => X"6ABFFFFFBEAB45A280155EF557FE8B55000428B55AAD168B55F7FFFDFEFFFAA9",
INIT_34 => X"000000007FEAB55A2D17FFEFFFD568B55A280021EF557FD755555042AB55AAD1",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000040000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(19),        -- Port A data input
DOA(0)   => data_read_a_hi_256(19),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(19),        -- Port B data input
DOB(0)   => data_read_b_hi_256(19),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_20_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000003",
INIT_01 => X"A65FF80000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000048002CC070000000000000000000000002FF86100200000000220002362",
INIT_03 => X"00000000000203D80025DC18004DC3D01E000000000000000000000000000000",
INIT_04 => X"07E5DF808071026F87C4191DD8005080679800000F300002998058068002C000",
INIT_05 => X"C205F23A2100557F70000004390021F61E1E87C3FD0CFBF80880072042000044",
INIT_06 => X"1209244C2000100006800000020010000008407FC800B0000000100600040000",
INIT_07 => X"8802000009FFBFE51886018002040020000800000554003E0000000002800000",
INIT_08 => X"30801F5780259FB0000000F7DF78020004011FEFE00000000020031502000083",
INIT_09 => X"00000000001000000000000000000056F8000001000000040000040141800802",
INIT_0A => X"0000000000000008000800000000000000000000000000000010010014800000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"00010240001721214E000004000000080000008000001000040080FFDB000000",
INIT_0D => X"0000000F3008001E00000000001803FF14FFC006000000008010200000000000",
INIT_0E => X"0000000F3040200000020000000026A70C0008020000200000000F3002000020",
INIT_0F => X"000030B86000400080000200000000004A58F0020000200000000F3002000020",
INIT_10 => X"0000000002183E61E6000040200001000000000019B140000800800000020000",
INIT_11 => X"C00010080000000000525801000000000014AC08000000508001030A0A400100",
INIT_12 => X"000002BC360020000000000292C0100000000000A56000090100000000001F86",
INIT_13 => X"8010000000000000574500001001060600000000001716800000803102020000",
INIT_14 => X"00000000000040040040002000080506049CDF70C08040100000706707600000",
INIT_15 => X"00000000000000000000000000802040200200604040000000000024FB7FE008",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"060070400020112240209A408004000000000000000000000000000000000000",
INIT_19 => X"65965965965965965965965965965861861861861860D30424343CF3CF340E00",
INIT_1A => X"90C86432190C86432190C86432190C86432190C86432190C8643219659659659",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000086432190C86432190C864321",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974AA55040201008000000000000000000000000",
INIT_1F => X"4AA550002000007BFFFFFFFFFFFFFFFFFFFFFFFFFAA954BA5500020BA5D7FFFF",
INIT_20 => X"FFFFFFFFFFFEFF7AE954BA5D04174AA00003FFFFFFFFFFFFFFFFFFFFFFF7AA97",
INIT_21 => X"7FFFF087FFFFFFFFFFFFFFFFFFFFDFEFFFAE974AA5D003FE005D043FFFFFFFFF",
INIT_22 => X"BFDFFFAA84000105D556AB55557BFFFFFFFFFFFFFFFFFBFDFEFFFAA974BA5D51",
INIT_23 => X"043FFFFFFFFFFFFFF7FBFDF55A28402000F7D56ABFF55003FFFFFFFFFFFFFF7F",
INIT_24 => X"A8002000F7D5575455D2EBFFFFFFFFFFFEFF7FBEAB55A28000010F7D16ABEF08",
INIT_25 => X"000000000000000000000000000000000000007BFFFFFFFFFFFFEFF7D16AB45A",
INIT_26 => X"A550000082557FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550400028000000000",
INIT_27 => X"FFFFFFFDFEFF7AE974BA5500050380071FFFFFFFFFFFFFFFFFFFFFFFF7AA954B",
INIT_28 => X"E285D0E3FFFFFFFFFFFFFFFFBFDFEFFFAE954AA55041549214043FFFFFFFFFFF",
INIT_29 => X"AFD7E3A4954BA555B7AFC70871FFFFFFFFFFFFFFF7FBFDFFFFFAA974BA550038",
INIT_2A => X"3FFFFFFFFFDFEFF7F1FAFC7A28002028555F6FB7D5D75FFFFFFFFFFFFEFF7FBF",
INIT_2B => X"402010FFDB6ABEF140A3FFFFFFFFFDFEFE3F5FAF45AA8000038F7DB6FBD7490E",
INIT_2C => X"FBF8FC7EBD568B55A28000000FFDF525455524BFFFFFFFBFDFC7E3F5E8B45A28",
INIT_2D => X"504000BA080000000000000000000000000000000000000000000007FFFFFFF7",
INIT_2E => X"FFFFFFFEFF7AA974AA550002000557FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5",
INIT_2F => X"055043FFFFFFFFFFFFFF7FBFDFEFFFAE954BA5500174AA08517FFFFFFFFFFFFF",
INIT_30 => X"EFF7AE974AA550028AAA5D2ABFFFFFFFFFFFEFF7FBFDFFFF7AA974BA55041541",
INIT_31 => X"FFFFFFBFDFEFFFFFEAB45AA80154AA557BEAB4500557FFFFFFFFFDFEFF7FFFFF",
INIT_32 => X"00BAF7FFFDF55002EBFFFFF7FBFDFEFFFD568B55A284020BA557FFFFFF5D517F",
INIT_33 => X"FFF55A2D16AB45AA8402000F7FBEABEF5D2ABFFEFF7FBFDFFFAAD168B55AA800",
INIT_34 => X"000000007BFDFEFF7FBEAB55A2D56AB55A28002000F7FFC215555043DFEFF7FB",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000007FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(20),        -- Port A data input
DOA(0)   => data_read_a_hi_256(20),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(20),        -- Port B data input
DOB(0)   => data_read_b_hi_256(20),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_21_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"4A302428B824900A128C090A5C1800261500213C005FE812D10420054085A202",
INIT_01 => X"081FFE3440B609703B0427F801A40B8115BC4F655300340288A40D30040E4DD8",
INIT_02 => X"04CA478082CC1740002019824E0203100640303FF8C0B31061096E21A1840814",
INIT_03 => X"230CA7A4810083F80095DE00102DC3823EA821094EC68248923200013290C800",
INIT_04 => X"07CFFFC04904AA7F8780409DF84A0202879800000F3000029980780EA2C3C002",
INIT_05 => X"DE87F0280000407FF900D914382091FE1E1C0FC3E01EFFF8000480200008D062",
INIT_06 => X"010E2182002BC107A03448808F0D7C002822987FC830F40134CC74D002016612",
INIT_07 => X"0401000011FBFFE00520000200422033025C4209104500000012004C004D8C0B",
INIT_08 => X"00EF1F5FA0041FF080AC70FFDF78220010841EFFE7116E144071268DFD3E4C24",
INIT_09 => X"FC8BFE18008083B4443151462A28C6DFF80010002605302248088950484550A3",
INIT_0A => X"10018C241102068006C620C03882019480E631A0855E924E2598038938404037",
INIT_0B => X"A641165448C80C103648A3648A3648A3648A3648A3648A3648A366451B2451B2",
INIT_0C => X"011100841200D001000624000100C002804A08221890004806A310FFDF000454",
INIT_0D => X"5004D8158809C86065941840B1014FFF56FFC0281280080180B2948004400220",
INIT_0E => X"5004D815810D42E04A08A80098C02450025360694101816002D41A4068C10181",
INIT_0F => X"134160C8125B0B271802242880A04482418A0068C101816002D41A4069410181",
INIT_10 => X"10080E05C0B06AA8B12CFD0D42E0441A300012682960828F05C96A001B029010",
INIT_11 => X"00010362A8A20826A88660D86B202049F115100920C54E8EA256ECF078BA081C",
INIT_12 => X"064802C0081B0D64040936443306C55144104F30A8801406D002900062803201",
INIT_13 => X"4581BA0038005A706680012280506A8010602011819E290048A2118EC8140C08",
INIT_14 => X"CC158092C044600466208CC5091011C322A4C40A0300600C0A80509F41800880",
INIT_15 => X"80200802008020080200802008020412002001000000381C02004000FBFFF80D",
INIT_16 => X"0200802008020080200802008020080200802008020080200802008020080200",
INIT_17 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_18 => X"FDDFEFFFBEFFE7C7BFBEFC000000000000000000000000080200802008020080",
INIT_19 => X"F7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7FFBFBFFF9E79E7FFFDF3",
INIT_1A => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFDFEFF7FBFDFEFF7FBFDF7DF7DF7D",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00001FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D000200008000000000000000000000000",
INIT_1F => X"4AA5D00020AA5D7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550402010087FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAA954BA5500020BA5D7FFFFFFFFFFFFFFFFFFFFFFFFFFAE95",
INIT_21 => X"0200000003FFFFFFFFFFFFFFFFFFFFFFF7AA974BA5D0402000557BFFFFFFFFFF",
INIT_22 => X"FFFFEFF7AE974BA5D00174BA00003FFFFFFFFFFFFFFFFFFFFFFF7AA974AA5500",
INIT_23 => X"043FFFFFFFFFFFFFFFFFFFFEFF7AE954BA5D04174AA00003FFFFFFFFFFFFFFFF",
INIT_24 => X"FAE974AA5D003FE005D2EBFFFFFFFFFFFFFFFFFFDFEFF7AE954AA5500174BA5D",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFDFEFF",
INIT_26 => X"A550400028007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0000010000000000",
INIT_27 => X"FFFFFFFFFFFFFAA954BA5D00000BA557FFFFFFFFFFFFFFFFFFFFFFFFFFAE974A",
INIT_28 => X"0005571FFFFFFFFFFFFFFFFFFFFFFFF7AA954BA550000082557BFFFFFFFFFFFF",
INIT_29 => X"DFEFF7AE974BA55000503800003FFFFFFFFFFFFFFFFFFFFEFF7AA974AA5D0405",
INIT_2A => X"3FFFFFFFFFFFFFFFFFFDFEFF7AE954BA5D00154AA00043FFFFFFFFFFFFFFFFFF",
INIT_2B => X"A974BA5D00104925D0E3FFFFFFFFFFFFFFFFBFDFEFFFAE954AA550415492140E",
INIT_2C => X"FFFFFFFF7FBFDFFFFFAA974BA550038E285D2ABFFFFFFFFFFFFFFFFBFDFEFFFA",
INIT_2D => X"D00000100000000000000000000000000000000000000000000000071FFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE954AA5504000BA087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0557BFFFFFFFFFFFFFFFFFFFFFFFF7AA954BA5D00000BA5D7FFFFFFFFFFFFFFF",
INIT_30 => X"EFF7AE954AA5D041740055517FFFFFFFFFFFFFFFFFFFFEFF7AA974AA55000200",
INIT_31 => X"FFFFFFFFFFFFF7FBFDFEFFFAE954BA5500174AA08043FFFFFFFFFFFFFFFFBFDF",
INIT_32 => X"74BA550415410552ABFFFFFFFFFFFFFF7FBFDFFFFFAA974AA5D00174BA08043F",
INIT_33 => X"FDFEFF7FBFFFFFF7AE954BA5D0000010552ABFFFFFFFFFFFEFF7FBFDFFFF7AA9",
INIT_34 => X"00000000557FFFFFFFFFDFEFF7FFFFFEFF7AE974AA550028AAA5D2EBFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(21),        -- Port A data input
DOA(0)   => data_read_a_hi_256(21),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(21),        -- Port B data input
DOB(0)   => data_read_b_hi_256(21),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_22_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"5290F4CDE914905A14A43D33F488243E17122300F55FEB189B343A1140548380",
INIT_01 => X"A94007B259F6A975386262000C344BA9573C6FF57B18A5FB0ABFCD3C2C5F4F0C",
INIT_02 => X"D56B4302AC01005111011BD506AA5205274056900596A539584E2E6DFE4B2418",
INIT_03 => X"9AC0FCBD854688207C90007A1000047A00E588632CA213C8903AD6B55AD0EB5A",
INIT_04 => X"30002047A6FCA110086C402022F2124A8022492580040440002021C922D9109B",
INIT_05 => X"14A206B6838151008D95DD1847811C08002380041F1104002205AC4140DAD060",
INIT_06 => X"1727FF2EB9EF113A10BD32F44289D1F840C1710010344DB9A808FDFF3DE03130",
INIT_07 => X"050700154A00401D00495A06A8D464C5F6B54AA8551040818F4C997AC80CBE05",
INIT_08 => X"0141008801018040E48D50080002B00A0C00801014541E9504703680017F6CB4",
INIT_09 => X"02680000010937986481514E2A29CE010708C0804C6A033F7FCFF9426A41F1AB",
INIT_0A => X"00500001840000C80B410014088040F4A944B1AA313C004554002381B8000500",
INIT_0B => X"A004D1594832824A070AA070AA070AA070AA070AA070AA070AA0725503855038",
INIT_0C => X"501428054278142151262CA50343854E506A2C6898B2950AA6A35B0004284058",
INIT_0D => X"90078E1F840A2B0114020104022460002200050F60E220A06880D2A14050A028",
INIT_0E => X"90078E1F891C239F8908003099C1ACF06273612B3482C0C0078E1F412B1582C0",
INIT_0F => X"1BA1B0FD16770236A4091621C08055C2C0DB012B1582C0C0078E1F412B3482C0",
INIT_10 => X"00101F09C030AB28B03C111C239F870828041BA859F213AFC14AA38043006018",
INIT_11 => X"10E8822A984B0025B0DE6089462660095337B08AA600CA88B143AB11880C2806",
INIT_12 => X"055412D4481128C4CC012A66F304553096004B61BD8068B92400D0004E303689",
INIT_13 => X"589C48082C006A9057CA4385809520F07830001AC2173B00E162563454C40804",
INIT_14 => X"00460848952220592745AC11A544B1BF006850840180A00E1C81900C4190E160",
INIT_15 => X"22088220882208822088220882208CD888088D940D2A3A9D5002001300800C8C",
INIT_16 => X"0080200882208822088220882208822088220882208822088220882208822088",
INIT_17 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_18 => X"FBDFD1FE3EFBD7BBEFBEFA0A245120000000007FFFFFFFF20080200802008020",
INIT_19 => X"F3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF7FFBFAFBBBEFBEFBEFBF7",
INIT_1A => X"CFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCF3CF3CF3C",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000007F3F9FCFE7F3F9FCFE7F3F9F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040000000000000000000000000000000",
INIT_1F => X"4BA550000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0002000087FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974AA550402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"020AA5D7FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5D00000AA007FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAA954BA5504000AA557FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5D00",
INIT_23 => X"7BFFFFFFFFFFFFFFFFFFFFFFFFFAA954BA5500020BA5D7FFFFFFFFFFFFFFFFFF",
INIT_24 => X"7AA974BA5D040200055517FFFFFFFFFFFFFFFFFFFFFFFFAA954BA5500000BA5D",
INIT_25 => X"00000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000080000000",
INIT_27 => X"FFFFFFFFFFFFFAE974AA550002010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"0BA087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550400028007FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAA954BA5D00000BA557FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5D0002",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAA954BA5504020AA5D7BFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"A974AA5D00070925D71FFFFFFFFFFFFFFFFFFFFFFFF7AA954BA5500000825571",
INIT_2C => X"FFFFFFFFFFFFFFEFF7AA974AA5D040500055517FFFFFFFFFFFFFFFFFFFFFFF7A",
INIT_2D => X"D040200008000000000000000000000000000000000000000000000003FFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"A087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550002000087FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAA954AA5D00020AA007FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5504000B",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFF7AA954BA5D00000BA5D7BFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"74AA55000200055517FFFFFFFFFFFFFFFFFFFFEFF7AA974BA5504020BA557BFF",
INIT_33 => X"FFFFFFFFFFDFEFF7AE974AA5D00154105D517FFFFFFFFFFFFFFFFFFFFEFF7AA9",
INIT_34 => X"00000000043FFFFFFFFFFFFFFFFBFDFEFF7AE954AA5D041740055557FFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000007FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(22),        -- Port A data input
DOA(0)   => data_read_a_hi_256(22),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(22),        -- Port B data input
DOB(0)   => data_read_b_hi_256(22),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_23_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"EF20906D902424807BC8241BC81801B97D38AD3C0800103362A6741C80A12A02",
INIT_01 => X"001FFF8409F089003B4422000D80C80106804A7951C5B9D1C828043EA28838F9",
INIT_02 => X"028406A002DC176444683862400003111001303FFC00F240D50146013B300500",
INIT_03 => X"0006C90C010203F80005DC00C52FC380BEAC25886C02034800200200A1008008",
INIT_04 => X"17DFFF8049000BFF878314BFF8488890979800002F702002BB807A068403C280",
INIT_05 => X"DA07F0000000007FF020C814380011FE5E1C2FC3E05FFFF90020000808900010",
INIT_06 => X"10004C9690A8CA008024685184097E81E872C8FFE900FC31348EFDF03BE15E22",
INIT_07 => X"402000001FFBFFFD00080200B8140011F0D8C108155542018D1A302193E94004",
INIT_08 => X"41BE1F5F80003FF0002023FFDF79000000000EFFE309606020008005FC000000",
INIT_09 => X"FC83FE1840C0902400300000000000DFFD4004040C4D32BF7C0EE860003CE680",
INIT_0A => X"10018C24110A860006C620C0312241C482B20420CC56924E2199000C00415037",
INIT_0B => X"4669070510C90C14304043040430404304043040430404304043040218202182",
INIT_0C => X"008000105400C00400100000A018000801000C024000004A940000FFDF820604",
INIT_0D => X"100152100801C17E61841950B1C10FFF57FFC02812F00429DC92C40002000100",
INIT_0E => X"10015210088528E00E02C8200A430A424202A1CAF13F214001521001CBF03F21",
INIT_0F => X"01C1C044006D0C94FB94320880603C420B8001CBF03F214001521001CAF13F21",
INIT_10 => X"30182800A018D9CA8000648528E00D12480202C86040902AC60BACDF0E02D020",
INIT_11 => X"0445C19960A00026880C006739000009B00300010AF5052419D1964419028014",
INIT_12 => X"01844068880CE72000013600600332C140004D101808458A5602E00089202911",
INIT_13 => X"41D0B9023402085020825132C8CB5B4040301009408021144CB042F880100C06",
INIT_14 => X"8E17C0D240406519400500840A9524EE38A1F80E02120018390320F050144CB2",
INIT_15 => X"01004010040100401004010040100100040040000000000001000900FBFFE000",
INIT_16 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_17 => X"0040100401004010040100401004010040100401004010040100401004010040",
INIT_18 => X"0000000000000000000000000000000000000000000000001004010040100401",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000000000000000000000000",
INIT_1F => X"4BA5D0400010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000007FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974BA5D0002000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"00010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA550002000007FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAE974AA550400000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5500",
INIT_23 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550402010087FFFFFFFFFFFFFFFFFF",
INIT_24 => X"FAE954AA5D00000AA007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA55040200008",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010000000000",
INIT_27 => X"FFFFFFFFFFFFFAE974BA5D0400010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0000010007FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAE974AA550002010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA550002",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550400010087FFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"E954AA5D0402038007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550400028007F",
INIT_2C => X"FFFFFFFFFFFFFFFFFFAE954AA5D00020BA087FFFFFFFFFFFFFFFFFFFFFFFFFFA",
INIT_2D => X"D0402010000000000000000000000000000000000000000000000007FFFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000087FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAE974BA550002010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D000001",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFFFAE974AA550002000087FFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"54AA5504000BA087FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA550400010007FFF",
INIT_33 => X"FFFFFFFFFFFFFFFFAA954AA5D04000AA087FFFFFFFFFFFFFFFFFFFFFFFFFFAE9",
INIT_34 => X"000000007BFFFFFFFFFFFFFFFFFFFFFFFFFAA954AA5D00020AA007BFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000007FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(23),        -- Port A data input
DOA(0)   => data_read_a_hi_256(23),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(23),        -- Port B data input
DOB(0)   => data_read_b_hi_256(23),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_24_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100600007FFF000080108004000800020000840041000080808",
INIT_02 => X"0000068002CC07400000090C080002000000103FF811F150231000520ABE4404",
INIT_03 => X"210A0600000203F80005DC00000DC3801EA000000745C4010220000000008000",
INIT_04 => X"07C5FF804900026F8780001DF8000000079800000F300002998078068003C080",
INIT_05 => X"C207F0000000007FF0000004380001FE1E1C07C3E00CFFF80000000000000000",
INIT_06 => X"0002648240F20035A0102000BD0000002802C87FC800FCAA035400001B918600",
INIT_07 => X"0000000001FBFFEC4D2B4AD0B8129063B2CC0000100042018408142F16C01848",
INIT_08 => X"008E1F5F80001FF0000000FFDF78000000000EFFE001600000000005FC000000",
INIT_09 => X"E883FE180000000000300000000000DFFD0000002A80D500000671000004A000",
INIT_0A => X"10018C0411020600048620C030020502000200000400920A2198000800404037",
INIT_0B => X"0641060400C00C00304003040030400304003040030400304003040018200182",
INIT_0C => X"000000001000C00000000000000240058000000000000000000000FFDF000404",
INIT_0D => X"E00880104809C1666594584031010FFF56FFC000104000000010440000000000",
INIT_0E => X"E0088010492064206100E81084200048C0804012500021B00880108012500021",
INIT_0F => X"04100144800803419043064900C0020501840012500021B00880108012500021",
INIT_10 => X"1018140F02C0000809408D206420530270040410004C840041A0D80054109038",
INIT_11 => X"110002C9E8010C00010480B35A0300400041020902F60002260D65B361BAA104",
INIT_12 => X"0228204300166B4060080008240593D0021800020818B06D9802F00030C02060",
INIT_13 => X"143B62023C00142800B04400095DFF90203020042108603100061516EE800C06",
INIT_14 => X"DC1180C7804400044029208301040214AE4C7C02000040206602C10B48110006",
INIT_15 => X"00000000000000000000000000000000000000000000000000000000FBFFE000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"DD5EDCF9822659B6888332000000000000000000000000000000000000000000",
INIT_19 => X"F3CF3CF3CF3CF3DF7DF7DF7DF7DF7DF3DF3DF3DF3DF4D30C2432AEBAEBFE5A15",
INIT_1A => X"C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783DF7DF7DF7C",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000F0783C1E0F0783C1E0F0783",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201008000000000000000000000000",
INIT_1F => X"4BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974BA5D0400000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"00010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000007FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAE974BA5D0000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_23 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0002000087FFFFFFFFFFFFFFFFFF",
INIT_24 => X"FAE974BA550002000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D000200000",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010080000000",
INIT_27 => X"FFFFFFFFFFFFFAE974BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000087FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAE974BA5D0400010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0000010007FFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"E974BA550002000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0000010007F",
INIT_2C => X"FFFFFFFFFFFFFFFFFFAE974BA550002000007FFFFFFFFFFFFFFFFFFFFFFFFFFA",
INIT_2D => X"D0402010080000000000000000000000000000000000000000000007FFFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAE974BA5D0400000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040200",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000087FFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"74BA5D0000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0000010087FFF",
INIT_33 => X"FFFFFFFFFFFFFFFFAE974BA550000010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE9",
INIT_34 => X"000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA550002010087FFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(24),        -- Port A data input
DOA(0)   => data_read_a_hi_256(24),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(24),        -- Port B data input
DOB(0)   => data_read_b_hi_256(24),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_25_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100200002000000080100004000000020000800041000080808",
INIT_02 => X"0000068002CC474000000800000002000000103FFCE302008000000880844A04",
INIT_03 => X"00000040700803FC0105DE00020DC3801EA00000040000000020000000008000",
INIT_04 => X"47C5FFC04904026F8780081DFC040000079C92484F30499299837C168003E400",
INIT_05 => X"C207F0382004407FF0000004382281FF1E1C07C3E00CFFFC090004B05000200A",
INIT_06 => X"1009015C4000000020000000390C10002802C87FC800F8000000000019810600",
INIT_07 => X"0501000001FBFFFD480A0280A816002010800001000054018408102000000002",
INIT_08 => X"0C8E1F5FA21C9FF8004000FFDF7C062031863EFFF75D78004001010DFC000020",
INIT_09 => X"E883FE180C00000000300000000000DFFF00180800000000000660100000A000",
INIT_0A => X"1001DCCC31222730A49620C030020100000200000400921A21D8000804404037",
INIT_0B => X"0641062400C00C00304003040030400304003040030400304003040018200182",
INIT_0C => X"C11160845004D04820000000000000000000000000000000940000FFDF000404",
INIT_0D => X"000800000801C0786184185031810FFF56FFC02812E0182000F2C48304418220",
INIT_0E => X"0008000000002020000008000000000800800002400001000800000002400001",
INIT_0F => X"0000010000000000900000080000000400000002400001000800000002400001",
INIT_10 => X"1000000002002000004000002020000200000000000404000000880000001000",
INIT_11 => X"010000082000000001000001080000000040000100C600800001040000040009",
INIT_12 => X"0000000100002100000000080000104000000002000000081001000000000040",
INIT_13 => X"0010200000000000001004000001080000400080000040010000001080001008",
INIT_14 => X"8C11808200400000400000C20000000420000000030280000000010000010000",
INIT_15 => X"82208822088220882208822088A20C52082081A30080000002005008FBFFF001",
INIT_16 => X"2208822088220882208822088220882208822088220882208822088220882208",
INIT_17 => X"2088220882208822088220882208822088220882208822088220882208822088",
INIT_18 => X"29432D518B45265D82BB4101000005FFFFFFFFFFFFFFFFF82208822088220882",
INIT_19 => X"24924924924924820820820820820820924820924824000A6242B4D34D7F7451",
INIT_1A => X"AC562B158AC562B158AC562B158AC562B1188C46231188C46231189249249249",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000162B158AC562B158AC562B158",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000000000000000000000000",
INIT_1F => X"4BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"02000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAE974BA5D0402000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_23 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000007FFFFFFFFFFFFFFFFFF",
INIT_24 => X"FAE974BA5D0400000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040000008",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010000000000",
INIT_27 => X"FFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAE974BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000007FFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"E974BA5D0400000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000087F",
INIT_2C => X"FFFFFFFFFFFFFFFFFFAE974BA5D0400000007FFFFFFFFFFFFFFFFFFFFFFFFFFA",
INIT_2D => X"D0402010000000000000000000000000000000000000000000000007FFFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"74BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000007FFF",
INIT_33 => X"FFFFFFFFFFFFFFFFAE974BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE9",
INIT_34 => X"000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000007FFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000007FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(25),        -- Port A data input
DOA(0)   => data_read_a_hi_256(25),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(25),        -- Port B data input
DOB(0)   => data_read_b_hi_256(25),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_26_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"E9264EAB20190CA3BA4997AA9002AE9C001006B0778015CFA17E0811039879C7",
INIT_01 => X"F1FFF9BB1F773C7F9BB07DFFFDD863FC5FFF3FEFFBBF9FFB22FFFBC7B9F30686",
INIT_02 => X"9B3184F8AFDEAF300029E4E300FC78A6258548EFFA71C00172082400003A2161",
INIT_03 => X"0084F0FF7FFF1FDD3FEFDCDE981DC3FF5F0D294A7B2B18A0001B9CE6CC606E73",
INIT_04 => X"0FC5DFD7EDFFD66F87FE605DDDBFF3690F9EDB7F5F7AFF639BD7DE37C2FEF591",
INIT_05 => X"F205F0F8E9D199FF76DFEE1C3FCC3FF7BE1FD7C3FFACFBFFDFF7B4FEFFDAA10E",
INIT_06 => X"042648C40179912406C1830639AFBEC14489737FDC00B13BB79DFDB83BF4112A",
INIT_07 => X"763A844769FFBFE4398E4390BB9C28B1D0F049080414583F9468D1AEFC000060",
INIT_08 => X"02C05FD7BC471FBD13D981F7DF7D7E6171AF3FEFE8A3E679FAC1FD1FFFBEB000",
INIT_09 => X"F8CFFE38FF7F6BD928F1ABB47476B5FEF9F59F5FCEEDE73FEE0EFC53B079F5CC",
INIT_0A => X"315BDDCC3B336F7C548667D47B7737AF3FD62601EDC2B66A67B9D60FE4C4427F",
INIT_0B => X"06E19F4DA0E80E903DE3035E3035E3035E3035E3035E3035E3035E981AF181AE",
INIT_0C => X"EBFBF7FEBD66DBFCA3F87501AE7B080607307DCFE1D4077B4D026FFFFBFFAFCD",
INIT_0D => X"0007E010084BCD7FF1B61B5C33813FFFFCFFC7D7D51D6F5FDCB935D7AFEBD7F5",
INIT_0E => X"0007E01001BD8020500008001F010040520201F45EC0010007E01001F45EC001",
INIT_0F => X"1DC0004600400F781429C0080000770001A001F45EC0010007E01001F45EC001",
INIT_10 => X"10003C064000E408010081BD8020600200001EC00040B02007EC09A0E0001000",
INIT_11 => X"360403E434588007200D00F88C84C081C203404B3BFD0402346235408402C080",
INIT_12 => X"07B00040091F1190982038406807C868B1000E401A08FE0012040000FC002001",
INIT_13 => X"7D00212000007C400082D81009FC08281D00001F010021560406758091454000",
INIT_14 => X"FFBFF5FA1040076065F730FC08043A903A80008320C0403C3400008860160406",
INIT_15 => X"D7F5FD7F5FD7F5FD7F5FD7F5FDFF7F7F7F77F9F761FFBFDFFDE5BFFFFF7FF005",
INIT_16 => X"7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5F",
INIT_17 => X"F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD",
INIT_18 => X"B79E923C2CD990AA7F0DDB6B910C8DFFFFFFFFFFFFFFFFFD7F5FD7F5FD7F5FD7",
INIT_19 => X"30C30C30C30C30C30C30C30C30C30C30D34D34C30C35F7AA9ABF0E38E3A8EB62",
INIT_1A => X"C26130984C26130984C26130984C26130984C26130984C26130984C30C30C30C",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000130984C26130984C26130984",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000000000000000000000000",
INIT_1F => X"4BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"02010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_23 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFF",
INIT_24 => X"FAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010000000000",
INIT_27 => X"FFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"E974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007F",
INIT_2C => X"FFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFA",
INIT_2D => X"D0402010000000000000000000000000000000000000000000000007FFFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"74BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFF",
INIT_33 => X"FFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE9",
INIT_34 => X"000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(26),        -- Port A data input
DOA(0)   => data_read_a_hi_256(26),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(26),        -- Port B data input
DOB(0)   => data_read_b_hi_256(26),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_27_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"00080A40000A41248002029000050A088000008242A0004404480002000A1155",
INIT_01 => X"F1FFF1C11F781C129C107DFFFE0860941E81258CA2B71C2220EC1B86E1A00002",
INIT_02 => X"183080988B2EAE00002BE001117C78C6848140CFFA0000800042008000011081",
INIT_03 => X"000000FF7CF91F1D3DEF3CDA881D23FB5C0C21085B0B0820001318C60C204C63",
INIT_04 => X"8FC51FD7EDFDD66E47EE205D1DB7F1490E5EDB7D5CBADB2385D79C3643D4E580",
INIT_05 => X"E001F0C0C991BBFC76DFEA1A3F8C3BC7391F9723FF2CE3FCD6D13096B79C8106",
INIT_06 => X"40000001000000084041830600A40C415004637FC4003021259CFDB01BF80028",
INIT_07 => X"3158954761FA3FE402088220AC1108001080400A400041018468D1A060000050",
INIT_08 => X"02005F0784411E390A4881C7BEFC5F6171CE2F8FE823E778DAC16C1FFBBC9000",
INIT_09 => X"F0C7FEBABF3F6BD108F40E04C0C084F0F8B58B5B8849673F6C0E7A01B00914C4",
INIT_0A => X"B51BFDCC39732F3554866AD57C37BEAF1C152201A4C0B6EA63AAD60B60D4427F",
INIT_0B => X"06F18FC5A0E00F0038D1030D1030D1030D1030D1030D1030D1030F0818688186",
INIT_0C => X"AB6AD7EAB962CBD8A3A83101F47E08040510768EA0C406630D0226FFE375ADE5",
INIT_0D => X"000760000843C561E5C55C42B9011FFF48FFCC57550D63564D1D2556ADAB56D5",
INIT_0E => X"0007600004BD8020100008001F010000130201E44A40010007600005E44A4001",
INIT_0F => X"1DC0000208400D781020C00800007700002005E44A40010007600005E44A4001",
INIT_10 => X"10003C064000C400018080BD8020200200001EC00000382006EC0820A0001000",
INIT_11 => X"3E0403A424108007200102E888808081C20040431BC504021462354004004080",
INIT_12 => X"07B00000015D1110102038400817484821000E400204FE0010040000FC000000",
INIT_13 => X"7D00202000007C400000F81001FC08080500001F0100005E0404758081014000",
INIT_14 => X"8DBBB5FA10400360649310FC08003A903A8000012040403C34000080201E0404",
INIT_15 => X"56D5B56D5B56D5B56D5B56D5B56D7E3D7B57B1C4E17F0944B8D596EEFC7FF001",
INIT_16 => X"6D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B",
INIT_17 => X"D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B5",
INIT_18 => X"2D0200903950C080420948E2D10E8FFFFFFFFFFFFFFFFFF56D5B56D5B56D5B56",
INIT_19 => X"00000000000000000000000000000104000000000004000E5E420000002921C4",
INIT_1A => X"28140A05028140A05028140A05028140A0100804020100804020100000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000140A05028140A05028140A050",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000000000000000000000000",
INIT_1F => X"4BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_23 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFF",
INIT_24 => X"FAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201008",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010000000000",
INIT_27 => X"FFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"E974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087F",
INIT_2C => X"FFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFA",
INIT_2D => X"D0402010000000000000000000000000000000000000000000000007FFFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"74BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFF",
INIT_33 => X"FFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE9",
INIT_34 => X"000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000007FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(27),        -- Port A data input
DOA(0)   => data_read_a_hi_256(27),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(27),        -- Port B data input
DOB(0)   => data_read_b_hi_256(27),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_28_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"02200AA400180030808802A900002A08001280A08A801044104A1000001818C3",
INIT_01 => X"50A00011460214428114180000882214413D0A71592A01D92213D28005210202",
INIT_02 => X"8A54800A210200111100C2110054289220810440030404010844000444410001",
INIT_03 => X"1080010208B51400007800000A000001000108C21008092000018C6295200631",
INIT_04 => X"0008000000017000000028000001610300000010000802202040012040040011",
INIT_05 => X"2000044440048880026A22000026A20000000000000000004994140203000064",
INIT_06 => X"1400922401041008004891224228810080010200040001020800000004000008",
INIT_07 => X"150B001328000001404010040084088404200020455514000224489028492201",
INIT_08 => X"00414000201800004080A0000002480B04008100011000088800081002C19020",
INIT_09 => X"000400001036584108415B4A6A694A0000100101C08200000001000190200044",
INIT_0A => X"004800210C19808400500010009110091500020B408820000200400040811600",
INIT_0B => X"40000800B00100040D8140581405814058140581405814058140580A02C0A02C",
INIT_0C => X"00200248010201008298150006210802043058C46054032981002D00201C8081",
INIT_0D => X"0000A00000400600841041108280300008000140000401028008330000800040",
INIT_0E => X"0000A000000080001000000000000000500000040A40000000A00000040A4000",
INIT_0F => X"00000006000000080020C00000000000012000040A40000000A00000040A4000",
INIT_10 => X"00000000000024000000000080002000000000000000A00000040020A0000000",
INIT_11 => X"2200000404108000000900008080808000024040152000000020000004004080",
INIT_12 => X"0000000009001010102000004800080821000000120002000004000000000001",
INIT_13 => X"2000002000000000000288000020000805000000000001420000200001014000",
INIT_14 => X"408010000000022000D610280000080000000001204000000000000820020000",
INIT_15 => X"00401004010040100401004010042024210218734CD52150A840827504000000",
INIT_16 => X"0401004010040100401004010040100401004010040100401004010040100401",
INIT_17 => X"4010040100401004010040100401004010040100401004010040100401004010",
INIT_18 => X"05822140048D2E57B1348141845C200000000000000000000401004010040100",
INIT_19 => X"04104104104104104104104104104104104104104101A6A0A0EB1861863BC422",
INIT_1A => X"2C160B0582C160B0582C160B0582C160B0180C06030180C06030181041041041",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000160B0582C160B0582C160B058",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000000000000000000000000",
INIT_1F => X"4BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_23 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFF",
INIT_24 => X"FAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010000000000",
INIT_27 => X"FFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"E974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007F",
INIT_2C => X"FFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFA",
INIT_2D => X"D0402010000000000000000000000000000000000000000000000007FFFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"74BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFF",
INIT_33 => X"FFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE9",
INIT_34 => X"000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000007FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(28),        -- Port A data input
DOA(0)   => data_read_a_hi_256(28),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(28),        -- Port B data input
DOB(0)   => data_read_b_hi_256(28),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_29_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"79964E4BA01DACAB9E659792D00AAE160002829C7FDFEFCEE97C2815039D70C3",
INIT_01 => X"50BFF9AB0775343F9AB01DF80D5821FC0FFF3FEFD1AF9FF1207FFBC7B9720586",
INIT_02 => X"0D15846807D207200021C4E200D428A2018408600271C000720A0000003A2161",
INIT_03 => X"0000B0027BBF17C43E6DC05E1A0DC07D1F0000803B2819A00019084345606421",
INIT_04 => X"07CDC047A4FB526F807C681DC4B97369078249370F482E62BA414627C2FE3000",
INIT_05 => X"F204007861C088FF0EFF260407C427F19E03C7C01F8CF80749B390EA4BCA202C",
INIT_06 => X"000248C00079800406C081023B233E804488527FDC008019968D74982C94110A",
INIT_07 => X"5229000221FF8000398641903B082831D05000200000083F942850AEB4000221",
INIT_08 => X"00805FD0180E1F8C1111A0F041056A0100A11FE000916249A800B915FE82B020",
INIT_09 => X"F80C000055FF7C492840AAB45456B55E015015058665A31DA603A4539058F54C",
INIT_0A => X"000850400A11414C005005000B51158936D20601A98A204006114005C4800217",
INIT_0B => X"40201948B029029409A3401A3401A3401A3401A3401A3401A3401A9A00D1A00C",
INIT_0C => X"40B1225C1506512C83E85500AC3A080406305587A154023141006DFFF89E82C9",
INIT_0D => X"0000A01008480D3EB4A24A0C910037FFFC0007C7C0140D0B50A8218102C08160",
INIT_0E => X"0000A010010080005000000000000040520000141EC0000000A01000141EC000",
INIT_0F => X"00000046000002080429C0000000000001A000141EC0000000A01000141EC000",
INIT_10 => X"00000000000024080100010080006000000000000040B000010401A0E0000000",
INIT_11 => X"3600004414588000000D00108484C080000340483B590000202000008402C080",
INIT_12 => X"00000040090210909820000068008828B10000001A0802000204000000002001",
INIT_13 => X"20000120000000000082D800082000281D000000000021560002200011454000",
INIT_14 => X"B29450580000066021F6303C000408000000008320C000000000000860160002",
INIT_15 => X"816058160581605816058160589625662522506344FF9FCFFF62EB6DFF001004",
INIT_16 => X"1605816058160581605816058160581605816058160581605816058160581605",
INIT_17 => X"6058160581605816058160581605816058160581605816058160581605816058",
INIT_18 => X"F2DDCFFFBEFFCF07FFBFFD41800C05FFFFFFFFFFFFFFFFF81605816058160581",
INIT_19 => X"7DF7DF7DF7DF7DF7DF7DF7DF7DF7DD75D75D75D75D77FFBF3F7DFFFFFFD779F3",
INIT_1A => X"FEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDF7DF7DF7DF",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00001F7FBFDFEFF7FBFDFEFF7FBFD",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000000000000000000000000",
INIT_1F => X"4BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_23 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFF",
INIT_24 => X"FAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010000000000",
INIT_27 => X"FFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"E974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007F",
INIT_2C => X"FFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFA",
INIT_2D => X"D0402010000000000000000000000000000000000000000000000007FFFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"74BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFF",
INIT_33 => X"FFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE9",
INIT_34 => X"000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(29),        -- Port A data input
DOA(0)   => data_read_a_hi_256(29),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(29),        -- Port B data input
DOB(0)   => data_read_b_hi_256(29),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_30_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"FFDFF3FC3EFFF7FFFFBFFA000000000000000000000000000000000000000000",
INIT_19 => X"F3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF5F7AEBEBFBEFBEFFEFFF7",
INIT_1A => X"CFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCF3CF3CF3C",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000007F3F9FCFE7F3F9FCFE7F3F9F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000000000000000000000000",
INIT_1F => X"4BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_23 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFF",
INIT_24 => X"FAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010000000000",
INIT_27 => X"FFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"E974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007F",
INIT_2C => X"FFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFA",
INIT_2D => X"D0402010000000000000000000000000000000000000000000000007FFFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"74BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFF",
INIT_33 => X"FFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE9",
INIT_34 => X"000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(30),        -- Port A data input
DOA(0)   => data_read_a_hi_256(30),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(30),        -- Port B data input
DOB(0)   => data_read_b_hi_256(30),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_31_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"129000008004A00804A40000400800020000000C005FEA005800200400050100",
INIT_01 => X"A15FF18019700810180065FFFC0040801E80258CA2951C2200EC0906A0804140",
INIT_02 => X"146000808A0C060444692000402850040400408FF80000000010000000004000",
INIT_03 => X"000000FD74480B1C3D951C5A800D03FA1C0C21084B0300000012108518004842",
INIT_04 => X"07C51FC7EDFCA26E07EE001D1CB6904A061EDB6D4C30490281831C1602D0E480",
INIT_05 => X"C001F0808181117C7C95C8183FA099C7181F8703FF0CE3FC0201209010988002",
INIT_06 => X"00000000000000010001020400840C41C000617FC0003021259CFDB01BF00020",
INIT_07 => X"0000000441FA3FE400080200A810000010804008100040018448912040000040",
INIT_08 => X"00011F0780011E38004801C79E7C162231862E8FE00166704041240DF93D0000",
INIT_09 => X"F0C3FE180D89279000B00000000000D0F80088080849673F6C0E780020091480",
INIT_0A => X"1011DCCC31222730048620C4382204A608142002A440924A6188020920404437",
INIT_0B => X"0661874500E00E00304003040030400304003040030400304003060018200182",
INIT_0C => X"810040801060C04821202001A05A00040100240A80800442040202FFC3200444",
INIT_0D => X"000740000803C0616184184031010FFF40FFC407500020004C10060204010200",
INIT_0E => X"0007400000BD0020000008001F010000020201E04000010007400001E0400001",
INIT_0F => X"1DC0000000400D701000000800007700000001E04000010007400001E0400001",
INIT_10 => X"10003C064000C000010080BD0020000200001EC00000102006E8080000001000",
INIT_11 => X"140403A020000007200000E808000001C200000308C504021442354000000000",
INIT_12 => X"07B00000001D0100000038400007404000000E400000FC0010000000FC000000",
INIT_13 => X"5D00200000007C400000501001DC08000000001F010000140404558080000000",
INIT_14 => X"8C1380DA10400140640100D4080032903A8000000000403C3400008000140404",
INIT_15 => X"02008020080200802008020080200C1808008184012A08041202500AF87FF001",
INIT_16 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_17 => X"0080200802008020080200802008020080200802008020080200802008020080",
INIT_18 => X"000000000000000000000002001005FFFFFFFFFFFFFFFFF02008020080200802",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000000000000000000000000",
INIT_1F => X"4BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_23 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFF",
INIT_24 => X"FAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010000000000",
INIT_27 => X"FFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"E974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007F",
INIT_2C => X"FFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFA",
INIT_2D => X"D0402010000000000000000000000000000000000000000000000007FFFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"74BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFF",
INIT_33 => X"FFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE9",
INIT_34 => X"000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(31),        -- Port A data input
DOA(0)   => data_read_a_hi_256(31),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(31),        -- Port B data input
DOB(0)   => data_read_b_hi_256(31),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_0_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"ED39BA795990D275FB4A6E96ACC4731DEA4598B0AFB54867F6EE4618C3749807",
INIT_01 => X"58A0047D8607944AC7DA180001ECA2444042106208408208C20022E9173734B3",
INIT_02 => X"8B1E49562021F8051500147A0E162923024F28000415F5787B09FBF999BB1EFC",
INIT_03 => X"1013BF028A959403C06A23A147723C01E140088280C4CF6996088862C7922221",
INIT_04 => X"781A003802015D9078011DE20340699198600000B08694916434804825241311",
INIT_05 => X"2CA000587E10C880036A3103C00F2000E1E0383C00730002B4409845E4425171",
INIT_06 => X"179B48CFF95DCF9EF730E1C3BB731138AF7B888025340C0888430047040FEE18",
INIT_07 => X"AF155113160400185F87C1F05707D415E664A6E7C5551EBE783060CEB164833F",
INIT_08 => X"4D7E40002B7AE005FDB47600208229010C6101001EFE198C96B0528202C0DCB4",
INIT_09 => X"062400608234D864444081048A80CC00062D42D30222108091C107A1DA040267",
INIT_0A => X"204A21008E514844EB5145000255DA599581D3A9583C24351240B58298011308",
INIT_0B => X"E08C4830F81380CE0F89E07A9E0789E07A9E0789E07A9E0789E070CF0184F038",
INIT_0C => X"3A4E9D63EA180EB150CA1CA45C254D4AF4AA414568729139F2A12C0000016110",
INIT_0D => X"F0009E0FC048211E9C11C31F82E4A000890022B827EB52F52347F174E93A749D",
INIT_0E => X"F0009E0FCC42EFDFBF0AE03080E2AEB2E0F1F80FA97FE0F0009E0FC40FA97FE0",
INIT_0F => X"0231F0BD9E3FC08FEBD6F661C0E008C3CB5F040FAB3FE0F0009E0FC40FAB3FE0",
INIT_10 => X"20180309A0F83BE2B87C7C42EFDFBF187806013879BA878FE807F65FBF12E038",
INIT_11 => X"0BE9F01FC8B38C2098DAE007F323A0C83136B248831ACBFC8BBDCAB779BC699F",
INIT_12 => X"004C72BEC800FE7464290626D7003F9947184131B59003FFEC07F00003F01FB9",
INIT_13 => X"A0FFDA2A3C0202B8776A2FA7F023F7D065703080E29F1B2BE9F8A27E6E915C0E",
INIT_14 => X"016C2D25E52630BB1AE49C2BA7F98D6F846DFC0C2352A0024B83F07F198BE9F8",
INIT_15 => X"749D2749D2749D2749D2749D2749F285F25D2C500815A5522CB5A4B400000CD4",
INIT_16 => X"49D2749D2749D2749D2749D2749D2749D2749D2749D2749D2749D2749D2749D2",
INIT_17 => X"9D2749D2749D2749D2749D2749D2749D2749D2749D2749D2749D2749D2749D27",
INIT_18 => X"31C136AD8E9B562BA39E2600654BA800000000000000000749D2749D2749D274",
INIT_19 => X"4104104104104104104104104104104104104104104104109C83B8E38E2ABE71",
INIT_1A => X"0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0410410410",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000007C3E1F0F87C3E1F0F87C3E1F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000187FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"BAF7FFD55EF007FD75EFFFAE97555557BD75EF5D000000000000000000000000",
INIT_1F => X"000AA843FE00AAFBE8B45AA803DFEFA28428B455D0017410A28428AAAA2FBD54",
INIT_20 => X"FEBAA2D5401450051401555D7FC0145F7AEBFFFF08002AA10A2AABFEAAA2FFC0",
INIT_21 => X"D755555517FFEFA280021FF082E974AA5D7BFFE000804000BAAAAAAAB45557FF",
INIT_22 => X"EA8B45005168A10AA8028A10087FD7410557FC21555D51574AAA2FFE8B455D7B",
INIT_23 => X"AE95410AA80000005D003FEAAFFAEBFE00A2803FEBA002A820AA0800174BA5D2",
INIT_24 => X"2AEA8A10000417410A2FFE8BEFF7FFE8B45FFFBC00005D003FF45557FC01FFFF",
INIT_25 => X"00000000000000000000000000000000000000557DF5500003DFEFFF84175EFA",
INIT_26 => X"5F524AFE38B780154BAFFF1D54AF0075D75EFEBAE9554540754717F1F8000000",
INIT_27 => X"50B6AABDE12BEA0AF010B7D1F8F47E00A2DB45AA8A3AFD7B68E2AB78550E1255",
INIT_28 => X"E9257F1E816D557095EAAA2D1401D500002A150038038E285D7F78FD7000B6AB",
INIT_29 => X"5A87AAD178A8002D1D21C5E8257D5C7AA854008700249243A412EBFF5542A43F",
INIT_2A => X"52A82000E3A5D2150AB8F401471EDBC0B680900AAF52B474385D75C502D15754",
INIT_2B => X"FD7E9541242FE920AD082E10A28F6A150012A2F02AFFDF40E85F475451D502D1",
INIT_2C => X"0550E87B7A405B52AAD152BD00151EAFEDB52E3F1EFFFF485A2DA3D5D24BD417",
INIT_2D => X"57F40545850000000000000000000000000000000000000000000005AAF55508",
INIT_2E => X"F7AEAABFF5D2A81151FB8635A02FA69574BAF7D5555AF0D79D55FFA2AC974450",
INIT_2F => X"8D46F6ABE7082AAAAF2FAC77FE00FF16565B2FA9075F4F7B3EBDF50FEAEAAB55",
INIT_30 => X"56803CE3AEB038662E5D81406014D5D51F5E08A394003A908B8410E707EF34A0",
INIT_31 => X"4AF0151555AF58794040077D774FAE8C798A11A0EAEF75F7AA84001A7052C952",
INIT_32 => X"4E1870108B11020AD4AA05542A0A05051023F9A9D57B63BFBF906CB45FABC095",
INIT_33 => X"F5F0DA6BC9525688C1A2A0C06E9FEE5555BE48AB2A2AE0A0F20C43EAC562245B",
INIT_34 => X"000000FF80F55E25C00A0BA7FBED407A97F6F35F498B96BEB12DAAB77558ABD5",
INIT_35 => X"8000000FF8000000FF8000000FF8000000FF8000000FF8000000FF8000000FF8",
INIT_36 => X"00000000000000000000000000FF8000000FF8000000FF8000000FF8000000FF",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000008000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(0),               -- Port A write enable input
DIA(0)   => data_write_a(0),        -- Port A data input
DOA(0)   => data_read_a_lo_512(0),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(0),               -- Port B write enable input
DIB(0)   => data_write_b(0),        -- Port B data input
DOB(0)   => data_read_b_lo_512(0),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_1_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"212C001411984004084D000508C53810A03D1450E839B003342114428A000803",
INIT_01 => X"08000010400A0008010600000084005000400002000000000000000000140000",
INIT_02 => X"C084484000002014400205851002007030450E0000A606C8C44CB4C6666C00E0",
INIT_03 => X"CCF7CE0002058001000000800240200001018CA1800001091408463061120118",
INIT_04 => X"082800100000000040000900010000100040000000008411600401C02100000C",
INIT_05 => X"10800202080422000020012200000000810000200000000004020C00200011A0",
INIT_06 => X"56BDBFBC48C315A8660C18305750C008940D8000011000820001000104050004",
INIT_07 => X"8B4344400004000150248912154404C6060A2FE24555013E13060C158AC97F01",
INIT_08 => X"00082080087A000559102400200281000469000008B000000090108000400430",
INIT_09 => X"0000000000001004140545402820020000010010208000008041060008200001",
INIT_0A => X"2102210182004840007845004044020000200080080844200000048088000000",
INIT_0B => X"48800000190191064620646A06468064680646A0646A06468064690321503234",
INIT_0C => X"02008100200800A1100707040101E20BE0B002605C1C110848200C0000000800",
INIT_0D => X"F000A000C0000012187087010AE4B00000000810010040108104100408020401",
INIT_0E => X"F000A000CC4200002F08E03080000010F18058000003C0F000A000C4000003C0",
INIT_0F => X"000000078808C00000023461C0E00000012704000003C0F000A000C4000003C0",
INIT_10 => X"201803000000240218C0044200001E1878060000000AAC00680000001F10E038",
INIT_11 => X"2100B00048230C200009A0001303204800025200040A00D000000202090C281F",
INIT_12 => X"00000002C9000260640900004D0000904618400012900001EC03F00000000039",
INIT_13 => X"80025A0A3C020000002A8400B00007806070308000000961002880204A901C0E",
INIT_14 => X"000801046004308A185000020128000904285C0C0312A0020000000838810028",
INIT_15 => X"0401004010040100401004010040100010410C002000040280100000000008D0",
INIT_16 => X"4010040100401004010040100401004010040100401004010040100401004010",
INIT_17 => X"0100401004010040100401004010040100401004010040100401004010040100",
INIT_18 => X"48D757DF8A9410218E8A56085142020000000000000000004010040100401004",
INIT_19 => X"555555555555555555555555555554514514514514550431A581924924B02651",
INIT_1A => X"4BA5D2E974BA5D2E974BA5D2E974BA5D2EB75BADD6EB75BADD6EB75555555555",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800005D2E974BA5D2E974BA5D2E97",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000607FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"10AAAABFFFFFF803FE10F7D17FEBA55556AAAAAA800000000000000000000000",
INIT_1F => X"EBAFFD555400557BD54BA5D7FFDF45A2FBD75EFA2AE97555F7FBFFF45FFAE800",
INIT_20 => X"ABEFA2D568A005D5157400AA8028AAAF7FBD54AA002A955555D7FE8ABA082EBF",
INIT_21 => X"FDF55AAFBC0010555540010550417555AA8028BEFAAAE97555082A80000AA802",
INIT_22 => X"BD7410550428ABA5D5168ABA552EBDFEF5D7FEAA00AAAABFEAA007BC0145FFFF",
INIT_23 => X"FFEAB55557FFFEBAAAD568B45A2D5575555D7FC2155F7AEA8BEFAAAA954BA557",
INIT_24 => X"D7BD74000804154BA082ABFF55FFD57DF45F7D568ABAF7AABFFFF082ABFFFFFF",
INIT_25 => X"000000000000000000000000000000000000002EBFFEFA280021FF082E974AA5",
INIT_26 => X"5E175EFF57BF8FC2000BEA4BAE97F78A3FE28E3D17DEAA485FE8E02B50000000",
INIT_27 => X"455571E8A2A087BF8EAAEB8E0016D5D75D54BA5D7BFFF7DA2FFD55EFAAA49554",
INIT_28 => X"157428145A00AA8A2FBD7B6DF6AA28550E10405F7A4AFE38EAA0924921C2FD55",
INIT_29 => X"8E971471C7010B7D168F47400A07A28415A001684104155C5B6DF6DBEFBFAA07",
INIT_2A => X"BFBD7B6A0BF492415FC20105D24AAABF1FFBC7010FF8A38FEF557FEAB78B6AAB",
INIT_2B => X"017EBA4A8EB8F6FFD5FE8B7D557495EAAA2D16D1FDBED56A55557A43DE385FD4",
INIT_2C => X"854008700249243A417FFF41542F5D717FE2AAAA56DEBD17FE3DF7FB7FEBFE38",
INIT_2D => X"07DFCA127B8000000000000000000000000000000000000000000002A3D5C7AA",
INIT_2E => X"AAFBD55FFAA8416545A6FB60F47AF2A00010F78028B15F7823FEAAA2D57DFBA0",
INIT_2F => X"22A38C20B2552E975F758516AAAA0869AAAB8A7C19C55550E8574BA557BFFFEF",
INIT_30 => X"55FFEFBCEE5FBAACB10085EE5DE10A2AEBFF55F7BAAA8565DBAC1112FFAC21A0",
INIT_31 => X"BEA097BEAAFAF2863FA00DD574201E7AD1FFF5575841DE08007FC20480028957",
INIT_32 => X"54FF57EFBFA18D4FBFFF40FF809D4000D7FC00FC5D062BBA05ED5034472A02EA",
INIT_33 => X"7DFBFF6963FCAAA2283CF14050062B0A2F7AE8B5D5D51F5E18ABD5EAFFF2AF95",
INIT_34 => X"000000002CB75F7AA84001A7052C95256807DC31AA8114DE55F5BED201FFFED1",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000008000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(0),               -- Port A write enable input
DIA(0)   => data_write_a(1),        -- Port A data input
DOA(0)   => data_read_a_lo_512(1),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(0),               -- Port B write enable input
DIB(0)   => data_write_b(1),        -- Port B data input
DOB(0)   => data_read_b_lo_512(1),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_2_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10E44660018259B2843913100062C98004802322D3E030235201006009B2813",
INIT_01 => X"000AC188084900481C8024A542400340404000720885800802000906E4910204",
INIT_02 => X"82040072AC248C31010204880000007401044C0550200000480E0080001300E0",
INIT_03 => X"0080812C130D0A0D1193088802182142494D218220021100001A8020C1004A00",
INIT_04 => X"090D0AD62824A44A428408540D1610020C6E510818923441A4908B0503404201",
INIT_05 => X"5000A004081122242420480A14A99C428908122144244150906124248C002168",
INIT_06 => X"1400088400450000460000001308890094082015800011012D41D518044C1100",
INIT_07 => X"26731111491C1541324C1114BD880004002040204050413F1400100480000201",
INIT_08 => X"02410582881E0C1511D02082AAAB016A2463288549B044605201D10AE11B0020",
INIT_09 => X"E80394280E40158020B591000800481051241A4A404B5035C60904502054E000",
INIT_0A => X"0102C9E12202EA6014D027C418428E220A5500024808922801A0900A84454458",
INIT_0B => X"4600070110C10D04340043400434A043420434A04342043480434102184021A0",
INIT_0C => X"E9CA34328E44CA1401306100A246000402100C088104010AC8005C5681812B04",
INIT_0D => X"0000A0000801487334E34C1A980001550055481204090A4C01351253A728D194",
INIT_0E => X"0000A000013800004000080000000000500000B01480010000A0000150148001",
INIT_0F => X"0000000608000A500409000800000000012001501480010000A00000B0148001",
INIT_10 => X"1000000000002400000001A100004002000000000000A0000360018040001000",
INIT_11 => X"380001C01048000000090298040440000002400008C400022042004080028000",
INIT_12 => X"0000000009530080880000004813802090000000120C94000200000000000001",
INIT_13 => X"4C000100000000000002E0000950002018000000000001580002508010440000",
INIT_14 => X"7120642000000400015020500004221018000082008000000000000820180002",
INIT_15 => X"5094A5294A5294A52942509425094209461468000822241A03835D88482AB001",
INIT_16 => X"09465094A5294A5294A5294250942509425094A5294A5294A529425094250942",
INIT_17 => X"94650946509465294E5294E5294E5094650946509465294E5294E5294E509465",
INIT_18 => X"080271AE180616A38A18FA204452A7F03F03F07E07E07E05294E5294E5294E50",
INIT_19 => X"20820820820820820820820820820820820820820820490C04102CB2CB2EB2C0",
INIT_1A => X"8944A25128944A25128944A25128944A25128944A25128944A25128208208208",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF1F804A25128944A25128944A2512",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000787FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"AAAA843DFFFAAD1554005D7FD74AA00040015500000000000000000000000000",
INIT_1F => X"F45AAAAA8A10A2AE80010A2AA975FF5D003FE10F7D17FEBAF7D5420AA0855420",
INIT_20 => X"FF45A2AA975EFA2FFD7555FFFBFFF45AAFBC20AAF7D1575EF55517DF555D2EBF",
INIT_21 => X"95555552E974105D517DF55AAAAAABEFAAD1575EFAAAE974AA5D51554BA5D7FF",
INIT_22 => X"E82010F7AABFE10FFD542145FFD5554AA555555555557FE8ABA082EBFFFFAAAE",
INIT_23 => X"FBC0010AA802ABEFAAD540000FFD540000AA802AABAF7FFC2010AAAE821EF552",
INIT_24 => X"A8028BEFAAAE821550851420AA002E800AA08042AB45007FC00BAFFD168BEFF7",
INIT_25 => X"000000000000000000000000000000000000002E80010555540010550417555A",
INIT_26 => X"AE95F40002157F470AABE803AE97A2DF55400557FD54AA1D04001C5150000000",
INIT_27 => X"EF55517DFC5552ABDF45B6AEAFFD5F7A482000BEAE905C755003FE28E3D17DEA",
INIT_28 => X"0BA5FD0154BA5D7BFAF7DA2AE955EFAAA495545E3F5EFF57F7FE80082FFDE105",
INIT_29 => X"8AAF082AB8EAAEB8E0016D5D2A924105D5B7FF7DB6AAAABC7BEDB505EFBEA407",
INIT_2A => X"95038AAAEAF1D7410E80000FF8438E00B6DF68FEF4871D24BA495B5556D5571E",
INIT_2B => X"1ED1EFEAF1EFFFDEAD1C5010AA8E2FBD7B6DF47A00EBDB50000A380AAE28E804",
INIT_2C => X"5A001684104155C5B68E2DBEFBFFBC703AE2DF42AAA002A851C214003FF68007",
INIT_2D => X"50002155510000000000000000000000000000000000000000000002087A2841",
INIT_2E => X"55003FEAAAAD57DEBAA2FDDC01051FBD74BAF7802AB05AAFBD5400557BD54AA5",
INIT_2F => X"7AF7FC20B2F7FBC015D58517FF555D2ABDF55F782BEB47AFAD00010F7AA82155",
INIT_30 => X"55FFFFC20FFF3AE544108410174BA557BEABEFAAEBD55FFAA1456547A2D360F4",
INIT_31 => X"0BA547FD75FF58516AAAA0828AAAB4A78016545540400010557BFDFFFF7822A9",
INIT_32 => X"550AAFACAAA122AA8954BAA2AE9D545002A800A8FF862BA00F2F9E8F0050D442",
INIT_33 => X"954505C417FFFF08555555BAAD335B57AB5155400A2AEBFF45FFFB404007FFBD",
INIT_34 => X"00000000061DE08007FC2048002895755FFAEBCFE57BBA57002DF3C4AAAA002E",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000010000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(0),               -- Port A write enable input
DIA(0)   => data_write_a(2),        -- Port A data input
DOA(0)   => data_read_a_lo_512(2),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(0),               -- Port B write enable input
DIB(0)   => data_write_b(2),        -- Port B data input
DOB(0)   => data_read_b_lo_512(2),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_3_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"210C44A20020248B08431120001604B8156023104C40771B3430400A02380206",
INIT_01 => X"015A2A4050B009683C0422C992000B61404040028804A0080A000C16A8990A0C",
INIT_02 => X"C0A406500CE0A95011000D1501005274B5041AB330860281CC08008222170060",
INIT_03 => X"AB488054270F08E1289084C8020420E005A48DA16C021100003A46B06900C91A",
INIT_04 => X"848966150DA0A02941A4080C612A104201C689044382FD403C17E491829B259B",
INIT_05 => X"D006620608843116942508120A208D18A5050160C600D4C894600094B49CA068",
INIT_06 => X"12002D9401C70008060408141788E2C094887033080071913209CC8004640100",
INIT_07 => X"221111454874CCC4122C0932155400C2023940284000003E15020525CE805E11",
INIT_08 => X"020103C9984A0AC511102029869D974214EDBA132891000052C1750B48290020",
INIT_09 => X"60808C8A2E41351020004148A289428730A51E5E644C8233A0090E1020208100",
INIT_0A => X"A4000041A600417914506F955D6422000934000A090A94A020229603A414144D",
INIT_0B => X"469100841001000406D04065040650406D0406D04065040670406C8201782032",
INIT_0C => X"6A4AF532A8040AF821042D01F14084030070262810340402C0000CCE4CC12520",
INIT_0D => X"000800000401C333494594532980733302CCC81300094E5C91200257AD2AD795",
INIT_0E => X"00080000051C0000400000000000000800000190148000000800000450148000",
INIT_0F => X"0000010000000B100409000000000004000005101480000008000004F0148000",
INIT_10 => X"0000000002000000000001B00000400000000000000400000168018040000000",
INIT_11 => X"1000034010480000010002D804044000004000812E4400002440014080028000",
INIT_12 => X"0000000100570080880000080015C02090000002000CCC000200000000000040",
INIT_13 => X"1C0001000000000000104000094C002018000000000040100006418010440000",
INIT_14 => X"4128652000004404010E20500004208018800082008000000000010000100006",
INIT_15 => X"5795A5595A5595A5595A5595A5595E1152556D008028341B13924D80C2E67009",
INIT_16 => X"69565795A5595A5595A5595A5595A5595A559525795257952579525795257952",
INIT_17 => X"95256956579525495E5595A5495E5595A5495E5595A569565795256956579525",
INIT_18 => X"7818F18E0C8514298B0C52A0115009AA9556AAD552AAD5556956579525695657",
INIT_19 => X"24924924924924924924924924924820820820820825042C0000249249202A60",
INIT_1A => X"8D46A351A8D46A351A8D46A351A8D46A353A9D4EA753A9D4EA753A9249249249",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF248086A351A8D46A351A8D46A351A",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"EFAAFFD54AAF7D168B45AAAABDF5500002AA1000000000000000000000000000",
INIT_1F => X"F45FFD168AAA0855420AAAA843DFFFAAD1554005D7FD74AAA284001550055421",
INIT_20 => X"55FF5D003FE10F7803FEBAFFD5420AA080400155AAD5554AAF7802AB4500043D",
INIT_21 => X"28B45A2AE82155A2FBFFEBA0800021550855555FFAA84001FFAAAE80010A2AA9",
INIT_22 => X"168ABAFFFBD54BAAAAE97400A2FBC20AAA284175EF55517DF555D2EBFE00AA80",
INIT_23 => X"AA954AA5D7FFFF45AAAA975EF007BD7555FFFBFDF55AAFBD55EF5D2EBFE10085",
INIT_24 => X"AD1575EFAAAE974AA5D00175555D0015410F7AAAAAAA55043DE00FFFFD5555AA",
INIT_25 => X"0000000000000000000000000000000000000004174105D517DF55AAAAAABEFA",
INIT_26 => X"ABC04001C51551471D7AAF1D05D2EBD56DB7DBEAEBFF551C042AA101D0000000",
INIT_27 => X"92EB842FB5508043FF55EBD56ABD75D5B470AABE8A3AFD7A2DF55400557FD54A",
INIT_28 => X"557FD2082000BEAE905C755003FE28E3D17DEAAEBDF40002550F47155AADB504",
INIT_29 => X"DF40552ABDF45B6AEAFFD5F7A48017DAAFFFAE821C0A0717D1C5B575FFB68E82",
INIT_2A => X"C55D7492E90E3808756DA92EBFFD74BAE3AE85480FFFFC00AABE8E105C755517",
INIT_2B => X"43AE10EAF5C5547FF80954AA5D7FFAF7DA2AE905EF0075D5545E3F5EFF57F7D5",
INIT_2C => X"5B7FF7DB6AAAABC7BEDB505EFBEF5C7092FF801756D490A10438EBA4B8E92410",
INIT_2D => X"D0028A00510000000000000000000000000000000000000000000000E124105D",
INIT_2E => X"AAFBD54005D7BD54AAF78002155515157555AAD142040A2D57FFFFFFAEBFF555",
INIT_2F => X"051AE955F7AAFBC0000AF843FF5500003FF55AAFD6AB455157D74BAF7AAA8B45",
INIT_30 => X"FF557BD74EFFBACD41577B8400010F7AA8215555003FEAAAAC53DEB8A2FDDC01",
INIT_31 => X"0BAF7AA8015558517FF555D2ABDF51F782BCB47ABAE801FFAAFBEAA105D2E955",
INIT_32 => X"214FA2D3EAF57AFFDD7555082AA0AAA00557FEA8A2FDD64BAAF8282012AFFEC2",
INIT_33 => X"820AAAB842AA00000028AB0AAFF48547AE04174BA557BEABEFA2AA951FF88554",
INIT_34 => X"000000002A80010557BFDFFFF7822A955FFFFC21FFF3BE40412DE02955FF082A",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000008000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(0),               -- Port A write enable input
DIA(0)   => data_write_a(3),        -- Port A data input
DOA(0)   => data_read_a_lo_512(3),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(0),               -- Port B write enable input
DIB(0)   => data_write_b(3),        -- Port B data input
DOB(0)   => data_read_b_lo_512(3),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_4_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A108400020612C80284210081034849800A000303100048B3432C82904204006",
INIT_01 => X"210668000008004C1C20250E12100368403008418984014902030906A8910200",
INIT_02 => X"120404C0024C0600000206100008402404040C00F104008040080080001310E0",
INIT_03 => X"7728805052470B5C1B873C04121D03845D0020CA0822018000080084C1000002",
INIT_04 => X"0B899E43891686690790485D5C3E02000E9892201D306D03A9835C16029AC186",
INIT_05 => X"C001E080005030767434C0003C8A01D6B81C5703C82CDBC000072400089C8120",
INIT_06 => X"1000088100410000460002041300004084080070D00030032009700024641102",
INIT_07 => X"4261950408CCBC2012048310951000000003402A4000143E1008912480000211",
INIT_08 => X"00811007AC0A1EB5131120C79E7D176251E53E80E8B361604041340838452020",
INIT_09 => X"C08360820C0912800035F1801630A8260900180C00C8021C800FEE522020A108",
INIT_0A => X"8400F88C166262E940D00D410D62AD02091704024D0A02882192020DA0544043",
INIT_0B => X"4011078510C90D143142430C243042430C24304243042430C24305121A612186",
INIT_0C => X"C08060101000C00401008800F004140009400E4002A0010240000DC3C080002C",
INIT_0D => X"000800100001C07261C51C42390240F050C3C000950008088130040100018000",
INIT_0E => X"00080010003510004000000000000048010002E0100000000800100220100000",
INIT_0F => X"0000014008001550000800000000000400800280100000000800100360100000",
INIT_10 => X"00000000020000080080009410004000000000000044080000D8008000000000",
INIT_11 => X"000005800008000001040168000040000041000100EC00004002214000008000",
INIT_12 => X"00000041003C000008000008200D00001000000208050C000200000000002040",
INIT_13 => X"17000100000000000090000002C8000008000000000060000004480000400000",
INIT_14 => X"8400C00208004844C00800000000528008000000008000000000010040000000",
INIT_15 => X"0100800004030080000C010000A00D1804404912802A261B53104810DB1E0028",
INIT_16 => X"000C030000200C01000020040300800004030000000C03000000040100802004",
INIT_17 => X"008020040100C010000200800004010040300800000020040100C03000020000",
INIT_18 => X"40C700FC0A000280C68A08A950520E964C3269B2C9864D30000C030040100800",
INIT_19 => X"555555555555555555555555555554514514514514526991A199A28A28981451",
INIT_1A => X"41A0D068341A0D068341A0D068341A0D06A351A8D46A351A8D46A35555555555",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF771F60D068341A0D068341A0D0683",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FF087FFDF5508003FEBA087FD54BAAA841540055000000000000000000000000",
INIT_1F => X"F5500003DF455555421EFAAFFD54AAF7D168B45AAAABDF55A2802AA1000002AB",
INIT_20 => X"DFFFAAD1554005D7FD74AAAA840015500002AABA082E954005500021FF5D2EBF",
INIT_21 => X"68BEF080028BFF0855555455500174BAA2AABDE0055517FF555555420AAAA843",
INIT_22 => X"168ABA0055574BA5555554BA5D0400155AAD1554AAF7802AB4500043DF45FFD1",
INIT_23 => X"0400010A2AA955FF55003FE10F7803FEBAFFD5420BA085168A00007BFDE10085",
INIT_24 => X"855555FFAA84001FFAAFBEAB45002A97545F7D1555EF55043DF5555517DEAA5D",
INIT_25 => X"000000000000000000000000000000000000002A82155A2FBFFEBA0800021550",
INIT_26 => X"5BC042AA101D0A28BC7007FFDF45080A3AEAA007BD2482BE84124285C0000000",
INIT_27 => X"004100021FF492AB8F7D1C0438E381451471D7AAFBD0492EBD56DB7DBEAEBFF5",
INIT_28 => X"FED1C5F470AABE8A3AFD7A2DF55400557FD54AABE84001C5550A28ABA1424974",
INIT_29 => X"FB5508043FF55EBD56ABD75D0428BEF005557545490012482B6A0BAE2849557A",
INIT_2A => X"6DA101475FDE10145F68A921C55504924955524AA140E0717DAADB50492EB842",
INIT_2B => X"43AF6D405F78E3A1C2002000BEAA905C755003FE28E3803DEAAEBDF40002557F",
INIT_2C => X"FFFAE821C0A0717D1C5B575FFB6DF425575D7BEFB55002097555FFD5401EF5D0",
INIT_2D => X"784000AA59000000000000000000000000000000000000000000000208017DAA",
INIT_2E => X"A2D57FFFFF7AEBFF55FF8028A00512EAAB45007FFFF55082EA8AAA087FC2010F",
INIT_2F => X"5512AAAA085D04174100800021FF002EA8BEF5D0428ABA595557555AAFBC2000",
INIT_30 => X"00FF802ABAA04552ABFF597FD74BAF7AAA8B45AAFBD54005D7BD54AAF7800215",
INIT_31 => X"5FFAAFBC0000AF843FF5500003FF55AAFD6AB4551002ABEF0055555550004020",
INIT_32 => X"DEB0A2FD5600051537DE005D557DE005D7BE8AA85555400100879560AA592F95",
INIT_33 => X"17545FFD5421FF5D0428BEF0079FCABA598400010F7AA8215555003FEAAAA843",
INIT_34 => X"0000000004001FFAAFBEAA105D2E955FF557BD75EFFBBCD415521FBFDF450004",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000010000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(0),               -- Port A write enable input
DIA(0)   => data_write_a(4),        -- Port A data input
DOA(0)   => data_read_a_lo_512(4),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(0),               -- Port B write enable input
DIB(0)   => data_write_b(4),        -- Port B data input
DOB(0)   => data_read_b_lo_512(4),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_5_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50DB0A0791B1B41694368283C81F9996A091A32152007AB36B20E03C040C002",
INIT_01 => X"880015C49830884C446A40000C34C24841280A00084000C8C212892EEA953231",
INIT_02 => X"408F417400B1D9100002171C1FA20171124E6AA00D8633F8CD09DBFBBB972F7C",
INIT_03 => X"88538F0182058082D800C3314722DC08A34084A100C4D7C99208521063D00148",
INIT_04 => X"F45E41AFAF420996B8411CA282F80A9091224800A2C61490363080C8A4000308",
INIT_05 => X"0EA416069640420901A01505C4410020C6E228DC30532839B043289D9C005031",
INIT_06 => X"13992D9AF8C74E92B7B568D19708C038AFFA89F0B9348C9204C389672407EF12",
INIT_07 => X"6255000016053C18162589725146F442222CE6AF844012BE795224458BA4DE0F",
INIT_08 => X"4F3F00503B4AE104B5347230418190420821006016FC18843630D285FC416CB4",
INIT_09 => X"EEA33E700340902C4424C442B0344724066C56C2248130A2D9C185B24A24832B",
INIT_0A => X"315325008348CC40AB570500204462508135D5AA593E043731E9B18A98440137",
INIT_0B => X"E0CD463C5813804E0258E0358E02D8E03D8E0258E03D8E02D8E03447012C701E",
INIT_0C => X"F8DE3C27CA181E5D710664A5F140C14BD32A2E281992940AFAA15C3FC0836310",
INIT_0D => X"F000BE0FC80020130841840308653FF0313FE92C23FB1EECB367C0F3E378F0BC",
INIT_0E => X"F000BE0FCD806FFFAF0AE83080E2AEB2F0F1E01BE53FE1F000BE0FC41BE53FE1",
INIT_0F => X"0231F0BF9E3F02A7FFD63669C0E008C3CB7F041BE1BFE1F000BE0FC41BE1BFE1",
INIT_10 => X"30180309A0F83FE2B87C7D006FFF9F1A7806013879BAA78FC103FF5F1F12F038",
INIT_11 => X"39E9C1DBF8A30C2098DBE2FF7F2320483136F200A822CBACAB9DDEB7F9BC291F",
INIT_12 => X"004C72BEC95FEF64E4090626DF15B7D1C6184131B7980DFFFC03F00003F01FB9",
INIT_13 => X"1DFFFA0A3C0202B8776AE7A7C9CBFFF060703080E29F1B79E9F6427EFE901C0E",
INIT_14 => X"2B716CA5C56620590350ACD3A7D5B7EFAC6DFC8C0312A0024B83F07F3999E9F2",
INIT_15 => X"F0BCAF3BC2F3BC6F0BCEF2BC2F3BC6DBC67C251104A2261253904580207E1C81",
INIT_16 => X"1BCEF0BC2F3BC2F1BCEF0BC6F2BC2F1BCAF1BC6F2BC6F2BCAF1BC2F3BC6F2BCE",
INIT_17 => X"BCEF0BC2F3BC2F1BCAF1BCAF3BC6F0BCEF0BCEF2BC6F2BCAF1BCAF1BC2F3BCAF",
INIT_18 => X"69CFEF73B6FFE7436DB6FD0831518424965B4D2492CB69AF1BCEF0BC6F2BC6F0",
INIT_19 => X"F7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF3EF9FBFBB9E79E7BEBCB7",
INIT_1A => X"DEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDF7DF7DF7D",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF29FDAF77BBDDEEF77BBDDEEF77BBD",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"AAA2802AA10FFFFFDE0008556AABA5D2ABFFEFFF800000000000000000000000",
INIT_1F => X"ABAF7AAA8BFFAA802ABFF087FFDF5508003FEBA087FD54BA0804154005555574",
INIT_20 => X"54AAF7D168B45AAAABDF55AA802AA1000003FEBA00002AABA5D2EBFEBAAAD16A",
INIT_21 => X"3DE005555575EFA2D142145A2FFE8B45FF80001555D2E955FFFFD5421EFAAFFD",
INIT_22 => X"FC00BA5D5568AAAF7AAAAAAAAA802AABA082E954005500021FF5D2EBFF550000",
INIT_23 => X"D5420AAAA843DFFFAAD1554005D7FD74AAAA840014500517FFEF007BEABFF5D7",
INIT_24 => X"2AABDE0055517FF555504154BAA2FBEAA105D2E97410FFD16AAAA5D2ABDEBAFF",
INIT_25 => X"000000000000000000000000000000000000000028BFF0855555455500174BAA",
INIT_26 => X"21E84124285C51574BAB68A2DA00FFFFFFE38085F6FA92552AB8FEFF78000000",
INIT_27 => X"925D2AB8EBABEDB6AA92F7AAA8BC7B68A28BC70075FDF45080A3AEAA007BD248",
INIT_28 => X"5FFFFD1471D7AAFBD0492EBD56DB7DBEAEBFF55BE842AA105D0A38EBA1C0428A",
INIT_29 => X"21FF492AB8F7D1C0438E38145B575EFA2DB45145B6F5EFB6DF78E05145552A92",
INIT_2A => X"7DFC70875EABC7557FC20AA415F68AAAF7AAAAA82BE8A28A9214249740041000",
INIT_2B => X"B6FABA542ABAE2AF7DF470AABE8A3AFD7A2DF55400557FD54AABE84001C55551",
INIT_2C => X"5557545490012482B6A0BAE2849043AFED1C0E10492B6FFEFA105D2A95410FFD",
INIT_2D => X"D2AAABEFFB8000000000000000000000000000000000000000000000428BEF00",
INIT_2E => X"082EA8AAA087FC20105504000AA5955554BAFFAEBDE10F7FBFDEBA007BFDE005",
INIT_2F => X"0512AA8AAA5D0028A005D2AA8ABAF7FBE8A00FFAEAAB45F3AAAAB4500557FF55",
INIT_30 => X"EFFFAA97545552A821EFFBD557555AAFBC2000A2D57FFFFF7AEBFF55FF8028A0",
INIT_31 => X"A005D04174100800021FF002EA8BEF5D0428ABA597FD55FFA2FFD5555FFD57FF",
INIT_32 => X"54AAF7800015551517DF45005168B55557FC0012087FEAABAF7AAAAA10F3AAAA",
INIT_33 => X"FFE005D2A95410F7FFFFEBA5D2EA8ABAFBFFD74BAF7AAA8B45AAFBD54005D7BD",
INIT_34 => X"00000000002ABEF005555555000402000FF802AAAA04452ABFF592E80010FFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000060000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(0),               -- Port A write enable input
DIA(0)   => data_write_a(5),        -- Port A data input
DOA(0)   => data_read_a_lo_512(5),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(0),               -- Port B write enable input
DIB(0)   => data_write_b(5),        -- Port B data input
DOB(0)   => data_read_b_lo_512(5),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_6_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10800B0061A01002840002C030028180004003220200403312301C4389B2082",
INIT_01 => X"060009C838394848188160000C42426041000000090800090210090000510200",
INIT_02 => X"00043040009001100000061000018070002408000000000648080000001210E0",
INIT_03 => X"0000800002054081020080801200A0000300008000201184681A0000410C4800",
INIT_04 => X"0808801040000001401048008100022401400002024024053200020089000100",
INIT_05 => X"0240040408402202002000C200400020A50000A0000010010001260808000520",
INIT_06 => X"44000881064500004600000013088002840C240F5048011200010000440C0146",
INIT_07 => X"0241914041FE83E010040110110003040020402A0000003E1000000488000201",
INIT_08 => X"8001BF002C4A01041B112020200110024029006FE09081002004902000012068",
INIT_09 => X"0083FE38A040100281353150ACB645AEF8C01404448000008011061204200108",
INIT_0A => X"3103AD0413424E4014D627C470462200011504420C0A962A2189002881404060",
INIT_0B => X"46C1060C16C96D15B0425B0425B1425B1425B0C25B0C25B1C25B1512D8212D82",
INIT_0C => X"009000140401100601016600A040220203A004480598010248000D0010420C0C",
INIT_0D => X"0000A01033A00013000000000018800F2400091081100C0090A5008200410020",
INIT_0E => X"0000A0103142000000000000000000455D0018100000000000A0103410000000",
INIT_0F => X"000000466800C200000000000000000001A0F4100000000000A0103410000000",
INIT_10 => X"00000000000024094680014200000000000000000041E8002900000000000000",
INIT_11 => X"F000322000000000000D1A000000000000034D240C2000502000000000000000",
INIT_12 => X"000000403F4000000000000068D24000000000001A60F0000000000000002007",
INIT_13 => X"C0000000000000000087C0003014000000000000000025D00008958000000000",
INIT_14 => X"02000000000814C219500150002800101280000000000000000000086670000C",
INIT_15 => X"8120C82208812048120882208892055A0060011280222413130449010301F051",
INIT_16 => X"3200802008320C82200802048320C82200812048320880200812048220880204",
INIT_17 => X"20C83208812048020883204802048120882204812008220C8220081204822088",
INIT_18 => X"79CFF1FE1E9F52ABEF9EFE8150120EC718638E38E30C71C812088220C8120080",
INIT_19 => X"71C71C71C71C71C71C71C71C71C71C71C71C71C71C736D9DBD9BBEFBEFBEBEF1",
INIT_1A => X"CFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FC71C71C71C",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCF29A7F3F9FCFE7F3F9FCFE7F3F9F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000607FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"EFA2FBD54BA5555554BAAAFBC20BA5D7BEAAAAFF800000000000000000000000",
INIT_1F => X"EBA0855421455555574AAA2802AA10FFFFFDE0008556AABA5D2ABFFEFFF843DF",
INIT_20 => X"DF5508003FEBA087FD54BA000415400550428AAAAA84021FF007BD54BAAAD17D",
INIT_21 => X"A8BFFAAD1554BA002A95555A28417400AAFBE8ABAF7FFD54AAAA802ABFF087FF",
INIT_22 => X"BD5545080417555A2D17FE1000003FEBA00002AABA5D2EBFEBAAAD16AABAF7AA",
INIT_23 => X"D5421EFAAFFD54AAF7D168B45AAAABDF55AA802AA100000001EF087FEAA00FFF",
INIT_24 => X"F80001555D2E955FFFF843DEAAA2803DFEF0855401FF082EA8B555D7FC21FFFF",
INIT_25 => X"0000000000000000000000000000000000000055575EFA2D142145A2FFE8B45F",
INIT_26 => X"2552AB8FEFF78E3DFFFAAFFD04AA415B52492B6F5C20825D7FE8A92FF8000000",
INIT_27 => X"EF147BD2482BED57AE921451421555551574BAB68A2DA00FFFFFFE38085F6FA9",
INIT_28 => X"4BAB68A28BC70075FDF45080A3AEAA007BD24821C04124281C0E2DA82BE8E001",
INIT_29 => X"8EBABEDB6AA92F7AAA8BC7B6D5524AA14209557DA28E15400BEF1EFA92FFFFD2",
INIT_2A => X"071FF0071EDA38F7F1D5555000417545B6D178E281C0A38EBA1C0428A925D2AB",
INIT_2B => X"4A8B555C7FC2147F7D1471D7AAFBD0492EBD56DB7DBEAEBFF55BE842AA105D0E",
INIT_2C => X"DB45145B6F5EFB6DF78E05145552A925FFFF8E3DE82BE8E38FFF0851401C7082",
INIT_2D => X"57FE8A00F38000000000000000000000000000000000000000000005B575EFA2",
INIT_2E => X"F7FBFDEBA007BFDE005D2AAABEFFBAABDFEFAAFBC00BA007BC0000FFD5420005",
INIT_2F => X"A592ABFE00F7AA821FF557FC0010F7D168A105D55421455155554BAFFAEBDE10",
INIT_30 => X"10F7D57DE00FFFBC00AAFBAAAAB4500557FF55082EA8AAA087FC20105504000A",
INIT_31 => X"AAA5D0028A005D2AA8ABAF7FBE8A00FFAEAAB45F3D5400BA5504155EFAAAE954",
INIT_32 => X"FF55FF8028A00512E975FF08557FEAAF7D157545080417545F7D56AAAA592AA8",
INIT_33 => X"AABEF005542155000028B555D7FC2145F3D557555AAFBC2000A2D57FFFFF7AEB",
INIT_34 => X"000000007FD55FFA2FFD5555FFD57FFEFFFAA97545552A821EFFBAABDE00F7AA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000048000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(0),               -- Port A write enable input
DIA(0)   => data_write_a(6),        -- Port A data input
DOA(0)   => data_read_a_lo_512(6),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(0),               -- Port B write enable input
DIB(0)   => data_write_b(6),        -- Port B data input
DOB(0)   => data_read_b_lo_512(6),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_7_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10844B00482258A2842112C02450418800002300500030B313300C418992002",
INIT_01 => X"020009C23838684D1C20E0000E11424840000000080000080200000000110204",
INIT_02 => X"000520700CA08910000206101180803081144880010400044808000000122160",
INIT_03 => X"000080040305208000008000328080040304008020303194289A000041484800",
INIT_04 => X"08088000000000010000CA008008060441000000028234493410820191000000",
INIT_05 => X"03500404000022020020044000000C208400408000001000984005949C002928",
INIT_06 => X"54000881044500004680000013008002940C24001A4A010200018920646410C7",
INIT_07 => X"22510040400500011204813015012204002040280000013E1000000488000201",
INIT_08 => X"9001A0602C4A01051B132820208001024069004008908002120851420001226A",
INIT_09 => X"01100020A2401008A20404E08200A05000A4264640800022C8198C4E05200018",
INIT_0A => X"20002000024040400050450440C48A0041140C420B0904208800904286000008",
INIT_0B => X"50822002120D2134800648006480064800648106481064810648193240432404",
INIT_0C => X"284A142288042A5C24202451505E00A621A5220A8091444040188C001B41210A",
INIT_0D => X"00F001F021141A12004104020810B000100000000109064C80010050A3285194",
INIT_0E => X"00F001F027420000400004C3201C514408081C1014800000F001F02810148000",
INIT_0F => X"E00E0E404100E200040900000B0380383480C81014800000F001F02810148000",
INIT_10 => X"4160C0301D07001D0402034200004000019860078641004039000180400002C0",
INIT_11 => X"08103BA0104810C8462416E8040446120C890814600010512000000080028400",
INIT_12 => X"98038D4030DD008088C2419120B740209021908C4846FC000200030F000FE006",
INIT_13 => X"DD000100411C81078884204035DC00201804C3201C60A408100DD58010440130",
INIT_14 => X"412024202211148019064200402A32901A8000B2048902C0807C0E00C448100D",
INIT_15 => X"50942509425194651946519465894619421421102000269243854D8002000250",
INIT_16 => X"19465194E50942509425094E51946519465094A50942509425194E5194651942",
INIT_17 => X"9425094251946539465094250946539465194250942509465194650942509425",
INIT_18 => X"0000000000000000000000080150890820800041041000052942509465194653",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF21E6C000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"AAF7D5575455D557DFEF002AAAB55002E820AAAA800000000000000000000000",
INIT_1F => X"B55007FD74AAAA843DFEFA2FBD54BA5555554BAAAFBC20BA5D7BEAAAAFFFBC00",
INIT_20 => X"AA10FFFFFDE0008556AABA5D2ABFFEFFFAAAAAAAF7D57FFEFF7D555555A2AEAA",
INIT_21 => X"42145552ABDFEFFFAA801EFFFFBFDF550000175555504175450055574AAA2802",
INIT_22 => X"A975EF00003DF55555168A00000428AAAAA84021FF007BD54BAAAD17DEBA0855",
INIT_23 => X"802ABFF087FFDF5508003FEBA087FD54BA000415400557BD74BAFFD140000082",
INIT_24 => X"AFBE8ABAF7FFD54AAAAAEA8ABA55557FEAAA2843FF55A2AEA8B55AAAABDEAAFF",
INIT_25 => X"0000000000000000000000000000000000000051554BA002A95555A28417400A",
INIT_26 => X"25D7FE8A92FFFFC70BAE3D155555415178FD7082EAAB550820870BAAA8000000",
INIT_27 => X"FFEBD55557DBEA4AFB550871D7482AA8E3DFFFAAFFD04AA415B52492B6F5C208",
INIT_28 => X"5550051574BAB68A2DA00FFFFFFE38085F6FA92552AB8FEFF7A0ADABAEBD578F",
INIT_29 => X"2482BED57AE921451421555524BDFD7FFA4801D7F7F5FDF55000E17545410E17",
INIT_2A => X"D2482E3D1450381C20905EF08003AF55415F6DA38080E2DA82BE8E001EF147BD",
INIT_2B => X"AAFB55ABA0BDE02EB8A28BC70075FDF45080A3AEAA007BD24821C04124281C7B",
INIT_2C => X"209557DA28E15400BEF1EFA92FFFFD24BAB6A4A8A82495F78E92AA843DF45BEA",
INIT_2D => X"800174BAA680000000000000000000000000000000000000000000055524AA14",
INIT_2E => X"007BC0000FFD542000557FE8A00F3FFD54BAAAD15754508556AB45002AA8B450",
INIT_2F => X"FFB803DEAAAAD56ABEFAAD5575EFF7803DF45085557410AEAABDFEFAAFBC00BA",
INIT_30 => X"55082E97555002E955550C55554BAFFAEBDE10F7FBFDEBA007BFDE005D2AAABE",
INIT_31 => X"E00F7AA821FF557FC0010F7D168A105D554214551003FF45FF8400145FFD57FF",
INIT_32 => X"20105504000AA597FC2010A2D1554AA5500021EF000028B55087BFDEBA042ABF",
INIT_33 => X"E8A00A2803FF45F7AABDF55AA843FE10AEAAAAB4500557FF55082EA8AAA087FC",
INIT_34 => X"0000000055400BA5504155EFAAAE95410F7D57DE00FFFBC00AAFB8028A00007F",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000007FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(0),               -- Port A write enable input
DIA(0)   => data_write_a(7),        -- Port A data input
DOA(0)   => data_read_a_lo_512(7),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(0),               -- Port B write enable input
DIB(0)   => data_write_b(7),        -- Port B data input
DOB(0)   => data_read_b_lo_512(7),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_8_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000B0000040042840002C0000001800000070000000033022000000000086",
INIT_01 => X"000009C21838284D1C2160000E12426840000000180800080200080040510200",
INIT_02 => X"0001004000900110000006100080003000240800014400004808000000122160",
INIT_03 => X"00008000020440810002A0801010A0044300000000200086011A000040404800",
INIT_04 => X"8000801000020401400040408108022029400000124004041200000089000100",
INIT_05 => X"02080424085022020000040200480020850010A0002010010120060800040400",
INIT_06 => X"50000880006500000680000011008006840C200018C1010200018920E0640102",
INIT_07 => X"426000404005000112048130150120240020400A0000013E1000000488000010",
INIT_08 => X"220100402C42010413110020200100024029004000A200002004902200012141",
INIT_09 => X"0000000080400008010410A2940A45240040140440800022C8388E1200A00008",
INIT_0A => X"00420100020048405000070440C0000001140412090000000021002081000048",
INIT_0B => X"0000000800000100011000010000100001000010000100001000010000880008",
INIT_0C => X"001000040001100008012008004020102180800804802000C0080D00100A0008",
INIT_0D => X"0FF0000002200A1200410402080080003000091085100C008124008000400020",
INIT_0E => X"0FF000000140000040F517CF600000000104081010001E0FF00000001010001E",
INIT_0F => X"E000000000804200000809963F1F80000000001010001E0FF00000001010001E",
INIT_10 => X"CFE7C0F00000000000810140000040E587F9E000000008100900008000ED0FC7",
INIT_11 => X"00021040030C73D80000021000585F3600000020240020102000000802419660",
INIT_12 => X"F80000000042000B0BD6C0000010800618E7B000000C000003F80FFF00000000",
INIT_13 => X"800005D5C3FD800000000008180000078A8FCF600000000002028001006AA3F1",
INIT_14 => X"020000000008808219002100100C000041120370DCAD1FC18000000000000202",
INIT_15 => X"8020080200812048120481204812055A04604930A02026934215410102000110",
INIT_16 => X"0200802008020080200802048120481204812048120481204802008020080200",
INIT_17 => X"2008020081204812048120481200802008020080200802048120481204812048",
INIT_18 => X"414A87D78AF42143CEBAC88151120A0000000000000000081204812008020080",
INIT_19 => X"F3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF7E799B1BEB65B65948051",
INIT_1A => X"C3E9F0FA7C3E9F0FA7C3E9F0FA7C3E9F0F87C3E1F0F87C3E1F0F87CF3CF3CF3C",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF1B5DA9F0FA7C3E9F0FA7C3E9F0FA7",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"0000043DF55087BC01EF007FD75FFFF84000AAFF800000000000000000000000",
INIT_1F => X"E10A28028AAAAAFBC00AAF7D5575455D557DFEF002AAAB55002E820AAAA84000",
INIT_20 => X"54BA5555554BAAAFBC20BA5D7BEAAAAFFAA95545552ABFE00087BC00AA082EBF",
INIT_21 => X"D74AAAAD57FF45002A975FF007BE8BFFA2FBFFFFFAAD5400AAFF843DFEFA2FBD",
INIT_22 => X"BE8A00082A97410F7D5555EFAAAAAAAAAF7D57FFEFF7D555555A2AEAAB55007F",
INIT_23 => X"55574AAA2802AA10FFFFFDE0008556AABA5D2ABFFEFFFAA82000555555545AAF",
INIT_24 => X"00017555550417545000015545087BC2010AAD54014500516ABFFA2AABDF4500",
INIT_25 => X"000000000000000000000000000000000000002ABDFEFFFAA801EFFFFBFDF550",
INIT_26 => X"50820870BAAA8407000140038F450075C71FF087BD75D7FF84050BAEB8000000",
INIT_27 => X"10007FC50BA002ABFE00AA8A2AABABEFFC70BAE3D155555415178FD7082EAAB5",
INIT_28 => X"082EB8E3DFFFAAFFD04AA415B52492B6F5C20825D7FE8A92FFA497545552AB8E",
INIT_29 => X"557DBEA4AFB550871D7482AAD17DF451C24955EF0875EFBD7B6F1FFFC7BEDB45",
INIT_2A => X"87000415B5057DAAFBE8A10082092410EBD5505EFB6A0ADABAEBD578FFFEBD55",
INIT_2B => X"B6ABC7B6AABFFED0051574BAB68A2DA00FFFFFFE38085F6FA92552AB8FEFF7AA",
INIT_2C => X"A4801D7F7F5FDF55000E17545410E17555000E17545007BC0000BED14217D005",
INIT_2D => X"784174AAA280000000000000000000000000000000000000000000024BDFD7FF",
INIT_2E => X"08556AB45002AA8B450800174BAA684174105D042AB550055555FF007BD7555F",
INIT_2F => X"0F384175555D2EA8A00087BD74BA082EBDE10AAAEA8ABAF7FFD54BAAAD157545",
INIT_30 => X"55FFD57DF55FFFBD5400A2AABDFEFAAFBC00BA007BC0000FFD542000557FE8A0",
INIT_31 => X"EAAAAD56ABEFAAD5575EFF7803DF45085557410AED17FF455D04155FF00557DF",
INIT_32 => X"DE005D2AAABEFFBAE97410087BC21EFA2FFEAA00000002010A2D5421FFFF803D",
INIT_33 => X"C0010FFD1401EF087FE8B55FFAEBDFEF0855554BAFFAEBDE10F7FBFDEBA007BF",
INIT_34 => X"00000000003FF45FF8400145FFD57FF55082E97555002E955550C2E95555087B",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000020000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(1),               -- Port A write enable input
DIA(0)   => data_write_a(8),        -- Port A data input
DOA(0)   => data_read_a_lo_512(8),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(1),               -- Port B write enable input
DIB(0)   => data_write_b(8),        -- Port B data input
DOB(0)   => data_read_b_lo_512(8),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_9_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00018248A2840112C00002C18000002300500030B3132000400812002",
INIT_01 => X"A140098218302849180060000C004240413C0A61590001D90213C90008510204",
INIT_02 => X"102008700CB089100002061031285074810448800104008048080080001210E2",
INIT_03 => X"00008015074608840390A0040040800203140000A00010800408108448020042",
INIT_04 => X"082080400004A00100000100840602020100000002C2344156108201811801C0",
INIT_05 => X"0200048480011502049500280020CC2084000080008010019161249C9C002188",
INIT_06 => X"70000881004500004E01020411D08000940C00001800010200018B20206C0102",
INIT_07 => X"EA70C0040005000312048130150100040020404A0000017E10408104C8000110",
INIT_08 => X"000000402C220104131004202081120050A5104000A204617201D10801002000",
INIT_09 => X"000800002F4924003085E51420A0100400641E4E40800022C8088C1220200908",
INIT_0A => X"20102000024040484028450001648C2229150400080244000401900284000440",
INIT_0B => X"0880110901081110411204112040120411204012041120401204111020090208",
INIT_0C => X"685B34A688841A5C21200101A01A0004009024028004044248404D00104B2100",
INIT_0D => X"0000A01000000213000000000000B0001000010000190E44802002D1A168D0B4",
INIT_0E => X"0000A010014000000000000000000040500008100400000000A0100410040000",
INIT_0F => X"0000004608004200040000000000000001A004100080000000A0100410008000",
INIT_10 => X"00000000000024080000014000000000000000000040A0000900010000000000",
INIT_11 => X"300013E010000000000D00F804000000000340000C0000102000000080000000",
INIT_12 => X"00000040091F0000800000006807C000800000001A0CFC000000000000002001",
INIT_13 => X"DD000000000000000082C00019DC002000000000000021500006D58010000000",
INIT_14 => X"03206420000000C019502050000C32901A800080000000000000000860100006",
INIT_15 => X"D1B46D1B46D0B42D0B42D0B42D8B424342342832002A24921082158802001011",
INIT_16 => X"0B42D0B42D0B42D0B42D0B46D1B46D1B46D1B46D1B46D1B46D1B46D1B46D1B46",
INIT_17 => X"B42D0B42D1B46D1B46D1B46D1B46D1B46D1B46D1B46D1B42D0B42D0B42D0B42D",
INIT_18 => X"89999E91BCD1512B871C4A0100000000000000000000000D0B42D0B42D0B42D0",
INIT_19 => X"A28A28A28A28A28A28A28A28A28A29A69A69A69A69A51C200807249041202AE6",
INIT_1A => X"8349A4D068341A0D269341A0D269341A0D068341A0D068341A0D068A28A28A28",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF2DA921A0D269341A0D068349A4D06",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"45A280154BA5555401EFFFD5421EFA2FFFFF555D000000000000000000000000",
INIT_1F => X"5EF00557DF555D040000000043DF55087BC01EF007FD75FFFF84000AAFFD57DF",
INIT_20 => X"75455D557DFEF002AAAB55002E820AAAA843DFEF00517DEBA007BFDFEFFFD157",
INIT_21 => X"28AAAAAAABDF45F7803FFEF555568AAAF7802AA00FFFBD7555087BC00AAF7D55",
INIT_22 => X"BD54BA550417400085155555082A95545552ABFE00087BC00AA082EBFE10A280",
INIT_23 => X"043DFEFA2FBD54BA5555554BAAAFBC20BA5D7BEAAAAFFFBC00AA552E95545087",
INIT_24 => X"2FBFFFFFAAD5400AAFF8402000A2FFFDF555D7BE8BFF5D51575EFA280175555D",
INIT_25 => X"00000000000000000000000000000000000000557FF45002A975FF007BE8BFFA",
INIT_26 => X"7FF84050BAEBDF78F45B68010482415B471C7E3DF451EFBEFBFAF45490000000",
INIT_27 => X"82007FFAFEFE3DB505EF1C5B7AF45490407000140038F450075C71FF087BD75D",
INIT_28 => X"5451C7FC70BAE3D155555415178FD7082EAAB550820870BAAA8438FFF00517DE",
INIT_29 => X"50BA002ABFE00AA8A2AABABEAEB8F45F78A3DFD741516DAAAE38E2DA28EBFFD5",
INIT_2A => X"C20BA5D2E905550071D54825D0A1543808515756D1C2497545552AB8E10007FC",
INIT_2B => X"5505FFBE801256D490E3DFFFAAFFD04AA415B52492B6F5C20825D7FE8A92FFFF",
INIT_2C => X"24955EF0875EFBD7B6F1FFFC7BEDB45082EB8002000AAFFFDF6D417FEABEF5D5",
INIT_2D => X"7FBE8B5500000000000000000000000000000000000000000000000517DF451C",
INIT_2E => X"0055555FF007BD7555F784174AAA2FBEAB45F78402010007BD5545AAFFD55EFF",
INIT_2F => X"AA68028BEF00517FE10007BE8BFFAAFFC01FF557FE8B550004174105D042AB55",
INIT_30 => X"AAAAAEBFEAAAAFFD5545557FD54BAAAD15754508556AB45002AA8B450800174B",
INIT_31 => X"5555D2EA8A00087BD74BA082EBDE10AAAEA8ABAF7AAAAB45F7AEBFF4508557FE",
INIT_32 => X"2000557FE8A00F3FFC00BA552E80145005557400552A954BA0051575EF550417",
INIT_33 => X"FDFFF007FE8BFF5551401EFF784021FF002ABDFEFAAFBC00BA007BC0000FFD54",
INIT_34 => X"00000000517FF455D04155FF00557DF55FFD57DF55FFFBD5400A28400010A2FB",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000040000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(1),               -- Port A write enable input
DIA(0)   => data_write_a(9),        -- Port A data input
DOA(0)   => data_read_a_lo_512(9),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(1),               -- Port B write enable input
DIB(0)   => data_write_b(9),        -- Port B data input
DOB(0)   => data_read_b_lo_512(9),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_10_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00018248A2840112C00002C18000202300500030B3132000400992006",
INIT_01 => X"A140098218302849180060000C00424040000000080000080200090008510204",
INIT_02 => X"102100400C8001100000061000A8503401044880010400004808000000122160",
INIT_03 => X"000080150746088401908000100080020304000020201080001A108448404842",
INIT_04 => X"800080400004A001000040008406020201000000020004401000000180180080",
INIT_05 => X"02000484800133020495040800208C20A4000080000010000001249010042008",
INIT_06 => X"50000881004500004681020411808000940C20001800010200018920206C0102",
INIT_07 => X"024084044005000112048130150120040020400A0000013E10408104C8000010",
INIT_08 => X"000100402C020105131100200000124250A51040088084614001110801012000",
INIT_09 => X"00080082CD09240820800000000000040000180840800022C8088C1220200108",
INIT_0A => X"841201000200484910000F050560262229140402080200A00402000484140400",
INIT_0B => X"0010118900080010000200102001020000200002001020010200001000010008",
INIT_0C => X"408120900404004821202001F05E00040180260A8080044240004C0010800228",
INIT_0D => X"0000A01000000813004104020800800030000800010008088124020102008100",
INIT_0E => X"0000A010014000004000000000000040500008101480000000A0100410148000",
INIT_0F => X"0000004608004200040900000000000001A004101480000000A0100410148000",
INIT_10 => X"00000000000024080000014000004000000000000040A0000900018040000000",
INIT_11 => X"3800100010480000000D00000404400000034000282000102000000080028000",
INIT_12 => X"00000040090000808800000068000020900000001A0000000200000000002001",
INIT_13 => X"80000100000000000082E0001000002018000000000021580000800010440000",
INIT_14 => X"00004000000004C0195000500008000000000082008000000000000860180000",
INIT_15 => X"0100401004010040100401004090055804404110802A24921317580802001011",
INIT_16 => X"0000000000000000000000040100401004010040100401004010040100401004",
INIT_17 => X"0040100400000000000000000000000000000000000000000000000000000000",
INIT_18 => X"215281FC1A72E2486AAA40A85052020000000000000000001004010040100401",
INIT_19 => X"51451451451451451451451451451451451451451452AA83330A8A28A29EA8D1",
INIT_1A => X"5CA6532994CA6532B95CAE572994CA6532994CA6532994CA6532994514514514",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF31CE2E572994CA6532994CAE572B9",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"10AAFBE8AAAA2D540000F7D57DF55A2AABFFEF08000000000000000000000000",
INIT_1F => X"F45FFFBC2010AAD57DF45A280154BA5555401EFFFD5421EFA2FFFFF555D003FE",
INIT_20 => X"DF55087BC01EF007FD75FFFF84000AAFF8002155AAFFE8B45AAD540000087FFD",
INIT_21 => X"7DF555D517FEBA082A801EFF7FBD5400FFD568B555D00155EF08040000000043",
INIT_22 => X"BFDE00A2FBC0145005168A10AA843DFEF00517DEBA007BFDFEFFFD1575EF0055",
INIT_23 => X"7BC00AAF7D5575455D557DFEF002AAAB55002E820AAAA803FEBA082AAAAAAF7F",
INIT_24 => X"7802AA00FFFBD7555082E82155FFAEAAB55AAD568B455D00154BAFFFBD75EF5D",
INIT_25 => X"000000000000000000000000000000000000002ABDF45F7803FFEF555568AAAF",
INIT_26 => X"FBEFBFAF4549003DE10BEF5EDAAAAAD547038EBD57DF7DA2AEB8FC7000000000",
INIT_27 => X"6DAADF470280075FFF45E3F1C7038A2DF78F45B68010482415B471C7E3DF451E",
INIT_28 => X"5C7000407000140038F450075C71FF087BD75D7FF84050BAEB8002155BEF5EDB",
INIT_29 => X"AFEFE3DB505EF1C5B7AF45495B7DEAA0824851EFEBFBD2410EBD168B7D410A17",
INIT_2A => X"38EAA0824A8AAAEBF5FAE28AAF1C2155005F68A10A28438FFF00517DE82007FF",
INIT_2B => X"4104AAF7F1D75EF557FC70BAE3D155555415178FD7082EAAB550820870BAAA80",
INIT_2C => X"8A3DFD741516DAAAE38E2DA28EBFFD55451C2087155EBA4A8B7DAADF68B7D410",
INIT_2D => X"2AEAAB55000000000000000000000000000000000000000000000002EB8F45F7",
INIT_2E => X"007BD5545AAFFD55EFF7FBE8B5500043FE00F7D17FEBAA2D5574BAAAD17DFEFA",
INIT_2F => X"AA28002155FFD17FFFFA2FBD74BA00557FF45A2D5554AAA2FBEAB45F78402010",
INIT_30 => X"00AAD16ABFF002A975450004174105D042AB550055555FF007BD7555F784174A",
INIT_31 => X"BEF00517FE10007BE8BFFAAFFC01FF557FE8B55007FFDEAA0004175FFA2FBC20",
INIT_32 => X"8B450800174BAA68428AAA08042AABAAAD56AABAAAD140155087FEAA10A28028",
INIT_33 => X"2ABEFAAFBE8BFF0004020AAFFD5555EF557FD54BAAAD15754508556AB45002AA",
INIT_34 => X"000000002AAAB45F7AEBFF4508557FEAAAAAEBFEAAAAFFD5545550015555A284",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000047FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(1),               -- Port A write enable input
DIA(0)   => data_write_a(10),        -- Port A data input
DOA(0)   => data_read_a_lo_512(10),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(1),               -- Port B write enable input
DIB(0)   => data_write_b(10),        -- Port B data input
DOB(0)   => data_read_b_lo_512(10),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_11_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10180B05A0010402840602C2D001019000000300000000330A20080EC180002",
INIT_01 => X"AB400984B830084C1820E0000C36424840000000080000088200000802112220",
INIT_02 => X"102A68440080011000000618062AD03502640800010410424908136019920868",
INIT_03 => X"001282118644C88481908001106088022300000080F4925CDC9A10844A9A4842",
INIT_04 => X"401280480004A1011000418084460002E12000000200040010000040A8000000",
INIT_05 => X"0FC8048484011502059511488020802084400888001110000000050000005400",
INIT_06 => X"1011088AE24500001631024511C08004A70AA40008B90D0200018B60A0650D45",
INIT_07 => X"020011005405000910040150110041040024400D800002BE18408104C9205908",
INIT_08 => X"89390040280241041D175820000001020061004004800567403512A801014C46",
INIT_09 => X"050800E20D09A424C5840400808000040680180840800022D8288E946CA00833",
INIT_0A => X"85002000024040410A000D0504408C32E915D9C208050084840201A099100400",
INIT_0B => X"B01011934A005101431CA821CA831CA821CA831CA831CA821CA83165410E5410",
INIT_0C => X"00010080028000010402214850444091019B02080885200042A9CC001000003A",
INIT_0D => X"5A5018C5A0A00812004104020808B00030000808024008008325820000000000",
INIT_0E => X"5A5018C5AB0062C38A4DB680A0D8241500D5761B011986695014A96E1A811986",
INIT_0F => X"42056A289A1BB2078A922DA2A8B180A2600AAE1A811986695014A96E1B011986",
INIT_10 => X"05AA429189B60AC43C6C7F0272C3841DB528802CAB18468F4101621B1BAC8455",
INIT_11 => X"C003104289A668B8CAB270106338317A3D94392020224ACDE215883078681B5C",
INIT_12 => X"804B020A06020C67061BC785938085134CD551BCA1C90006C0C2958502861120",
INIT_13 => X"80819A5539D503336D61056ABA006282806CA64090B89E015AAA880E48382EB8",
INIT_14 => X"40000000E808989003066E03513E41470126C6284B2D20410AB4503089C00A82",
INIT_15 => X"0000000000000000000000000000041800400110200026124202500802000800",
INIT_16 => X"1004010040100401004010000000000000000000000000000000000000000000",
INIT_17 => X"0040100401004010040100401004010040100401004010040100401004010040",
INIT_18 => X"C110083018162148420840280050800000000000000000001004010040100401",
INIT_19 => X"000000000000000000000000000001041041041041003882928E0000000AA0C4",
INIT_1A => X"0000000000008040000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3E0FC000000000000020100000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"EFAA842ABEFA280155EFFFFBC01EF08554000055000000000000000000000000",
INIT_1F => X"F4508514000000003FE10AAFBE8AAAA2D540000F7D57DF55A2AABFFEF0804155",
INIT_20 => X"54BA5555401EFFFD5421EFA2FFFFF555D51575FFA2FFD75FF550015400FFFBFF",
INIT_21 => X"C2010AAD568AAAAAD142145FF80155EF0051555FF0804155FFF7D57DF45A2801",
INIT_22 => X"01540008514215555003DFFFA28002155AAFFE8B45AAD540000087FFDF45FFFB",
INIT_23 => X"040000000043DF55087BC01EF007FD75FFFF84000AAFF802ABFFA2AABFE10080",
INIT_24 => X"FD568B555D00155EF085168B45085142010FFAE800AA5D7BFDF45F7FFEAA0000",
INIT_25 => X"00000000000000000000000000000000000000517FEBA082A801EFF7FBD5400F",
INIT_26 => X"DA2AEB8FC70000175EFB6802DBC7BE8A155EFE3FBC71FF145B42038550000000",
INIT_27 => X"EF550E15400E3F1FFF7D085B420381C003DE10BEF5EDAAAAAD547038EBD57DF7",
INIT_28 => X"5C7F7DF78F45B68010482415B471C7E3DF451EFBEFBFAF45495F575FFBEF5D05",
INIT_29 => X"70280075FFF45E3F1C7038A2DB68ABAB6D145145FF84155D7085B555C7140410",
INIT_2A => X"28BEFBEA4BDE28140A1543800514515549003FFC7BE8002155BEF5EDB6DAADF4",
INIT_2B => X"FFFF7DE3F1EFA10140407000140038F450075C71FF087BD75D7FF84050BAEB84",
INIT_2C => X"24851EFEBFBD2410EBD168B7D410A175C7005B6DB55145140000FFAE85082417",
INIT_2D => X"57BC20AA5D0000000000000000000000000000000000000000000005B7DEAA08",
INIT_2E => X"A2D5574BAAAD17DFEFA2AEAAB550004175FFF7803DF45FFAE955EFAAFBD55EF5",
INIT_2F => X"5007FD75FFF7D5401EF5D2E97410AAD17DFEF007FC20AA5D043FE00F7D17FEBA",
INIT_30 => X"55007FD5545550400145FFFBEAB45F78402010007BD5545AAFFD55EFF7FBE8B5",
INIT_31 => X"155FFD17FFFFA2FBD74BA00557FF45A2D5554AAA2FBEAAAAFFD555545FF80155",
INIT_32 => X"7555F784174AAA2842ABEFFF803DEAA5D2E974AA00515754500003FF55FF8002",
INIT_33 => X"40000FFAE97410007BFFFFFA2D57FE105D04174105D042AB550055555FF007BD",
INIT_34 => X"000000007FFDEAA0004175FFA2FBC2000AAD16ABFF002A97545007FFFF455555",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000040000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(1),               -- Port A write enable input
DIA(0)   => data_write_a(11),        -- Port A data input
DOA(0)   => data_read_a_lo_512(11),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(1),               -- Port B write enable input
DIB(0)   => data_write_b(11),        -- Port B data input
DOB(0)   => data_read_b_lo_512(11),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_12_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50080B01BC002006940202C0DE041196A83183000000023322287E0FC000006",
INIT_01 => X"0E000C068000E04D40238000001702484000000008000008820009280A553231",
INIT_02 => X"400B71440C8001100000171C0283813013766A800586235ECC09C8423B962966",
INIT_03 => X"CC618E048306E082000081000040900003548421A080025EDF08421042DC0108",
INIT_04 => X"00028020000000812000012080080000E100001002000448100000C1BC18008C",
INIT_05 => X"0FF8060610000402010015E100004C2084800090000310000000079010007C19",
INIT_06 => X"33992D98DEC74A003EA468D01510C03E8F580C800A3F018200418927E0668645",
INIT_07 => X"0204000406050013142409121142F746222EE2498000007E111204058B84C50C",
INIT_08 => X"E826A0602902A10491165C200000820018A5104010C01086003C13E000004EDF",
INIT_09 => X"023000000000000867000000000000040000600060801022C9F88D244FA40133",
INIT_0A => X"00100000820040482B28050001600010C13499F01B334015980001E09F000000",
INIT_0B => X"B80460124F16F06BC20CBC30CBC20CBC20CBC30CBC20CBC20CBC3065E1865E10",
INIT_0C => X"00000000029D204B7C0382FD0100F3F9F80FA0200E0BF40063F99C0010000012",
INIT_0D => X"93900F6EE230301208008001007A80001100002002801000A042000000000000",
INIT_0E => X"93900F6EEC421392C96B1237E0D8BD9629F97E0B348EDAC3900F6EFA0B158EDA",
INIT_0F => X"622DBC31D73F6006A5891533EF9500EAE64BCA0B158EDAC3900F6EFA0B348EDA",
INIT_10 => X"C2B083798D341B10DEFE14400392C74CAEAD412EDD2B4FCFF812A383430C669E",
INIT_11 => X"49FAB442994B3238D4E2FB104636652E19B8BA30C022DAD8C100CA39E8CEBE66",
INIT_12 => X"30469392526208C6CC95C33717D88532966471A9C5DD00B12728D5360234D62A",
INIT_13 => X"828C4999AF580395542D27CDBA0020F0FABAC800DA550C29F36A8A2554E48A64",
INIT_14 => X"40000000873FB80B8A00EF03F56CC12B416A51B60585A5C28895962502E9F36A",
INIT_15 => X"0000000000000000000000000000008000000410802A26924010000002000EE0",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"28C1111026C152A121960A884042020000000000000000000000000000000000",
INIT_19 => X"2082082082082082082082082082092492492492492400200005A8A28A200A37",
INIT_1A => X"964B2592C964B2592C964B2592C964B2590C86432190C86432190C8208208208",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF400FEB2592C964B2592C964B2592C",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FF00042ABEFFF8400010082EAABFF55002ABEF08000000000000000000000000",
INIT_1F => X"BEFFFFBD54000004155EFAA842ABEFA280155EFFFFBC01EF0855400005555421",
INIT_20 => X"8AAAA2D540000F7D57DF55A2AABFFEF08556AA10000028AAAFFD15541000002A",
INIT_21 => X"40000005168AAA087BFFFFF5D04001FF00041554555557FE005D003FE10AAFBE",
INIT_22 => X"1555FF082AA8B55F7AEA8BEF5551575FFA2FFD75FF550015400FFFBFFF450851",
INIT_23 => X"D57DF45A280154BA5555401EFFFD5421EFA2FFFFF555D0000145082E955FF085",
INIT_24 => X"051555FF0804155FFF7842AA100000020BAAA801541055042ABEFFFFBD5410AA",
INIT_25 => X"000000000000000000000000000000000000005568AAAAAD142145FF80155EF0",
INIT_26 => X"F145B42038555F401D71C0A2DBC7EB80000280824ADBD7490E28BEF080000000",
INIT_27 => X"82FFDB5243800002FBD7EBFBD24101C00175EFB6802DBC7BE8A155EFE3FBC71F",
INIT_28 => X"E1041003DE10BEF5EDAAAAAD547038EBD57DF7DA2AEB8FC7005F6AA381C0A2DA",
INIT_29 => X"5400E3F1FFF7D085B420381C5B6AA82147FF8FEF410E001FF000E17555555B7A",
INIT_2A => X"0017D142E905EF1451525C7082AADB45F7AEA8BEF555F575FFBEF5D05EF550E1",
INIT_2B => X"02FBEFEBFBD2410AADF78F45B68010482415B471C7E3DF451EFBEFBFAF454900",
INIT_2C => X"D145145FF84155D7085B555C71404105C7F7842FA381C0A00082AA8A10410410",
INIT_2D => X"02AA8BEF000000000000000000000000000000000000000000000005B68ABAB6",
INIT_2E => X"FFAE955EFAAFBD55EF557BC20AA5D7BC01555D2EBFF55A284000AA08003FF550",
INIT_2F => X"5007BE8AAA5D2EBDE00FFFFC00AA08003FF55A2FBC00105D04175FFF7803DF45",
INIT_30 => X"FF082A97555557FE8A0000043FE00F7D17FEBAA2D5574BAAAD17DFEFA2AEAAB5",
INIT_31 => X"5FFF7D5401EF5D2E97410AAD17DFEF007FC20AA5D7BE8A005D7FEABFF002E821",
INIT_32 => X"55EFF7FBE8B550004001FF5D2A801EF5D5142145082EBFF55F7AAAABEF5D7FD7",
INIT_33 => X"82010A2AA8000008043FFFFA2FBC2010A2FBEAB45F78402010007BD5545AAFFD",
INIT_34 => X"000000007BEAAAAFFD555545FF8015555007FD5545550400145FF843DEAA552A",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000007FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(1),               -- Port A write enable input
DIA(0)   => data_write_a(12),        -- Port A data input
DOA(0)   => data_read_a_lo_512(12),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(1),               -- Port B write enable input
DIB(0)   => data_write_b(12),        -- Port B data input
DOB(0)   => data_read_b_lo_512(12),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_13_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10110A0441812402840402822007818000E00700000000330A3000000008042",
INIT_01 => X"A1400986B830E84D182260000C1042484001000008220008A20019080A510200",
INIT_02 => X"10A108600C9141100000C6180CA85035010E4880010431004908135980122D60",
INIT_03 => X"0013881507460886C190832175809C02030400002020124C441A108468424842",
INIT_04 => X"203080680204A0113801D600864E0C96C12000008244244052200201801802C0",
INIT_05 => X"030004849601110204950409C0208C2084E0009C0000100120A00C9918002098",
INIT_06 => X"10000882804544921681428591908000AF28A8002BC00D020003896020658FC4",
INIT_07 => X"CA20400450050009100501501102E0042020448D0000023E10408144C800D800",
INIT_08 => X"1D2B00402B220104B53100200001020218A5104016CC1C616401910801010100",
INIT_09 => X"050800404D49A42EB08000000000000406481C8C408000A2D8088D1820200B00",
INIT_0A => X"0010000002004048AA08050401604462E9144002090740148441200484000500",
INIT_0B => X"000A112100000000010000000001000000000000001000000000000000800000",
INIT_0C => X"509528954404144C200425010040000001B020081094040072005C0030864208",
INIT_0D => X"1C10B3831034081200000000000430003000206822F20CA8826AC2A14250A128",
INIT_0E => X"1C10B383110218CB0E54C2EA404A4F03D404A41AA5B7344C10B383081BA4B734",
INIT_0F => X"8001CE3E20A5B284ED1132909C72885A2B2C381BA4B7344C10B383081AA5B734",
INIT_10 => X"AC3CC0C0B8182597A801610218CB0C3548B3A008E730A01AB113A5524E6ACA67",
INIT_11 => X"A151EC5952E44128CA194517354C180A3C066430202021252991C22C99731014",
INIT_12 => X"1804C8A0ADA2E6A983014780CA28B2A5C8825194332B018A444AEA2701288A15",
INIT_13 => X"02D09852745F80112C428562EE0353635232D50048A411C158BB0A7910142C77",
INIT_14 => X"4240480068001C9B9150A0000297046E4023F8BE8E3E1E0109472C3EB50158BB",
INIT_15 => X"A1284A1284A1284A1284A1284A12851A84284110406A26924302590806000110",
INIT_16 => X"1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284",
INIT_17 => X"284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A",
INIT_18 => X"7DDFE7EFBEFFE7D3EFBEFC48A0550000000000000000000A1284A1284A1284A1",
INIT_19 => X"D75D75D75D75D75D75D75D75D75D75D75D75D75D75D7EFBFBFBBAAAAAABEFDF7",
INIT_1A => X"5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5D75D75D75",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000FEFD7EBF5FAFD7EBF5FAFD7EBF",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"AA5D043FFFFAAAABDEAA557BFDE00FFD140155F7800000000000000000000000",
INIT_1F => X"400AAD540155A2D5421FF00042ABEFFF8400010082EAABFF55002ABEF08556AA",
INIT_20 => X"ABEFA280155EFFFFBC01EF08554000055043DEBAF7843FFFFF7AABDF55A2AA97",
INIT_21 => X"D5400005568A1055043DEBAAAFFE8B45557FD7410552EAAABAAA84155EFAA842",
INIT_22 => X"FE8ABAAA8428A00087BD7555FFD56AA10000028AAAFFD15541000002ABEFFFFB",
INIT_23 => X"803FE10AAFBE8AAAA2D540000F7D57DF55A2AABFFEF085557545FFD17DEBAA2F",
INIT_24 => X"0041554555557FE005D0000155557BEAABA5D2ABDF450851420AA5D7FD5555A2",
INIT_25 => X"000000000000000000000000000000000000005168AAA087BFFFFF5D04001FF0",
INIT_26 => X"7490E28BEF08516DA82410A3FFD7AAA4B8E824971F8E38E3DF45155EB8000000",
INIT_27 => X"D7EBA4BDF45AAAA90410BEDF45155A2DF401D71C0A2DBC7EB80000280824ADBD",
INIT_28 => X"A82B680175EFB6802DBC7BE8A155EFE3FBC71FF145B42038550E38E92EB803FF",
INIT_29 => X"243800002FBD7EBFBD24101C556FA38490A3FE92BEFFEAB45417FD24385D2AAF",
INIT_2A => X"5056DE3D17FE92BEF1EFA92AA8428A10007FD557DFFDF6AA381C0A2DA82FFDB5",
INIT_2B => X"B400925D7FD557DA2803DE10BEF5EDAAAAAD547038EBD57DF7DA2AEB8FC70051",
INIT_2C => X"7FF8FEF410E001FF000E17555555B7AE10410E00155497FEFABA4120B8F55085",
INIT_2D => X"2FBD7545AA8000000000000000000000000000000000000000000005B6AA8214",
INIT_2E => X"A284000AA08003FF55002AA8BEF00517FE00082EBDF45AA8428A10085568ABAA",
INIT_2F => X"A5D2EA8A00A2803DF45AA843DF55AAAE82000F7FBD5545AAFBC01555D2EBFF55",
INIT_30 => X"55087FC00BA552ABFE10F784175FFF7803DF45FFAE955EFAAFBD55EF557BC20A",
INIT_31 => X"AAA5D2EBDE00FFFFC00AA08003FF55A2FBC00105D517FEAA082EBFE10F7FFE8B",
INIT_32 => X"DFEFA2AEAAB550051401FFA2D57FE10F7D57DE00AA842AA00007FD75FFF7FBE8",
INIT_33 => X"FDEAA08042AB45087FC0010557FD55FFAA843FE00F7D17FEBAA2D5574BAAAD17",
INIT_34 => X"000000007BE8A005D7FEABFF002E821FF082A97555557FE8A00002E82155007B",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000067FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(1),               -- Port A write enable input
DIA(0)   => data_write_a(13),        -- Port A data input
DOA(0)   => data_read_a_lo_512(13),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(1),               -- Port B write enable input
DIB(0)   => data_write_b(13),        -- Port B data input
DOB(0)   => data_read_b_lo_512(13),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_14_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10020A000180000284008280000281800000030000000033022000000580002",
INIT_01 => X"A14009821830284D186860000C30C24840000000084000084200090008510200",
INIT_02 => X"102100600C9001100000061020A8503401044880010400204908012018122F64",
INIT_03 => X"00008015074608840190800010008002030400002074F401209A108448404842",
INIT_04 => X"000080400004A00100004000840E000201000000024024401200020180180080",
INIT_05 => X"0A000484800111020495040800208C2084000080000010010020049818002008",
INIT_06 => X"1000088020450402B6A1420511C080008468A80008000D0200018B202067AF10",
INIT_07 => X"422000044005000910040110510260040024400C800000BE3850A144C924080E",
INIT_08 => X"000B004028020104111100200001020210A51040008004616001910801010000",
INIT_09 => X"000800004D492408208000000000000406401C0C40800022C8088DB420200900",
INIT_0A => X"0010000002004048000005040160042229140002090200000401000484000400",
INIT_0B => X"0000110100000000010000100000000000000100000000000000100000000000",
INIT_0C => X"409120940404104C2000210100400000011020080084040040005C0010820208",
INIT_0D => X"E0E0A0000190081200000000000000003000000000100C088020028102408120",
INIT_0E => X"E0E0A0000B02740421A0E5D1A024002050805210040000B0E0A0000210040000",
INIT_0F => X"E01200860008920106460D4501CB000111300210008000B0E0A0000210008000",
INIT_10 => X"0ABBC00905C33C6000400F02740412C0715C40110080A4006110510C14D18178",
INIT_11 => X"20000041DB011CC000090012565306500002411420220080220C0093C3892324",
INIT_12 => X"5809240C09024A4AE0CA00004800839682398000120800658992F3C700C30181",
INIT_13 => X"002B46867DBC002A830280000800F7B7A0B1E240240A8340000200067EAA8CB6",
INIT_14 => X"42004005800004801150A00341244000845C7DB0D0200900422ACA4B28000002",
INIT_15 => X"8120481204812048120481204812051A04204110002A26924302590802000000",
INIT_16 => X"1204812048120481204812048120481204812048120481204812048120481204",
INIT_17 => X"2048120481204812048120481204812048120481204812048120481204812048",
INIT_18 => X"69CB91FE1EF7D3ABEFBECA080050000000000000000000081204812048120481",
INIT_19 => X"F3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF7EFBBBBBF9E79E7BEAAF3",
INIT_1A => X"CFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCF3CF3CF3C",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FF007F3F9FCFE7F3F9FCFE7F3F9F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"45AAD157400007BEAAAAAAAE955555D5568A105D000000000000000000000000",
INIT_1F => X"0AAF784020AAF7D56AAAA5D043FFFFAAAABDEAA557BFDE00FFD140155F7D17DF",
INIT_20 => X"ABEFFF8400010082EAABFF55002ABEF085155400FFD1420100055574AAA2AA80",
INIT_21 => X"40155A28028B550051574005D7FFFE105D7BD7545A284020BA0055421FF00042",
INIT_22 => X"1421FF5D7FFDEBA085168B45FF843DEBAF7843FFFFF7AABDF55A2AA97400AAD5",
INIT_23 => X"04155EFAA842ABEFA280155EFFFFBC01EF08554000055002AB455D5142010085",
INIT_24 => X"57FD7410552EAAABAAA8017400AAD140000002EBFFEFA2AAA8BEFF780021FF55",
INIT_25 => X"000000000000000000000000000000000000005568A1055043DEBAAAFFE8B455",
INIT_26 => X"8E3DF45155EBD17FF6DAADB504001C71EDA82AAA0955455D556DA00490000000",
INIT_27 => X"101C55554AAAAA480082FF84000BAEBD16DA82410A3FFD7AAA4B8E824971F8E3",
INIT_28 => X"092085F401D71C0A2DBC7EB80000280824ADBD7490E28BEF085157428FFDB420",
INIT_29 => X"DF45AAAA90410BEDF45155A28E2AB7D0051504005D71F8E004975D556DB68405",
INIT_2A => X"28B6D5D51420101C5B401EF417BFAEAA08516AB45E38E38E92EB803FFD7EBA4B",
INIT_2B => X"EAFBC7EB80071FF5500175EFB6802DBC7BE8A155EFE3FBC71FF145B420385500",
INIT_2C => X"0A3FE92BEFFEAB45417FD24385D2AAFA82B68015400AADB40000082EBFFC7A2A",
INIT_2D => X"5557FE1000000000000000000000000000000000000000000000000556FA3849",
INIT_2E => X"AA8428A10085568ABAA2FBD7545AAD17DFFFAAFFC200055557DE00A280155455",
INIT_2F => X"F0051554AAFFFFC00105D55554BAA28400000F784020BAAAD17FE00082EBDF45",
INIT_30 => X"000051575FFF78415410087BC01555D2EBFF55A284000AA08003FF55002AA8BE",
INIT_31 => X"A00A2803DF45AA843DF55AAAE82000F7FBD5545AAAEAABFF0051400105D5568A",
INIT_32 => X"55EF557BC20AA5D042ABFF555142000557FC01EF007FEAABA00556AB55A2AEA8",
INIT_33 => X"C0010082EBDF55A2AABDF45A284175FF5D04175FFF7803DF45FFAE955EFAAFBD",
INIT_34 => X"00000000517FEAA082EBFE10F7FFE8B55087FC00BA552ABFE10F78415400A2FB",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000007FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(1),               -- Port A write enable input
DIA(0)   => data_write_a(14),        -- Port A data input
DOA(0)   => data_read_a_lo_512(14),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(1),               -- Port B write enable input
DIB(0)   => data_write_b(14),        -- Port B data input
DOB(0)   => data_read_b_lo_512(14),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_15_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000A000000000284000280000001800020030000000033022000000180002",
INIT_01 => X"A140098018300848180060000C00426040000000080000080200000000110200",
INIT_02 => X"1020004000801110000006100028503400040800010430004808000180120278",
INIT_03 => X"00008011064408840190800000228002A3000000000010000008108448000042",
INIT_04 => X"701280400004A991000000A28406000211000000220004941000000880000000",
INIT_05 => X"02000484800155020495000800218020C4002880005310000000040000000001",
INIT_06 => X"10000880004540000711224491C08000850A880008000D020001892020656300",
INIT_07 => X"8A04000016050009140501505100000420204008000000BE70408104C8000000",
INIT_08 => X"001F004028026104111002200000000200210040008004614001100801010000",
INIT_09 => X"000800000D09240000800000000000040600180840800022C8088C1020200000",
INIT_0A => X"0000000002004040000105000040042229140002080000000400000080000400",
INIT_0B => X"0000110100000000010000100001000010000000000000000000100000800008",
INIT_0C => X"0001008000000000000025000040000001300008009400006200580010000000",
INIT_0D => X"0000000002300012000000000004200030000000000008008020020000000000",
INIT_0E => X"0000000001000000400000000000000000000010108000000000000010108000",
INIT_0F => X"0000000000000200000900000000000000000010140000000000000010140000",
INIT_10 => X"0140000000000000000001000000400000000000000000000100008040000000",
INIT_11 => X"0000004000480000000000100004400000000030002000406000000000068409",
INIT_12 => X"8000000000020080080000000000802010000000000800000201000800000000",
INIT_13 => X"00000100000000000000000008000000184400A0000000000002000000441108",
INIT_14 => X"4000000000000000010620000004000000000242038B82800000000000000002",
INIT_15 => X"0000000000000000000000000000041800000110000024130202500802000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000080050000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"000804154AA5D00001EFF78428AAA007BC2145F7800000000000000000000000",
INIT_1F => X"0AA007FC2000F7D17DF45AAD157400007BEAAAAAAAE955555D5568A105D7FC00",
INIT_20 => X"FFFFAAAABDEAA557BFDE00FFD140155F7FBD74AAAAD17DF45F7D1421EF005540",
INIT_21 => X"020AAF7FFFDF45FF84000BA552ABDFEF08517DF55A2FBEAB555D556AAAA5D043",
INIT_22 => X"FEAB45F7843FF45082A801FF005155400FFD1420100055574AAA2AA800AAF784",
INIT_23 => X"D5421FF00042ABEFFF8400010082EAABFF55002ABEF087BE8ABA555168B55AAF",
INIT_24 => X"D7BD7545A284020BA007FFFE10A284000AA0055401550055574005D2E800AAA2",
INIT_25 => X"000000000000000000000000000000000000000028B550051574005D7FFFE105",
INIT_26 => X"55D556DA004971C7038140012482550E021C7EB8028A821C7BC516DFF8000000",
INIT_27 => X"45E3DF471C70851400BA0071C5028FFD17FF6DAADB504001C71EDA82AAA09554",
INIT_28 => X"B555D516DA82410A3FFD7AAA4B8E824971F8E38E3DF45155EBF1D5492BED17FF",
INIT_29 => X"54AAAAA480082FF84000BAEBF1FFF7DEB8000092552ABFFEF08517DF6DB6FBE8",
INIT_2A => X"EFA8241516DB55A2FFEAB6DEB843DF551C20801C71C5157428FFDB420101C555",
INIT_2B => X"550428412A85082BEDF401D71C0A2DBC7EB80000280824ADBD7490E28BEF087F",
INIT_2C => X"51504005D71F8E004975D556DB68405092087FF8E00BE8A02082005F47145085",
INIT_2D => X"57BD75EFF78000000000000000000000000000000000000000000000E2AB7D00",
INIT_2E => X"55557DE00A2801554555557FE100055554BA5504000105D2A80145AA842AA005",
INIT_2F => X"5AAD557410F7D57DF55AAFBD55450055420BA0055574BAF7D17DFFFAAFFC2000",
INIT_30 => X"FF08517FFFFF7FBEAB455D517FE00082EBDF45AA8428A10085568ABAA2FBD754",
INIT_31 => X"4AAFFFFC00105D55554BAA28400000F784020BAAAD57FFEFA28402010552ABDF",
INIT_32 => X"FF55002AA8BEF007FFDE1000557DF45AAFBE8BEFA2803FF45550400155555155",
INIT_33 => X"80000087BD55450855400BA002A95400F7FBC01555D2EBFF55A284000AA08003",
INIT_34 => X"000000002EAABFF0051400105D5568A000051575FFF78415410087FEAA10F7AE",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000060000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(1),               -- Port A write enable input
DIA(0)   => data_write_a(15),        -- Port A data input
DOA(0)   => data_read_a_lo_512(15),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(1),               -- Port B write enable input
DIB(0)   => data_write_b(15),        -- Port B data input
DOB(0)   => data_read_b_lo_512(15),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_16_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"DA22C618B1000482B688B186588884862A400438255FC38381441205BA803003",
INIT_01 => X"264AC80028404C211203A952A90341080B173340412000E1005D628000820484",
INIT_02 => X"400034C206C405000001A48202084004003008255040826EE008B440200E2042",
INIT_03 => X"2916704900606AC82B49CC56DF8CC1E50E4800202115005760010010000C0400",
INIT_04 => X"052DCA856DC7504B82BF6614C86D2B7F85AAD17F4B100000B88148C4804A428A",
INIT_05 => X"373CB02A00C0502F301180141A42A5720E0F43C17A8479580001AC20000000E2",
INIT_06 => X"303E2094282B85242C85001038D5710E8410D5959BC4800015001219D0550077",
INIT_07 => X"880100000159954501280B0080146F7112D949A0015018220540000382805001",
INIT_08 => X"30015452880C8D90409A05B2CB2CA400200209E5601044A24000000462A60018",
INIT_09 => X"452D54000C0907000330000000000096480050000685400005FC014743E0DC92",
INIT_0A => X"00014808A02004200E540480212000A448C0080024AEA00C9688000000000005",
INIT_0B => X"000D58460018F6D3D84400044000440004400044000440004400042000220002",
INIT_0C => X"0001004010A8812831605DA0000A054052E40000817680220040025699200002",
INIT_0D => X"AAADA0C343F1AC1B01040A002024895514554485D00000012400240000000000",
INIT_0E => X"AAADA0CC421CA003B694B68018FAAA708E2CB5320018CAC99BA0A3B9320018CA",
INIT_0F => X"B1443A1891E4A928C29020E6A8524CE7A3EE59320018CAC99BA0ACB9320018CA",
INIT_10 => X"04B2A5A40B1E6644AF0F021EA003AC24352AB2449A3FF2FA04E5E09B128834AD",
INIT_11 => X"60ED838E890B703C6260D8E3A21275714C902375B801324301AB0067622E5E54",
INIT_12 => X"064F70DBDB1C74424E91E1C194C71D1216F50A8C241815FEB6A9158863F638FB",
INIT_13 => X"45FDF9D364DBD9435A6D45C9E81BED555E4C15F11133D171727A2550EE2F1BA0",
INIT_14 => X"08150013F162119014204373517700ACCC59432A2B2D001F803471A9A960E572",
INIT_15 => X"000000000000000000000000000000880002054000229088542210206B2AB015",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"2A898D21B4C98389ED146C080000000000000000000000000000000000000000",
INIT_19 => X"A29A29A29A29A29A29A29A29A29A28A28A28A28A28A53CBF0F0D3CF3CF0AB1A2",
INIT_1A => X"8F47A3D1E8F4FA7D3E9F4FA7D3E9F4FA7D3E8F4FA3D3E8F4FA3D3E9A29A29A29",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000FA7D3E9F4FA7D1E8F47A3D1E",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFF7FBE8B45AAD568BFFFFAA975FF00003FE0055000000000000000000000000",
INIT_1F => X"0005D2A95410FFFFC00000804154AA5D00001EFF78428AAA007BC2145F7843FF",
INIT_20 => X"7400007BEAAAAAAAE955555D5568A105D2E974BAF7FBEAB45FFFFC00BAF78002",
INIT_21 => X"C2000F78000010552E800AA002E821FFA2AAAAA00000417555FFD17DF45AAD15",
INIT_22 => X"43FEBA5D55575FFF7AABFE00557BD74AAAAD17DF45F7D1421EF0055400AA007F",
INIT_23 => X"D56AAAA5D043FFFFAAAABDEAA557BFDE00FFD140155F7AABDF55F7AE820AA080",
INIT_24 => X"8517DF55A2FBEAB555D04154BAA2FBE8B55FFFFD55FF557FC2000FF8015410FF",
INIT_25 => X"000000000000000000000000000000000000007FFDF45FF84000BA552ABDFEF0",
INIT_26 => X"21C7BC516DFF8438FC7E3F1EAB55B6DF6DBFFF7AA955C71C043FE10490000000",
INIT_27 => X"55FFF1C70BAF78A000005D2097438FFF1C7038140012482550E021C7EB8028A8",
INIT_28 => X"57DEBD17FF6DAADB504001C71EDA82AAA0955455D556DA00492490492F7FBE8B",
INIT_29 => X"71C70851400BA0071C5028FF84020285D2085092002A801FFB6AAA8A10080E17",
INIT_2A => X"BAF6DE3AA8709208043FEBA555B555FFE3AABFE005D71D5492BED17FF45E3DF4",
INIT_2B => X"BC0028E38412428EBD16DA82410A3FFD7AAA4B8E824971F8E38E3DF45155EBA4",
INIT_2C => X"8000092552ABFFEF08517DF6DB6FBE8B555D04124BAB6FBE8B45E3FBD55D7557",
INIT_2D => X"5003DE000000000000000000000000000000000000000000000000071FFF7DEB",
INIT_2E => X"5D2A80145AA842AA00557BD75EFF78428B55AAD168B55F7FFFDFEFFFAA955555",
INIT_2F => X"0000000010F7FBEAB45FFD1554AAFFAE820105500154AAF7D5554BA550400010",
INIT_30 => X"EFF7AEA8A10002E955FFA2D17DFFFAAFFC200055557DE00A2801554555557FE1",
INIT_31 => X"410F7D57DF55AAFBD55450055420BA0055574BAF784000BA5D0017410082E801",
INIT_32 => X"8ABAA2FBD7545AA802ABEFA2AA9541000003DEBA557BD75EFA2AEBDE105D5557",
INIT_33 => X"EAB45AAFFD55555D7FC20AAA280000AAAAD17FE00082EBDF45AA8428A1008556",
INIT_34 => X"00000000557FFEFA28402010552ABDFFF08517FFFFF7FBEAB455D04020AAFFFB",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000020000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(2),               -- Port A write enable input
DIA(0)   => data_write_a(16),        -- Port A data input
DOA(0)   => data_read_a_lo_512(16),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(2),               -- Port B write enable input
DIB(0)   => data_write_b(16),        -- Port B data input
DOB(0)   => data_read_b_lo_512(16),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_17_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"5284CE4FB7BD2C8994A13392DBD02E14006B82AC7E800D44D3DD2FD5F9B961C0",
INIT_01 => X"F9BA301F7E03FC6793F2199B39FC233C11D93AE6F3BB92B32091DBC339B24542",
INIT_02 => X"1D5FC0C08F040404446965C0607FB8A217C400C33A908078551BD04222186338",
INIT_03 => X"A14124C28DFD960832C90446DF8400A5055C25295B695FF97E1B5AC757F06D6B",
INIT_04 => X"04A106866DA3D02A01FB660C08A4AB7F840EDB6F48100DFC8081081D78AC7402",
INIT_05 => X"51E072F0C0C58D9C125EBFC00A46CF0388054100F680E0CE0107B8D040DAFCDA",
INIT_06 => X"019A4D00786B048112C58B16307F15DE8408B233661C10BBA5DAAFA9DDA1194D",
INIT_07 => X"8E00001660700CE170284A00891C7C03D29DE26814515835902AC089A2801540",
INIT_08 => X"C009F3A1B0120A1C51DFF881861CBE0305A12A0321810217C01D34EDC98FFA1C",
INIT_09 => X"747E6610052CDEE97FF1F9F63E3EF790380078002CE976AB6BF769769E4D437D",
INIT_0A => X"00185C44B91BC1740B7605040BE0018CFC7429F326B9D045FF8000E9AB415606",
INIT_0B => X"3A28FC1AAF5CF6F3D3EF3D3EF3D3EF3D3EF3D3EF3D3EF3D3EF3D3EF9E9F79E9E",
INIT_0C => X"0000020012E9E10A31EB5FF9296A67F5B4FFBD2FAD7FE653C3FBFF33E10C001B",
INIT_0D => X"333EA16031F2BD47BDA2CA5D8164FCCFE833C5C3D00018006C68170000000000",
INIT_0E => X"333EA160391BEFF2C32FB695F919110D5ECE542A6FEEB2533EA160782A6FEEB2",
INIT_0F => X"D18C0D06638A207CFDE1F7DDAD76D5282400F82A6FEEB2533EA160782A6FEEB2",
INIT_10 => X"E6E43E59AFE4A59B57679D19EFF2C7573FAD5A86840354D1706FFFA3EF6E24B6",
INIT_11 => X"F7D7A0ABD6DAAAB96529382B74E4E1FE4ACA4D77FAAB77CE3AF3EE78F58DB737",
INIT_12 => X"2D1281017F056E9C9C3FC95949C157ADB55572CA52606DFED6CA55334C04C04F",
INIT_13 => X"59FDEB974F486905001FDF5FA0D719F9956EAA1A184045D5D7A870D2F5A5D752",
INIT_14 => X"60158015177F916A039EF41FDB34A91F432EA58949D5B5C85F97871876F7D7E8",
INIT_15 => X"000000000000000000000000000004DC200005E705B7B3D9FC22F00BE419FB55",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"06013DB9880A5D22E229F3030018000000000000000000000000000000000000",
INIT_19 => X"D35D74D35D74D34D35D74D35D74D34D34D34D34D34D0D30D0D303AEBAE886E40",
INIT_1A => X"51A8D46A351A0D068341A0D068341A0D068341A8D468341A8D46834D35D74D34",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000008D46A351A8D46A351A8D46A3",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFF7FBFDF55A28402000F7D56ABFF55000000000000000000000000",
INIT_1F => X"A00F7843FEBA55043FFFFF7FBE8B45AAD568BFFFFAA975FF00003FE0055043FF",
INIT_20 => X"54AA5D00001EFF78428AAA007BC2145F7D568B45000002010552EBDF45A28028",
INIT_21 => X"95410FFAE800105D2A95410002A95410AAAEBFF55AAFFC00BAF7FFC000008041",
INIT_22 => X"57DE00F7AE800AAAAAABDFEF5D2E974BAF7FBEAB45FFFFC00BAF780020005D2A",
INIT_23 => X"517DF45AAD157400007BEAAAAAAAE955555D5568A105D7FFFFEFA2D568BFFFFD",
INIT_24 => X"2AAAAA00000417555FF8028B55082A974105D003FF55F7802AAAAAAD168AAA5D",
INIT_25 => X"000000000000000000000000000000000000000000010552E800AA002E821FFA",
INIT_26 => X"71C043FE10490A3FFFFFFFFFDFEFE3F5FAF45AA8000038F7DB6FBD7490000000",
INIT_27 => X"384124BFF7DB68A28A38F7803DE82490438FC7E3F1EAB55B6DF6DBFFF7AA955C",
INIT_28 => X"0BAFFF1C7038140012482550E021C7EB8028A821C7BC516DFFDF68B551C0E050",
INIT_29 => X"70BAF78A000005D2097438FFAA85000492495428082E95400AAA0BDF7DB6F5C7",
INIT_2A => X"FAFFFB6D56FBFFEBDB78E38F7AA800BAB6AEBDFD75D2490492F7FBE8B55FFF1C",
INIT_2B => X"028AAAB6D16FA8249517FF6DAADB504001C71EDA82AAA0955455D556DA00497F",
INIT_2C => X"2085092002A801FFB6AAA8A10080E1757DEB8A2DB5514249243841003FF6DEB8",
INIT_2D => X"7FFFDF550000000000000000000000000000000000000000000000004020285D",
INIT_2E => X"F7FFFDFEFFFAA9555555003DE00002ABFFEFF7FBFDFFFAAD168B55AA80000BAF",
INIT_2F => X"FF7FBEAB45552E954BA08003DFFFFFAAA8AAAF7843FE10000428B55AAD168B55",
INIT_30 => X"10AA843FFFFF7D5554BAF7D5554BA5504000105D2A80145AA842AA00557BD75E",
INIT_31 => X"010F7FBEAB45FFD1554AAFFAE820105500154AAF7AE974000800154AA002E954",
INIT_32 => X"554555557FE10007FEABEFFFD57FFEFAAFFE8ABAFFAA820BAF7AEBFF55550000",
INIT_33 => X"020AA08003DFFFA28028AAAF7D17DE0000517DFFFAAFFC200055557DE00A2801",
INIT_34 => X"0000000004000BA5D0017410082E801EFF7AEA8A10002E955FFA2AABFF455500",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000067FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(2),               -- Port A write enable input
DIA(0)   => data_write_a(17),        -- Port A data input
DOA(0)   => data_read_a_lo_512(17),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(2),               -- Port B write enable input
DIB(0)   => data_write_b(17),        -- Port B data input
DOB(0)   => data_read_b_lo_512(17),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_18_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"69844019080000A21A611406840014122A641074155FC28A2024001001801003",
INIT_01 => X"01067920034004180005E9E3C90360C0041C0181002001602025800008440084",
INIT_02 => X"40AC3CAA22D605200000856E2481902400344A20F802C22054001000021E2379",
INIT_03 => X"A95308ECD3207AC81D91C4002004C08A06008080BA868007E58040102B0E0100",
INIT_04 => X"044CC183800CA00780808004C8DB841405A80A100B586200FAC24AE4805242CA",
INIT_05 => X"771C10000000000B1135883C08A115320E0401C0200038394230070A19000020",
INIT_06 => X"3001499C602A8A003E800A042D8132A00098408F79E3901218050018024110D6",
INIT_07 => X"5029401000C983E60004010030400353C05806800104004E0000042E52800E20",
INIT_08 => X"0000117088080990419005B0C309402030060860E01004A828408800440405E3",
INIT_09 => X"6B8186185C42900693A002004040001E1950850C848601008708114A2030B480",
INIT_0A => X"100180A8062026000DC425C0301311324AA237108857220BA089420440000030",
INIT_0B => X"C44703657083080C2800C2000C2000C2000C2000C2000C2000C2000610006100",
INIT_0C => X"C1B0609C05013065CC042004040808084001E000108010230400800FD9B286C4",
INIT_0D => X"CCC15F9CBA45505640000A402019003F140FC2060014250B9080008306C18360",
INIT_0E => X"CCC15F9FB1962FCB69E08AAAEAEBCDDF7C728582081483ACC15F9C3982081483",
INIT_0F => X"EBF1CFFF7670ACC3811A28AB57523CDFEBFBF982081483ACC15F9F3982081483",
INIT_10 => X"C9002BF05800D875E63CC9962FCB52CAA02FE3F8E7F5E3AC3620805298B15A3F",
INIT_11 => X"F1B72A8A800B7546DB9F1CA320037F01BD67DC4041D4CF03138DD865103EFEEA",
INIT_12 => X"81CCFAFDBF9464006FD037AEFAE5150016EA8DB7BFE25208E8F46A228BF8A757",
INIT_13 => X"641256EC844B8AF92FD7CEDC24A9E181A8A29509EAAE7FD3B749471C48F8A459",
INIT_14 => X"0297D086E00036D2440E0880AAD62BEFF5778802A3AF8E8FB0440CE78773B709",
INIT_15 => X"8360D8360D8360D8360D8360D83609220D20D00000080C0601400B402307E480",
INIT_16 => X"360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D",
INIT_17 => X"60D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8",
INIT_18 => X"D9D701DC2E784601EFBE2C00000000000000000000000008360D8360D8360D83",
INIT_19 => X"5155555545145145155555545145145145145145145220B22A0B820820965177",
INIT_1A => X"44A25128944A25128944A25128944A25128944AA552A954A2512895554514514",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000025128944A25128944A251289",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFEFF7AE954BA5D04174AA00000000000000000000000000",
INIT_1F => X"145AA801741000043FFFFFFFFFFFFFF7FBFDF55A28402000F7D56ABFF55043FF",
INIT_20 => X"8B45AAD568BFFFFAA975FF00003FE0055043FFFFFFFFFDFEFA2D56AB45AA8400",
INIT_21 => X"3FEBA55557FFEFA2D168B55AAFBFFFFFFF80021EF0855421EF00043FFFFF7FBE",
INIT_22 => X"A82155F7AEBFEBAFFD56AA00A2D568B45000002010552EBDF45A28028A00F784",
INIT_23 => X"FFC00000804154AA5D00001EFF78428AAA007BC2145F7D5400000004020AA5D2",
INIT_24 => X"AAEBFF55AAFFC00BAF7AE80010082E954BA0004174AAAA8428B45082ABFEBAA2",
INIT_25 => X"000000000000000000000000000000000000002E800105D2A95410002A95410A",
INIT_26 => X"8F7DB6FBD7490E3FFFFFFFFFFFFFFFFBFDFEFFFAE954AA550415492140000000",
INIT_27 => X"D7AAD16FB6DBE8E00155BE8015410140A3FFFFFFFFFDFEFE3F5FAF45AA800003",
INIT_28 => X"1C7140438FC7E3F1EAB55B6DF6DBFFF7AA955C71C043FE1049043FFEFE3F1F8F",
INIT_29 => X"FF7DB68A28A38F7803DE82495B78FC7AAD56FB6DBEF1FAFD7E384001EF145B47",
INIT_2A => X"420381C0A02082492A85155E3A4BDE92FFD56FA28B6DF68B551C0E050384124B",
INIT_2B => X"E28B7D1420BDEAAA2F1C7038140012482550E021C7EB8028A821C7BC516DFFD1",
INIT_2C => X"2495428082E95400AAA0BDF7DB6F5C70BAFFAE870280024904BA1400174AABE8",
INIT_2D => X"50415410550000000000000000000000000000000000000000000002A8500049",
INIT_2E => X"AAD168B55AA80000BAF7FFFDF55002ABFFFFFFFFFFFEFF7FBFDFFFF7AA974BA5",
INIT_2F => X"000043DFEFA2D56AB45AAD57DFEFF7AA82155F78015400552ABFFEFF7FBFDFFF",
INIT_30 => X"55A280021EF557FD7555550428B55AAD168B55F7FFFDFEFFFAA9555555003DE0",
INIT_31 => X"B45552E954BA08003DFFFFFAAA8AAAF7843FE10007FEAB55A2D17FFEFFFD568B",
INIT_32 => X"AA00557BD75EFF7D1400AA5D2A82000002A95545A2843FE00F7D17FEAAF7FBEA",
INIT_33 => X"020AA5D04154BAF7AEA8BEF55003DEAAA2D5554BA5504000105D2A80145AA842",
INIT_34 => X"000000002E974000800154AA002E95410AA843FFFFF7D5554BAF7AE974BA0004",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000020000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(2),               -- Port A write enable input
DIA(0)   => data_write_a(18),        -- Port A data input
DOA(0)   => data_read_a_lo_512(18),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(2),               -- Port B write enable input
DIB(0)   => data_write_b(18),        -- Port B data input
DOB(0)   => data_read_b_lo_512(18),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_19_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"042200000000000041088001001AA00000000000000000000000500802000003",
INIT_01 => X"074018000024000000000404000000000A22000800000800004A200000000001",
INIT_02 => X"0000048002C405000000000006A84000000000200893C246A20000000020031A",
INIT_03 => X"020A9639044012C80001C4000004C08006000000001025000000000000000000",
INIT_04 => X"0400C0800000000380800004C8000000058800000B1000009880480480024200",
INIT_05 => X"420410000000000B10804004080001320E0401C0200038080000000000000000",
INIT_06 => X"2002409006F00A8428050A000280493104004500480090080A01120220140020",
INIT_07 => X"0000000000418026090240923240002190400000000000C0054A912054004021",
INIT_08 => X"0000115080000990000000B0C308000000000860200160000000000038380000",
INIT_09 => X"8000F80001012590001000000000001618000000020280008180810200000000",
INIT_0A => X"0000000000000000000000000000000100008000110000000000000000000017",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000840007600000000000000000800259000000",
INIT_0D => X"0008A0034078104B41A41000000000031400C002000000000000000000000000",
INIT_0E => X"0008A0004263C0343EDD414004042228DC0D385598035D0008A003B05598035D",
INIT_0F => X"040231068187C39F5A4F985C008902041124505598035D0008A000B05598035D",
INIT_10 => X"1BFBD406451B02000E033263C0343CB740500401180DE053A98F6ECC739D8140",
INIT_11 => X"420851546B2400000040D8549B5800000010227848D4303807FC8CC5508AEAED",
INIT_12 => X"52210402120A936B0000000004C2A8D6480000000018A700FCF980CC300318A2",
INIT_13 => X"B1427ED430B41402D025082359700181C21140E40511802208D6B30C48F8A8A4",
INIT_14 => X"9C000018440021011821B35254E99AF9E9410006362A2B6424287B08286208D6",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000023006000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"7747E18E0218CC18E88324000000000000000000000000000000000000000000",
INIT_19 => X"34C30C30C30C30D34C30C30C30C30C30C30C30C30C3504118982A69A6980E411",
INIT_1A => X"C26130984C26130984C26130984C261309A4D26130984C26130984C30C30C30D",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000130984C26130984C26130984",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAA954BA5500020BA5D000000000000000000000000",
INIT_1F => X"4BA5D517FFFF08043FFFFFFFFFFFFFFFFFFFFEFF7AE954BA5D04174AA007BFFF",
INIT_20 => X"FFFFF7FBFDF55A28402000F7D56ABFF557BFFFFFFFFFFFFFFFFFBFDFEFFFAA97",
INIT_21 => X"17410007BFFFFFFFFFFFFEFF7D16AB45AA8002000F7D5575455D043FFFFFFFFF",
INIT_22 => X"568B55F7AE955FFAA840201008043FFFFFFFFFDFEFA2D56AB45AA8400145AA80",
INIT_23 => X"043FFFFF7FBE8B45AAD568BFFFFAA975FF00003FE00557BFFFFFFFFBFDF45AAD",
INIT_24 => X"F80021EF0855421EF002ABFFEFF7D168B55AAD17FFEFF7AE975FF00557FFFF5D",
INIT_25 => X"00000000000000000000000000000000000000557FFEFA2D168B55AAFBFFFFFF",
INIT_26 => X"A5504154921471FFFFFFFFFFFFFFFFFFFFFFFF7AA954BA550000082550000000",
INIT_27 => X"EFF7FBFAFD7E3A4954BA555B7AFC7080E3FFFFFFFFFFFFFFFFBFDFEFFFAE954A",
INIT_28 => X"545550A3FFFFFFFFFDFEFE3F5FAF45AA8000038F7DB6FBD74975FFFFFFFFFFFF",
INIT_29 => X"FB6DBE8E00155BE8015410147FFFFFFF7FBF8FC7EBD568B55A28000000FFDF52",
INIT_2A => X"FDFC7E3F1FAF55A2DB6FB7DF7AE955C7BE800000008043FFEFE3F1F8FD7AAD16",
INIT_2B => X"0955FF145B7AFC7410438FC7E3F1EAB55B6DF6DBFFF7AA955C71C043FE10497B",
INIT_2C => X"D56FB6DBEF1FAFD7E384001EF145B471C71424B8FC7E3D56AB6DB6DF7AFC7EBA",
INIT_2D => X"50002000550000000000000000000000000000000000000000000005B78FC7AA",
INIT_2E => X"F7FBFDFFFF7AA974BA55041541055517FFFFFFFFFFFFFFFFFFFFEFF7AA974AA5",
INIT_2F => X"500517FFFFFFFBFDFEFFFFFEAB45AA80154AA557BEAB45002ABFFFFFFFFFFFEF",
INIT_30 => X"55A28002000F7FFC2155552ABFFEFF7FBFDFFFAAD168B55AA80000BAF7FFFDF5",
INIT_31 => X"FEFA2D56AB45AAD57DFEFF7AA82155F78015400557BFDFEFF7FBEAB55A2D56AB",
INIT_32 => X"555555003DE00007FFDF45AAD568B45AAFBFFFFFFFAA95545F7840201000043D",
INIT_33 => X"6ABFFFFFBEAB45A280155EF557FE8B55000428B55AAD168B55F7FFFDFEFFFAA9",
INIT_34 => X"000000007FEAB55A2D17FFEFFFD568B55A280021EF557FD755555042AB55AAD1",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000040000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(2),               -- Port A write enable input
DIA(0)   => data_write_a(19),        -- Port A data input
DOA(0)   => data_read_a_lo_512(19),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(2),               -- Port B write enable input
DIB(0)   => data_write_b(19),        -- Port B data input
DOB(0)   => data_read_b_lo_512(19),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_20_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000003",
INIT_01 => X"A65FF80000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000048002CC070000000000000000000000002FF86100200000000220002362",
INIT_03 => X"00000000000203D80025DC18004DC3D01E000000000000000000000000000000",
INIT_04 => X"07E5DF808071026F87C4191DD8005080679800000F300002998058068002C000",
INIT_05 => X"C205F23A2100557F70000004390021F61E1E87C3FD0CFBF80880072042000044",
INIT_06 => X"1209244C2000100006800000020010000008407FC800B0000000100600040000",
INIT_07 => X"8802000009FFBFE51886018002040020000800000554003E0000000002800000",
INIT_08 => X"30801F5780259FB0000000F7DF78020004011FEFE00000000020031502000083",
INIT_09 => X"00000000001000000000000000000056F8000001000000040000040141800802",
INIT_0A => X"0000000000000008000800000000000000000000000000000010010014800000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"00010240001721214E000004000000080000008000001000040080FFDB000000",
INIT_0D => X"0000000F3008001E00000000001803FF14FFC006000000008010200000000000",
INIT_0E => X"0000000F3040200000020000000026A70C0008020000200000000F3002000020",
INIT_0F => X"000030B86000400080000200000000004A58F0020000200000000F3002000020",
INIT_10 => X"0000000002183E61E6000040200001000000000019B140000800800000020000",
INIT_11 => X"C00010080000000000525801000000000014AC08000000508001030A0A400100",
INIT_12 => X"000002BC360020000000000292C0100000000000A56000090100000000001F86",
INIT_13 => X"8010000000000000574500001001060600000000001716800000803102020000",
INIT_14 => X"00000000000040040040002000080506049CDF70C08040100000706707600000",
INIT_15 => X"00000000000000000000000000802040200200604040000000000024FB7FE008",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"060070400020112240209A408004000000000000000000000000000000000000",
INIT_19 => X"65965965965965965965965965965861861861861860D30424343CF3CF340E00",
INIT_1A => X"90C86432190C86432190C86432190C86432190C86432190C8643219659659659",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000086432190C86432190C864321",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974AA55040201008000000000000000000000000",
INIT_1F => X"4AA550002000007BFFFFFFFFFFFFFFFFFFFFFFFFFAA954BA5500020BA5D7FFFF",
INIT_20 => X"FFFFFFFFFFFEFF7AE954BA5D04174AA00003FFFFFFFFFFFFFFFFFFFFFFF7AA97",
INIT_21 => X"7FFFF087FFFFFFFFFFFFFFFFFFFFDFEFFFAE974AA5D003FE005D043FFFFFFFFF",
INIT_22 => X"BFDFFFAA84000105D556AB55557BFFFFFFFFFFFFFFFFFBFDFEFFFAA974BA5D51",
INIT_23 => X"043FFFFFFFFFFFFFF7FBFDF55A28402000F7D56ABFF55003FFFFFFFFFFFFFF7F",
INIT_24 => X"A8002000F7D5575455D2EBFFFFFFFFFFFEFF7FBEAB55A28000010F7D16ABEF08",
INIT_25 => X"000000000000000000000000000000000000007BFFFFFFFFFFFFEFF7D16AB45A",
INIT_26 => X"A550000082557FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550400028000000000",
INIT_27 => X"FFFFFFFDFEFF7AE974BA5500050380071FFFFFFFFFFFFFFFFFFFFFFFF7AA954B",
INIT_28 => X"E285D0E3FFFFFFFFFFFFFFFFBFDFEFFFAE954AA55041549214043FFFFFFFFFFF",
INIT_29 => X"AFD7E3A4954BA555B7AFC70871FFFFFFFFFFFFFFF7FBFDFFFFFAA974BA550038",
INIT_2A => X"3FFFFFFFFFDFEFF7F1FAFC7A28002028555F6FB7D5D75FFFFFFFFFFFFEFF7FBF",
INIT_2B => X"402010FFDB6ABEF140A3FFFFFFFFFDFEFE3F5FAF45AA8000038F7DB6FBD7490E",
INIT_2C => X"FBF8FC7EBD568B55A28000000FFDF525455524BFFFFFFFBFDFC7E3F5E8B45A28",
INIT_2D => X"504000BA080000000000000000000000000000000000000000000007FFFFFFF7",
INIT_2E => X"FFFFFFFEFF7AA974AA550002000557FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5",
INIT_2F => X"055043FFFFFFFFFFFFFF7FBFDFEFFFAE954BA5500174AA08517FFFFFFFFFFFFF",
INIT_30 => X"EFF7AE974AA550028AAA5D2ABFFFFFFFFFFFEFF7FBFDFFFF7AA974BA55041541",
INIT_31 => X"FFFFFFBFDFEFFFFFEAB45AA80154AA557BEAB4500557FFFFFFFFFDFEFF7FFFFF",
INIT_32 => X"00BAF7FFFDF55002EBFFFFF7FBFDFEFFFD568B55A284020BA557FFFFFF5D517F",
INIT_33 => X"FFF55A2D16AB45AA8402000F7FBEABEF5D2ABFFEFF7FBFDFFFAAD168B55AA800",
INIT_34 => X"000000007BFDFEFF7FBEAB55A2D56AB55A28002000F7FFC215555043DFEFF7FB",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000007FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(2),               -- Port A write enable input
DIA(0)   => data_write_a(20),        -- Port A data input
DOA(0)   => data_read_a_lo_512(20),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(2),               -- Port B write enable input
DIB(0)   => data_write_b(20),        -- Port B data input
DOB(0)   => data_read_b_lo_512(20),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_21_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"4A302428B824900A128C090A5C1800261500213C005FE812D10420054085A202",
INIT_01 => X"081FFE3440B609703B0427F801A40B8115BC4F655300340288A40D30040E4DD8",
INIT_02 => X"04CA478082CC1740002019824E0203100640303FF8C0B31061096E21A1840814",
INIT_03 => X"230CA7A4810083F80095DE00102DC3823EA821094EC68248923200013290C800",
INIT_04 => X"07CFFFC04904AA7F8780409DF84A0202879800000F3000029980780EA2C3C002",
INIT_05 => X"DE87F0280000407FF900D914382091FE1E1C0FC3E01EFFF8000480200008D062",
INIT_06 => X"010E2182002BC107A03448808F0D7C002822987FC830F40134CC74D002016612",
INIT_07 => X"0401000011FBFFE00520000200422033025C4209104500000012004C004D8C0B",
INIT_08 => X"00EF1F5FA0041FF080AC70FFDF78220010841EFFE7116E144071268DFD3E4C24",
INIT_09 => X"FC8BFE18008083B4443151462A28C6DFF80010002605302248088950484550A3",
INIT_0A => X"10018C241102068006C620C03882019480E631A0855E924E2598038938404037",
INIT_0B => X"A641165448C80C103648A3648A3648A3648A3648A3648A3648A366451B2451B2",
INIT_0C => X"011100841200D001000624000100C002804A08221890004806A310FFDF000454",
INIT_0D => X"5004D8158809C86065941840B1014FFF56FFC0281280080180B2948004400220",
INIT_0E => X"5004D815810D42E04A08A80098C02450025360694101816002D41A4068C10181",
INIT_0F => X"134160C8125B0B271802242880A04482418A0068C101816002D41A4069410181",
INIT_10 => X"10080E05C0B06AA8B12CFD0D42E0441A300012682960828F05C96A001B029010",
INIT_11 => X"00010362A8A20826A88660D86B202049F115100920C54E8EA256ECF078BA081C",
INIT_12 => X"064802C0081B0D64040936443306C55144104F30A8801406D002900062803201",
INIT_13 => X"4581BA0038005A706680012280506A8010602011819E290048A2118EC8140C08",
INIT_14 => X"CC158092C044600466208CC5091011C322A4C40A0300600C0A80509F41800880",
INIT_15 => X"80200802008020080200802008020412002001000000381C02004000FBFFF80D",
INIT_16 => X"0200802008020080200802008020080200802008020080200802008020080200",
INIT_17 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_18 => X"FDDFEFFFBEFFE7C7BFBEFC000000000000000000000000080200802008020080",
INIT_19 => X"F7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7FFBFBFFF9E79E7FFFDF3",
INIT_1A => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFDFEFF7FBFDFEFF7FBFDF7DF7DF7D",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00001FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D000200008000000000000000000000000",
INIT_1F => X"4AA5D00020AA5D7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550402010087FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAA954BA5500020BA5D7FFFFFFFFFFFFFFFFFFFFFFFFFFAE95",
INIT_21 => X"0200000003FFFFFFFFFFFFFFFFFFFFFFF7AA974BA5D0402000557BFFFFFFFFFF",
INIT_22 => X"FFFFEFF7AE974BA5D00174BA00003FFFFFFFFFFFFFFFFFFFFFFF7AA974AA5500",
INIT_23 => X"043FFFFFFFFFFFFFFFFFFFFEFF7AE954BA5D04174AA00003FFFFFFFFFFFFFFFF",
INIT_24 => X"FAE974AA5D003FE005D2EBFFFFFFFFFFFFFFFFFFDFEFF7AE954AA5500174BA5D",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFDFEFF",
INIT_26 => X"A550400028007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0000010000000000",
INIT_27 => X"FFFFFFFFFFFFFAA954BA5D00000BA557FFFFFFFFFFFFFFFFFFFFFFFFFFAE974A",
INIT_28 => X"0005571FFFFFFFFFFFFFFFFFFFFFFFF7AA954BA550000082557BFFFFFFFFFFFF",
INIT_29 => X"DFEFF7AE974BA55000503800003FFFFFFFFFFFFFFFFFFFFEFF7AA974AA5D0405",
INIT_2A => X"3FFFFFFFFFFFFFFFFFFDFEFF7AE954BA5D00154AA00043FFFFFFFFFFFFFFFFFF",
INIT_2B => X"A974BA5D00104925D0E3FFFFFFFFFFFFFFFFBFDFEFFFAE954AA550415492140E",
INIT_2C => X"FFFFFFFF7FBFDFFFFFAA974BA550038E285D2ABFFFFFFFFFFFFFFFFBFDFEFFFA",
INIT_2D => X"D00000100000000000000000000000000000000000000000000000071FFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE954AA5504000BA087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0557BFFFFFFFFFFFFFFFFFFFFFFFF7AA954BA5D00000BA5D7FFFFFFFFFFFFFFF",
INIT_30 => X"EFF7AE954AA5D041740055517FFFFFFFFFFFFFFFFFFFFEFF7AA974AA55000200",
INIT_31 => X"FFFFFFFFFFFFF7FBFDFEFFFAE954BA5500174AA08043FFFFFFFFFFFFFFFFBFDF",
INIT_32 => X"74BA550415410552ABFFFFFFFFFFFFFF7FBFDFFFFFAA974AA5D00174BA08043F",
INIT_33 => X"FDFEFF7FBFFFFFF7AE954BA5D0000010552ABFFFFFFFFFFFEFF7FBFDFFFF7AA9",
INIT_34 => X"00000000557FFFFFFFFFDFEFF7FFFFFEFF7AE974AA550028AAA5D2EBFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(2),               -- Port A write enable input
DIA(0)   => data_write_a(21),        -- Port A data input
DOA(0)   => data_read_a_lo_512(21),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(2),               -- Port B write enable input
DIB(0)   => data_write_b(21),        -- Port B data input
DOB(0)   => data_read_b_lo_512(21),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_22_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"5290F4CDE914905A14A43D33F488243E17122300F55FEB189B343A1140548380",
INIT_01 => X"A94007B259F6A975386262000C344BA9573C6FF57B18A5FB0ABFCD3C2C5F4F0C",
INIT_02 => X"D56B4302AC01005111011BD506AA5205274056900596A539584E2E6DFE4B2418",
INIT_03 => X"9AC0FCBD854688207C90007A1000047A00E588632CA213C8903AD6B55AD0EB5A",
INIT_04 => X"30002047A6FCA110086C402022F2124A8022492580040440002021C922D9109B",
INIT_05 => X"14A206B6838151008D95DD1847811C08002380041F1104002205AC4140DAD060",
INIT_06 => X"1727FF2EB9EF113A10BD32F44289D1F840C1710010344DB9A808FDFF3DE03130",
INIT_07 => X"050700154A00401D00495A06A8D464C5F6B54AA8551040818F4C997AC80CBE05",
INIT_08 => X"0141008801018040E48D50080002B00A0C00801014541E9504703680017F6CB4",
INIT_09 => X"02680000010937986481514E2A29CE010708C0804C6A033F7FCFF9426A41F1AB",
INIT_0A => X"00500001840000C80B410014088040F4A944B1AA313C004554002381B8000500",
INIT_0B => X"A004D1594832824A070AA070AA070AA070AA070AA070AA070AA0725503855038",
INIT_0C => X"501428054278142151262CA50343854E506A2C6898B2950AA6A35B0004284058",
INIT_0D => X"90078E1F840A2B0114020104022460002200050F60E220A06880D2A14050A028",
INIT_0E => X"90078E1F891C239F8908003099C1ACF06273612B3482C0C0078E1F412B1582C0",
INIT_0F => X"1BA1B0FD16770236A4091621C08055C2C0DB012B1582C0C0078E1F412B3482C0",
INIT_10 => X"00101F09C030AB28B03C111C239F870828041BA859F213AFC14AA38043006018",
INIT_11 => X"10E8822A984B0025B0DE6089462660095337B08AA600CA88B143AB11880C2806",
INIT_12 => X"055412D4481128C4CC012A66F304553096004B61BD8068B92400D0004E303689",
INIT_13 => X"589C48082C006A9057CA4385809520F07830001AC2173B00E162563454C40804",
INIT_14 => X"00460848952220592745AC11A544B1BF006850840180A00E1C81900C4190E160",
INIT_15 => X"22088220882208822088220882208CD888088D940D2A3A9D5002001300800C8C",
INIT_16 => X"0080200882208822088220882208822088220882208822088220882208822088",
INIT_17 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_18 => X"FBDFD1FE3EFBD7BBEFBEFA0A245120000000007FFFFFFFF20080200802008020",
INIT_19 => X"F3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF7FFBFAFBBBEFBEFBEFBF7",
INIT_1A => X"CFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCF3CF3CF3C",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000007F3F9FCFE7F3F9FCFE7F3F9F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040000000000000000000000000000000",
INIT_1F => X"4BA550000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0002000087FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974AA550402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"020AA5D7FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5D00000AA007FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAA954BA5504000AA557FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5D00",
INIT_23 => X"7BFFFFFFFFFFFFFFFFFFFFFFFFFAA954BA5500020BA5D7FFFFFFFFFFFFFFFFFF",
INIT_24 => X"7AA974BA5D040200055517FFFFFFFFFFFFFFFFFFFFFFFFAA954BA5500000BA5D",
INIT_25 => X"00000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000080000000",
INIT_27 => X"FFFFFFFFFFFFFAE974AA550002010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"0BA087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550400028007FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAA954BA5D00000BA557FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5D0002",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAA954BA5504020AA5D7BFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"A974AA5D00070925D71FFFFFFFFFFFFFFFFFFFFFFFF7AA954BA5500000825571",
INIT_2C => X"FFFFFFFFFFFFFFEFF7AA974AA5D040500055517FFFFFFFFFFFFFFFFFFFFFFF7A",
INIT_2D => X"D040200008000000000000000000000000000000000000000000000003FFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"A087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550002000087FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAA954AA5D00020AA007FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5504000B",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFF7AA954BA5D00000BA5D7BFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"74AA55000200055517FFFFFFFFFFFFFFFFFFFFEFF7AA974BA5504020BA557BFF",
INIT_33 => X"FFFFFFFFFFDFEFF7AE974AA5D00154105D517FFFFFFFFFFFFFFFFFFFFEFF7AA9",
INIT_34 => X"00000000043FFFFFFFFFFFFFFFFBFDFEFF7AE954AA5D041740055557FFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000007FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(2),               -- Port A write enable input
DIA(0)   => data_write_a(22),        -- Port A data input
DOA(0)   => data_read_a_lo_512(22),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(2),               -- Port B write enable input
DIB(0)   => data_write_b(22),        -- Port B data input
DOB(0)   => data_read_b_lo_512(22),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_23_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"EF20906D902424807BC8241BC81801B97D38AD3C0800103362A6741C80A12A02",
INIT_01 => X"001FFF8409F089003B4422000D80C80106804A7951C5B9D1C828043EA28838F9",
INIT_02 => X"028406A002DC176444683862400003111001303FFC00F240D50146013B300500",
INIT_03 => X"0006C90C010203F80005DC00C52FC380BEAC25886C02034800200200A1008008",
INIT_04 => X"17DFFF8049000BFF878314BFF8488890979800002F702002BB807A068403C280",
INIT_05 => X"DA07F0000000007FF020C814380011FE5E1C2FC3E05FFFF90020000808900010",
INIT_06 => X"10004C9690A8CA008024685184097E81E872C8FFE900FC31348EFDF03BE15E22",
INIT_07 => X"402000001FFBFFFD00080200B8140011F0D8C108155542018D1A302193E94004",
INIT_08 => X"41BE1F5F80003FF0002023FFDF79000000000EFFE309606020008005FC000000",
INIT_09 => X"FC83FE1840C0902400300000000000DFFD4004040C4D32BF7C0EE860003CE680",
INIT_0A => X"10018C24110A860006C620C0312241C482B20420CC56924E2199000C00415037",
INIT_0B => X"4669070510C90C14304043040430404304043040430404304043040218202182",
INIT_0C => X"008000105400C00400100000A018000801000C024000004A940000FFDF820604",
INIT_0D => X"100152100801C17E61841950B1C10FFF57FFC02812F00429DC92C40002000100",
INIT_0E => X"10015210088528E00E02C8200A430A424202A1CAF13F214001521001CBF03F21",
INIT_0F => X"01C1C044006D0C94FB94320880603C420B8001CBF03F214001521001CAF13F21",
INIT_10 => X"30182800A018D9CA8000648528E00D12480202C86040902AC60BACDF0E02D020",
INIT_11 => X"0445C19960A00026880C006739000009B00300010AF5052419D1964419028014",
INIT_12 => X"01844068880CE72000013600600332C140004D101808458A5602E00089202911",
INIT_13 => X"41D0B9023402085020825132C8CB5B4040301009408021144CB042F880100C06",
INIT_14 => X"8E17C0D240406519400500840A9524EE38A1F80E02120018390320F050144CB2",
INIT_15 => X"01004010040100401004010040100100040040000000000001000900FBFFE000",
INIT_16 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_17 => X"0040100401004010040100401004010040100401004010040100401004010040",
INIT_18 => X"0000000000000000000000000000000000000000000000001004010040100401",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000000000000000000000000",
INIT_1F => X"4BA5D0400010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000007FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974BA5D0002000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"00010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA550002000007FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAE974AA550400000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5500",
INIT_23 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550402010087FFFFFFFFFFFFFFFFFF",
INIT_24 => X"FAE954AA5D00000AA007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA55040200008",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010000000000",
INIT_27 => X"FFFFFFFFFFFFFAE974BA5D0400010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0000010007FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAE974AA550002010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA550002",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550400010087FFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"E954AA5D0402038007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550400028007F",
INIT_2C => X"FFFFFFFFFFFFFFFFFFAE954AA5D00020BA087FFFFFFFFFFFFFFFFFFFFFFFFFFA",
INIT_2D => X"D0402010000000000000000000000000000000000000000000000007FFFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000087FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAE974BA550002010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D000001",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFFFAE974AA550002000087FFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"54AA5504000BA087FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA550400010007FFF",
INIT_33 => X"FFFFFFFFFFFFFFFFAA954AA5D04000AA087FFFFFFFFFFFFFFFFFFFFFFFFFFAE9",
INIT_34 => X"000000007BFFFFFFFFFFFFFFFFFFFFFFFFFAA954AA5D00020AA007BFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000007FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(2),               -- Port A write enable input
DIA(0)   => data_write_a(23),        -- Port A data input
DOA(0)   => data_read_a_lo_512(23),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(2),               -- Port B write enable input
DIB(0)   => data_write_b(23),        -- Port B data input
DOB(0)   => data_read_b_lo_512(23),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_24_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100600007FFF000080108004000800020000840041000080808",
INIT_02 => X"0000068002CC07400000090C080002000000103FF811F150231000520ABE4404",
INIT_03 => X"210A0600000203F80005DC00000DC3801EA000000745C4010220000000008000",
INIT_04 => X"07C5FF804900026F8780001DF8000000079800000F300002998078068003C080",
INIT_05 => X"C207F0000000007FF0000004380001FE1E1C07C3E00CFFF80000000000000000",
INIT_06 => X"0002648240F20035A0102000BD0000002802C87FC800FCAA035400001B918600",
INIT_07 => X"0000000001FBFFEC4D2B4AD0B8129063B2CC0000100042018408142F16C01848",
INIT_08 => X"008E1F5F80001FF0000000FFDF78000000000EFFE001600000000005FC000000",
INIT_09 => X"E883FE180000000000300000000000DFFD0000002A80D500000671000004A000",
INIT_0A => X"10018C0411020600048620C030020502000200000400920A2198000800404037",
INIT_0B => X"0641060400C00C00304003040030400304003040030400304003040018200182",
INIT_0C => X"000000001000C00000000000000240058000000000000000000000FFDF000404",
INIT_0D => X"E00880104809C1666594584031010FFF56FFC000104000000010440000000000",
INIT_0E => X"E0088010492064206100E81084200048C0804012500021B00880108012500021",
INIT_0F => X"04100144800803419043064900C0020501840012500021B00880108012500021",
INIT_10 => X"1018140F02C0000809408D206420530270040410004C840041A0D80054109038",
INIT_11 => X"110002C9E8010C00010480B35A0300400041020902F60002260D65B361BAA104",
INIT_12 => X"0228204300166B4060080008240593D0021800020818B06D9802F00030C02060",
INIT_13 => X"143B62023C00142800B04400095DFF90203020042108603100061516EE800C06",
INIT_14 => X"DC1180C7804400044029208301040214AE4C7C02000040206602C10B48110006",
INIT_15 => X"00000000000000000000000000000000000000000000000000000000FBFFE000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"DD5EDCF9822659B6888332000000000000000000000000000000000000000000",
INIT_19 => X"F3CF3CF3CF3CF3DF7DF7DF7DF7DF7DF3DF3DF3DF3DF4D30C2432AEBAEBFE5A15",
INIT_1A => X"C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783DF7DF7DF7C",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000F0783C1E0F0783C1E0F0783",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201008000000000000000000000000",
INIT_1F => X"4BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974BA5D0400000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"00010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000007FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAE974BA5D0000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_23 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0002000087FFFFFFFFFFFFFFFFFF",
INIT_24 => X"FAE974BA550002000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D000200000",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010080000000",
INIT_27 => X"FFFFFFFFFFFFFAE974BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000087FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAE974BA5D0400010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0000010007FFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"E974BA550002000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0000010007F",
INIT_2C => X"FFFFFFFFFFFFFFFFFFAE974BA550002000007FFFFFFFFFFFFFFFFFFFFFFFFFFA",
INIT_2D => X"D0402010080000000000000000000000000000000000000000000007FFFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAE974BA5D0400000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040200",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000087FFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"74BA5D0000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0000010087FFF",
INIT_33 => X"FFFFFFFFFFFFFFFFAE974BA550000010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE9",
INIT_34 => X"000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA550002010087FFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(3),               -- Port A write enable input
DIA(0)   => data_write_a(24),        -- Port A data input
DOA(0)   => data_read_a_lo_512(24),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(3),               -- Port B write enable input
DIB(0)   => data_write_b(24),        -- Port B data input
DOB(0)   => data_read_b_lo_512(24),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_25_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100200002000000080100004000000020000800041000080808",
INIT_02 => X"0000068002CC474000000800000002000000103FFCE302008000000880844A04",
INIT_03 => X"00000040700803FC0105DE00020DC3801EA00000040000000020000000008000",
INIT_04 => X"47C5FFC04904026F8780081DFC040000079C92484F30499299837C168003E400",
INIT_05 => X"C207F0382004407FF0000004382281FF1E1C07C3E00CFFFC090004B05000200A",
INIT_06 => X"1009015C4000000020000000390C10002802C87FC800F8000000000019810600",
INIT_07 => X"0501000001FBFFFD480A0280A816002010800001000054018408102000000002",
INIT_08 => X"0C8E1F5FA21C9FF8004000FFDF7C062031863EFFF75D78004001010DFC000020",
INIT_09 => X"E883FE180C00000000300000000000DFFF00180800000000000660100000A000",
INIT_0A => X"1001DCCC31222730A49620C030020100000200000400921A21D8000804404037",
INIT_0B => X"0641062400C00C00304003040030400304003040030400304003040018200182",
INIT_0C => X"C11160845004D04820000000000000000000000000000000940000FFDF000404",
INIT_0D => X"000800000801C0786184185031810FFF56FFC02812E0182000F2C48304418220",
INIT_0E => X"0008000000002020000008000000000800800002400001000800000002400001",
INIT_0F => X"0000010000000000900000080000000400000002400001000800000002400001",
INIT_10 => X"1000000002002000004000002020000200000000000404000000880000001000",
INIT_11 => X"010000082000000001000001080000000040000100C600800001040000040009",
INIT_12 => X"0000000100002100000000080000104000000002000000081001000000000040",
INIT_13 => X"0010200000000000001004000001080000400080000040010000001080001008",
INIT_14 => X"8C11808200400000400000C20000000420000000030280000000010000010000",
INIT_15 => X"82208822088220882208822088A20C52082081A30080000002005008FBFFF001",
INIT_16 => X"2208822088220882208822088220882208822088220882208822088220882208",
INIT_17 => X"2088220882208822088220882208822088220882208822088220882208822088",
INIT_18 => X"29432D518B45265D82BB4101000005FFFFFFFFFFFFFFFFF82208822088220882",
INIT_19 => X"24924924924924820820820820820820924820924824000A6242B4D34D7F7451",
INIT_1A => X"AC562B158AC562B158AC562B158AC562B1188C46231188C46231189249249249",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000162B158AC562B158AC562B158",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000000000000000000000000",
INIT_1F => X"4BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"02000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAE974BA5D0402000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_23 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000007FFFFFFFFFFFFFFFFFF",
INIT_24 => X"FAE974BA5D0400000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040000008",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010000000000",
INIT_27 => X"FFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAE974BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000007FFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"E974BA5D0400000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000087F",
INIT_2C => X"FFFFFFFFFFFFFFFFFFAE974BA5D0400000007FFFFFFFFFFFFFFFFFFFFFFFFFFA",
INIT_2D => X"D0402010000000000000000000000000000000000000000000000007FFFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"74BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000007FFF",
INIT_33 => X"FFFFFFFFFFFFFFFFAE974BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE9",
INIT_34 => X"000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000007FFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000007FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(3),               -- Port A write enable input
DIA(0)   => data_write_a(25),        -- Port A data input
DOA(0)   => data_read_a_lo_512(25),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(3),               -- Port B write enable input
DIB(0)   => data_write_b(25),        -- Port B data input
DOB(0)   => data_read_b_lo_512(25),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_26_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"E9264EAB20190CA3BA4997AA9002AE9C001006B0778015CFA17E0811039879C7",
INIT_01 => X"F1FFF9BB1F773C7F9BB07DFFFDD863FC5FFF3FEFFBBF9FFB22FFFBC7B9F30686",
INIT_02 => X"9B3184F8AFDEAF300029E4E300FC78A6258548EFFA71C00172082400003A2161",
INIT_03 => X"0084F0FF7FFF1FDD3FEFDCDE981DC3FF5F0D294A7B2B18A0001B9CE6CC606E73",
INIT_04 => X"0FC5DFD7EDFFD66F87FE605DDDBFF3690F9EDB7F5F7AFF639BD7DE37C2FEF591",
INIT_05 => X"F205F0F8E9D199FF76DFEE1C3FCC3FF7BE1FD7C3FFACFBFFDFF7B4FEFFDAA10E",
INIT_06 => X"042648C40179912406C1830639AFBEC14489737FDC00B13BB79DFDB83BF4112A",
INIT_07 => X"763A844769FFBFE4398E4390BB9C28B1D0F049080414583F9468D1AEFC000060",
INIT_08 => X"02C05FD7BC471FBD13D981F7DF7D7E6171AF3FEFE8A3E679FAC1FD1FFFBEB000",
INIT_09 => X"F8CFFE38FF7F6BD928F1ABB47476B5FEF9F59F5FCEEDE73FEE0EFC53B079F5CC",
INIT_0A => X"315BDDCC3B336F7C548667D47B7737AF3FD62601EDC2B66A67B9D60FE4C4427F",
INIT_0B => X"06E19F4DA0E80E903DE3035E3035E3035E3035E3035E3035E3035E981AF181AE",
INIT_0C => X"EBFBF7FEBD66DBFCA3F87501AE7B080607307DCFE1D4077B4D026FFFFBFFAFCD",
INIT_0D => X"0007E010084BCD7FF1B61B5C33813FFFFCFFC7D7D51D6F5FDCB935D7AFEBD7F5",
INIT_0E => X"0007E01001BD8020500008001F010040520201F45EC0010007E01001F45EC001",
INIT_0F => X"1DC0004600400F781429C0080000770001A001F45EC0010007E01001F45EC001",
INIT_10 => X"10003C064000E408010081BD8020600200001EC00040B02007EC09A0E0001000",
INIT_11 => X"360403E434588007200D00F88C84C081C203404B3BFD0402346235408402C080",
INIT_12 => X"07B00040091F1190982038406807C868B1000E401A08FE0012040000FC002001",
INIT_13 => X"7D00212000007C400082D81009FC08281D00001F010021560406758091454000",
INIT_14 => X"FFBFF5FA1040076065F730FC08043A903A80008320C0403C3400008860160406",
INIT_15 => X"D7F5FD7F5FD7F5FD7F5FD7F5FDFF7F7F7F77F9F761FFBFDFFDE5BFFFFF7FF005",
INIT_16 => X"7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5F",
INIT_17 => X"F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD",
INIT_18 => X"B79E923C2CD990AA7F0DDB6B910C8DFFFFFFFFFFFFFFFFFD7F5FD7F5FD7F5FD7",
INIT_19 => X"30C30C30C30C30C30C30C30C30C30C30D34D34C30C35F7AA9ABF0E38E3A8EB62",
INIT_1A => X"C26130984C26130984C26130984C26130984C26130984C26130984C30C30C30C",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000130984C26130984C26130984",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000000000000000000000000",
INIT_1F => X"4BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"02010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_23 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFF",
INIT_24 => X"FAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010000000000",
INIT_27 => X"FFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"E974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007F",
INIT_2C => X"FFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFA",
INIT_2D => X"D0402010000000000000000000000000000000000000000000000007FFFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"74BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFF",
INIT_33 => X"FFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE9",
INIT_34 => X"000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(3),               -- Port A write enable input
DIA(0)   => data_write_a(26),        -- Port A data input
DOA(0)   => data_read_a_lo_512(26),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(3),               -- Port B write enable input
DIB(0)   => data_write_b(26),        -- Port B data input
DOB(0)   => data_read_b_lo_512(26),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_27_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"00080A40000A41248002029000050A088000008242A0004404480002000A1155",
INIT_01 => X"F1FFF1C11F781C129C107DFFFE0860941E81258CA2B71C2220EC1B86E1A00002",
INIT_02 => X"183080988B2EAE00002BE001117C78C6848140CFFA0000800042008000011081",
INIT_03 => X"000000FF7CF91F1D3DEF3CDA881D23FB5C0C21085B0B0820001318C60C204C63",
INIT_04 => X"8FC51FD7EDFDD66E47EE205D1DB7F1490E5EDB7D5CBADB2385D79C3643D4E580",
INIT_05 => X"E001F0C0C991BBFC76DFEA1A3F8C3BC7391F9723FF2CE3FCD6D13096B79C8106",
INIT_06 => X"40000001000000084041830600A40C415004637FC4003021259CFDB01BF80028",
INIT_07 => X"3158954761FA3FE402088220AC1108001080400A400041018468D1A060000050",
INIT_08 => X"02005F0784411E390A4881C7BEFC5F6171CE2F8FE823E778DAC16C1FFBBC9000",
INIT_09 => X"F0C7FEBABF3F6BD108F40E04C0C084F0F8B58B5B8849673F6C0E7A01B00914C4",
INIT_0A => X"B51BFDCC39732F3554866AD57C37BEAF1C152201A4C0B6EA63AAD60B60D4427F",
INIT_0B => X"06F18FC5A0E00F0038D1030D1030D1030D1030D1030D1030D1030F0818688186",
INIT_0C => X"AB6AD7EAB962CBD8A3A83101F47E08040510768EA0C406630D0226FFE375ADE5",
INIT_0D => X"000760000843C561E5C55C42B9011FFF48FFCC57550D63564D1D2556ADAB56D5",
INIT_0E => X"0007600004BD8020100008001F010000130201E44A40010007600005E44A4001",
INIT_0F => X"1DC0000208400D781020C00800007700002005E44A40010007600005E44A4001",
INIT_10 => X"10003C064000C400018080BD8020200200001EC00000382006EC0820A0001000",
INIT_11 => X"3E0403A424108007200102E888808081C20040431BC504021462354004004080",
INIT_12 => X"07B00000015D1110102038400817484821000E400204FE0010040000FC000000",
INIT_13 => X"7D00202000007C400000F81001FC08080500001F0100005E0404758081014000",
INIT_14 => X"8DBBB5FA10400360649310FC08003A903A8000012040403C34000080201E0404",
INIT_15 => X"56D5B56D5B56D5B56D5B56D5B56D7E3D7B57B1C4E17F0944B8D596EEFC7FF001",
INIT_16 => X"6D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B",
INIT_17 => X"D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B5",
INIT_18 => X"2D0200903950C080420948E2D10E8FFFFFFFFFFFFFFFFFF56D5B56D5B56D5B56",
INIT_19 => X"00000000000000000000000000000104000000000004000E5E420000002921C4",
INIT_1A => X"28140A05028140A05028140A05028140A0100804020100804020100000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000140A05028140A05028140A050",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000000000000000000000000",
INIT_1F => X"4BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_23 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFF",
INIT_24 => X"FAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201008",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010000000000",
INIT_27 => X"FFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"E974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087F",
INIT_2C => X"FFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFA",
INIT_2D => X"D0402010000000000000000000000000000000000000000000000007FFFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"74BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFF",
INIT_33 => X"FFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE9",
INIT_34 => X"000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000007FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(3),               -- Port A write enable input
DIA(0)   => data_write_a(27),        -- Port A data input
DOA(0)   => data_read_a_lo_512(27),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(3),               -- Port B write enable input
DIB(0)   => data_write_b(27),        -- Port B data input
DOB(0)   => data_read_b_lo_512(27),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_28_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"02200AA400180030808802A900002A08001280A08A801044104A1000001818C3",
INIT_01 => X"50A00011460214428114180000882214413D0A71592A01D92213D28005210202",
INIT_02 => X"8A54800A210200111100C2110054289220810440030404010844000444410001",
INIT_03 => X"1080010208B51400007800000A000001000108C21008092000018C6295200631",
INIT_04 => X"0008000000017000000028000001610300000010000802202040012040040011",
INIT_05 => X"2000044440048880026A22000026A20000000000000000004994140203000064",
INIT_06 => X"1400922401041008004891224228810080010200040001020800000004000008",
INIT_07 => X"150B001328000001404010040084088404200020455514000224489028492201",
INIT_08 => X"00414000201800004080A0000002480B04008100011000088800081002C19020",
INIT_09 => X"000400001036584108415B4A6A694A0000100101C08200000001000190200044",
INIT_0A => X"004800210C19808400500010009110091500020B408820000200400040811600",
INIT_0B => X"40000800B00100040D8140581405814058140581405814058140580A02C0A02C",
INIT_0C => X"00200248010201008298150006210802043058C46054032981002D00201C8081",
INIT_0D => X"0000A00000400600841041108280300008000140000401028008330000800040",
INIT_0E => X"0000A000000080001000000000000000500000040A40000000A00000040A4000",
INIT_0F => X"00000006000000080020C00000000000012000040A40000000A00000040A4000",
INIT_10 => X"00000000000024000000000080002000000000000000A00000040020A0000000",
INIT_11 => X"2200000404108000000900008080808000024040152000000020000004004080",
INIT_12 => X"0000000009001010102000004800080821000000120002000004000000000001",
INIT_13 => X"2000002000000000000288000020000805000000000001420000200001014000",
INIT_14 => X"408010000000022000D610280000080000000001204000000000000820020000",
INIT_15 => X"00401004010040100401004010042024210218734CD52150A840827504000000",
INIT_16 => X"0401004010040100401004010040100401004010040100401004010040100401",
INIT_17 => X"4010040100401004010040100401004010040100401004010040100401004010",
INIT_18 => X"05822140048D2E57B1348141845C200000000000000000000401004010040100",
INIT_19 => X"04104104104104104104104104104104104104104101A6A0A0EB1861863BC422",
INIT_1A => X"2C160B0582C160B0582C160B0582C160B0180C06030180C06030181041041041",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000160B0582C160B0582C160B058",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000000000000000000000000",
INIT_1F => X"4BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_23 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFF",
INIT_24 => X"FAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010000000000",
INIT_27 => X"FFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"E974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007F",
INIT_2C => X"FFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFA",
INIT_2D => X"D0402010000000000000000000000000000000000000000000000007FFFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"74BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFF",
INIT_33 => X"FFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE9",
INIT_34 => X"000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000007FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(3),               -- Port A write enable input
DIA(0)   => data_write_a(28),        -- Port A data input
DOA(0)   => data_read_a_lo_512(28),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(3),               -- Port B write enable input
DIB(0)   => data_write_b(28),        -- Port B data input
DOB(0)   => data_read_b_lo_512(28),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_29_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"79964E4BA01DACAB9E659792D00AAE160002829C7FDFEFCEE97C2815039D70C3",
INIT_01 => X"50BFF9AB0775343F9AB01DF80D5821FC0FFF3FEFD1AF9FF1207FFBC7B9720586",
INIT_02 => X"0D15846807D207200021C4E200D428A2018408600271C000720A0000003A2161",
INIT_03 => X"0000B0027BBF17C43E6DC05E1A0DC07D1F0000803B2819A00019084345606421",
INIT_04 => X"07CDC047A4FB526F807C681DC4B97369078249370F482E62BA414627C2FE3000",
INIT_05 => X"F204007861C088FF0EFF260407C427F19E03C7C01F8CF80749B390EA4BCA202C",
INIT_06 => X"000248C00079800406C081023B233E804488527FDC008019968D74982C94110A",
INIT_07 => X"5229000221FF8000398641903B082831D05000200000083F942850AEB4000221",
INIT_08 => X"00805FD0180E1F8C1111A0F041056A0100A11FE000916249A800B915FE82B020",
INIT_09 => X"F80C000055FF7C492840AAB45456B55E015015058665A31DA603A4539058F54C",
INIT_0A => X"000850400A11414C005005000B51158936D20601A98A204006114005C4800217",
INIT_0B => X"40201948B029029409A3401A3401A3401A3401A3401A3401A3401A9A00D1A00C",
INIT_0C => X"40B1225C1506512C83E85500AC3A080406305587A154023141006DFFF89E82C9",
INIT_0D => X"0000A01008480D3EB4A24A0C910037FFFC0007C7C0140D0B50A8218102C08160",
INIT_0E => X"0000A010010080005000000000000040520000141EC0000000A01000141EC000",
INIT_0F => X"00000046000002080429C0000000000001A000141EC0000000A01000141EC000",
INIT_10 => X"00000000000024080100010080006000000000000040B000010401A0E0000000",
INIT_11 => X"3600004414588000000D00108484C080000340483B590000202000008402C080",
INIT_12 => X"00000040090210909820000068008828B10000001A0802000204000000002001",
INIT_13 => X"20000120000000000082D800082000281D000000000021560002200011454000",
INIT_14 => X"B29450580000066021F6303C000408000000008320C000000000000860160002",
INIT_15 => X"816058160581605816058160589625662522506344FF9FCFFF62EB6DFF001004",
INIT_16 => X"1605816058160581605816058160581605816058160581605816058160581605",
INIT_17 => X"6058160581605816058160581605816058160581605816058160581605816058",
INIT_18 => X"F2DDCFFFBEFFCF07FFBFFD41800C05FFFFFFFFFFFFFFFFF81605816058160581",
INIT_19 => X"7DF7DF7DF7DF7DF7DF7DF7DF7DF7DD75D75D75D75D77FFBF3F7DFFFFFFD779F3",
INIT_1A => X"FEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDF7DF7DF7DF",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00001F7FBFDFEFF7FBFDFEFF7FBFD",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000000000000000000000000",
INIT_1F => X"4BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_23 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFF",
INIT_24 => X"FAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010000000000",
INIT_27 => X"FFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"E974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007F",
INIT_2C => X"FFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFA",
INIT_2D => X"D0402010000000000000000000000000000000000000000000000007FFFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"74BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFF",
INIT_33 => X"FFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE9",
INIT_34 => X"000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(3),               -- Port A write enable input
DIA(0)   => data_write_a(29),        -- Port A data input
DOA(0)   => data_read_a_lo_512(29),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(3),               -- Port B write enable input
DIB(0)   => data_write_b(29),        -- Port B data input
DOB(0)   => data_read_b_lo_512(29),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_30_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"FFDFF3FC3EFFF7FFFFBFFA000000000000000000000000000000000000000000",
INIT_19 => X"F3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF5F7AEBEBFBEFBEFFEFFF7",
INIT_1A => X"CFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCF3CF3CF3C",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000007F3F9FCFE7F3F9FCFE7F3F9F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000000000000000000000000",
INIT_1F => X"4BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_23 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFF",
INIT_24 => X"FAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010000000000",
INIT_27 => X"FFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"E974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007F",
INIT_2C => X"FFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFA",
INIT_2D => X"D0402010000000000000000000000000000000000000000000000007FFFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"74BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFF",
INIT_33 => X"FFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE9",
INIT_34 => X"000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(3),               -- Port A write enable input
DIA(0)   => data_write_a(30),        -- Port A data input
DOA(0)   => data_read_a_lo_512(30),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(3),               -- Port B write enable input
DIB(0)   => data_write_b(30),        -- Port B data input
DOB(0)   => data_read_b_lo_512(30),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_31_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"129000008004A00804A40000400800020000000C005FEA005800200400050100",
INIT_01 => X"A15FF18019700810180065FFFC0040801E80258CA2951C2200EC0906A0804140",
INIT_02 => X"146000808A0C060444692000402850040400408FF80000000010000000004000",
INIT_03 => X"000000FD74480B1C3D951C5A800D03FA1C0C21084B0300000012108518004842",
INIT_04 => X"07C51FC7EDFCA26E07EE001D1CB6904A061EDB6D4C30490281831C1602D0E480",
INIT_05 => X"C001F0808181117C7C95C8183FA099C7181F8703FF0CE3FC0201209010988002",
INIT_06 => X"00000000000000010001020400840C41C000617FC0003021259CFDB01BF00020",
INIT_07 => X"0000000441FA3FE400080200A810000010804008100040018448912040000040",
INIT_08 => X"00011F0780011E38004801C79E7C162231862E8FE00166704041240DF93D0000",
INIT_09 => X"F0C3FE180D89279000B00000000000D0F80088080849673F6C0E780020091480",
INIT_0A => X"1011DCCC31222730048620C4382204A608142002A440924A6188020920404437",
INIT_0B => X"0661874500E00E00304003040030400304003040030400304003060018200182",
INIT_0C => X"810040801060C04821202001A05A00040100240A80800442040202FFC3200444",
INIT_0D => X"000740000803C0616184184031010FFF40FFC407500020004C10060204010200",
INIT_0E => X"0007400000BD0020000008001F010000020201E04000010007400001E0400001",
INIT_0F => X"1DC0000000400D701000000800007700000001E04000010007400001E0400001",
INIT_10 => X"10003C064000C000010080BD0020000200001EC00000102006E8080000001000",
INIT_11 => X"140403A020000007200000E808000001C200000308C504021442354000000000",
INIT_12 => X"07B00000001D0100000038400007404000000E400000FC0010000000FC000000",
INIT_13 => X"5D00200000007C400000501001DC08000000001F010000140404558080000000",
INIT_14 => X"8C1380DA10400140640100D4080032903A8000000000403C3400008000140404",
INIT_15 => X"02008020080200802008020080200C1808008184012A08041202500AF87FF001",
INIT_16 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_17 => X"0080200802008020080200802008020080200802008020080200802008020080",
INIT_18 => X"000000000000000000000002001005FFFFFFFFFFFFFFFFF02008020080200802",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000000000000000000000000",
INIT_1F => X"4BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_23 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFF",
INIT_24 => X"FAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010000000000",
INIT_27 => X"FFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"E974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007F",
INIT_2C => X"FFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFA",
INIT_2D => X"D0402010000000000000000000000000000000000000000000000007FFFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"74BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFF",
INIT_33 => X"FFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE9",
INIT_34 => X"000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(3),               -- Port A write enable input
DIA(0)   => data_write_a(31),        -- Port A data input
DOA(0)   => data_read_a_lo_512(31),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(3),               -- Port B write enable input
DIB(0)   => data_write_b(31),        -- Port B data input
DOB(0)   => data_read_b_lo_512(31),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_0_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"ED39BA795990D275FB4A6E96ACC4731DEA4598B0AFB54867F6EE4618C3749807",
INIT_01 => X"58A0047D8607944AC7DA180001ECA2444042106208408208C20022E9173734B3",
INIT_02 => X"8B1E49562021F8051500147A0E162923024F28000415F5787B09FBF999BB1EFC",
INIT_03 => X"1013BF028A959403C06A23A147723C01E140088280C4CF6996088862C7922221",
INIT_04 => X"781A003802015D9078011DE20340699198600000B08694916434804825241311",
INIT_05 => X"2CA000587E10C880036A3103C00F2000E1E0383C00730002B4409845E4425171",
INIT_06 => X"179B48CFF95DCF9EF730E1C3BB731138AF7B888025340C0888430047040FEE18",
INIT_07 => X"AF155113160400185F87C1F05707D415E664A6E7C5551EBE783060CEB164833F",
INIT_08 => X"4D7E40002B7AE005FDB47600208229010C6101001EFE198C96B0528202C0DCB4",
INIT_09 => X"062400608234D864444081048A80CC00062D42D30222108091C107A1DA040267",
INIT_0A => X"204A21008E514844EB5145000255DA599581D3A9583C24351240B58298011308",
INIT_0B => X"E08C4830F81380CE0F89E07A9E0789E07A9E0789E07A9E0789E070CF0184F038",
INIT_0C => X"3A4E9D63EA180EB150CA1CA45C254D4AF4AA414568729139F2A12C0000016110",
INIT_0D => X"F0009E0FC048211E9C11C31F82E4A000890022B827EB52F52347F174E93A749D",
INIT_0E => X"F0009E0FCC42EFDFBF0AE03080E2AEB2E0F1F80FA97FE0F0009E0FC40FA97FE0",
INIT_0F => X"0231F0BD9E3FC08FEBD6F661C0E008C3CB5F040FAB3FE0F0009E0FC40FAB3FE0",
INIT_10 => X"20180309A0F83BE2B87C7C42EFDFBF187806013879BA878FE807F65FBF12E038",
INIT_11 => X"0BE9F01FC8B38C2098DAE007F323A0C83136B248831ACBFC8BBDCAB779BC699F",
INIT_12 => X"004C72BEC800FE7464290626D7003F9947184131B59003FFEC07F00003F01FB9",
INIT_13 => X"A0FFDA2A3C0202B8776A2FA7F023F7D065703080E29F1B2BE9F8A27E6E915C0E",
INIT_14 => X"016C2D25E52630BB1AE49C2BA7F98D6F846DFC0C2352A0024B83F07F198BE9F8",
INIT_15 => X"749D2749D2749D2749D2749D2749F285F25D2C500815A5522CB5A4B400000CD4",
INIT_16 => X"49D2749D2749D2749D2749D2749D2749D2749D2749D2749D2749D2749D2749D2",
INIT_17 => X"9D2749D2749D2749D2749D2749D2749D2749D2749D2749D2749D2749D2749D27",
INIT_18 => X"31C136AD8E9B562BA39E2600654BA800000000000000000749D2749D2749D274",
INIT_19 => X"4104104104104104104104104104104104104104104104109C83B8E38E2ABE71",
INIT_1A => X"0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0410410410",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000007C3E1F0F87C3E1F0F87C3E1F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000187FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"BAF7FFD55EF007FD75EFFFAE97555557BD75EF5D000000000000000000000000",
INIT_1F => X"000AA843FE00AAFBE8B45AA803DFEFA28428B455D0017410A28428AAAA2FBD54",
INIT_20 => X"FEBAA2D5401450051401555D7FC0145F7AEBFFFF08002AA10A2AABFEAAA2FFC0",
INIT_21 => X"D755555517FFEFA280021FF082E974AA5D7BFFE000804000BAAAAAAAB45557FF",
INIT_22 => X"EA8B45005168A10AA8028A10087FD7410557FC21555D51574AAA2FFE8B455D7B",
INIT_23 => X"AE95410AA80000005D003FEAAFFAEBFE00A2803FEBA002A820AA0800174BA5D2",
INIT_24 => X"2AEA8A10000417410A2FFE8BEFF7FFE8B45FFFBC00005D003FF45557FC01FFFF",
INIT_25 => X"00000000000000000000000000000000000000557DF5500003DFEFFF84175EFA",
INIT_26 => X"5F524AFE38B780154BAFFF1D54AF0075D75EFEBAE9554540754717F1F8000000",
INIT_27 => X"50B6AABDE12BEA0AF010B7D1F8F47E00A2DB45AA8A3AFD7B68E2AB78550E1255",
INIT_28 => X"E9257F1E816D557095EAAA2D1401D500002A150038038E285D7F78FD7000B6AB",
INIT_29 => X"5A87AAD178A8002D1D21C5E8257D5C7AA854008700249243A412EBFF5542A43F",
INIT_2A => X"52A82000E3A5D2150AB8F401471EDBC0B680900AAF52B474385D75C502D15754",
INIT_2B => X"FD7E9541242FE920AD082E10A28F6A150012A2F02AFFDF40E85F475451D502D1",
INIT_2C => X"0550E87B7A405B52AAD152BD00151EAFEDB52E3F1EFFFF485A2DA3D5D24BD417",
INIT_2D => X"57F40545850000000000000000000000000000000000000000000005AAF55508",
INIT_2E => X"F7AEAABFF5D2A81151FB8635A02FA69574BAF7D5555AF0D79D55FFA2AC974450",
INIT_2F => X"8D46F6ABE7082AAAAF2FAC77FE00FF16565B2FA9075F4F7B3EBDF50FEAEAAB55",
INIT_30 => X"56803CE3AEB038662E5D81406014D5D51F5E08A394003A908B8410E707EF34A0",
INIT_31 => X"4AF0151555AF58794040077D774FAE8C798A11A0EAEF75F7AA84001A7052C952",
INIT_32 => X"4E1870108B11020AD4AA05542A0A05051023F9A9D57B63BFBF906CB45FABC095",
INIT_33 => X"F5F0DA6BC9525688C1A2A0C06E9FEE5555BE48AB2A2AE0A0F20C43EAC562245B",
INIT_34 => X"000000FF80F55E25C00A0BA7FBED407A97F6F35F498B96BEB12DAAB77558ABD5",
INIT_35 => X"8000000FF8000000FF8000000FF8000000FF8000000FF8000000FF8000000FF8",
INIT_36 => X"00000000000000000000000000FF8000000FF8000000FF8000000FF8000000FF",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000008000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(0),               -- Port A write enable input
DIA(0)   => data_write_a(0),        -- Port A data input
DOA(0)   => data_read_a_hi_512(0),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(0),               -- Port B write enable input
DIB(0)   => data_write_b(0),        -- Port B data input
DOB(0)   => data_read_b_hi_512(0),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_1_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"212C001411984004084D000508C53810A03D1450E839B003342114428A000803",
INIT_01 => X"08000010400A0008010600000084005000400002000000000000000000140000",
INIT_02 => X"C084484000002014400205851002007030450E0000A606C8C44CB4C6666C00E0",
INIT_03 => X"CCF7CE0002058001000000800240200001018CA1800001091408463061120118",
INIT_04 => X"082800100000000040000900010000100040000000008411600401C02100000C",
INIT_05 => X"10800202080422000020012200000000810000200000000004020C00200011A0",
INIT_06 => X"56BDBFBC48C315A8660C18305750C008940D8000011000820001000104050004",
INIT_07 => X"8B4344400004000150248912154404C6060A2FE24555013E13060C158AC97F01",
INIT_08 => X"00082080087A000559102400200281000469000008B000000090108000400430",
INIT_09 => X"0000000000001004140545402820020000010010208000008041060008200001",
INIT_0A => X"2102210182004840007845004044020000200080080844200000048088000000",
INIT_0B => X"48800000190191064620646A06468064680646A0646A06468064690321503234",
INIT_0C => X"02008100200800A1100707040101E20BE0B002605C1C110848200C0000000800",
INIT_0D => X"F000A000C0000012187087010AE4B00000000810010040108104100408020401",
INIT_0E => X"F000A000CC4200002F08E03080000010F18058000003C0F000A000C4000003C0",
INIT_0F => X"000000078808C00000023461C0E00000012704000003C0F000A000C4000003C0",
INIT_10 => X"201803000000240218C0044200001E1878060000000AAC00680000001F10E038",
INIT_11 => X"2100B00048230C200009A0001303204800025200040A00D000000202090C281F",
INIT_12 => X"00000002C9000260640900004D0000904618400012900001EC03F00000000039",
INIT_13 => X"80025A0A3C020000002A8400B00007806070308000000961002880204A901C0E",
INIT_14 => X"000801046004308A185000020128000904285C0C0312A0020000000838810028",
INIT_15 => X"0401004010040100401004010040100010410C002000040280100000000008D0",
INIT_16 => X"4010040100401004010040100401004010040100401004010040100401004010",
INIT_17 => X"0100401004010040100401004010040100401004010040100401004010040100",
INIT_18 => X"48D757DF8A9410218E8A56085142020000000000000000004010040100401004",
INIT_19 => X"555555555555555555555555555554514514514514550431A581924924B02651",
INIT_1A => X"4BA5D2E974BA5D2E974BA5D2E974BA5D2EB75BADD6EB75BADD6EB75555555555",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800005D2E974BA5D2E974BA5D2E97",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000607FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"10AAAABFFFFFF803FE10F7D17FEBA55556AAAAAA800000000000000000000000",
INIT_1F => X"EBAFFD555400557BD54BA5D7FFDF45A2FBD75EFA2AE97555F7FBFFF45FFAE800",
INIT_20 => X"ABEFA2D568A005D5157400AA8028AAAF7FBD54AA002A955555D7FE8ABA082EBF",
INIT_21 => X"FDF55AAFBC0010555540010550417555AA8028BEFAAAE97555082A80000AA802",
INIT_22 => X"BD7410550428ABA5D5168ABA552EBDFEF5D7FEAA00AAAABFEAA007BC0145FFFF",
INIT_23 => X"FFEAB55557FFFEBAAAD568B45A2D5575555D7FC2155F7AEA8BEFAAAA954BA557",
INIT_24 => X"D7BD74000804154BA082ABFF55FFD57DF45F7D568ABAF7AABFFFF082ABFFFFFF",
INIT_25 => X"000000000000000000000000000000000000002EBFFEFA280021FF082E974AA5",
INIT_26 => X"5E175EFF57BF8FC2000BEA4BAE97F78A3FE28E3D17DEAA485FE8E02B50000000",
INIT_27 => X"455571E8A2A087BF8EAAEB8E0016D5D75D54BA5D7BFFF7DA2FFD55EFAAA49554",
INIT_28 => X"157428145A00AA8A2FBD7B6DF6AA28550E10405F7A4AFE38EAA0924921C2FD55",
INIT_29 => X"8E971471C7010B7D168F47400A07A28415A001684104155C5B6DF6DBEFBFAA07",
INIT_2A => X"BFBD7B6A0BF492415FC20105D24AAABF1FFBC7010FF8A38FEF557FEAB78B6AAB",
INIT_2B => X"017EBA4A8EB8F6FFD5FE8B7D557495EAAA2D16D1FDBED56A55557A43DE385FD4",
INIT_2C => X"854008700249243A417FFF41542F5D717FE2AAAA56DEBD17FE3DF7FB7FEBFE38",
INIT_2D => X"07DFCA127B8000000000000000000000000000000000000000000002A3D5C7AA",
INIT_2E => X"AAFBD55FFAA8416545A6FB60F47AF2A00010F78028B15F7823FEAAA2D57DFBA0",
INIT_2F => X"22A38C20B2552E975F758516AAAA0869AAAB8A7C19C55550E8574BA557BFFFEF",
INIT_30 => X"55FFEFBCEE5FBAACB10085EE5DE10A2AEBFF55F7BAAA8565DBAC1112FFAC21A0",
INIT_31 => X"BEA097BEAAFAF2863FA00DD574201E7AD1FFF5575841DE08007FC20480028957",
INIT_32 => X"54FF57EFBFA18D4FBFFF40FF809D4000D7FC00FC5D062BBA05ED5034472A02EA",
INIT_33 => X"7DFBFF6963FCAAA2283CF14050062B0A2F7AE8B5D5D51F5E18ABD5EAFFF2AF95",
INIT_34 => X"000000002CB75F7AA84001A7052C95256807DC31AA8114DE55F5BED201FFFED1",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000008000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(0),               -- Port A write enable input
DIA(0)   => data_write_a(1),        -- Port A data input
DOA(0)   => data_read_a_hi_512(1),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(0),               -- Port B write enable input
DIB(0)   => data_write_b(1),        -- Port B data input
DOB(0)   => data_read_b_hi_512(1),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_2_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10E44660018259B2843913100062C98004802322D3E030235201006009B2813",
INIT_01 => X"000AC188084900481C8024A542400340404000720885800802000906E4910204",
INIT_02 => X"82040072AC248C31010204880000007401044C0550200000480E0080001300E0",
INIT_03 => X"0080812C130D0A0D1193088802182142494D218220021100001A8020C1004A00",
INIT_04 => X"090D0AD62824A44A428408540D1610020C6E510818923441A4908B0503404201",
INIT_05 => X"5000A004081122242420480A14A99C428908122144244150906124248C002168",
INIT_06 => X"1400088400450000460000001308890094082015800011012D41D518044C1100",
INIT_07 => X"26731111491C1541324C1114BD880004002040204050413F1400100480000201",
INIT_08 => X"02410582881E0C1511D02082AAAB016A2463288549B044605201D10AE11B0020",
INIT_09 => X"E80394280E40158020B591000800481051241A4A404B5035C60904502054E000",
INIT_0A => X"0102C9E12202EA6014D027C418428E220A5500024808922801A0900A84454458",
INIT_0B => X"4600070110C10D04340043400434A043420434A04342043480434102184021A0",
INIT_0C => X"E9CA34328E44CA1401306100A246000402100C088104010AC8005C5681812B04",
INIT_0D => X"0000A0000801487334E34C1A980001550055481204090A4C01351253A728D194",
INIT_0E => X"0000A000013800004000080000000000500000B01480010000A0000150148001",
INIT_0F => X"0000000608000A500409000800000000012001501480010000A00000B0148001",
INIT_10 => X"1000000000002400000001A100004002000000000000A0000360018040001000",
INIT_11 => X"380001C01048000000090298040440000002400008C400022042004080028000",
INIT_12 => X"0000000009530080880000004813802090000000120C94000200000000000001",
INIT_13 => X"4C000100000000000002E0000950002018000000000001580002508010440000",
INIT_14 => X"7120642000000400015020500004221018000082008000000000000820180002",
INIT_15 => X"5094A5294A5294A52942509425094209461468000822241A03835D88482AB001",
INIT_16 => X"09465094A5294A5294A5294250942509425094A5294A5294A529425094250942",
INIT_17 => X"94650946509465294E5294E5294E5094650946509465294E5294E5294E509465",
INIT_18 => X"080271AE180616A38A18FA204452A7F03F03F07E07E07E05294E5294E5294E50",
INIT_19 => X"20820820820820820820820820820820820820820820490C04102CB2CB2EB2C0",
INIT_1A => X"8944A25128944A25128944A25128944A25128944A25128944A25128208208208",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF1F804A25128944A25128944A2512",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000787FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"AAAA843DFFFAAD1554005D7FD74AA00040015500000000000000000000000000",
INIT_1F => X"F45AAAAA8A10A2AE80010A2AA975FF5D003FE10F7D17FEBAF7D5420AA0855420",
INIT_20 => X"FF45A2AA975EFA2FFD7555FFFBFFF45AAFBC20AAF7D1575EF55517DF555D2EBF",
INIT_21 => X"95555552E974105D517DF55AAAAAABEFAAD1575EFAAAE974AA5D51554BA5D7FF",
INIT_22 => X"E82010F7AABFE10FFD542145FFD5554AA555555555557FE8ABA082EBFFFFAAAE",
INIT_23 => X"FBC0010AA802ABEFAAD540000FFD540000AA802AABAF7FFC2010AAAE821EF552",
INIT_24 => X"A8028BEFAAAE821550851420AA002E800AA08042AB45007FC00BAFFD168BEFF7",
INIT_25 => X"000000000000000000000000000000000000002E80010555540010550417555A",
INIT_26 => X"AE95F40002157F470AABE803AE97A2DF55400557FD54AA1D04001C5150000000",
INIT_27 => X"EF55517DFC5552ABDF45B6AEAFFD5F7A482000BEAE905C755003FE28E3D17DEA",
INIT_28 => X"0BA5FD0154BA5D7BFAF7DA2AE955EFAAA495545E3F5EFF57F7FE80082FFDE105",
INIT_29 => X"8AAF082AB8EAAEB8E0016D5D2A924105D5B7FF7DB6AAAABC7BEDB505EFBEA407",
INIT_2A => X"95038AAAEAF1D7410E80000FF8438E00B6DF68FEF4871D24BA495B5556D5571E",
INIT_2B => X"1ED1EFEAF1EFFFDEAD1C5010AA8E2FBD7B6DF47A00EBDB50000A380AAE28E804",
INIT_2C => X"5A001684104155C5B68E2DBEFBFFBC703AE2DF42AAA002A851C214003FF68007",
INIT_2D => X"50002155510000000000000000000000000000000000000000000002087A2841",
INIT_2E => X"55003FEAAAAD57DEBAA2FDDC01051FBD74BAF7802AB05AAFBD5400557BD54AA5",
INIT_2F => X"7AF7FC20B2F7FBC015D58517FF555D2ABDF55F782BEB47AFAD00010F7AA82155",
INIT_30 => X"55FFFFC20FFF3AE544108410174BA557BEABEFAAEBD55FFAA1456547A2D360F4",
INIT_31 => X"0BA547FD75FF58516AAAA0828AAAB4A78016545540400010557BFDFFFF7822A9",
INIT_32 => X"550AAFACAAA122AA8954BAA2AE9D545002A800A8FF862BA00F2F9E8F0050D442",
INIT_33 => X"954505C417FFFF08555555BAAD335B57AB5155400A2AEBFF45FFFB404007FFBD",
INIT_34 => X"00000000061DE08007FC2048002895755FFAEBCFE57BBA57002DF3C4AAAA002E",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000010000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(0),               -- Port A write enable input
DIA(0)   => data_write_a(2),        -- Port A data input
DOA(0)   => data_read_a_hi_512(2),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(0),               -- Port B write enable input
DIB(0)   => data_write_b(2),        -- Port B data input
DOB(0)   => data_read_b_hi_512(2),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_3_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"210C44A20020248B08431120001604B8156023104C40771B3430400A02380206",
INIT_01 => X"015A2A4050B009683C0422C992000B61404040028804A0080A000C16A8990A0C",
INIT_02 => X"C0A406500CE0A95011000D1501005274B5041AB330860281CC08008222170060",
INIT_03 => X"AB488054270F08E1289084C8020420E005A48DA16C021100003A46B06900C91A",
INIT_04 => X"848966150DA0A02941A4080C612A104201C689044382FD403C17E491829B259B",
INIT_05 => X"D006620608843116942508120A208D18A5050160C600D4C894600094B49CA068",
INIT_06 => X"12002D9401C70008060408141788E2C094887033080071913209CC8004640100",
INIT_07 => X"221111454874CCC4122C0932155400C2023940284000003E15020525CE805E11",
INIT_08 => X"020103C9984A0AC511102029869D974214EDBA132891000052C1750B48290020",
INIT_09 => X"60808C8A2E41351020004148A289428730A51E5E644C8233A0090E1020208100",
INIT_0A => X"A4000041A600417914506F955D6422000934000A090A94A020229603A414144D",
INIT_0B => X"469100841001000406D04065040650406D0406D04065040670406C8201782032",
INIT_0C => X"6A4AF532A8040AF821042D01F14084030070262810340402C0000CCE4CC12520",
INIT_0D => X"000800000401C333494594532980733302CCC81300094E5C91200257AD2AD795",
INIT_0E => X"00080000051C0000400000000000000800000190148000000800000450148000",
INIT_0F => X"0000010000000B100409000000000004000005101480000008000004F0148000",
INIT_10 => X"0000000002000000000001B00000400000000000000400000168018040000000",
INIT_11 => X"1000034010480000010002D804044000004000812E4400002440014080028000",
INIT_12 => X"0000000100570080880000080015C02090000002000CCC000200000000000040",
INIT_13 => X"1C0001000000000000104000094C002018000000000040100006418010440000",
INIT_14 => X"4128652000004404010E20500004208018800082008000000000010000100006",
INIT_15 => X"5795A5595A5595A5595A5595A5595E1152556D008028341B13924D80C2E67009",
INIT_16 => X"69565795A5595A5595A5595A5595A5595A559525795257952579525795257952",
INIT_17 => X"95256956579525495E5595A5495E5595A5495E5595A569565795256956579525",
INIT_18 => X"7818F18E0C8514298B0C52A0115009AA9556AAD552AAD5556956579525695657",
INIT_19 => X"24924924924924924924924924924820820820820825042C0000249249202A60",
INIT_1A => X"8D46A351A8D46A351A8D46A351A8D46A353A9D4EA753A9D4EA753A9249249249",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF248086A351A8D46A351A8D46A351A",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"EFAAFFD54AAF7D168B45AAAABDF5500002AA1000000000000000000000000000",
INIT_1F => X"F45FFD168AAA0855420AAAA843DFFFAAD1554005D7FD74AAA284001550055421",
INIT_20 => X"55FF5D003FE10F7803FEBAFFD5420AA080400155AAD5554AAF7802AB4500043D",
INIT_21 => X"28B45A2AE82155A2FBFFEBA0800021550855555FFAA84001FFAAAE80010A2AA9",
INIT_22 => X"168ABAFFFBD54BAAAAE97400A2FBC20AAA284175EF55517DF555D2EBFE00AA80",
INIT_23 => X"AA954AA5D7FFFF45AAAA975EF007BD7555FFFBFDF55AAFBD55EF5D2EBFE10085",
INIT_24 => X"AD1575EFAAAE974AA5D00175555D0015410F7AAAAAAA55043DE00FFFFD5555AA",
INIT_25 => X"0000000000000000000000000000000000000004174105D517DF55AAAAAABEFA",
INIT_26 => X"ABC04001C51551471D7AAF1D05D2EBD56DB7DBEAEBFF551C042AA101D0000000",
INIT_27 => X"92EB842FB5508043FF55EBD56ABD75D5B470AABE8A3AFD7A2DF55400557FD54A",
INIT_28 => X"557FD2082000BEAE905C755003FE28E3D17DEAAEBDF40002550F47155AADB504",
INIT_29 => X"DF40552ABDF45B6AEAFFD5F7A48017DAAFFFAE821C0A0717D1C5B575FFB68E82",
INIT_2A => X"C55D7492E90E3808756DA92EBFFD74BAE3AE85480FFFFC00AABE8E105C755517",
INIT_2B => X"43AE10EAF5C5547FF80954AA5D7FFAF7DA2AE905EF0075D5545E3F5EFF57F7D5",
INIT_2C => X"5B7FF7DB6AAAABC7BEDB505EFBEF5C7092FF801756D490A10438EBA4B8E92410",
INIT_2D => X"D0028A00510000000000000000000000000000000000000000000000E124105D",
INIT_2E => X"AAFBD54005D7BD54AAF78002155515157555AAD142040A2D57FFFFFFAEBFF555",
INIT_2F => X"051AE955F7AAFBC0000AF843FF5500003FF55AAFD6AB455157D74BAF7AAA8B45",
INIT_30 => X"FF557BD74EFFBACD41577B8400010F7AA8215555003FEAAAAC53DEB8A2FDDC01",
INIT_31 => X"0BAF7AA8015558517FF555D2ABDF51F782BCB47ABAE801FFAAFBEAA105D2E955",
INIT_32 => X"214FA2D3EAF57AFFDD7555082AA0AAA00557FEA8A2FDD64BAAF8282012AFFEC2",
INIT_33 => X"820AAAB842AA00000028AB0AAFF48547AE04174BA557BEABEFA2AA951FF88554",
INIT_34 => X"000000002A80010557BFDFFFF7822A955FFFFC21FFF3BE40412DE02955FF082A",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000008000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(0),               -- Port A write enable input
DIA(0)   => data_write_a(3),        -- Port A data input
DOA(0)   => data_read_a_hi_512(3),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(0),               -- Port B write enable input
DIB(0)   => data_write_b(3),        -- Port B data input
DOB(0)   => data_read_b_hi_512(3),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_4_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A108400020612C80284210081034849800A000303100048B3432C82904204006",
INIT_01 => X"210668000008004C1C20250E12100368403008418984014902030906A8910200",
INIT_02 => X"120404C0024C0600000206100008402404040C00F104008040080080001310E0",
INIT_03 => X"7728805052470B5C1B873C04121D03845D0020CA0822018000080084C1000002",
INIT_04 => X"0B899E43891686690790485D5C3E02000E9892201D306D03A9835C16029AC186",
INIT_05 => X"C001E080005030767434C0003C8A01D6B81C5703C82CDBC000072400089C8120",
INIT_06 => X"1000088100410000460002041300004084080070D00030032009700024641102",
INIT_07 => X"4261950408CCBC2012048310951000000003402A4000143E1008912480000211",
INIT_08 => X"00811007AC0A1EB5131120C79E7D176251E53E80E8B361604041340838452020",
INIT_09 => X"C08360820C0912800035F1801630A8260900180C00C8021C800FEE522020A108",
INIT_0A => X"8400F88C166262E940D00D410D62AD02091704024D0A02882192020DA0544043",
INIT_0B => X"4011078510C90D143142430C243042430C24304243042430C24305121A612186",
INIT_0C => X"C08060101000C00401008800F004140009400E4002A0010240000DC3C080002C",
INIT_0D => X"000800100001C07261C51C42390240F050C3C000950008088130040100018000",
INIT_0E => X"00080010003510004000000000000048010002E0100000000800100220100000",
INIT_0F => X"0000014008001550000800000000000400800280100000000800100360100000",
INIT_10 => X"00000000020000080080009410004000000000000044080000D8008000000000",
INIT_11 => X"000005800008000001040168000040000041000100EC00004002214000008000",
INIT_12 => X"00000041003C000008000008200D00001000000208050C000200000000002040",
INIT_13 => X"17000100000000000090000002C8000008000000000060000004480000400000",
INIT_14 => X"8400C00208004844C00800000000528008000000008000000000010040000000",
INIT_15 => X"0100800004030080000C010000A00D1804404912802A261B53104810DB1E0028",
INIT_16 => X"000C030000200C01000020040300800004030000000C03000000040100802004",
INIT_17 => X"008020040100C010000200800004010040300800000020040100C03000020000",
INIT_18 => X"40C700FC0A000280C68A08A950520E964C3269B2C9864D30000C030040100800",
INIT_19 => X"555555555555555555555555555554514514514514526991A199A28A28981451",
INIT_1A => X"41A0D068341A0D068341A0D068341A0D06A351A8D46A351A8D46A35555555555",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF771F60D068341A0D068341A0D0683",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FF087FFDF5508003FEBA087FD54BAAA841540055000000000000000000000000",
INIT_1F => X"F5500003DF455555421EFAAFFD54AAF7D168B45AAAABDF55A2802AA1000002AB",
INIT_20 => X"DFFFAAD1554005D7FD74AAAA840015500002AABA082E954005500021FF5D2EBF",
INIT_21 => X"68BEF080028BFF0855555455500174BAA2AABDE0055517FF555555420AAAA843",
INIT_22 => X"168ABA0055574BA5555554BA5D0400155AAD1554AAF7802AB4500043DF45FFD1",
INIT_23 => X"0400010A2AA955FF55003FE10F7803FEBAFFD5420BA085168A00007BFDE10085",
INIT_24 => X"855555FFAA84001FFAAFBEAB45002A97545F7D1555EF55043DF5555517DEAA5D",
INIT_25 => X"000000000000000000000000000000000000002A82155A2FBFFEBA0800021550",
INIT_26 => X"5BC042AA101D0A28BC7007FFDF45080A3AEAA007BD2482BE84124285C0000000",
INIT_27 => X"004100021FF492AB8F7D1C0438E381451471D7AAFBD0492EBD56DB7DBEAEBFF5",
INIT_28 => X"FED1C5F470AABE8A3AFD7A2DF55400557FD54AABE84001C5550A28ABA1424974",
INIT_29 => X"FB5508043FF55EBD56ABD75D0428BEF005557545490012482B6A0BAE2849557A",
INIT_2A => X"6DA101475FDE10145F68A921C55504924955524AA140E0717DAADB50492EB842",
INIT_2B => X"43AF6D405F78E3A1C2002000BEAA905C755003FE28E3803DEAAEBDF40002557F",
INIT_2C => X"FFFAE821C0A0717D1C5B575FFB6DF425575D7BEFB55002097555FFD5401EF5D0",
INIT_2D => X"784000AA59000000000000000000000000000000000000000000000208017DAA",
INIT_2E => X"A2D57FFFFF7AEBFF55FF8028A00512EAAB45007FFFF55082EA8AAA087FC2010F",
INIT_2F => X"5512AAAA085D04174100800021FF002EA8BEF5D0428ABA595557555AAFBC2000",
INIT_30 => X"00FF802ABAA04552ABFF597FD74BAF7AAA8B45AAFBD54005D7BD54AAF7800215",
INIT_31 => X"5FFAAFBC0000AF843FF5500003FF55AAFD6AB4551002ABEF0055555550004020",
INIT_32 => X"DEB0A2FD5600051537DE005D557DE005D7BE8AA85555400100879560AA592F95",
INIT_33 => X"17545FFD5421FF5D0428BEF0079FCABA598400010F7AA8215555003FEAAAA843",
INIT_34 => X"0000000004001FFAAFBEAA105D2E955FF557BD75EFFBBCD415521FBFDF450004",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000010000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(0),               -- Port A write enable input
DIA(0)   => data_write_a(4),        -- Port A data input
DOA(0)   => data_read_a_hi_512(4),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(0),               -- Port B write enable input
DIB(0)   => data_write_b(4),        -- Port B data input
DOB(0)   => data_read_b_hi_512(4),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_5_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50DB0A0791B1B41694368283C81F9996A091A32152007AB36B20E03C040C002",
INIT_01 => X"880015C49830884C446A40000C34C24841280A00084000C8C212892EEA953231",
INIT_02 => X"408F417400B1D9100002171C1FA20171124E6AA00D8633F8CD09DBFBBB972F7C",
INIT_03 => X"88538F0182058082D800C3314722DC08A34084A100C4D7C99208521063D00148",
INIT_04 => X"F45E41AFAF420996B8411CA282F80A9091224800A2C61490363080C8A4000308",
INIT_05 => X"0EA416069640420901A01505C4410020C6E228DC30532839B043289D9C005031",
INIT_06 => X"13992D9AF8C74E92B7B568D19708C038AFFA89F0B9348C9204C389672407EF12",
INIT_07 => X"6255000016053C18162589725146F442222CE6AF844012BE795224458BA4DE0F",
INIT_08 => X"4F3F00503B4AE104B5347230418190420821006016FC18843630D285FC416CB4",
INIT_09 => X"EEA33E700340902C4424C442B0344724066C56C2248130A2D9C185B24A24832B",
INIT_0A => X"315325008348CC40AB570500204462508135D5AA593E043731E9B18A98440137",
INIT_0B => X"E0CD463C5813804E0258E0358E02D8E03D8E0258E03D8E02D8E03447012C701E",
INIT_0C => X"F8DE3C27CA181E5D710664A5F140C14BD32A2E281992940AFAA15C3FC0836310",
INIT_0D => X"F000BE0FC80020130841840308653FF0313FE92C23FB1EECB367C0F3E378F0BC",
INIT_0E => X"F000BE0FCD806FFFAF0AE83080E2AEB2F0F1E01BE53FE1F000BE0FC41BE53FE1",
INIT_0F => X"0231F0BF9E3F02A7FFD63669C0E008C3CB7F041BE1BFE1F000BE0FC41BE1BFE1",
INIT_10 => X"30180309A0F83FE2B87C7D006FFF9F1A7806013879BAA78FC103FF5F1F12F038",
INIT_11 => X"39E9C1DBF8A30C2098DBE2FF7F2320483136F200A822CBACAB9DDEB7F9BC291F",
INIT_12 => X"004C72BEC95FEF64E4090626DF15B7D1C6184131B7980DFFFC03F00003F01FB9",
INIT_13 => X"1DFFFA0A3C0202B8776AE7A7C9CBFFF060703080E29F1B79E9F6427EFE901C0E",
INIT_14 => X"2B716CA5C56620590350ACD3A7D5B7EFAC6DFC8C0312A0024B83F07F3999E9F2",
INIT_15 => X"F0BCAF3BC2F3BC6F0BCEF2BC2F3BC6DBC67C251104A2261253904580207E1C81",
INIT_16 => X"1BCEF0BC2F3BC2F1BCEF0BC6F2BC2F1BCAF1BC6F2BC6F2BCAF1BC2F3BC6F2BCE",
INIT_17 => X"BCEF0BC2F3BC2F1BCAF1BCAF3BC6F0BCEF0BCEF2BC6F2BCAF1BCAF1BC2F3BCAF",
INIT_18 => X"69CFEF73B6FFE7436DB6FD0831518424965B4D2492CB69AF1BCEF0BC6F2BC6F0",
INIT_19 => X"F7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF3EF9FBFBB9E79E7BEBCB7",
INIT_1A => X"DEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDF7DF7DF7D",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF29FDAF77BBDDEEF77BBDDEEF77BBD",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"AAA2802AA10FFFFFDE0008556AABA5D2ABFFEFFF800000000000000000000000",
INIT_1F => X"ABAF7AAA8BFFAA802ABFF087FFDF5508003FEBA087FD54BA0804154005555574",
INIT_20 => X"54AAF7D168B45AAAABDF55AA802AA1000003FEBA00002AABA5D2EBFEBAAAD16A",
INIT_21 => X"3DE005555575EFA2D142145A2FFE8B45FF80001555D2E955FFFFD5421EFAAFFD",
INIT_22 => X"FC00BA5D5568AAAF7AAAAAAAAA802AABA082E954005500021FF5D2EBFF550000",
INIT_23 => X"D5420AAAA843DFFFAAD1554005D7FD74AAAA840014500517FFEF007BEABFF5D7",
INIT_24 => X"2AABDE0055517FF555504154BAA2FBEAA105D2E97410FFD16AAAA5D2ABDEBAFF",
INIT_25 => X"000000000000000000000000000000000000000028BFF0855555455500174BAA",
INIT_26 => X"21E84124285C51574BAB68A2DA00FFFFFFE38085F6FA92552AB8FEFF78000000",
INIT_27 => X"925D2AB8EBABEDB6AA92F7AAA8BC7B68A28BC70075FDF45080A3AEAA007BD248",
INIT_28 => X"5FFFFD1471D7AAFBD0492EBD56DB7DBEAEBFF55BE842AA105D0A38EBA1C0428A",
INIT_29 => X"21FF492AB8F7D1C0438E38145B575EFA2DB45145B6F5EFB6DF78E05145552A92",
INIT_2A => X"7DFC70875EABC7557FC20AA415F68AAAF7AAAAA82BE8A28A9214249740041000",
INIT_2B => X"B6FABA542ABAE2AF7DF470AABE8A3AFD7A2DF55400557FD54AABE84001C55551",
INIT_2C => X"5557545490012482B6A0BAE2849043AFED1C0E10492B6FFEFA105D2A95410FFD",
INIT_2D => X"D2AAABEFFB8000000000000000000000000000000000000000000000428BEF00",
INIT_2E => X"082EA8AAA087FC20105504000AA5955554BAFFAEBDE10F7FBFDEBA007BFDE005",
INIT_2F => X"0512AA8AAA5D0028A005D2AA8ABAF7FBE8A00FFAEAAB45F3AAAAB4500557FF55",
INIT_30 => X"EFFFAA97545552A821EFFBD557555AAFBC2000A2D57FFFFF7AEBFF55FF8028A0",
INIT_31 => X"A005D04174100800021FF002EA8BEF5D0428ABA597FD55FFA2FFD5555FFD57FF",
INIT_32 => X"54AAF7800015551517DF45005168B55557FC0012087FEAABAF7AAAAA10F3AAAA",
INIT_33 => X"FFE005D2A95410F7FFFFEBA5D2EA8ABAFBFFD74BAF7AAA8B45AAFBD54005D7BD",
INIT_34 => X"00000000002ABEF005555555000402000FF802AAAA04452ABFF592E80010FFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000060000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(0),               -- Port A write enable input
DIA(0)   => data_write_a(5),        -- Port A data input
DOA(0)   => data_read_a_hi_512(5),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(0),               -- Port B write enable input
DIB(0)   => data_write_b(5),        -- Port B data input
DOB(0)   => data_read_b_hi_512(5),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_6_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10800B0061A01002840002C030028180004003220200403312301C4389B2082",
INIT_01 => X"060009C838394848188160000C42426041000000090800090210090000510200",
INIT_02 => X"00043040009001100000061000018070002408000000000648080000001210E0",
INIT_03 => X"0000800002054081020080801200A0000300008000201184681A0000410C4800",
INIT_04 => X"0808801040000001401048008100022401400002024024053200020089000100",
INIT_05 => X"0240040408402202002000C200400020A50000A0000010010001260808000520",
INIT_06 => X"44000881064500004600000013088002840C240F5048011200010000440C0146",
INIT_07 => X"0241914041FE83E010040110110003040020402A0000003E1000000488000201",
INIT_08 => X"8001BF002C4A01041B112020200110024029006FE09081002004902000012068",
INIT_09 => X"0083FE38A040100281353150ACB645AEF8C01404448000008011061204200108",
INIT_0A => X"3103AD0413424E4014D627C470462200011504420C0A962A2189002881404060",
INIT_0B => X"46C1060C16C96D15B0425B0425B1425B1425B0C25B0C25B1C25B1512D8212D82",
INIT_0C => X"009000140401100601016600A040220203A004480598010248000D0010420C0C",
INIT_0D => X"0000A01033A00013000000000018800F2400091081100C0090A5008200410020",
INIT_0E => X"0000A0103142000000000000000000455D0018100000000000A0103410000000",
INIT_0F => X"000000466800C200000000000000000001A0F4100000000000A0103410000000",
INIT_10 => X"00000000000024094680014200000000000000000041E8002900000000000000",
INIT_11 => X"F000322000000000000D1A000000000000034D240C2000502000000000000000",
INIT_12 => X"000000403F4000000000000068D24000000000001A60F0000000000000002007",
INIT_13 => X"C0000000000000000087C0003014000000000000000025D00008958000000000",
INIT_14 => X"02000000000814C219500150002800101280000000000000000000086670000C",
INIT_15 => X"8120C82208812048120882208892055A0060011280222413130449010301F051",
INIT_16 => X"3200802008320C82200802048320C82200812048320880200812048220880204",
INIT_17 => X"20C83208812048020883204802048120882204812008220C8220081204822088",
INIT_18 => X"79CFF1FE1E9F52ABEF9EFE8150120EC718638E38E30C71C812088220C8120080",
INIT_19 => X"71C71C71C71C71C71C71C71C71C71C71C71C71C71C736D9DBD9BBEFBEFBEBEF1",
INIT_1A => X"CFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FC71C71C71C",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCF29A7F3F9FCFE7F3F9FCFE7F3F9F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000607FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"EFA2FBD54BA5555554BAAAFBC20BA5D7BEAAAAFF800000000000000000000000",
INIT_1F => X"EBA0855421455555574AAA2802AA10FFFFFDE0008556AABA5D2ABFFEFFF843DF",
INIT_20 => X"DF5508003FEBA087FD54BA000415400550428AAAAA84021FF007BD54BAAAD17D",
INIT_21 => X"A8BFFAAD1554BA002A95555A28417400AAFBE8ABAF7FFD54AAAA802ABFF087FF",
INIT_22 => X"BD5545080417555A2D17FE1000003FEBA00002AABA5D2EBFEBAAAD16AABAF7AA",
INIT_23 => X"D5421EFAAFFD54AAF7D168B45AAAABDF55AA802AA100000001EF087FEAA00FFF",
INIT_24 => X"F80001555D2E955FFFF843DEAAA2803DFEF0855401FF082EA8B555D7FC21FFFF",
INIT_25 => X"0000000000000000000000000000000000000055575EFA2D142145A2FFE8B45F",
INIT_26 => X"2552AB8FEFF78E3DFFFAAFFD04AA415B52492B6F5C20825D7FE8A92FF8000000",
INIT_27 => X"EF147BD2482BED57AE921451421555551574BAB68A2DA00FFFFFFE38085F6FA9",
INIT_28 => X"4BAB68A28BC70075FDF45080A3AEAA007BD24821C04124281C0E2DA82BE8E001",
INIT_29 => X"8EBABEDB6AA92F7AAA8BC7B6D5524AA14209557DA28E15400BEF1EFA92FFFFD2",
INIT_2A => X"071FF0071EDA38F7F1D5555000417545B6D178E281C0A38EBA1C0428A925D2AB",
INIT_2B => X"4A8B555C7FC2147F7D1471D7AAFBD0492EBD56DB7DBEAEBFF55BE842AA105D0E",
INIT_2C => X"DB45145B6F5EFB6DF78E05145552A925FFFF8E3DE82BE8E38FFF0851401C7082",
INIT_2D => X"57FE8A00F38000000000000000000000000000000000000000000005B575EFA2",
INIT_2E => X"F7FBFDEBA007BFDE005D2AAABEFFBAABDFEFAAFBC00BA007BC0000FFD5420005",
INIT_2F => X"A592ABFE00F7AA821FF557FC0010F7D168A105D55421455155554BAFFAEBDE10",
INIT_30 => X"10F7D57DE00FFFBC00AAFBAAAAB4500557FF55082EA8AAA087FC20105504000A",
INIT_31 => X"AAA5D0028A005D2AA8ABAF7FBE8A00FFAEAAB45F3D5400BA5504155EFAAAE954",
INIT_32 => X"FF55FF8028A00512E975FF08557FEAAF7D157545080417545F7D56AAAA592AA8",
INIT_33 => X"AABEF005542155000028B555D7FC2145F3D557555AAFBC2000A2D57FFFFF7AEB",
INIT_34 => X"000000007FD55FFA2FFD5555FFD57FFEFFFAA97545552A821EFFBAABDE00F7AA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000048000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(0),               -- Port A write enable input
DIA(0)   => data_write_a(6),        -- Port A data input
DOA(0)   => data_read_a_hi_512(6),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(0),               -- Port B write enable input
DIB(0)   => data_write_b(6),        -- Port B data input
DOB(0)   => data_read_b_hi_512(6),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_7_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10844B00482258A2842112C02450418800002300500030B313300C418992002",
INIT_01 => X"020009C23838684D1C20E0000E11424840000000080000080200000000110204",
INIT_02 => X"000520700CA08910000206101180803081144880010400044808000000122160",
INIT_03 => X"000080040305208000008000328080040304008020303194289A000041484800",
INIT_04 => X"08088000000000010000CA008008060441000000028234493410820191000000",
INIT_05 => X"03500404000022020020044000000C208400408000001000984005949C002928",
INIT_06 => X"54000881044500004680000013008002940C24001A4A010200018920646410C7",
INIT_07 => X"22510040400500011204813015012204002040280000013E1000000488000201",
INIT_08 => X"9001A0602C4A01051B132820208001024069004008908002120851420001226A",
INIT_09 => X"01100020A2401008A20404E08200A05000A4264640800022C8198C4E05200018",
INIT_0A => X"20002000024040400050450440C48A0041140C420B0904208800904286000008",
INIT_0B => X"50822002120D2134800648006480064800648106481064810648193240432404",
INIT_0C => X"284A142288042A5C24202451505E00A621A5220A8091444040188C001B41210A",
INIT_0D => X"00F001F021141A12004104020810B000100000000109064C80010050A3285194",
INIT_0E => X"00F001F027420000400004C3201C514408081C1014800000F001F02810148000",
INIT_0F => X"E00E0E404100E200040900000B0380383480C81014800000F001F02810148000",
INIT_10 => X"4160C0301D07001D0402034200004000019860078641004039000180400002C0",
INIT_11 => X"08103BA0104810C8462416E8040446120C890814600010512000000080028400",
INIT_12 => X"98038D4030DD008088C2419120B740209021908C4846FC000200030F000FE006",
INIT_13 => X"DD000100411C81078884204035DC00201804C3201C60A408100DD58010440130",
INIT_14 => X"412024202211148019064200402A32901A8000B2048902C0807C0E00C448100D",
INIT_15 => X"50942509425194651946519465894619421421102000269243854D8002000250",
INIT_16 => X"19465194E50942509425094E51946519465094A50942509425194E5194651942",
INIT_17 => X"9425094251946539465094250946539465194250942509465194650942509425",
INIT_18 => X"0000000000000000000000080150890820800041041000052942509465194653",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF21E6C000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"AAF7D5575455D557DFEF002AAAB55002E820AAAA800000000000000000000000",
INIT_1F => X"B55007FD74AAAA843DFEFA2FBD54BA5555554BAAAFBC20BA5D7BEAAAAFFFBC00",
INIT_20 => X"AA10FFFFFDE0008556AABA5D2ABFFEFFFAAAAAAAF7D57FFEFF7D555555A2AEAA",
INIT_21 => X"42145552ABDFEFFFAA801EFFFFBFDF550000175555504175450055574AAA2802",
INIT_22 => X"A975EF00003DF55555168A00000428AAAAA84021FF007BD54BAAAD17DEBA0855",
INIT_23 => X"802ABFF087FFDF5508003FEBA087FD54BA000415400557BD74BAFFD140000082",
INIT_24 => X"AFBE8ABAF7FFD54AAAAAEA8ABA55557FEAAA2843FF55A2AEA8B55AAAABDEAAFF",
INIT_25 => X"0000000000000000000000000000000000000051554BA002A95555A28417400A",
INIT_26 => X"25D7FE8A92FFFFC70BAE3D155555415178FD7082EAAB550820870BAAA8000000",
INIT_27 => X"FFEBD55557DBEA4AFB550871D7482AA8E3DFFFAAFFD04AA415B52492B6F5C208",
INIT_28 => X"5550051574BAB68A2DA00FFFFFFE38085F6FA92552AB8FEFF7A0ADABAEBD578F",
INIT_29 => X"2482BED57AE921451421555524BDFD7FFA4801D7F7F5FDF55000E17545410E17",
INIT_2A => X"D2482E3D1450381C20905EF08003AF55415F6DA38080E2DA82BE8E001EF147BD",
INIT_2B => X"AAFB55ABA0BDE02EB8A28BC70075FDF45080A3AEAA007BD24821C04124281C7B",
INIT_2C => X"209557DA28E15400BEF1EFA92FFFFD24BAB6A4A8A82495F78E92AA843DF45BEA",
INIT_2D => X"800174BAA680000000000000000000000000000000000000000000055524AA14",
INIT_2E => X"007BC0000FFD542000557FE8A00F3FFD54BAAAD15754508556AB45002AA8B450",
INIT_2F => X"FFB803DEAAAAD56ABEFAAD5575EFF7803DF45085557410AEAABDFEFAAFBC00BA",
INIT_30 => X"55082E97555002E955550C55554BAFFAEBDE10F7FBFDEBA007BFDE005D2AAABE",
INIT_31 => X"E00F7AA821FF557FC0010F7D168A105D554214551003FF45FF8400145FFD57FF",
INIT_32 => X"20105504000AA597FC2010A2D1554AA5500021EF000028B55087BFDEBA042ABF",
INIT_33 => X"E8A00A2803FF45F7AABDF55AA843FE10AEAAAAB4500557FF55082EA8AAA087FC",
INIT_34 => X"0000000055400BA5504155EFAAAE95410F7D57DE00FFFBC00AAFB8028A00007F",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000007FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(0),               -- Port A write enable input
DIA(0)   => data_write_a(7),        -- Port A data input
DOA(0)   => data_read_a_hi_512(7),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(0),               -- Port B write enable input
DIB(0)   => data_write_b(7),        -- Port B data input
DOB(0)   => data_read_b_hi_512(7),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_8_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000B0000040042840002C0000001800000070000000033022000000000086",
INIT_01 => X"000009C21838284D1C2160000E12426840000000180800080200080040510200",
INIT_02 => X"0001004000900110000006100080003000240800014400004808000000122160",
INIT_03 => X"00008000020440810002A0801010A0044300000000200086011A000040404800",
INIT_04 => X"8000801000020401400040408108022029400000124004041200000089000100",
INIT_05 => X"02080424085022020000040200480020850010A0002010010120060800040400",
INIT_06 => X"50000880006500000680000011008006840C200018C1010200018920E0640102",
INIT_07 => X"426000404005000112048130150120240020400A0000013E1000000488000010",
INIT_08 => X"220100402C42010413110020200100024029004000A200002004902200012141",
INIT_09 => X"0000000080400008010410A2940A45240040140440800022C8388E1200A00008",
INIT_0A => X"00420100020048405000070440C0000001140412090000000021002081000048",
INIT_0B => X"0000000800000100011000010000100001000010000100001000010000880008",
INIT_0C => X"001000040001100008012008004020102180800804802000C0080D00100A0008",
INIT_0D => X"0FF0000002200A1200410402080080003000091085100C008124008000400020",
INIT_0E => X"0FF000000140000040F517CF600000000104081010001E0FF00000001010001E",
INIT_0F => X"E000000000804200000809963F1F80000000001010001E0FF00000001010001E",
INIT_10 => X"CFE7C0F00000000000810140000040E587F9E000000008100900008000ED0FC7",
INIT_11 => X"00021040030C73D80000021000585F3600000020240020102000000802419660",
INIT_12 => X"F80000000042000B0BD6C0000010800618E7B000000C000003F80FFF00000000",
INIT_13 => X"800005D5C3FD800000000008180000078A8FCF600000000002028001006AA3F1",
INIT_14 => X"020000000008808219002100100C000041120370DCAD1FC18000000000000202",
INIT_15 => X"8020080200812048120481204812055A04604930A02026934215410102000110",
INIT_16 => X"0200802008020080200802048120481204812048120481204802008020080200",
INIT_17 => X"2008020081204812048120481200802008020080200802048120481204812048",
INIT_18 => X"414A87D78AF42143CEBAC88151120A0000000000000000081204812008020080",
INIT_19 => X"F3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF7E799B1BEB65B65948051",
INIT_1A => X"C3E9F0FA7C3E9F0FA7C3E9F0FA7C3E9F0F87C3E1F0F87C3E1F0F87CF3CF3CF3C",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF1B5DA9F0FA7C3E9F0FA7C3E9F0FA7",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"0000043DF55087BC01EF007FD75FFFF84000AAFF800000000000000000000000",
INIT_1F => X"E10A28028AAAAAFBC00AAF7D5575455D557DFEF002AAAB55002E820AAAA84000",
INIT_20 => X"54BA5555554BAAAFBC20BA5D7BEAAAAFFAA95545552ABFE00087BC00AA082EBF",
INIT_21 => X"D74AAAAD57FF45002A975FF007BE8BFFA2FBFFFFFAAD5400AAFF843DFEFA2FBD",
INIT_22 => X"BE8A00082A97410F7D5555EFAAAAAAAAAF7D57FFEFF7D555555A2AEAAB55007F",
INIT_23 => X"55574AAA2802AA10FFFFFDE0008556AABA5D2ABFFEFFFAA82000555555545AAF",
INIT_24 => X"00017555550417545000015545087BC2010AAD54014500516ABFFA2AABDF4500",
INIT_25 => X"000000000000000000000000000000000000002ABDFEFFFAA801EFFFFBFDF550",
INIT_26 => X"50820870BAAA8407000140038F450075C71FF087BD75D7FF84050BAEB8000000",
INIT_27 => X"10007FC50BA002ABFE00AA8A2AABABEFFC70BAE3D155555415178FD7082EAAB5",
INIT_28 => X"082EB8E3DFFFAAFFD04AA415B52492B6F5C20825D7FE8A92FFA497545552AB8E",
INIT_29 => X"557DBEA4AFB550871D7482AAD17DF451C24955EF0875EFBD7B6F1FFFC7BEDB45",
INIT_2A => X"87000415B5057DAAFBE8A10082092410EBD5505EFB6A0ADABAEBD578FFFEBD55",
INIT_2B => X"B6ABC7B6AABFFED0051574BAB68A2DA00FFFFFFE38085F6FA92552AB8FEFF7AA",
INIT_2C => X"A4801D7F7F5FDF55000E17545410E17555000E17545007BC0000BED14217D005",
INIT_2D => X"784174AAA280000000000000000000000000000000000000000000024BDFD7FF",
INIT_2E => X"08556AB45002AA8B450800174BAA684174105D042AB550055555FF007BD7555F",
INIT_2F => X"0F384175555D2EA8A00087BD74BA082EBDE10AAAEA8ABAF7FFD54BAAAD157545",
INIT_30 => X"55FFD57DF55FFFBD5400A2AABDFEFAAFBC00BA007BC0000FFD542000557FE8A0",
INIT_31 => X"EAAAAD56ABEFAAD5575EFF7803DF45085557410AED17FF455D04155FF00557DF",
INIT_32 => X"DE005D2AAABEFFBAE97410087BC21EFA2FFEAA00000002010A2D5421FFFF803D",
INIT_33 => X"C0010FFD1401EF087FE8B55FFAEBDFEF0855554BAFFAEBDE10F7FBFDEBA007BF",
INIT_34 => X"00000000003FF45FF8400145FFD57FF55082E97555002E955550C2E95555087B",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000020000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(1),               -- Port A write enable input
DIA(0)   => data_write_a(8),        -- Port A data input
DOA(0)   => data_read_a_hi_512(8),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(1),               -- Port B write enable input
DIB(0)   => data_write_b(8),        -- Port B data input
DOB(0)   => data_read_b_hi_512(8),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_9_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00018248A2840112C00002C18000002300500030B3132000400812002",
INIT_01 => X"A140098218302849180060000C004240413C0A61590001D90213C90008510204",
INIT_02 => X"102008700CB089100002061031285074810448800104008048080080001210E2",
INIT_03 => X"00008015074608840390A0040040800203140000A00010800408108448020042",
INIT_04 => X"082080400004A00100000100840602020100000002C2344156108201811801C0",
INIT_05 => X"0200048480011502049500280020CC2084000080008010019161249C9C002188",
INIT_06 => X"70000881004500004E01020411D08000940C00001800010200018B20206C0102",
INIT_07 => X"EA70C0040005000312048130150100040020404A0000017E10408104C8000110",
INIT_08 => X"000000402C220104131004202081120050A5104000A204617201D10801002000",
INIT_09 => X"000800002F4924003085E51420A0100400641E4E40800022C8088C1220200908",
INIT_0A => X"20102000024040484028450001648C2229150400080244000401900284000440",
INIT_0B => X"0880110901081110411204112040120411204012041120401204111020090208",
INIT_0C => X"685B34A688841A5C21200101A01A0004009024028004044248404D00104B2100",
INIT_0D => X"0000A01000000213000000000000B0001000010000190E44802002D1A168D0B4",
INIT_0E => X"0000A010014000000000000000000040500008100400000000A0100410040000",
INIT_0F => X"0000004608004200040000000000000001A004100080000000A0100410008000",
INIT_10 => X"00000000000024080000014000000000000000000040A0000900010000000000",
INIT_11 => X"300013E010000000000D00F804000000000340000C0000102000000080000000",
INIT_12 => X"00000040091F0000800000006807C000800000001A0CFC000000000000002001",
INIT_13 => X"DD000000000000000082C00019DC002000000000000021500006D58010000000",
INIT_14 => X"03206420000000C019502050000C32901A800080000000000000000860100006",
INIT_15 => X"D1B46D1B46D0B42D0B42D0B42D8B424342342832002A24921082158802001011",
INIT_16 => X"0B42D0B42D0B42D0B42D0B46D1B46D1B46D1B46D1B46D1B46D1B46D1B46D1B46",
INIT_17 => X"B42D0B42D1B46D1B46D1B46D1B46D1B46D1B46D1B46D1B42D0B42D0B42D0B42D",
INIT_18 => X"89999E91BCD1512B871C4A0100000000000000000000000D0B42D0B42D0B42D0",
INIT_19 => X"A28A28A28A28A28A28A28A28A28A29A69A69A69A69A51C200807249041202AE6",
INIT_1A => X"8349A4D068341A0D269341A0D269341A0D068341A0D068341A0D068A28A28A28",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF2DA921A0D269341A0D068349A4D06",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"45A280154BA5555401EFFFD5421EFA2FFFFF555D000000000000000000000000",
INIT_1F => X"5EF00557DF555D040000000043DF55087BC01EF007FD75FFFF84000AAFFD57DF",
INIT_20 => X"75455D557DFEF002AAAB55002E820AAAA843DFEF00517DEBA007BFDFEFFFD157",
INIT_21 => X"28AAAAAAABDF45F7803FFEF555568AAAF7802AA00FFFBD7555087BC00AAF7D55",
INIT_22 => X"BD54BA550417400085155555082A95545552ABFE00087BC00AA082EBFE10A280",
INIT_23 => X"043DFEFA2FBD54BA5555554BAAAFBC20BA5D7BEAAAAFFFBC00AA552E95545087",
INIT_24 => X"2FBFFFFFAAD5400AAFF8402000A2FFFDF555D7BE8BFF5D51575EFA280175555D",
INIT_25 => X"00000000000000000000000000000000000000557FF45002A975FF007BE8BFFA",
INIT_26 => X"7FF84050BAEBDF78F45B68010482415B471C7E3DF451EFBEFBFAF45490000000",
INIT_27 => X"82007FFAFEFE3DB505EF1C5B7AF45490407000140038F450075C71FF087BD75D",
INIT_28 => X"5451C7FC70BAE3D155555415178FD7082EAAB550820870BAAA8438FFF00517DE",
INIT_29 => X"50BA002ABFE00AA8A2AABABEAEB8F45F78A3DFD741516DAAAE38E2DA28EBFFD5",
INIT_2A => X"C20BA5D2E905550071D54825D0A1543808515756D1C2497545552AB8E10007FC",
INIT_2B => X"5505FFBE801256D490E3DFFFAAFFD04AA415B52492B6F5C20825D7FE8A92FFFF",
INIT_2C => X"24955EF0875EFBD7B6F1FFFC7BEDB45082EB8002000AAFFFDF6D417FEABEF5D5",
INIT_2D => X"7FBE8B5500000000000000000000000000000000000000000000000517DF451C",
INIT_2E => X"0055555FF007BD7555F784174AAA2FBEAB45F78402010007BD5545AAFFD55EFF",
INIT_2F => X"AA68028BEF00517FE10007BE8BFFAAFFC01FF557FE8B550004174105D042AB55",
INIT_30 => X"AAAAAEBFEAAAAFFD5545557FD54BAAAD15754508556AB45002AA8B450800174B",
INIT_31 => X"5555D2EA8A00087BD74BA082EBDE10AAAEA8ABAF7AAAAB45F7AEBFF4508557FE",
INIT_32 => X"2000557FE8A00F3FFC00BA552E80145005557400552A954BA0051575EF550417",
INIT_33 => X"FDFFF007FE8BFF5551401EFF784021FF002ABDFEFAAFBC00BA007BC0000FFD54",
INIT_34 => X"00000000517FF455D04155FF00557DF55FFD57DF55FFFBD5400A28400010A2FB",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000040000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(1),               -- Port A write enable input
DIA(0)   => data_write_a(9),        -- Port A data input
DOA(0)   => data_read_a_hi_512(9),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(1),               -- Port B write enable input
DIB(0)   => data_write_b(9),        -- Port B data input
DOB(0)   => data_read_b_hi_512(9),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_10_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00018248A2840112C00002C18000202300500030B3132000400992006",
INIT_01 => X"A140098218302849180060000C00424040000000080000080200090008510204",
INIT_02 => X"102100400C8001100000061000A8503401044880010400004808000000122160",
INIT_03 => X"000080150746088401908000100080020304000020201080001A108448404842",
INIT_04 => X"800080400004A001000040008406020201000000020004401000000180180080",
INIT_05 => X"02000484800133020495040800208C20A4000080000010000001249010042008",
INIT_06 => X"50000881004500004681020411808000940C20001800010200018920206C0102",
INIT_07 => X"024084044005000112048130150120040020400A0000013E10408104C8000010",
INIT_08 => X"000100402C020105131100200000124250A51040088084614001110801012000",
INIT_09 => X"00080082CD09240820800000000000040000180840800022C8088C1220200108",
INIT_0A => X"841201000200484910000F050560262229140402080200A00402000484140400",
INIT_0B => X"0010118900080010000200102001020000200002001020010200001000010008",
INIT_0C => X"408120900404004821202001F05E00040180260A8080044240004C0010800228",
INIT_0D => X"0000A01000000813004104020800800030000800010008088124020102008100",
INIT_0E => X"0000A010014000004000000000000040500008101480000000A0100410148000",
INIT_0F => X"0000004608004200040900000000000001A004101480000000A0100410148000",
INIT_10 => X"00000000000024080000014000004000000000000040A0000900018040000000",
INIT_11 => X"3800100010480000000D00000404400000034000282000102000000080028000",
INIT_12 => X"00000040090000808800000068000020900000001A0000000200000000002001",
INIT_13 => X"80000100000000000082E0001000002018000000000021580000800010440000",
INIT_14 => X"00004000000004C0195000500008000000000082008000000000000860180000",
INIT_15 => X"0100401004010040100401004090055804404110802A24921317580802001011",
INIT_16 => X"0000000000000000000000040100401004010040100401004010040100401004",
INIT_17 => X"0040100400000000000000000000000000000000000000000000000000000000",
INIT_18 => X"215281FC1A72E2486AAA40A85052020000000000000000001004010040100401",
INIT_19 => X"51451451451451451451451451451451451451451452AA83330A8A28A29EA8D1",
INIT_1A => X"5CA6532994CA6532B95CAE572994CA6532994CA6532994CA6532994514514514",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF31CE2E572994CA6532994CAE572B9",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"10AAFBE8AAAA2D540000F7D57DF55A2AABFFEF08000000000000000000000000",
INIT_1F => X"F45FFFBC2010AAD57DF45A280154BA5555401EFFFD5421EFA2FFFFF555D003FE",
INIT_20 => X"DF55087BC01EF007FD75FFFF84000AAFF8002155AAFFE8B45AAD540000087FFD",
INIT_21 => X"7DF555D517FEBA082A801EFF7FBD5400FFD568B555D00155EF08040000000043",
INIT_22 => X"BFDE00A2FBC0145005168A10AA843DFEF00517DEBA007BFDFEFFFD1575EF0055",
INIT_23 => X"7BC00AAF7D5575455D557DFEF002AAAB55002E820AAAA803FEBA082AAAAAAF7F",
INIT_24 => X"7802AA00FFFBD7555082E82155FFAEAAB55AAD568B455D00154BAFFFBD75EF5D",
INIT_25 => X"000000000000000000000000000000000000002ABDF45F7803FFEF555568AAAF",
INIT_26 => X"FBEFBFAF4549003DE10BEF5EDAAAAAD547038EBD57DF7DA2AEB8FC7000000000",
INIT_27 => X"6DAADF470280075FFF45E3F1C7038A2DF78F45B68010482415B471C7E3DF451E",
INIT_28 => X"5C7000407000140038F450075C71FF087BD75D7FF84050BAEB8002155BEF5EDB",
INIT_29 => X"AFEFE3DB505EF1C5B7AF45495B7DEAA0824851EFEBFBD2410EBD168B7D410A17",
INIT_2A => X"38EAA0824A8AAAEBF5FAE28AAF1C2155005F68A10A28438FFF00517DE82007FF",
INIT_2B => X"4104AAF7F1D75EF557FC70BAE3D155555415178FD7082EAAB550820870BAAA80",
INIT_2C => X"8A3DFD741516DAAAE38E2DA28EBFFD55451C2087155EBA4A8B7DAADF68B7D410",
INIT_2D => X"2AEAAB55000000000000000000000000000000000000000000000002EB8F45F7",
INIT_2E => X"007BD5545AAFFD55EFF7FBE8B5500043FE00F7D17FEBAA2D5574BAAAD17DFEFA",
INIT_2F => X"AA28002155FFD17FFFFA2FBD74BA00557FF45A2D5554AAA2FBEAB45F78402010",
INIT_30 => X"00AAD16ABFF002A975450004174105D042AB550055555FF007BD7555F784174A",
INIT_31 => X"BEF00517FE10007BE8BFFAAFFC01FF557FE8B55007FFDEAA0004175FFA2FBC20",
INIT_32 => X"8B450800174BAA68428AAA08042AABAAAD56AABAAAD140155087FEAA10A28028",
INIT_33 => X"2ABEFAAFBE8BFF0004020AAFFD5555EF557FD54BAAAD15754508556AB45002AA",
INIT_34 => X"000000002AAAB45F7AEBFF4508557FEAAAAAEBFEAAAAFFD5545550015555A284",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000047FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(1),               -- Port A write enable input
DIA(0)   => data_write_a(10),        -- Port A data input
DOA(0)   => data_read_a_hi_512(10),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(1),               -- Port B write enable input
DIB(0)   => data_write_b(10),        -- Port B data input
DOB(0)   => data_read_b_hi_512(10),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_11_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10180B05A0010402840602C2D001019000000300000000330A20080EC180002",
INIT_01 => X"AB400984B830084C1820E0000C36424840000000080000088200000802112220",
INIT_02 => X"102A68440080011000000618062AD03502640800010410424908136019920868",
INIT_03 => X"001282118644C88481908001106088022300000080F4925CDC9A10844A9A4842",
INIT_04 => X"401280480004A1011000418084460002E12000000200040010000040A8000000",
INIT_05 => X"0FC8048484011502059511488020802084400888001110000000050000005400",
INIT_06 => X"1011088AE24500001631024511C08004A70AA40008B90D0200018B60A0650D45",
INIT_07 => X"020011005405000910040150110041040024400D800002BE18408104C9205908",
INIT_08 => X"89390040280241041D175820000001020061004004800567403512A801014C46",
INIT_09 => X"050800E20D09A424C5840400808000040680180840800022D8288E946CA00833",
INIT_0A => X"85002000024040410A000D0504408C32E915D9C208050084840201A099100400",
INIT_0B => X"B01011934A005101431CA821CA831CA821CA831CA831CA821CA83165410E5410",
INIT_0C => X"00010080028000010402214850444091019B02080885200042A9CC001000003A",
INIT_0D => X"5A5018C5A0A00812004104020808B00030000808024008008325820000000000",
INIT_0E => X"5A5018C5AB0062C38A4DB680A0D8241500D5761B011986695014A96E1A811986",
INIT_0F => X"42056A289A1BB2078A922DA2A8B180A2600AAE1A811986695014A96E1B011986",
INIT_10 => X"05AA429189B60AC43C6C7F0272C3841DB528802CAB18468F4101621B1BAC8455",
INIT_11 => X"C003104289A668B8CAB270106338317A3D94392020224ACDE215883078681B5C",
INIT_12 => X"804B020A06020C67061BC785938085134CD551BCA1C90006C0C2958502861120",
INIT_13 => X"80819A5539D503336D61056ABA006282806CA64090B89E015AAA880E48382EB8",
INIT_14 => X"40000000E808989003066E03513E41470126C6284B2D20410AB4503089C00A82",
INIT_15 => X"0000000000000000000000000000041800400110200026124202500802000800",
INIT_16 => X"1004010040100401004010000000000000000000000000000000000000000000",
INIT_17 => X"0040100401004010040100401004010040100401004010040100401004010040",
INIT_18 => X"C110083018162148420840280050800000000000000000001004010040100401",
INIT_19 => X"000000000000000000000000000001041041041041003882928E0000000AA0C4",
INIT_1A => X"0000000000008040000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3E0FC000000000000020100000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"EFAA842ABEFA280155EFFFFBC01EF08554000055000000000000000000000000",
INIT_1F => X"F4508514000000003FE10AAFBE8AAAA2D540000F7D57DF55A2AABFFEF0804155",
INIT_20 => X"54BA5555401EFFFD5421EFA2FFFFF555D51575FFA2FFD75FF550015400FFFBFF",
INIT_21 => X"C2010AAD568AAAAAD142145FF80155EF0051555FF0804155FFF7D57DF45A2801",
INIT_22 => X"01540008514215555003DFFFA28002155AAFFE8B45AAD540000087FFDF45FFFB",
INIT_23 => X"040000000043DF55087BC01EF007FD75FFFF84000AAFF802ABFFA2AABFE10080",
INIT_24 => X"FD568B555D00155EF085168B45085142010FFAE800AA5D7BFDF45F7FFEAA0000",
INIT_25 => X"00000000000000000000000000000000000000517FEBA082A801EFF7FBD5400F",
INIT_26 => X"DA2AEB8FC70000175EFB6802DBC7BE8A155EFE3FBC71FF145B42038550000000",
INIT_27 => X"EF550E15400E3F1FFF7D085B420381C003DE10BEF5EDAAAAAD547038EBD57DF7",
INIT_28 => X"5C7F7DF78F45B68010482415B471C7E3DF451EFBEFBFAF45495F575FFBEF5D05",
INIT_29 => X"70280075FFF45E3F1C7038A2DB68ABAB6D145145FF84155D7085B555C7140410",
INIT_2A => X"28BEFBEA4BDE28140A1543800514515549003FFC7BE8002155BEF5EDB6DAADF4",
INIT_2B => X"FFFF7DE3F1EFA10140407000140038F450075C71FF087BD75D7FF84050BAEB84",
INIT_2C => X"24851EFEBFBD2410EBD168B7D410A175C7005B6DB55145140000FFAE85082417",
INIT_2D => X"57BC20AA5D0000000000000000000000000000000000000000000005B7DEAA08",
INIT_2E => X"A2D5574BAAAD17DFEFA2AEAAB550004175FFF7803DF45FFAE955EFAAFBD55EF5",
INIT_2F => X"5007FD75FFF7D5401EF5D2E97410AAD17DFEF007FC20AA5D043FE00F7D17FEBA",
INIT_30 => X"55007FD5545550400145FFFBEAB45F78402010007BD5545AAFFD55EFF7FBE8B5",
INIT_31 => X"155FFD17FFFFA2FBD74BA00557FF45A2D5554AAA2FBEAAAAFFD555545FF80155",
INIT_32 => X"7555F784174AAA2842ABEFFF803DEAA5D2E974AA00515754500003FF55FF8002",
INIT_33 => X"40000FFAE97410007BFFFFFA2D57FE105D04174105D042AB550055555FF007BD",
INIT_34 => X"000000007FFDEAA0004175FFA2FBC2000AAD16ABFF002A97545007FFFF455555",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000040000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(1),               -- Port A write enable input
DIA(0)   => data_write_a(11),        -- Port A data input
DOA(0)   => data_read_a_hi_512(11),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(1),               -- Port B write enable input
DIB(0)   => data_write_b(11),        -- Port B data input
DOB(0)   => data_read_b_hi_512(11),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_12_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50080B01BC002006940202C0DE041196A83183000000023322287E0FC000006",
INIT_01 => X"0E000C068000E04D40238000001702484000000008000008820009280A553231",
INIT_02 => X"400B71440C8001100000171C0283813013766A800586235ECC09C8423B962966",
INIT_03 => X"CC618E048306E082000081000040900003548421A080025EDF08421042DC0108",
INIT_04 => X"00028020000000812000012080080000E100001002000448100000C1BC18008C",
INIT_05 => X"0FF8060610000402010015E100004C2084800090000310000000079010007C19",
INIT_06 => X"33992D98DEC74A003EA468D01510C03E8F580C800A3F018200418927E0668645",
INIT_07 => X"0204000406050013142409121142F746222EE2498000007E111204058B84C50C",
INIT_08 => X"E826A0602902A10491165C200000820018A5104010C01086003C13E000004EDF",
INIT_09 => X"023000000000000867000000000000040000600060801022C9F88D244FA40133",
INIT_0A => X"00100000820040482B28050001600010C13499F01B334015980001E09F000000",
INIT_0B => X"B80460124F16F06BC20CBC30CBC20CBC20CBC30CBC20CBC20CBC3065E1865E10",
INIT_0C => X"00000000029D204B7C0382FD0100F3F9F80FA0200E0BF40063F99C0010000012",
INIT_0D => X"93900F6EE230301208008001007A80001100002002801000A042000000000000",
INIT_0E => X"93900F6EEC421392C96B1237E0D8BD9629F97E0B348EDAC3900F6EFA0B158EDA",
INIT_0F => X"622DBC31D73F6006A5891533EF9500EAE64BCA0B158EDAC3900F6EFA0B348EDA",
INIT_10 => X"C2B083798D341B10DEFE14400392C74CAEAD412EDD2B4FCFF812A383430C669E",
INIT_11 => X"49FAB442994B3238D4E2FB104636652E19B8BA30C022DAD8C100CA39E8CEBE66",
INIT_12 => X"30469392526208C6CC95C33717D88532966471A9C5DD00B12728D5360234D62A",
INIT_13 => X"828C4999AF580395542D27CDBA0020F0FABAC800DA550C29F36A8A2554E48A64",
INIT_14 => X"40000000873FB80B8A00EF03F56CC12B416A51B60585A5C28895962502E9F36A",
INIT_15 => X"0000000000000000000000000000008000000410802A26924010000002000EE0",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"28C1111026C152A121960A884042020000000000000000000000000000000000",
INIT_19 => X"2082082082082082082082082082092492492492492400200005A8A28A200A37",
INIT_1A => X"964B2592C964B2592C964B2592C964B2590C86432190C86432190C8208208208",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF400FEB2592C964B2592C964B2592C",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FF00042ABEFFF8400010082EAABFF55002ABEF08000000000000000000000000",
INIT_1F => X"BEFFFFBD54000004155EFAA842ABEFA280155EFFFFBC01EF0855400005555421",
INIT_20 => X"8AAAA2D540000F7D57DF55A2AABFFEF08556AA10000028AAAFFD15541000002A",
INIT_21 => X"40000005168AAA087BFFFFF5D04001FF00041554555557FE005D003FE10AAFBE",
INIT_22 => X"1555FF082AA8B55F7AEA8BEF5551575FFA2FFD75FF550015400FFFBFFF450851",
INIT_23 => X"D57DF45A280154BA5555401EFFFD5421EFA2FFFFF555D0000145082E955FF085",
INIT_24 => X"051555FF0804155FFF7842AA100000020BAAA801541055042ABEFFFFBD5410AA",
INIT_25 => X"000000000000000000000000000000000000005568AAAAAD142145FF80155EF0",
INIT_26 => X"F145B42038555F401D71C0A2DBC7EB80000280824ADBD7490E28BEF080000000",
INIT_27 => X"82FFDB5243800002FBD7EBFBD24101C00175EFB6802DBC7BE8A155EFE3FBC71F",
INIT_28 => X"E1041003DE10BEF5EDAAAAAD547038EBD57DF7DA2AEB8FC7005F6AA381C0A2DA",
INIT_29 => X"5400E3F1FFF7D085B420381C5B6AA82147FF8FEF410E001FF000E17555555B7A",
INIT_2A => X"0017D142E905EF1451525C7082AADB45F7AEA8BEF555F575FFBEF5D05EF550E1",
INIT_2B => X"02FBEFEBFBD2410AADF78F45B68010482415B471C7E3DF451EFBEFBFAF454900",
INIT_2C => X"D145145FF84155D7085B555C71404105C7F7842FA381C0A00082AA8A10410410",
INIT_2D => X"02AA8BEF000000000000000000000000000000000000000000000005B68ABAB6",
INIT_2E => X"FFAE955EFAAFBD55EF557BC20AA5D7BC01555D2EBFF55A284000AA08003FF550",
INIT_2F => X"5007BE8AAA5D2EBDE00FFFFC00AA08003FF55A2FBC00105D04175FFF7803DF45",
INIT_30 => X"FF082A97555557FE8A0000043FE00F7D17FEBAA2D5574BAAAD17DFEFA2AEAAB5",
INIT_31 => X"5FFF7D5401EF5D2E97410AAD17DFEF007FC20AA5D7BE8A005D7FEABFF002E821",
INIT_32 => X"55EFF7FBE8B550004001FF5D2A801EF5D5142145082EBFF55F7AAAABEF5D7FD7",
INIT_33 => X"82010A2AA8000008043FFFFA2FBC2010A2FBEAB45F78402010007BD5545AAFFD",
INIT_34 => X"000000007BEAAAAFFD555545FF8015555007FD5545550400145FF843DEAA552A",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000007FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(1),               -- Port A write enable input
DIA(0)   => data_write_a(12),        -- Port A data input
DOA(0)   => data_read_a_hi_512(12),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(1),               -- Port B write enable input
DIB(0)   => data_write_b(12),        -- Port B data input
DOB(0)   => data_read_b_hi_512(12),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_13_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10110A0441812402840402822007818000E00700000000330A3000000008042",
INIT_01 => X"A1400986B830E84D182260000C1042484001000008220008A20019080A510200",
INIT_02 => X"10A108600C9141100000C6180CA85035010E4880010431004908135980122D60",
INIT_03 => X"0013881507460886C190832175809C02030400002020124C441A108468424842",
INIT_04 => X"203080680204A0113801D600864E0C96C12000008244244052200201801802C0",
INIT_05 => X"030004849601110204950409C0208C2084E0009C0000100120A00C9918002098",
INIT_06 => X"10000882804544921681428591908000AF28A8002BC00D020003896020658FC4",
INIT_07 => X"CA20400450050009100501501102E0042020448D0000023E10408144C800D800",
INIT_08 => X"1D2B00402B220104B53100200001020218A5104016CC1C616401910801010100",
INIT_09 => X"050800404D49A42EB08000000000000406481C8C408000A2D8088D1820200B00",
INIT_0A => X"0010000002004048AA08050401604462E9144002090740148441200484000500",
INIT_0B => X"000A112100000000010000000001000000000000001000000000000000800000",
INIT_0C => X"509528954404144C200425010040000001B020081094040072005C0030864208",
INIT_0D => X"1C10B3831034081200000000000430003000206822F20CA8826AC2A14250A128",
INIT_0E => X"1C10B383110218CB0E54C2EA404A4F03D404A41AA5B7344C10B383081BA4B734",
INIT_0F => X"8001CE3E20A5B284ED1132909C72885A2B2C381BA4B7344C10B383081AA5B734",
INIT_10 => X"AC3CC0C0B8182597A801610218CB0C3548B3A008E730A01AB113A5524E6ACA67",
INIT_11 => X"A151EC5952E44128CA194517354C180A3C066430202021252991C22C99731014",
INIT_12 => X"1804C8A0ADA2E6A983014780CA28B2A5C8825194332B018A444AEA2701288A15",
INIT_13 => X"02D09852745F80112C428562EE0353635232D50048A411C158BB0A7910142C77",
INIT_14 => X"4240480068001C9B9150A0000297046E4023F8BE8E3E1E0109472C3EB50158BB",
INIT_15 => X"A1284A1284A1284A1284A1284A12851A84284110406A26924302590806000110",
INIT_16 => X"1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284",
INIT_17 => X"284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A",
INIT_18 => X"7DDFE7EFBEFFE7D3EFBEFC48A0550000000000000000000A1284A1284A1284A1",
INIT_19 => X"D75D75D75D75D75D75D75D75D75D75D75D75D75D75D7EFBFBFBBAAAAAABEFDF7",
INIT_1A => X"5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5D75D75D75",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000FEFD7EBF5FAFD7EBF5FAFD7EBF",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"AA5D043FFFFAAAABDEAA557BFDE00FFD140155F7800000000000000000000000",
INIT_1F => X"400AAD540155A2D5421FF00042ABEFFF8400010082EAABFF55002ABEF08556AA",
INIT_20 => X"ABEFA280155EFFFFBC01EF08554000055043DEBAF7843FFFFF7AABDF55A2AA97",
INIT_21 => X"D5400005568A1055043DEBAAAFFE8B45557FD7410552EAAABAAA84155EFAA842",
INIT_22 => X"FE8ABAAA8428A00087BD7555FFD56AA10000028AAAFFD15541000002ABEFFFFB",
INIT_23 => X"803FE10AAFBE8AAAA2D540000F7D57DF55A2AABFFEF085557545FFD17DEBAA2F",
INIT_24 => X"0041554555557FE005D0000155557BEAABA5D2ABDF450851420AA5D7FD5555A2",
INIT_25 => X"000000000000000000000000000000000000005168AAA087BFFFFF5D04001FF0",
INIT_26 => X"7490E28BEF08516DA82410A3FFD7AAA4B8E824971F8E38E3DF45155EB8000000",
INIT_27 => X"D7EBA4BDF45AAAA90410BEDF45155A2DF401D71C0A2DBC7EB80000280824ADBD",
INIT_28 => X"A82B680175EFB6802DBC7BE8A155EFE3FBC71FF145B42038550E38E92EB803FF",
INIT_29 => X"243800002FBD7EBFBD24101C556FA38490A3FE92BEFFEAB45417FD24385D2AAF",
INIT_2A => X"5056DE3D17FE92BEF1EFA92AA8428A10007FD557DFFDF6AA381C0A2DA82FFDB5",
INIT_2B => X"B400925D7FD557DA2803DE10BEF5EDAAAAAD547038EBD57DF7DA2AEB8FC70051",
INIT_2C => X"7FF8FEF410E001FF000E17555555B7AE10410E00155497FEFABA4120B8F55085",
INIT_2D => X"2FBD7545AA8000000000000000000000000000000000000000000005B6AA8214",
INIT_2E => X"A284000AA08003FF55002AA8BEF00517FE00082EBDF45AA8428A10085568ABAA",
INIT_2F => X"A5D2EA8A00A2803DF45AA843DF55AAAE82000F7FBD5545AAFBC01555D2EBFF55",
INIT_30 => X"55087FC00BA552ABFE10F784175FFF7803DF45FFAE955EFAAFBD55EF557BC20A",
INIT_31 => X"AAA5D2EBDE00FFFFC00AA08003FF55A2FBC00105D517FEAA082EBFE10F7FFE8B",
INIT_32 => X"DFEFA2AEAAB550051401FFA2D57FE10F7D57DE00AA842AA00007FD75FFF7FBE8",
INIT_33 => X"FDEAA08042AB45087FC0010557FD55FFAA843FE00F7D17FEBAA2D5574BAAAD17",
INIT_34 => X"000000007BE8A005D7FEABFF002E821FF082A97555557FE8A00002E82155007B",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000067FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(1),               -- Port A write enable input
DIA(0)   => data_write_a(13),        -- Port A data input
DOA(0)   => data_read_a_hi_512(13),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(1),               -- Port B write enable input
DIB(0)   => data_write_b(13),        -- Port B data input
DOB(0)   => data_read_b_hi_512(13),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_14_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10020A000180000284008280000281800000030000000033022000000580002",
INIT_01 => X"A14009821830284D186860000C30C24840000000084000084200090008510200",
INIT_02 => X"102100600C9001100000061020A8503401044880010400204908012018122F64",
INIT_03 => X"00008015074608840190800010008002030400002074F401209A108448404842",
INIT_04 => X"000080400004A00100004000840E000201000000024024401200020180180080",
INIT_05 => X"0A000484800111020495040800208C2084000080000010010020049818002008",
INIT_06 => X"1000088020450402B6A1420511C080008468A80008000D0200018B202067AF10",
INIT_07 => X"422000044005000910040110510260040024400C800000BE3850A144C924080E",
INIT_08 => X"000B004028020104111100200001020210A51040008004616001910801010000",
INIT_09 => X"000800004D492408208000000000000406401C0C40800022C8088DB420200900",
INIT_0A => X"0010000002004048000005040160042229140002090200000401000484000400",
INIT_0B => X"0000110100000000010000100000000000000100000000000000100000000000",
INIT_0C => X"409120940404104C2000210100400000011020080084040040005C0010820208",
INIT_0D => X"E0E0A0000190081200000000000000003000000000100C088020028102408120",
INIT_0E => X"E0E0A0000B02740421A0E5D1A024002050805210040000B0E0A0000210040000",
INIT_0F => X"E01200860008920106460D4501CB000111300210008000B0E0A0000210008000",
INIT_10 => X"0ABBC00905C33C6000400F02740412C0715C40110080A4006110510C14D18178",
INIT_11 => X"20000041DB011CC000090012565306500002411420220080220C0093C3892324",
INIT_12 => X"5809240C09024A4AE0CA00004800839682398000120800658992F3C700C30181",
INIT_13 => X"002B46867DBC002A830280000800F7B7A0B1E240240A8340000200067EAA8CB6",
INIT_14 => X"42004005800004801150A00341244000845C7DB0D0200900422ACA4B28000002",
INIT_15 => X"8120481204812048120481204812051A04204110002A26924302590802000000",
INIT_16 => X"1204812048120481204812048120481204812048120481204812048120481204",
INIT_17 => X"2048120481204812048120481204812048120481204812048120481204812048",
INIT_18 => X"69CB91FE1EF7D3ABEFBECA080050000000000000000000081204812048120481",
INIT_19 => X"F3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF7EFBBBBBF9E79E7BEAAF3",
INIT_1A => X"CFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCF3CF3CF3C",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FF007F3F9FCFE7F3F9FCFE7F3F9F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"45AAD157400007BEAAAAAAAE955555D5568A105D000000000000000000000000",
INIT_1F => X"0AAF784020AAF7D56AAAA5D043FFFFAAAABDEAA557BFDE00FFD140155F7D17DF",
INIT_20 => X"ABEFFF8400010082EAABFF55002ABEF085155400FFD1420100055574AAA2AA80",
INIT_21 => X"40155A28028B550051574005D7FFFE105D7BD7545A284020BA0055421FF00042",
INIT_22 => X"1421FF5D7FFDEBA085168B45FF843DEBAF7843FFFFF7AABDF55A2AA97400AAD5",
INIT_23 => X"04155EFAA842ABEFA280155EFFFFBC01EF08554000055002AB455D5142010085",
INIT_24 => X"57FD7410552EAAABAAA8017400AAD140000002EBFFEFA2AAA8BEFF780021FF55",
INIT_25 => X"000000000000000000000000000000000000005568A1055043DEBAAAFFE8B455",
INIT_26 => X"8E3DF45155EBD17FF6DAADB504001C71EDA82AAA0955455D556DA00490000000",
INIT_27 => X"101C55554AAAAA480082FF84000BAEBD16DA82410A3FFD7AAA4B8E824971F8E3",
INIT_28 => X"092085F401D71C0A2DBC7EB80000280824ADBD7490E28BEF085157428FFDB420",
INIT_29 => X"DF45AAAA90410BEDF45155A28E2AB7D0051504005D71F8E004975D556DB68405",
INIT_2A => X"28B6D5D51420101C5B401EF417BFAEAA08516AB45E38E38E92EB803FFD7EBA4B",
INIT_2B => X"EAFBC7EB80071FF5500175EFB6802DBC7BE8A155EFE3FBC71FF145B420385500",
INIT_2C => X"0A3FE92BEFFEAB45417FD24385D2AAFA82B68015400AADB40000082EBFFC7A2A",
INIT_2D => X"5557FE1000000000000000000000000000000000000000000000000556FA3849",
INIT_2E => X"AA8428A10085568ABAA2FBD7545AAD17DFFFAAFFC200055557DE00A280155455",
INIT_2F => X"F0051554AAFFFFC00105D55554BAA28400000F784020BAAAD17FE00082EBDF45",
INIT_30 => X"000051575FFF78415410087BC01555D2EBFF55A284000AA08003FF55002AA8BE",
INIT_31 => X"A00A2803DF45AA843DF55AAAE82000F7FBD5545AAAEAABFF0051400105D5568A",
INIT_32 => X"55EF557BC20AA5D042ABFF555142000557FC01EF007FEAABA00556AB55A2AEA8",
INIT_33 => X"C0010082EBDF55A2AABDF45A284175FF5D04175FFF7803DF45FFAE955EFAAFBD",
INIT_34 => X"00000000517FEAA082EBFE10F7FFE8B55087FC00BA552ABFE10F78415400A2FB",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000007FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(1),               -- Port A write enable input
DIA(0)   => data_write_a(14),        -- Port A data input
DOA(0)   => data_read_a_hi_512(14),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(1),               -- Port B write enable input
DIB(0)   => data_write_b(14),        -- Port B data input
DOB(0)   => data_read_b_hi_512(14),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_15_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000A000000000284000280000001800020030000000033022000000180002",
INIT_01 => X"A140098018300848180060000C00426040000000080000080200000000110200",
INIT_02 => X"1020004000801110000006100028503400040800010430004808000180120278",
INIT_03 => X"00008011064408840190800000228002A3000000000010000008108448000042",
INIT_04 => X"701280400004A991000000A28406000211000000220004941000000880000000",
INIT_05 => X"02000484800155020495000800218020C4002880005310000000040000000001",
INIT_06 => X"10000880004540000711224491C08000850A880008000D020001892020656300",
INIT_07 => X"8A04000016050009140501505100000420204008000000BE70408104C8000000",
INIT_08 => X"001F004028026104111002200000000200210040008004614001100801010000",
INIT_09 => X"000800000D09240000800000000000040600180840800022C8088C1020200000",
INIT_0A => X"0000000002004040000105000040042229140002080000000400000080000400",
INIT_0B => X"0000110100000000010000100001000010000000000000000000100000800008",
INIT_0C => X"0001008000000000000025000040000001300008009400006200580010000000",
INIT_0D => X"0000000002300012000000000004200030000000000008008020020000000000",
INIT_0E => X"0000000001000000400000000000000000000010108000000000000010108000",
INIT_0F => X"0000000000000200000900000000000000000010140000000000000010140000",
INIT_10 => X"0140000000000000000001000000400000000000000000000100008040000000",
INIT_11 => X"0000004000480000000000100004400000000030002000406000000000068409",
INIT_12 => X"8000000000020080080000000000802010000000000800000201000800000000",
INIT_13 => X"00000100000000000000000008000000184400A0000000000002000000441108",
INIT_14 => X"4000000000000000010620000004000000000242038B82800000000000000002",
INIT_15 => X"0000000000000000000000000000041800000110000024130202500802000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000080050000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"000804154AA5D00001EFF78428AAA007BC2145F7800000000000000000000000",
INIT_1F => X"0AA007FC2000F7D17DF45AAD157400007BEAAAAAAAE955555D5568A105D7FC00",
INIT_20 => X"FFFFAAAABDEAA557BFDE00FFD140155F7FBD74AAAAD17DF45F7D1421EF005540",
INIT_21 => X"020AAF7FFFDF45FF84000BA552ABDFEF08517DF55A2FBEAB555D556AAAA5D043",
INIT_22 => X"FEAB45F7843FF45082A801FF005155400FFD1420100055574AAA2AA800AAF784",
INIT_23 => X"D5421FF00042ABEFFF8400010082EAABFF55002ABEF087BE8ABA555168B55AAF",
INIT_24 => X"D7BD7545A284020BA007FFFE10A284000AA0055401550055574005D2E800AAA2",
INIT_25 => X"000000000000000000000000000000000000000028B550051574005D7FFFE105",
INIT_26 => X"55D556DA004971C7038140012482550E021C7EB8028A821C7BC516DFF8000000",
INIT_27 => X"45E3DF471C70851400BA0071C5028FFD17FF6DAADB504001C71EDA82AAA09554",
INIT_28 => X"B555D516DA82410A3FFD7AAA4B8E824971F8E38E3DF45155EBF1D5492BED17FF",
INIT_29 => X"54AAAAA480082FF84000BAEBF1FFF7DEB8000092552ABFFEF08517DF6DB6FBE8",
INIT_2A => X"EFA8241516DB55A2FFEAB6DEB843DF551C20801C71C5157428FFDB420101C555",
INIT_2B => X"550428412A85082BEDF401D71C0A2DBC7EB80000280824ADBD7490E28BEF087F",
INIT_2C => X"51504005D71F8E004975D556DB68405092087FF8E00BE8A02082005F47145085",
INIT_2D => X"57BD75EFF78000000000000000000000000000000000000000000000E2AB7D00",
INIT_2E => X"55557DE00A2801554555557FE100055554BA5504000105D2A80145AA842AA005",
INIT_2F => X"5AAD557410F7D57DF55AAFBD55450055420BA0055574BAF7D17DFFFAAFFC2000",
INIT_30 => X"FF08517FFFFF7FBEAB455D517FE00082EBDF45AA8428A10085568ABAA2FBD754",
INIT_31 => X"4AAFFFFC00105D55554BAA28400000F784020BAAAD57FFEFA28402010552ABDF",
INIT_32 => X"FF55002AA8BEF007FFDE1000557DF45AAFBE8BEFA2803FF45550400155555155",
INIT_33 => X"80000087BD55450855400BA002A95400F7FBC01555D2EBFF55A284000AA08003",
INIT_34 => X"000000002EAABFF0051400105D5568A000051575FFF78415410087FEAA10F7AE",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000060000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(1),               -- Port A write enable input
DIA(0)   => data_write_a(15),        -- Port A data input
DOA(0)   => data_read_a_hi_512(15),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(1),               -- Port B write enable input
DIB(0)   => data_write_b(15),        -- Port B data input
DOB(0)   => data_read_b_hi_512(15),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_16_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"DA22C618B1000482B688B186588884862A400438255FC38381441205BA803003",
INIT_01 => X"264AC80028404C211203A952A90341080B173340412000E1005D628000820484",
INIT_02 => X"400034C206C405000001A48202084004003008255040826EE008B440200E2042",
INIT_03 => X"2916704900606AC82B49CC56DF8CC1E50E4800202115005760010010000C0400",
INIT_04 => X"052DCA856DC7504B82BF6614C86D2B7F85AAD17F4B100000B88148C4804A428A",
INIT_05 => X"373CB02A00C0502F301180141A42A5720E0F43C17A8479580001AC20000000E2",
INIT_06 => X"303E2094282B85242C85001038D5710E8410D5959BC4800015001219D0550077",
INIT_07 => X"880100000159954501280B0080146F7112D949A0015018220540000382805001",
INIT_08 => X"30015452880C8D90409A05B2CB2CA400200209E5601044A24000000462A60018",
INIT_09 => X"452D54000C0907000330000000000096480050000685400005FC014743E0DC92",
INIT_0A => X"00014808A02004200E540480212000A448C0080024AEA00C9688000000000005",
INIT_0B => X"000D58460018F6D3D84400044000440004400044000440004400042000220002",
INIT_0C => X"0001004010A8812831605DA0000A054052E40000817680220040025699200002",
INIT_0D => X"AAADA0C343F1AC1B01040A002024895514554485D00000012400240000000000",
INIT_0E => X"AAADA0CC421CA003B694B68018FAAA708E2CB5320018CAC99BA0A3B9320018CA",
INIT_0F => X"B1443A1891E4A928C29020E6A8524CE7A3EE59320018CAC99BA0ACB9320018CA",
INIT_10 => X"04B2A5A40B1E6644AF0F021EA003AC24352AB2449A3FF2FA04E5E09B128834AD",
INIT_11 => X"60ED838E890B703C6260D8E3A21275714C902375B801324301AB0067622E5E54",
INIT_12 => X"064F70DBDB1C74424E91E1C194C71D1216F50A8C241815FEB6A9158863F638FB",
INIT_13 => X"45FDF9D364DBD9435A6D45C9E81BED555E4C15F11133D171727A2550EE2F1BA0",
INIT_14 => X"08150013F162119014204373517700ACCC59432A2B2D001F803471A9A960E572",
INIT_15 => X"000000000000000000000000000000880002054000229088542210206B2AB015",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"2A898D21B4C98389ED146C080000000000000000000000000000000000000000",
INIT_19 => X"A29A29A29A29A29A29A29A29A29A28A28A28A28A28A53CBF0F0D3CF3CF0AB1A2",
INIT_1A => X"8F47A3D1E8F4FA7D3E9F4FA7D3E9F4FA7D3E8F4FA3D3E8F4FA3D3E9A29A29A29",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000FA7D3E9F4FA7D1E8F47A3D1E",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFF7FBE8B45AAD568BFFFFAA975FF00003FE0055000000000000000000000000",
INIT_1F => X"0005D2A95410FFFFC00000804154AA5D00001EFF78428AAA007BC2145F7843FF",
INIT_20 => X"7400007BEAAAAAAAE955555D5568A105D2E974BAF7FBEAB45FFFFC00BAF78002",
INIT_21 => X"C2000F78000010552E800AA002E821FFA2AAAAA00000417555FFD17DF45AAD15",
INIT_22 => X"43FEBA5D55575FFF7AABFE00557BD74AAAAD17DF45F7D1421EF0055400AA007F",
INIT_23 => X"D56AAAA5D043FFFFAAAABDEAA557BFDE00FFD140155F7AABDF55F7AE820AA080",
INIT_24 => X"8517DF55A2FBEAB555D04154BAA2FBE8B55FFFFD55FF557FC2000FF8015410FF",
INIT_25 => X"000000000000000000000000000000000000007FFDF45FF84000BA552ABDFEF0",
INIT_26 => X"21C7BC516DFF8438FC7E3F1EAB55B6DF6DBFFF7AA955C71C043FE10490000000",
INIT_27 => X"55FFF1C70BAF78A000005D2097438FFF1C7038140012482550E021C7EB8028A8",
INIT_28 => X"57DEBD17FF6DAADB504001C71EDA82AAA0955455D556DA00492490492F7FBE8B",
INIT_29 => X"71C70851400BA0071C5028FF84020285D2085092002A801FFB6AAA8A10080E17",
INIT_2A => X"BAF6DE3AA8709208043FEBA555B555FFE3AABFE005D71D5492BED17FF45E3DF4",
INIT_2B => X"BC0028E38412428EBD16DA82410A3FFD7AAA4B8E824971F8E38E3DF45155EBA4",
INIT_2C => X"8000092552ABFFEF08517DF6DB6FBE8B555D04124BAB6FBE8B45E3FBD55D7557",
INIT_2D => X"5003DE000000000000000000000000000000000000000000000000071FFF7DEB",
INIT_2E => X"5D2A80145AA842AA00557BD75EFF78428B55AAD168B55F7FFFDFEFFFAA955555",
INIT_2F => X"0000000010F7FBEAB45FFD1554AAFFAE820105500154AAF7D5554BA550400010",
INIT_30 => X"EFF7AEA8A10002E955FFA2D17DFFFAAFFC200055557DE00A2801554555557FE1",
INIT_31 => X"410F7D57DF55AAFBD55450055420BA0055574BAF784000BA5D0017410082E801",
INIT_32 => X"8ABAA2FBD7545AA802ABEFA2AA9541000003DEBA557BD75EFA2AEBDE105D5557",
INIT_33 => X"EAB45AAFFD55555D7FC20AAA280000AAAAD17FE00082EBDF45AA8428A1008556",
INIT_34 => X"00000000557FFEFA28402010552ABDFFF08517FFFFF7FBEAB455D04020AAFFFB",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000020000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(2),               -- Port A write enable input
DIA(0)   => data_write_a(16),        -- Port A data input
DOA(0)   => data_read_a_hi_512(16),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(2),               -- Port B write enable input
DIB(0)   => data_write_b(16),        -- Port B data input
DOB(0)   => data_read_b_hi_512(16),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_17_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"5284CE4FB7BD2C8994A13392DBD02E14006B82AC7E800D44D3DD2FD5F9B961C0",
INIT_01 => X"F9BA301F7E03FC6793F2199B39FC233C11D93AE6F3BB92B32091DBC339B24542",
INIT_02 => X"1D5FC0C08F040404446965C0607FB8A217C400C33A908078551BD04222186338",
INIT_03 => X"A14124C28DFD960832C90446DF8400A5055C25295B695FF97E1B5AC757F06D6B",
INIT_04 => X"04A106866DA3D02A01FB660C08A4AB7F840EDB6F48100DFC8081081D78AC7402",
INIT_05 => X"51E072F0C0C58D9C125EBFC00A46CF0388054100F680E0CE0107B8D040DAFCDA",
INIT_06 => X"019A4D00786B048112C58B16307F15DE8408B233661C10BBA5DAAFA9DDA1194D",
INIT_07 => X"8E00001660700CE170284A00891C7C03D29DE26814515835902AC089A2801540",
INIT_08 => X"C009F3A1B0120A1C51DFF881861CBE0305A12A0321810217C01D34EDC98FFA1C",
INIT_09 => X"747E6610052CDEE97FF1F9F63E3EF790380078002CE976AB6BF769769E4D437D",
INIT_0A => X"00185C44B91BC1740B7605040BE0018CFC7429F326B9D045FF8000E9AB415606",
INIT_0B => X"3A28FC1AAF5CF6F3D3EF3D3EF3D3EF3D3EF3D3EF3D3EF3D3EF3D3EF9E9F79E9E",
INIT_0C => X"0000020012E9E10A31EB5FF9296A67F5B4FFBD2FAD7FE653C3FBFF33E10C001B",
INIT_0D => X"333EA16031F2BD47BDA2CA5D8164FCCFE833C5C3D00018006C68170000000000",
INIT_0E => X"333EA160391BEFF2C32FB695F919110D5ECE542A6FEEB2533EA160782A6FEEB2",
INIT_0F => X"D18C0D06638A207CFDE1F7DDAD76D5282400F82A6FEEB2533EA160782A6FEEB2",
INIT_10 => X"E6E43E59AFE4A59B57679D19EFF2C7573FAD5A86840354D1706FFFA3EF6E24B6",
INIT_11 => X"F7D7A0ABD6DAAAB96529382B74E4E1FE4ACA4D77FAAB77CE3AF3EE78F58DB737",
INIT_12 => X"2D1281017F056E9C9C3FC95949C157ADB55572CA52606DFED6CA55334C04C04F",
INIT_13 => X"59FDEB974F486905001FDF5FA0D719F9956EAA1A184045D5D7A870D2F5A5D752",
INIT_14 => X"60158015177F916A039EF41FDB34A91F432EA58949D5B5C85F97871876F7D7E8",
INIT_15 => X"000000000000000000000000000004DC200005E705B7B3D9FC22F00BE419FB55",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"06013DB9880A5D22E229F3030018000000000000000000000000000000000000",
INIT_19 => X"D35D74D35D74D34D35D74D35D74D34D34D34D34D34D0D30D0D303AEBAE886E40",
INIT_1A => X"51A8D46A351A0D068341A0D068341A0D068341A8D468341A8D46834D35D74D34",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000008D46A351A8D46A351A8D46A3",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFF7FBFDF55A28402000F7D56ABFF55000000000000000000000000",
INIT_1F => X"A00F7843FEBA55043FFFFF7FBE8B45AAD568BFFFFAA975FF00003FE0055043FF",
INIT_20 => X"54AA5D00001EFF78428AAA007BC2145F7D568B45000002010552EBDF45A28028",
INIT_21 => X"95410FFAE800105D2A95410002A95410AAAEBFF55AAFFC00BAF7FFC000008041",
INIT_22 => X"57DE00F7AE800AAAAAABDFEF5D2E974BAF7FBEAB45FFFFC00BAF780020005D2A",
INIT_23 => X"517DF45AAD157400007BEAAAAAAAE955555D5568A105D7FFFFEFA2D568BFFFFD",
INIT_24 => X"2AAAAA00000417555FF8028B55082A974105D003FF55F7802AAAAAAD168AAA5D",
INIT_25 => X"000000000000000000000000000000000000000000010552E800AA002E821FFA",
INIT_26 => X"71C043FE10490A3FFFFFFFFFDFEFE3F5FAF45AA8000038F7DB6FBD7490000000",
INIT_27 => X"384124BFF7DB68A28A38F7803DE82490438FC7E3F1EAB55B6DF6DBFFF7AA955C",
INIT_28 => X"0BAFFF1C7038140012482550E021C7EB8028A821C7BC516DFFDF68B551C0E050",
INIT_29 => X"70BAF78A000005D2097438FFAA85000492495428082E95400AAA0BDF7DB6F5C7",
INIT_2A => X"FAFFFB6D56FBFFEBDB78E38F7AA800BAB6AEBDFD75D2490492F7FBE8B55FFF1C",
INIT_2B => X"028AAAB6D16FA8249517FF6DAADB504001C71EDA82AAA0955455D556DA00497F",
INIT_2C => X"2085092002A801FFB6AAA8A10080E1757DEB8A2DB5514249243841003FF6DEB8",
INIT_2D => X"7FFFDF550000000000000000000000000000000000000000000000004020285D",
INIT_2E => X"F7FFFDFEFFFAA9555555003DE00002ABFFEFF7FBFDFFFAAD168B55AA80000BAF",
INIT_2F => X"FF7FBEAB45552E954BA08003DFFFFFAAA8AAAF7843FE10000428B55AAD168B55",
INIT_30 => X"10AA843FFFFF7D5554BAF7D5554BA5504000105D2A80145AA842AA00557BD75E",
INIT_31 => X"010F7FBEAB45FFD1554AAFFAE820105500154AAF7AE974000800154AA002E954",
INIT_32 => X"554555557FE10007FEABEFFFD57FFEFAAFFE8ABAFFAA820BAF7AEBFF55550000",
INIT_33 => X"020AA08003DFFFA28028AAAF7D17DE0000517DFFFAAFFC200055557DE00A2801",
INIT_34 => X"0000000004000BA5D0017410082E801EFF7AEA8A10002E955FFA2AABFF455500",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000067FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(2),               -- Port A write enable input
DIA(0)   => data_write_a(17),        -- Port A data input
DOA(0)   => data_read_a_hi_512(17),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(2),               -- Port B write enable input
DIB(0)   => data_write_b(17),        -- Port B data input
DOB(0)   => data_read_b_hi_512(17),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_18_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"69844019080000A21A611406840014122A641074155FC28A2024001001801003",
INIT_01 => X"01067920034004180005E9E3C90360C0041C0181002001602025800008440084",
INIT_02 => X"40AC3CAA22D605200000856E2481902400344A20F802C22054001000021E2379",
INIT_03 => X"A95308ECD3207AC81D91C4002004C08A06008080BA868007E58040102B0E0100",
INIT_04 => X"044CC183800CA00780808004C8DB841405A80A100B586200FAC24AE4805242CA",
INIT_05 => X"771C10000000000B1135883C08A115320E0401C0200038394230070A19000020",
INIT_06 => X"3001499C602A8A003E800A042D8132A00098408F79E3901218050018024110D6",
INIT_07 => X"5029401000C983E60004010030400353C05806800104004E0000042E52800E20",
INIT_08 => X"0000117088080990419005B0C309402030060860E01004A828408800440405E3",
INIT_09 => X"6B8186185C42900693A002004040001E1950850C848601008708114A2030B480",
INIT_0A => X"100180A8062026000DC425C0301311324AA237108857220BA089420440000030",
INIT_0B => X"C44703657083080C2800C2000C2000C2000C2000C2000C2000C2000610006100",
INIT_0C => X"C1B0609C05013065CC042004040808084001E000108010230400800FD9B286C4",
INIT_0D => X"CCC15F9CBA45505640000A402019003F140FC2060014250B9080008306C18360",
INIT_0E => X"CCC15F9FB1962FCB69E08AAAEAEBCDDF7C728582081483ACC15F9C3982081483",
INIT_0F => X"EBF1CFFF7670ACC3811A28AB57523CDFEBFBF982081483ACC15F9F3982081483",
INIT_10 => X"C9002BF05800D875E63CC9962FCB52CAA02FE3F8E7F5E3AC3620805298B15A3F",
INIT_11 => X"F1B72A8A800B7546DB9F1CA320037F01BD67DC4041D4CF03138DD865103EFEEA",
INIT_12 => X"81CCFAFDBF9464006FD037AEFAE5150016EA8DB7BFE25208E8F46A228BF8A757",
INIT_13 => X"641256EC844B8AF92FD7CEDC24A9E181A8A29509EAAE7FD3B749471C48F8A459",
INIT_14 => X"0297D086E00036D2440E0880AAD62BEFF5778802A3AF8E8FB0440CE78773B709",
INIT_15 => X"8360D8360D8360D8360D8360D83609220D20D00000080C0601400B402307E480",
INIT_16 => X"360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D",
INIT_17 => X"60D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8",
INIT_18 => X"D9D701DC2E784601EFBE2C00000000000000000000000008360D8360D8360D83",
INIT_19 => X"5155555545145145155555545145145145145145145220B22A0B820820965177",
INIT_1A => X"44A25128944A25128944A25128944A25128944AA552A954A2512895554514514",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000025128944A25128944A251289",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFEFF7AE954BA5D04174AA00000000000000000000000000",
INIT_1F => X"145AA801741000043FFFFFFFFFFFFFF7FBFDF55A28402000F7D56ABFF55043FF",
INIT_20 => X"8B45AAD568BFFFFAA975FF00003FE0055043FFFFFFFFFDFEFA2D56AB45AA8400",
INIT_21 => X"3FEBA55557FFEFA2D168B55AAFBFFFFFFF80021EF0855421EF00043FFFFF7FBE",
INIT_22 => X"A82155F7AEBFEBAFFD56AA00A2D568B45000002010552EBDF45A28028A00F784",
INIT_23 => X"FFC00000804154AA5D00001EFF78428AAA007BC2145F7D5400000004020AA5D2",
INIT_24 => X"AAEBFF55AAFFC00BAF7AE80010082E954BA0004174AAAA8428B45082ABFEBAA2",
INIT_25 => X"000000000000000000000000000000000000002E800105D2A95410002A95410A",
INIT_26 => X"8F7DB6FBD7490E3FFFFFFFFFFFFFFFFBFDFEFFFAE954AA550415492140000000",
INIT_27 => X"D7AAD16FB6DBE8E00155BE8015410140A3FFFFFFFFFDFEFE3F5FAF45AA800003",
INIT_28 => X"1C7140438FC7E3F1EAB55B6DF6DBFFF7AA955C71C043FE1049043FFEFE3F1F8F",
INIT_29 => X"FF7DB68A28A38F7803DE82495B78FC7AAD56FB6DBEF1FAFD7E384001EF145B47",
INIT_2A => X"420381C0A02082492A85155E3A4BDE92FFD56FA28B6DF68B551C0E050384124B",
INIT_2B => X"E28B7D1420BDEAAA2F1C7038140012482550E021C7EB8028A821C7BC516DFFD1",
INIT_2C => X"2495428082E95400AAA0BDF7DB6F5C70BAFFAE870280024904BA1400174AABE8",
INIT_2D => X"50415410550000000000000000000000000000000000000000000002A8500049",
INIT_2E => X"AAD168B55AA80000BAF7FFFDF55002ABFFFFFFFFFFFEFF7FBFDFFFF7AA974BA5",
INIT_2F => X"000043DFEFA2D56AB45AAD57DFEFF7AA82155F78015400552ABFFEFF7FBFDFFF",
INIT_30 => X"55A280021EF557FD7555550428B55AAD168B55F7FFFDFEFFFAA9555555003DE0",
INIT_31 => X"B45552E954BA08003DFFFFFAAA8AAAF7843FE10007FEAB55A2D17FFEFFFD568B",
INIT_32 => X"AA00557BD75EFF7D1400AA5D2A82000002A95545A2843FE00F7D17FEAAF7FBEA",
INIT_33 => X"020AA5D04154BAF7AEA8BEF55003DEAAA2D5554BA5504000105D2A80145AA842",
INIT_34 => X"000000002E974000800154AA002E95410AA843FFFFF7D5554BAF7AE974BA0004",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000020000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(2),               -- Port A write enable input
DIA(0)   => data_write_a(18),        -- Port A data input
DOA(0)   => data_read_a_hi_512(18),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(2),               -- Port B write enable input
DIB(0)   => data_write_b(18),        -- Port B data input
DOB(0)   => data_read_b_hi_512(18),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_19_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"042200000000000041088001001AA00000000000000000000000500802000003",
INIT_01 => X"074018000024000000000404000000000A22000800000800004A200000000001",
INIT_02 => X"0000048002C405000000000006A84000000000200893C246A20000000020031A",
INIT_03 => X"020A9639044012C80001C4000004C08006000000001025000000000000000000",
INIT_04 => X"0400C0800000000380800004C8000000058800000B1000009880480480024200",
INIT_05 => X"420410000000000B10804004080001320E0401C0200038080000000000000000",
INIT_06 => X"2002409006F00A8428050A000280493104004500480090080A01120220140020",
INIT_07 => X"0000000000418026090240923240002190400000000000C0054A912054004021",
INIT_08 => X"0000115080000990000000B0C308000000000860200160000000000038380000",
INIT_09 => X"8000F80001012590001000000000001618000000020280008180810200000000",
INIT_0A => X"0000000000000000000000000000000100008000110000000000000000000017",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000840007600000000000000000800259000000",
INIT_0D => X"0008A0034078104B41A41000000000031400C002000000000000000000000000",
INIT_0E => X"0008A0004263C0343EDD414004042228DC0D385598035D0008A003B05598035D",
INIT_0F => X"040231068187C39F5A4F985C008902041124505598035D0008A000B05598035D",
INIT_10 => X"1BFBD406451B02000E033263C0343CB740500401180DE053A98F6ECC739D8140",
INIT_11 => X"420851546B2400000040D8549B5800000010227848D4303807FC8CC5508AEAED",
INIT_12 => X"52210402120A936B0000000004C2A8D6480000000018A700FCF980CC300318A2",
INIT_13 => X"B1427ED430B41402D025082359700181C21140E40511802208D6B30C48F8A8A4",
INIT_14 => X"9C000018440021011821B35254E99AF9E9410006362A2B6424287B08286208D6",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000023006000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"7747E18E0218CC18E88324000000000000000000000000000000000000000000",
INIT_19 => X"34C30C30C30C30D34C30C30C30C30C30C30C30C30C3504118982A69A6980E411",
INIT_1A => X"C26130984C26130984C26130984C261309A4D26130984C26130984C30C30C30D",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000130984C26130984C26130984",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAA954BA5500020BA5D000000000000000000000000",
INIT_1F => X"4BA5D517FFFF08043FFFFFFFFFFFFFFFFFFFFEFF7AE954BA5D04174AA007BFFF",
INIT_20 => X"FFFFF7FBFDF55A28402000F7D56ABFF557BFFFFFFFFFFFFFFFFFBFDFEFFFAA97",
INIT_21 => X"17410007BFFFFFFFFFFFFEFF7D16AB45AA8002000F7D5575455D043FFFFFFFFF",
INIT_22 => X"568B55F7AE955FFAA840201008043FFFFFFFFFDFEFA2D56AB45AA8400145AA80",
INIT_23 => X"043FFFFF7FBE8B45AAD568BFFFFAA975FF00003FE00557BFFFFFFFFBFDF45AAD",
INIT_24 => X"F80021EF0855421EF002ABFFEFF7D168B55AAD17FFEFF7AE975FF00557FFFF5D",
INIT_25 => X"00000000000000000000000000000000000000557FFEFA2D168B55AAFBFFFFFF",
INIT_26 => X"A5504154921471FFFFFFFFFFFFFFFFFFFFFFFF7AA954BA550000082550000000",
INIT_27 => X"EFF7FBFAFD7E3A4954BA555B7AFC7080E3FFFFFFFFFFFFFFFFBFDFEFFFAE954A",
INIT_28 => X"545550A3FFFFFFFFFDFEFE3F5FAF45AA8000038F7DB6FBD74975FFFFFFFFFFFF",
INIT_29 => X"FB6DBE8E00155BE8015410147FFFFFFF7FBF8FC7EBD568B55A28000000FFDF52",
INIT_2A => X"FDFC7E3F1FAF55A2DB6FB7DF7AE955C7BE800000008043FFEFE3F1F8FD7AAD16",
INIT_2B => X"0955FF145B7AFC7410438FC7E3F1EAB55B6DF6DBFFF7AA955C71C043FE10497B",
INIT_2C => X"D56FB6DBEF1FAFD7E384001EF145B471C71424B8FC7E3D56AB6DB6DF7AFC7EBA",
INIT_2D => X"50002000550000000000000000000000000000000000000000000005B78FC7AA",
INIT_2E => X"F7FBFDFFFF7AA974BA55041541055517FFFFFFFFFFFFFFFFFFFFEFF7AA974AA5",
INIT_2F => X"500517FFFFFFFBFDFEFFFFFEAB45AA80154AA557BEAB45002ABFFFFFFFFFFFEF",
INIT_30 => X"55A28002000F7FFC2155552ABFFEFF7FBFDFFFAAD168B55AA80000BAF7FFFDF5",
INIT_31 => X"FEFA2D56AB45AAD57DFEFF7AA82155F78015400557BFDFEFF7FBEAB55A2D56AB",
INIT_32 => X"555555003DE00007FFDF45AAD568B45AAFBFFFFFFFAA95545F7840201000043D",
INIT_33 => X"6ABFFFFFBEAB45A280155EF557FE8B55000428B55AAD168B55F7FFFDFEFFFAA9",
INIT_34 => X"000000007FEAB55A2D17FFEFFFD568B55A280021EF557FD755555042AB55AAD1",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000040000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(2),               -- Port A write enable input
DIA(0)   => data_write_a(19),        -- Port A data input
DOA(0)   => data_read_a_hi_512(19),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(2),               -- Port B write enable input
DIB(0)   => data_write_b(19),        -- Port B data input
DOB(0)   => data_read_b_hi_512(19),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_20_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000003",
INIT_01 => X"A65FF80000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000048002CC070000000000000000000000002FF86100200000000220002362",
INIT_03 => X"00000000000203D80025DC18004DC3D01E000000000000000000000000000000",
INIT_04 => X"07E5DF808071026F87C4191DD8005080679800000F300002998058068002C000",
INIT_05 => X"C205F23A2100557F70000004390021F61E1E87C3FD0CFBF80880072042000044",
INIT_06 => X"1209244C2000100006800000020010000008407FC800B0000000100600040000",
INIT_07 => X"8802000009FFBFE51886018002040020000800000554003E0000000002800000",
INIT_08 => X"30801F5780259FB0000000F7DF78020004011FEFE00000000020031502000083",
INIT_09 => X"00000000001000000000000000000056F8000001000000040000040141800802",
INIT_0A => X"0000000000000008000800000000000000000000000000000010010014800000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"00010240001721214E000004000000080000008000001000040080FFDB000000",
INIT_0D => X"0000000F3008001E00000000001803FF14FFC006000000008010200000000000",
INIT_0E => X"0000000F3040200000020000000026A70C0008020000200000000F3002000020",
INIT_0F => X"000030B86000400080000200000000004A58F0020000200000000F3002000020",
INIT_10 => X"0000000002183E61E6000040200001000000000019B140000800800000020000",
INIT_11 => X"C00010080000000000525801000000000014AC08000000508001030A0A400100",
INIT_12 => X"000002BC360020000000000292C0100000000000A56000090100000000001F86",
INIT_13 => X"8010000000000000574500001001060600000000001716800000803102020000",
INIT_14 => X"00000000000040040040002000080506049CDF70C08040100000706707600000",
INIT_15 => X"00000000000000000000000000802040200200604040000000000024FB7FE008",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"060070400020112240209A408004000000000000000000000000000000000000",
INIT_19 => X"65965965965965965965965965965861861861861860D30424343CF3CF340E00",
INIT_1A => X"90C86432190C86432190C86432190C86432190C86432190C8643219659659659",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000086432190C86432190C864321",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974AA55040201008000000000000000000000000",
INIT_1F => X"4AA550002000007BFFFFFFFFFFFFFFFFFFFFFFFFFAA954BA5500020BA5D7FFFF",
INIT_20 => X"FFFFFFFFFFFEFF7AE954BA5D04174AA00003FFFFFFFFFFFFFFFFFFFFFFF7AA97",
INIT_21 => X"7FFFF087FFFFFFFFFFFFFFFFFFFFDFEFFFAE974AA5D003FE005D043FFFFFFFFF",
INIT_22 => X"BFDFFFAA84000105D556AB55557BFFFFFFFFFFFFFFFFFBFDFEFFFAA974BA5D51",
INIT_23 => X"043FFFFFFFFFFFFFF7FBFDF55A28402000F7D56ABFF55003FFFFFFFFFFFFFF7F",
INIT_24 => X"A8002000F7D5575455D2EBFFFFFFFFFFFEFF7FBEAB55A28000010F7D16ABEF08",
INIT_25 => X"000000000000000000000000000000000000007BFFFFFFFFFFFFEFF7D16AB45A",
INIT_26 => X"A550000082557FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550400028000000000",
INIT_27 => X"FFFFFFFDFEFF7AE974BA5500050380071FFFFFFFFFFFFFFFFFFFFFFFF7AA954B",
INIT_28 => X"E285D0E3FFFFFFFFFFFFFFFFBFDFEFFFAE954AA55041549214043FFFFFFFFFFF",
INIT_29 => X"AFD7E3A4954BA555B7AFC70871FFFFFFFFFFFFFFF7FBFDFFFFFAA974BA550038",
INIT_2A => X"3FFFFFFFFFDFEFF7F1FAFC7A28002028555F6FB7D5D75FFFFFFFFFFFFEFF7FBF",
INIT_2B => X"402010FFDB6ABEF140A3FFFFFFFFFDFEFE3F5FAF45AA8000038F7DB6FBD7490E",
INIT_2C => X"FBF8FC7EBD568B55A28000000FFDF525455524BFFFFFFFBFDFC7E3F5E8B45A28",
INIT_2D => X"504000BA080000000000000000000000000000000000000000000007FFFFFFF7",
INIT_2E => X"FFFFFFFEFF7AA974AA550002000557FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5",
INIT_2F => X"055043FFFFFFFFFFFFFF7FBFDFEFFFAE954BA5500174AA08517FFFFFFFFFFFFF",
INIT_30 => X"EFF7AE974AA550028AAA5D2ABFFFFFFFFFFFEFF7FBFDFFFF7AA974BA55041541",
INIT_31 => X"FFFFFFBFDFEFFFFFEAB45AA80154AA557BEAB4500557FFFFFFFFFDFEFF7FFFFF",
INIT_32 => X"00BAF7FFFDF55002EBFFFFF7FBFDFEFFFD568B55A284020BA557FFFFFF5D517F",
INIT_33 => X"FFF55A2D16AB45AA8402000F7FBEABEF5D2ABFFEFF7FBFDFFFAAD168B55AA800",
INIT_34 => X"000000007BFDFEFF7FBEAB55A2D56AB55A28002000F7FFC215555043DFEFF7FB",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000007FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(2),               -- Port A write enable input
DIA(0)   => data_write_a(20),        -- Port A data input
DOA(0)   => data_read_a_hi_512(20),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(2),               -- Port B write enable input
DIB(0)   => data_write_b(20),        -- Port B data input
DOB(0)   => data_read_b_hi_512(20),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_21_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"4A302428B824900A128C090A5C1800261500213C005FE812D10420054085A202",
INIT_01 => X"081FFE3440B609703B0427F801A40B8115BC4F655300340288A40D30040E4DD8",
INIT_02 => X"04CA478082CC1740002019824E0203100640303FF8C0B31061096E21A1840814",
INIT_03 => X"230CA7A4810083F80095DE00102DC3823EA821094EC68248923200013290C800",
INIT_04 => X"07CFFFC04904AA7F8780409DF84A0202879800000F3000029980780EA2C3C002",
INIT_05 => X"DE87F0280000407FF900D914382091FE1E1C0FC3E01EFFF8000480200008D062",
INIT_06 => X"010E2182002BC107A03448808F0D7C002822987FC830F40134CC74D002016612",
INIT_07 => X"0401000011FBFFE00520000200422033025C4209104500000012004C004D8C0B",
INIT_08 => X"00EF1F5FA0041FF080AC70FFDF78220010841EFFE7116E144071268DFD3E4C24",
INIT_09 => X"FC8BFE18008083B4443151462A28C6DFF80010002605302248088950484550A3",
INIT_0A => X"10018C241102068006C620C03882019480E631A0855E924E2598038938404037",
INIT_0B => X"A641165448C80C103648A3648A3648A3648A3648A3648A3648A366451B2451B2",
INIT_0C => X"011100841200D001000624000100C002804A08221890004806A310FFDF000454",
INIT_0D => X"5004D8158809C86065941840B1014FFF56FFC0281280080180B2948004400220",
INIT_0E => X"5004D815810D42E04A08A80098C02450025360694101816002D41A4068C10181",
INIT_0F => X"134160C8125B0B271802242880A04482418A0068C101816002D41A4069410181",
INIT_10 => X"10080E05C0B06AA8B12CFD0D42E0441A300012682960828F05C96A001B029010",
INIT_11 => X"00010362A8A20826A88660D86B202049F115100920C54E8EA256ECF078BA081C",
INIT_12 => X"064802C0081B0D64040936443306C55144104F30A8801406D002900062803201",
INIT_13 => X"4581BA0038005A706680012280506A8010602011819E290048A2118EC8140C08",
INIT_14 => X"CC158092C044600466208CC5091011C322A4C40A0300600C0A80509F41800880",
INIT_15 => X"80200802008020080200802008020412002001000000381C02004000FBFFF80D",
INIT_16 => X"0200802008020080200802008020080200802008020080200802008020080200",
INIT_17 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_18 => X"FDDFEFFFBEFFE7C7BFBEFC000000000000000000000000080200802008020080",
INIT_19 => X"F7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7FFBFBFFF9E79E7FFFDF3",
INIT_1A => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFDFEFF7FBFDFEFF7FBFDF7DF7DF7D",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00001FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D000200008000000000000000000000000",
INIT_1F => X"4AA5D00020AA5D7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550402010087FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAA954BA5500020BA5D7FFFFFFFFFFFFFFFFFFFFFFFFFFAE95",
INIT_21 => X"0200000003FFFFFFFFFFFFFFFFFFFFFFF7AA974BA5D0402000557BFFFFFFFFFF",
INIT_22 => X"FFFFEFF7AE974BA5D00174BA00003FFFFFFFFFFFFFFFFFFFFFFF7AA974AA5500",
INIT_23 => X"043FFFFFFFFFFFFFFFFFFFFEFF7AE954BA5D04174AA00003FFFFFFFFFFFFFFFF",
INIT_24 => X"FAE974AA5D003FE005D2EBFFFFFFFFFFFFFFFFFFDFEFF7AE954AA5500174BA5D",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFDFEFF",
INIT_26 => X"A550400028007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0000010000000000",
INIT_27 => X"FFFFFFFFFFFFFAA954BA5D00000BA557FFFFFFFFFFFFFFFFFFFFFFFFFFAE974A",
INIT_28 => X"0005571FFFFFFFFFFFFFFFFFFFFFFFF7AA954BA550000082557BFFFFFFFFFFFF",
INIT_29 => X"DFEFF7AE974BA55000503800003FFFFFFFFFFFFFFFFFFFFEFF7AA974AA5D0405",
INIT_2A => X"3FFFFFFFFFFFFFFFFFFDFEFF7AE954BA5D00154AA00043FFFFFFFFFFFFFFFFFF",
INIT_2B => X"A974BA5D00104925D0E3FFFFFFFFFFFFFFFFBFDFEFFFAE954AA550415492140E",
INIT_2C => X"FFFFFFFF7FBFDFFFFFAA974BA550038E285D2ABFFFFFFFFFFFFFFFFBFDFEFFFA",
INIT_2D => X"D00000100000000000000000000000000000000000000000000000071FFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE954AA5504000BA087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0557BFFFFFFFFFFFFFFFFFFFFFFFF7AA954BA5D00000BA5D7FFFFFFFFFFFFFFF",
INIT_30 => X"EFF7AE954AA5D041740055517FFFFFFFFFFFFFFFFFFFFEFF7AA974AA55000200",
INIT_31 => X"FFFFFFFFFFFFF7FBFDFEFFFAE954BA5500174AA08043FFFFFFFFFFFFFFFFBFDF",
INIT_32 => X"74BA550415410552ABFFFFFFFFFFFFFF7FBFDFFFFFAA974AA5D00174BA08043F",
INIT_33 => X"FDFEFF7FBFFFFFF7AE954BA5D0000010552ABFFFFFFFFFFFEFF7FBFDFFFF7AA9",
INIT_34 => X"00000000557FFFFFFFFFDFEFF7FFFFFEFF7AE974AA550028AAA5D2EBFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(2),               -- Port A write enable input
DIA(0)   => data_write_a(21),        -- Port A data input
DOA(0)   => data_read_a_hi_512(21),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(2),               -- Port B write enable input
DIB(0)   => data_write_b(21),        -- Port B data input
DOB(0)   => data_read_b_hi_512(21),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_22_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"5290F4CDE914905A14A43D33F488243E17122300F55FEB189B343A1140548380",
INIT_01 => X"A94007B259F6A975386262000C344BA9573C6FF57B18A5FB0ABFCD3C2C5F4F0C",
INIT_02 => X"D56B4302AC01005111011BD506AA5205274056900596A539584E2E6DFE4B2418",
INIT_03 => X"9AC0FCBD854688207C90007A1000047A00E588632CA213C8903AD6B55AD0EB5A",
INIT_04 => X"30002047A6FCA110086C402022F2124A8022492580040440002021C922D9109B",
INIT_05 => X"14A206B6838151008D95DD1847811C08002380041F1104002205AC4140DAD060",
INIT_06 => X"1727FF2EB9EF113A10BD32F44289D1F840C1710010344DB9A808FDFF3DE03130",
INIT_07 => X"050700154A00401D00495A06A8D464C5F6B54AA8551040818F4C997AC80CBE05",
INIT_08 => X"0141008801018040E48D50080002B00A0C00801014541E9504703680017F6CB4",
INIT_09 => X"02680000010937986481514E2A29CE010708C0804C6A033F7FCFF9426A41F1AB",
INIT_0A => X"00500001840000C80B410014088040F4A944B1AA313C004554002381B8000500",
INIT_0B => X"A004D1594832824A070AA070AA070AA070AA070AA070AA070AA0725503855038",
INIT_0C => X"501428054278142151262CA50343854E506A2C6898B2950AA6A35B0004284058",
INIT_0D => X"90078E1F840A2B0114020104022460002200050F60E220A06880D2A14050A028",
INIT_0E => X"90078E1F891C239F8908003099C1ACF06273612B3482C0C0078E1F412B1582C0",
INIT_0F => X"1BA1B0FD16770236A4091621C08055C2C0DB012B1582C0C0078E1F412B3482C0",
INIT_10 => X"00101F09C030AB28B03C111C239F870828041BA859F213AFC14AA38043006018",
INIT_11 => X"10E8822A984B0025B0DE6089462660095337B08AA600CA88B143AB11880C2806",
INIT_12 => X"055412D4481128C4CC012A66F304553096004B61BD8068B92400D0004E303689",
INIT_13 => X"589C48082C006A9057CA4385809520F07830001AC2173B00E162563454C40804",
INIT_14 => X"00460848952220592745AC11A544B1BF006850840180A00E1C81900C4190E160",
INIT_15 => X"22088220882208822088220882208CD888088D940D2A3A9D5002001300800C8C",
INIT_16 => X"0080200882208822088220882208822088220882208822088220882208822088",
INIT_17 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_18 => X"FBDFD1FE3EFBD7BBEFBEFA0A245120000000007FFFFFFFF20080200802008020",
INIT_19 => X"F3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF7FFBFAFBBBEFBEFBEFBF7",
INIT_1A => X"CFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCF3CF3CF3C",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000007F3F9FCFE7F3F9FCFE7F3F9F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040000000000000000000000000000000",
INIT_1F => X"4BA550000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0002000087FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974AA550402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"020AA5D7FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5D00000AA007FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAA954BA5504000AA557FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5D00",
INIT_23 => X"7BFFFFFFFFFFFFFFFFFFFFFFFFFAA954BA5500020BA5D7FFFFFFFFFFFFFFFFFF",
INIT_24 => X"7AA974BA5D040200055517FFFFFFFFFFFFFFFFFFFFFFFFAA954BA5500000BA5D",
INIT_25 => X"00000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000080000000",
INIT_27 => X"FFFFFFFFFFFFFAE974AA550002010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"0BA087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550400028007FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAA954BA5D00000BA557FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5D0002",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAA954BA5504020AA5D7BFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"A974AA5D00070925D71FFFFFFFFFFFFFFFFFFFFFFFF7AA954BA5500000825571",
INIT_2C => X"FFFFFFFFFFFFFFEFF7AA974AA5D040500055517FFFFFFFFFFFFFFFFFFFFFFF7A",
INIT_2D => X"D040200008000000000000000000000000000000000000000000000003FFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"A087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550002000087FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAA954AA5D00020AA007FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5504000B",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFF7AA954BA5D00000BA5D7BFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"74AA55000200055517FFFFFFFFFFFFFFFFFFFFEFF7AA974BA5504020BA557BFF",
INIT_33 => X"FFFFFFFFFFDFEFF7AE974AA5D00154105D517FFFFFFFFFFFFFFFFFFFFEFF7AA9",
INIT_34 => X"00000000043FFFFFFFFFFFFFFFFBFDFEFF7AE954AA5D041740055557FFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000007FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(2),               -- Port A write enable input
DIA(0)   => data_write_a(22),        -- Port A data input
DOA(0)   => data_read_a_hi_512(22),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(2),               -- Port B write enable input
DIB(0)   => data_write_b(22),        -- Port B data input
DOB(0)   => data_read_b_hi_512(22),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_23_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"EF20906D902424807BC8241BC81801B97D38AD3C0800103362A6741C80A12A02",
INIT_01 => X"001FFF8409F089003B4422000D80C80106804A7951C5B9D1C828043EA28838F9",
INIT_02 => X"028406A002DC176444683862400003111001303FFC00F240D50146013B300500",
INIT_03 => X"0006C90C010203F80005DC00C52FC380BEAC25886C02034800200200A1008008",
INIT_04 => X"17DFFF8049000BFF878314BFF8488890979800002F702002BB807A068403C280",
INIT_05 => X"DA07F0000000007FF020C814380011FE5E1C2FC3E05FFFF90020000808900010",
INIT_06 => X"10004C9690A8CA008024685184097E81E872C8FFE900FC31348EFDF03BE15E22",
INIT_07 => X"402000001FFBFFFD00080200B8140011F0D8C108155542018D1A302193E94004",
INIT_08 => X"41BE1F5F80003FF0002023FFDF79000000000EFFE309606020008005FC000000",
INIT_09 => X"FC83FE1840C0902400300000000000DFFD4004040C4D32BF7C0EE860003CE680",
INIT_0A => X"10018C24110A860006C620C0312241C482B20420CC56924E2199000C00415037",
INIT_0B => X"4669070510C90C14304043040430404304043040430404304043040218202182",
INIT_0C => X"008000105400C00400100000A018000801000C024000004A940000FFDF820604",
INIT_0D => X"100152100801C17E61841950B1C10FFF57FFC02812F00429DC92C40002000100",
INIT_0E => X"10015210088528E00E02C8200A430A424202A1CAF13F214001521001CBF03F21",
INIT_0F => X"01C1C044006D0C94FB94320880603C420B8001CBF03F214001521001CAF13F21",
INIT_10 => X"30182800A018D9CA8000648528E00D12480202C86040902AC60BACDF0E02D020",
INIT_11 => X"0445C19960A00026880C006739000009B00300010AF5052419D1964419028014",
INIT_12 => X"01844068880CE72000013600600332C140004D101808458A5602E00089202911",
INIT_13 => X"41D0B9023402085020825132C8CB5B4040301009408021144CB042F880100C06",
INIT_14 => X"8E17C0D240406519400500840A9524EE38A1F80E02120018390320F050144CB2",
INIT_15 => X"01004010040100401004010040100100040040000000000001000900FBFFE000",
INIT_16 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_17 => X"0040100401004010040100401004010040100401004010040100401004010040",
INIT_18 => X"0000000000000000000000000000000000000000000000001004010040100401",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000000000000000000000000",
INIT_1F => X"4BA5D0400010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000007FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974BA5D0002000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"00010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA550002000007FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAE974AA550400000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5500",
INIT_23 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550402010087FFFFFFFFFFFFFFFFFF",
INIT_24 => X"FAE954AA5D00000AA007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA55040200008",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010000000000",
INIT_27 => X"FFFFFFFFFFFFFAE974BA5D0400010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0000010007FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAE974AA550002010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA550002",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550400010087FFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"E954AA5D0402038007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550400028007F",
INIT_2C => X"FFFFFFFFFFFFFFFFFFAE954AA5D00020BA087FFFFFFFFFFFFFFFFFFFFFFFFFFA",
INIT_2D => X"D0402010000000000000000000000000000000000000000000000007FFFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000087FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAE974BA550002010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D000001",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFFFAE974AA550002000087FFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"54AA5504000BA087FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA550400010007FFF",
INIT_33 => X"FFFFFFFFFFFFFFFFAA954AA5D04000AA087FFFFFFFFFFFFFFFFFFFFFFFFFFAE9",
INIT_34 => X"000000007BFFFFFFFFFFFFFFFFFFFFFFFFFAA954AA5D00020AA007BFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000007FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(2),               -- Port A write enable input
DIA(0)   => data_write_a(23),        -- Port A data input
DOA(0)   => data_read_a_hi_512(23),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(2),               -- Port B write enable input
DIB(0)   => data_write_b(23),        -- Port B data input
DOB(0)   => data_read_b_hi_512(23),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_24_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100600007FFF000080108004000800020000840041000080808",
INIT_02 => X"0000068002CC07400000090C080002000000103FF811F150231000520ABE4404",
INIT_03 => X"210A0600000203F80005DC00000DC3801EA000000745C4010220000000008000",
INIT_04 => X"07C5FF804900026F8780001DF8000000079800000F300002998078068003C080",
INIT_05 => X"C207F0000000007FF0000004380001FE1E1C07C3E00CFFF80000000000000000",
INIT_06 => X"0002648240F20035A0102000BD0000002802C87FC800FCAA035400001B918600",
INIT_07 => X"0000000001FBFFEC4D2B4AD0B8129063B2CC0000100042018408142F16C01848",
INIT_08 => X"008E1F5F80001FF0000000FFDF78000000000EFFE001600000000005FC000000",
INIT_09 => X"E883FE180000000000300000000000DFFD0000002A80D500000671000004A000",
INIT_0A => X"10018C0411020600048620C030020502000200000400920A2198000800404037",
INIT_0B => X"0641060400C00C00304003040030400304003040030400304003040018200182",
INIT_0C => X"000000001000C00000000000000240058000000000000000000000FFDF000404",
INIT_0D => X"E00880104809C1666594584031010FFF56FFC000104000000010440000000000",
INIT_0E => X"E0088010492064206100E81084200048C0804012500021B00880108012500021",
INIT_0F => X"04100144800803419043064900C0020501840012500021B00880108012500021",
INIT_10 => X"1018140F02C0000809408D206420530270040410004C840041A0D80054109038",
INIT_11 => X"110002C9E8010C00010480B35A0300400041020902F60002260D65B361BAA104",
INIT_12 => X"0228204300166B4060080008240593D0021800020818B06D9802F00030C02060",
INIT_13 => X"143B62023C00142800B04400095DFF90203020042108603100061516EE800C06",
INIT_14 => X"DC1180C7804400044029208301040214AE4C7C02000040206602C10B48110006",
INIT_15 => X"00000000000000000000000000000000000000000000000000000000FBFFE000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"DD5EDCF9822659B6888332000000000000000000000000000000000000000000",
INIT_19 => X"F3CF3CF3CF3CF3DF7DF7DF7DF7DF7DF3DF3DF3DF3DF4D30C2432AEBAEBFE5A15",
INIT_1A => X"C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783DF7DF7DF7C",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000F0783C1E0F0783C1E0F0783",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201008000000000000000000000000",
INIT_1F => X"4BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974BA5D0400000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"00010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000007FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAE974BA5D0000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_23 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0002000087FFFFFFFFFFFFFFFFFF",
INIT_24 => X"FAE974BA550002000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D000200000",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010080000000",
INIT_27 => X"FFFFFFFFFFFFFAE974BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000087FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAE974BA5D0400010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0000010007FFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"E974BA550002000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0000010007F",
INIT_2C => X"FFFFFFFFFFFFFFFFFFAE974BA550002000007FFFFFFFFFFFFFFFFFFFFFFFFFFA",
INIT_2D => X"D0402010080000000000000000000000000000000000000000000007FFFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAE974BA5D0400000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040200",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000087FFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"74BA5D0000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0000010087FFF",
INIT_33 => X"FFFFFFFFFFFFFFFFAE974BA550000010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE9",
INIT_34 => X"000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA550002010087FFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(3),               -- Port A write enable input
DIA(0)   => data_write_a(24),        -- Port A data input
DOA(0)   => data_read_a_hi_512(24),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(3),               -- Port B write enable input
DIB(0)   => data_write_b(24),        -- Port B data input
DOB(0)   => data_read_b_hi_512(24),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_25_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100200002000000080100004000000020000800041000080808",
INIT_02 => X"0000068002CC474000000800000002000000103FFCE302008000000880844A04",
INIT_03 => X"00000040700803FC0105DE00020DC3801EA00000040000000020000000008000",
INIT_04 => X"47C5FFC04904026F8780081DFC040000079C92484F30499299837C168003E400",
INIT_05 => X"C207F0382004407FF0000004382281FF1E1C07C3E00CFFFC090004B05000200A",
INIT_06 => X"1009015C4000000020000000390C10002802C87FC800F8000000000019810600",
INIT_07 => X"0501000001FBFFFD480A0280A816002010800001000054018408102000000002",
INIT_08 => X"0C8E1F5FA21C9FF8004000FFDF7C062031863EFFF75D78004001010DFC000020",
INIT_09 => X"E883FE180C00000000300000000000DFFF00180800000000000660100000A000",
INIT_0A => X"1001DCCC31222730A49620C030020100000200000400921A21D8000804404037",
INIT_0B => X"0641062400C00C00304003040030400304003040030400304003040018200182",
INIT_0C => X"C11160845004D04820000000000000000000000000000000940000FFDF000404",
INIT_0D => X"000800000801C0786184185031810FFF56FFC02812E0182000F2C48304418220",
INIT_0E => X"0008000000002020000008000000000800800002400001000800000002400001",
INIT_0F => X"0000010000000000900000080000000400000002400001000800000002400001",
INIT_10 => X"1000000002002000004000002020000200000000000404000000880000001000",
INIT_11 => X"010000082000000001000001080000000040000100C600800001040000040009",
INIT_12 => X"0000000100002100000000080000104000000002000000081001000000000040",
INIT_13 => X"0010200000000000001004000001080000400080000040010000001080001008",
INIT_14 => X"8C11808200400000400000C20000000420000000030280000000010000010000",
INIT_15 => X"82208822088220882208822088A20C52082081A30080000002005008FBFFF001",
INIT_16 => X"2208822088220882208822088220882208822088220882208822088220882208",
INIT_17 => X"2088220882208822088220882208822088220882208822088220882208822088",
INIT_18 => X"29432D518B45265D82BB4101000005FFFFFFFFFFFFFFFFF82208822088220882",
INIT_19 => X"24924924924924820820820820820820924820924824000A6242B4D34D7F7451",
INIT_1A => X"AC562B158AC562B158AC562B158AC562B1188C46231188C46231189249249249",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000162B158AC562B158AC562B158",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000000000000000000000000",
INIT_1F => X"4BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"02000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAE974BA5D0402000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_23 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000007FFFFFFFFFFFFFFFFFF",
INIT_24 => X"FAE974BA5D0400000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040000008",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010000000000",
INIT_27 => X"FFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAE974BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000007FFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"E974BA5D0400000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000087F",
INIT_2C => X"FFFFFFFFFFFFFFFFFFAE974BA5D0400000007FFFFFFFFFFFFFFFFFFFFFFFFFFA",
INIT_2D => X"D0402010000000000000000000000000000000000000000000000007FFFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"74BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000007FFF",
INIT_33 => X"FFFFFFFFFFFFFFFFAE974BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE9",
INIT_34 => X"000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000007FFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000007FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(3),               -- Port A write enable input
DIA(0)   => data_write_a(25),        -- Port A data input
DOA(0)   => data_read_a_hi_512(25),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(3),               -- Port B write enable input
DIB(0)   => data_write_b(25),        -- Port B data input
DOB(0)   => data_read_b_hi_512(25),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_26_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"E9264EAB20190CA3BA4997AA9002AE9C001006B0778015CFA17E0811039879C7",
INIT_01 => X"F1FFF9BB1F773C7F9BB07DFFFDD863FC5FFF3FEFFBBF9FFB22FFFBC7B9F30686",
INIT_02 => X"9B3184F8AFDEAF300029E4E300FC78A6258548EFFA71C00172082400003A2161",
INIT_03 => X"0084F0FF7FFF1FDD3FEFDCDE981DC3FF5F0D294A7B2B18A0001B9CE6CC606E73",
INIT_04 => X"0FC5DFD7EDFFD66F87FE605DDDBFF3690F9EDB7F5F7AFF639BD7DE37C2FEF591",
INIT_05 => X"F205F0F8E9D199FF76DFEE1C3FCC3FF7BE1FD7C3FFACFBFFDFF7B4FEFFDAA10E",
INIT_06 => X"042648C40179912406C1830639AFBEC14489737FDC00B13BB79DFDB83BF4112A",
INIT_07 => X"763A844769FFBFE4398E4390BB9C28B1D0F049080414583F9468D1AEFC000060",
INIT_08 => X"02C05FD7BC471FBD13D981F7DF7D7E6171AF3FEFE8A3E679FAC1FD1FFFBEB000",
INIT_09 => X"F8CFFE38FF7F6BD928F1ABB47476B5FEF9F59F5FCEEDE73FEE0EFC53B079F5CC",
INIT_0A => X"315BDDCC3B336F7C548667D47B7737AF3FD62601EDC2B66A67B9D60FE4C4427F",
INIT_0B => X"06E19F4DA0E80E903DE3035E3035E3035E3035E3035E3035E3035E981AF181AE",
INIT_0C => X"EBFBF7FEBD66DBFCA3F87501AE7B080607307DCFE1D4077B4D026FFFFBFFAFCD",
INIT_0D => X"0007E010084BCD7FF1B61B5C33813FFFFCFFC7D7D51D6F5FDCB935D7AFEBD7F5",
INIT_0E => X"0007E01001BD8020500008001F010040520201F45EC0010007E01001F45EC001",
INIT_0F => X"1DC0004600400F781429C0080000770001A001F45EC0010007E01001F45EC001",
INIT_10 => X"10003C064000E408010081BD8020600200001EC00040B02007EC09A0E0001000",
INIT_11 => X"360403E434588007200D00F88C84C081C203404B3BFD0402346235408402C080",
INIT_12 => X"07B00040091F1190982038406807C868B1000E401A08FE0012040000FC002001",
INIT_13 => X"7D00212000007C400082D81009FC08281D00001F010021560406758091454000",
INIT_14 => X"FFBFF5FA1040076065F730FC08043A903A80008320C0403C3400008860160406",
INIT_15 => X"D7F5FD7F5FD7F5FD7F5FD7F5FDFF7F7F7F77F9F761FFBFDFFDE5BFFFFF7FF005",
INIT_16 => X"7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5F",
INIT_17 => X"F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD",
INIT_18 => X"B79E923C2CD990AA7F0DDB6B910C8DFFFFFFFFFFFFFFFFFD7F5FD7F5FD7F5FD7",
INIT_19 => X"30C30C30C30C30C30C30C30C30C30C30D34D34C30C35F7AA9ABF0E38E3A8EB62",
INIT_1A => X"C26130984C26130984C26130984C26130984C26130984C26130984C30C30C30C",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000130984C26130984C26130984",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000000000000000000000000",
INIT_1F => X"4BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"02010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_23 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFF",
INIT_24 => X"FAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010000000000",
INIT_27 => X"FFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"E974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007F",
INIT_2C => X"FFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFA",
INIT_2D => X"D0402010000000000000000000000000000000000000000000000007FFFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"74BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFF",
INIT_33 => X"FFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE9",
INIT_34 => X"000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(3),               -- Port A write enable input
DIA(0)   => data_write_a(26),        -- Port A data input
DOA(0)   => data_read_a_hi_512(26),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(3),               -- Port B write enable input
DIB(0)   => data_write_b(26),        -- Port B data input
DOB(0)   => data_read_b_hi_512(26),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_27_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"00080A40000A41248002029000050A088000008242A0004404480002000A1155",
INIT_01 => X"F1FFF1C11F781C129C107DFFFE0860941E81258CA2B71C2220EC1B86E1A00002",
INIT_02 => X"183080988B2EAE00002BE001117C78C6848140CFFA0000800042008000011081",
INIT_03 => X"000000FF7CF91F1D3DEF3CDA881D23FB5C0C21085B0B0820001318C60C204C63",
INIT_04 => X"8FC51FD7EDFDD66E47EE205D1DB7F1490E5EDB7D5CBADB2385D79C3643D4E580",
INIT_05 => X"E001F0C0C991BBFC76DFEA1A3F8C3BC7391F9723FF2CE3FCD6D13096B79C8106",
INIT_06 => X"40000001000000084041830600A40C415004637FC4003021259CFDB01BF80028",
INIT_07 => X"3158954761FA3FE402088220AC1108001080400A400041018468D1A060000050",
INIT_08 => X"02005F0784411E390A4881C7BEFC5F6171CE2F8FE823E778DAC16C1FFBBC9000",
INIT_09 => X"F0C7FEBABF3F6BD108F40E04C0C084F0F8B58B5B8849673F6C0E7A01B00914C4",
INIT_0A => X"B51BFDCC39732F3554866AD57C37BEAF1C152201A4C0B6EA63AAD60B60D4427F",
INIT_0B => X"06F18FC5A0E00F0038D1030D1030D1030D1030D1030D1030D1030F0818688186",
INIT_0C => X"AB6AD7EAB962CBD8A3A83101F47E08040510768EA0C406630D0226FFE375ADE5",
INIT_0D => X"000760000843C561E5C55C42B9011FFF48FFCC57550D63564D1D2556ADAB56D5",
INIT_0E => X"0007600004BD8020100008001F010000130201E44A40010007600005E44A4001",
INIT_0F => X"1DC0000208400D781020C00800007700002005E44A40010007600005E44A4001",
INIT_10 => X"10003C064000C400018080BD8020200200001EC00000382006EC0820A0001000",
INIT_11 => X"3E0403A424108007200102E888808081C20040431BC504021462354004004080",
INIT_12 => X"07B00000015D1110102038400817484821000E400204FE0010040000FC000000",
INIT_13 => X"7D00202000007C400000F81001FC08080500001F0100005E0404758081014000",
INIT_14 => X"8DBBB5FA10400360649310FC08003A903A8000012040403C34000080201E0404",
INIT_15 => X"56D5B56D5B56D5B56D5B56D5B56D7E3D7B57B1C4E17F0944B8D596EEFC7FF001",
INIT_16 => X"6D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B",
INIT_17 => X"D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B5",
INIT_18 => X"2D0200903950C080420948E2D10E8FFFFFFFFFFFFFFFFFF56D5B56D5B56D5B56",
INIT_19 => X"00000000000000000000000000000104000000000004000E5E420000002921C4",
INIT_1A => X"28140A05028140A05028140A05028140A0100804020100804020100000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000140A05028140A05028140A050",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000000000000000000000000",
INIT_1F => X"4BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_23 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFF",
INIT_24 => X"FAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201008",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010000000000",
INIT_27 => X"FFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"E974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087F",
INIT_2C => X"FFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFA",
INIT_2D => X"D0402010000000000000000000000000000000000000000000000007FFFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"74BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFF",
INIT_33 => X"FFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE9",
INIT_34 => X"000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000007FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(3),               -- Port A write enable input
DIA(0)   => data_write_a(27),        -- Port A data input
DOA(0)   => data_read_a_hi_512(27),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(3),               -- Port B write enable input
DIB(0)   => data_write_b(27),        -- Port B data input
DOB(0)   => data_read_b_hi_512(27),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_28_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"02200AA400180030808802A900002A08001280A08A801044104A1000001818C3",
INIT_01 => X"50A00011460214428114180000882214413D0A71592A01D92213D28005210202",
INIT_02 => X"8A54800A210200111100C2110054289220810440030404010844000444410001",
INIT_03 => X"1080010208B51400007800000A000001000108C21008092000018C6295200631",
INIT_04 => X"0008000000017000000028000001610300000010000802202040012040040011",
INIT_05 => X"2000044440048880026A22000026A20000000000000000004994140203000064",
INIT_06 => X"1400922401041008004891224228810080010200040001020800000004000008",
INIT_07 => X"150B001328000001404010040084088404200020455514000224489028492201",
INIT_08 => X"00414000201800004080A0000002480B04008100011000088800081002C19020",
INIT_09 => X"000400001036584108415B4A6A694A0000100101C08200000001000190200044",
INIT_0A => X"004800210C19808400500010009110091500020B408820000200400040811600",
INIT_0B => X"40000800B00100040D8140581405814058140581405814058140580A02C0A02C",
INIT_0C => X"00200248010201008298150006210802043058C46054032981002D00201C8081",
INIT_0D => X"0000A00000400600841041108280300008000140000401028008330000800040",
INIT_0E => X"0000A000000080001000000000000000500000040A40000000A00000040A4000",
INIT_0F => X"00000006000000080020C00000000000012000040A40000000A00000040A4000",
INIT_10 => X"00000000000024000000000080002000000000000000A00000040020A0000000",
INIT_11 => X"2200000404108000000900008080808000024040152000000020000004004080",
INIT_12 => X"0000000009001010102000004800080821000000120002000004000000000001",
INIT_13 => X"2000002000000000000288000020000805000000000001420000200001014000",
INIT_14 => X"408010000000022000D610280000080000000001204000000000000820020000",
INIT_15 => X"00401004010040100401004010042024210218734CD52150A840827504000000",
INIT_16 => X"0401004010040100401004010040100401004010040100401004010040100401",
INIT_17 => X"4010040100401004010040100401004010040100401004010040100401004010",
INIT_18 => X"05822140048D2E57B1348141845C200000000000000000000401004010040100",
INIT_19 => X"04104104104104104104104104104104104104104101A6A0A0EB1861863BC422",
INIT_1A => X"2C160B0582C160B0582C160B0582C160B0180C06030180C06030181041041041",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000160B0582C160B0582C160B058",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000000000000000000000000",
INIT_1F => X"4BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_23 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFF",
INIT_24 => X"FAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010000000000",
INIT_27 => X"FFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"E974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007F",
INIT_2C => X"FFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFA",
INIT_2D => X"D0402010000000000000000000000000000000000000000000000007FFFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"74BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFF",
INIT_33 => X"FFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE9",
INIT_34 => X"000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000007FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(3),               -- Port A write enable input
DIA(0)   => data_write_a(28),        -- Port A data input
DOA(0)   => data_read_a_hi_512(28),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(3),               -- Port B write enable input
DIB(0)   => data_write_b(28),        -- Port B data input
DOB(0)   => data_read_b_hi_512(28),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_29_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"79964E4BA01DACAB9E659792D00AAE160002829C7FDFEFCEE97C2815039D70C3",
INIT_01 => X"50BFF9AB0775343F9AB01DF80D5821FC0FFF3FEFD1AF9FF1207FFBC7B9720586",
INIT_02 => X"0D15846807D207200021C4E200D428A2018408600271C000720A0000003A2161",
INIT_03 => X"0000B0027BBF17C43E6DC05E1A0DC07D1F0000803B2819A00019084345606421",
INIT_04 => X"07CDC047A4FB526F807C681DC4B97369078249370F482E62BA414627C2FE3000",
INIT_05 => X"F204007861C088FF0EFF260407C427F19E03C7C01F8CF80749B390EA4BCA202C",
INIT_06 => X"000248C00079800406C081023B233E804488527FDC008019968D74982C94110A",
INIT_07 => X"5229000221FF8000398641903B082831D05000200000083F942850AEB4000221",
INIT_08 => X"00805FD0180E1F8C1111A0F041056A0100A11FE000916249A800B915FE82B020",
INIT_09 => X"F80C000055FF7C492840AAB45456B55E015015058665A31DA603A4539058F54C",
INIT_0A => X"000850400A11414C005005000B51158936D20601A98A204006114005C4800217",
INIT_0B => X"40201948B029029409A3401A3401A3401A3401A3401A3401A3401A9A00D1A00C",
INIT_0C => X"40B1225C1506512C83E85500AC3A080406305587A154023141006DFFF89E82C9",
INIT_0D => X"0000A01008480D3EB4A24A0C910037FFFC0007C7C0140D0B50A8218102C08160",
INIT_0E => X"0000A010010080005000000000000040520000141EC0000000A01000141EC000",
INIT_0F => X"00000046000002080429C0000000000001A000141EC0000000A01000141EC000",
INIT_10 => X"00000000000024080100010080006000000000000040B000010401A0E0000000",
INIT_11 => X"3600004414588000000D00108484C080000340483B590000202000008402C080",
INIT_12 => X"00000040090210909820000068008828B10000001A0802000204000000002001",
INIT_13 => X"20000120000000000082D800082000281D000000000021560002200011454000",
INIT_14 => X"B29450580000066021F6303C000408000000008320C000000000000860160002",
INIT_15 => X"816058160581605816058160589625662522506344FF9FCFFF62EB6DFF001004",
INIT_16 => X"1605816058160581605816058160581605816058160581605816058160581605",
INIT_17 => X"6058160581605816058160581605816058160581605816058160581605816058",
INIT_18 => X"F2DDCFFFBEFFCF07FFBFFD41800C05FFFFFFFFFFFFFFFFF81605816058160581",
INIT_19 => X"7DF7DF7DF7DF7DF7DF7DF7DF7DF7DD75D75D75D75D77FFBF3F7DFFFFFFD779F3",
INIT_1A => X"FEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDF7DF7DF7DF",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00001F7FBFDFEFF7FBFDFEFF7FBFD",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000000000000000000000000",
INIT_1F => X"4BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_23 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFF",
INIT_24 => X"FAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010000000000",
INIT_27 => X"FFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"E974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007F",
INIT_2C => X"FFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFA",
INIT_2D => X"D0402010000000000000000000000000000000000000000000000007FFFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"74BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFF",
INIT_33 => X"FFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE9",
INIT_34 => X"000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(3),               -- Port A write enable input
DIA(0)   => data_write_a(29),        -- Port A data input
DOA(0)   => data_read_a_hi_512(29),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(3),               -- Port B write enable input
DIB(0)   => data_write_b(29),        -- Port B data input
DOB(0)   => data_read_b_hi_512(29),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_30_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"FFDFF3FC3EFFF7FFFFBFFA000000000000000000000000000000000000000000",
INIT_19 => X"F3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF5F7AEBEBFBEFBEFFEFFF7",
INIT_1A => X"CFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCF3CF3CF3C",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000007F3F9FCFE7F3F9FCFE7F3F9F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000000000000000000000000",
INIT_1F => X"4BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_23 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFF",
INIT_24 => X"FAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010000000000",
INIT_27 => X"FFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"E974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007F",
INIT_2C => X"FFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFA",
INIT_2D => X"D0402010000000000000000000000000000000000000000000000007FFFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"74BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFF",
INIT_33 => X"FFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE9",
INIT_34 => X"000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(3),               -- Port A write enable input
DIA(0)   => data_write_a(30),        -- Port A data input
DOA(0)   => data_read_a_hi_512(30),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(3),               -- Port B write enable input
DIB(0)   => data_write_b(30),        -- Port B data input
DOB(0)   => data_read_b_hi_512(30),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_31_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"129000008004A00804A40000400800020000000C005FEA005800200400050100",
INIT_01 => X"A15FF18019700810180065FFFC0040801E80258CA2951C2200EC0906A0804140",
INIT_02 => X"146000808A0C060444692000402850040400408FF80000000010000000004000",
INIT_03 => X"000000FD74480B1C3D951C5A800D03FA1C0C21084B0300000012108518004842",
INIT_04 => X"07C51FC7EDFCA26E07EE001D1CB6904A061EDB6D4C30490281831C1602D0E480",
INIT_05 => X"C001F0808181117C7C95C8183FA099C7181F8703FF0CE3FC0201209010988002",
INIT_06 => X"00000000000000010001020400840C41C000617FC0003021259CFDB01BF00020",
INIT_07 => X"0000000441FA3FE400080200A810000010804008100040018448912040000040",
INIT_08 => X"00011F0780011E38004801C79E7C162231862E8FE00166704041240DF93D0000",
INIT_09 => X"F0C3FE180D89279000B00000000000D0F80088080849673F6C0E780020091480",
INIT_0A => X"1011DCCC31222730048620C4382204A608142002A440924A6188020920404437",
INIT_0B => X"0661874500E00E00304003040030400304003040030400304003060018200182",
INIT_0C => X"810040801060C04821202001A05A00040100240A80800442040202FFC3200444",
INIT_0D => X"000740000803C0616184184031010FFF40FFC407500020004C10060204010200",
INIT_0E => X"0007400000BD0020000008001F010000020201E04000010007400001E0400001",
INIT_0F => X"1DC0000000400D701000000800007700000001E04000010007400001E0400001",
INIT_10 => X"10003C064000C000010080BD0020000200001EC00000102006E8080000001000",
INIT_11 => X"140403A020000007200000E808000001C200000308C504021442354000000000",
INIT_12 => X"07B00000001D0100000038400007404000000E400000FC0010000000FC000000",
INIT_13 => X"5D00200000007C400000501001DC08000000001F010000140404558080000000",
INIT_14 => X"8C1380DA10400140640100D4080032903A8000000000403C3400008000140404",
INIT_15 => X"02008020080200802008020080200C1808008184012A08041202500AF87FF001",
INIT_16 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_17 => X"0080200802008020080200802008020080200802008020080200802008020080",
INIT_18 => X"000000000000000000000002001005FFFFFFFFFFFFFFFFF02008020080200802",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000000000000000000000000",
INIT_1F => X"4BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_23 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFF",
INIT_24 => X"FAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010000000000",
INIT_27 => X"FFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"E974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007F",
INIT_2C => X"FFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFA",
INIT_2D => X"D0402010000000000000000000000000000000000000000000000007FFFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"74BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFF",
INIT_33 => X"FFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE9",
INIT_34 => X"000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(3),               -- Port A write enable input
DIA(0)   => data_write_a(31),        -- Port A data input
DOA(0)   => data_read_a_hi_512(31),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(3),               -- Port B write enable input
DIB(0)   => data_write_b(31),        -- Port B data input
DOB(0)   => data_read_b_hi_512(31),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_0_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"ED39BA795990D275FB4A6E96ACC4731DEA4598B0AFB54867F6EE4618C3749807",
INIT_01 => X"58A0047D8607944AC7DA180001ECA2444042106208408208C20022E9173734B3",
INIT_02 => X"8B1E49562021F8051500147A0E162923024F28000415F5787B09FBF999BB1EFC",
INIT_03 => X"1013BF028A959403C06A23A147723C01E140088280C4CF6996088862C7922221",
INIT_04 => X"781A003802015D9078011DE20340699198600000B08694916434804825241311",
INIT_05 => X"2CA000587E10C880036A3103C00F2000E1E0383C00730002B4409845E4425171",
INIT_06 => X"179B48CFF95DCF9EF730E1C3BB731138AF7B888025340C0888430047040FEE18",
INIT_07 => X"AF155113160400185F87C1F05707D415E664A6E7C5551EBE783060CEB164833F",
INIT_08 => X"4D7E40002B7AE005FDB47600208229010C6101001EFE198C96B0528202C0DCB4",
INIT_09 => X"062400608234D864444081048A80CC00062D42D30222108091C107A1DA040267",
INIT_0A => X"204A21008E514844EB5145000255DA599581D3A9583C24351240B58298011308",
INIT_0B => X"E08C4830F81380CE0F89E07A9E0789E07A9E0789E07A9E0789E070CF0184F038",
INIT_0C => X"3A4E9D63EA180EB150CA1CA45C254D4AF4AA414568729139F2A12C0000016110",
INIT_0D => X"F0009E0FC048211E9C11C31F82E4A000890022B827EB52F52347F174E93A749D",
INIT_0E => X"F0009E0FCC42EFDFBF0AE03080E2AEB2E0F1F80FA97FE0F0009E0FC40FA97FE0",
INIT_0F => X"0231F0BD9E3FC08FEBD6F661C0E008C3CB5F040FAB3FE0F0009E0FC40FAB3FE0",
INIT_10 => X"20180309A0F83BE2B87C7C42EFDFBF187806013879BA878FE807F65FBF12E038",
INIT_11 => X"0BE9F01FC8B38C2098DAE007F323A0C83136B248831ACBFC8BBDCAB779BC699F",
INIT_12 => X"004C72BEC800FE7464290626D7003F9947184131B59003FFEC07F00003F01FB9",
INIT_13 => X"A0FFDA2A3C0202B8776A2FA7F023F7D065703080E29F1B2BE9F8A27E6E915C0E",
INIT_14 => X"016C2D25E52630BB1AE49C2BA7F98D6F846DFC0C2352A0024B83F07F198BE9F8",
INIT_15 => X"749D2749D2749D2749D2749D2749F285F25D2C500815A5522CB5A4B400000CD4",
INIT_16 => X"49D2749D2749D2749D2749D2749D2749D2749D2749D2749D2749D2749D2749D2",
INIT_17 => X"9D2749D2749D2749D2749D2749D2749D2749D2749D2749D2749D2749D2749D27",
INIT_18 => X"31C136AD8E9B562BA39E2600654BA800000000000000000749D2749D2749D274",
INIT_19 => X"4104104104104104104104104104104104104104104104109C83B8E38E2ABE71",
INIT_1A => X"0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0410410410",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000007C3E1F0F87C3E1F0F87C3E1F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000187FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"BAF7FFD55EF007FD75EFFFAE97555557BD75EF5D000000000000000000000000",
INIT_1F => X"000AA843FE00AAFBE8B45AA803DFEFA28428B455D0017410A28428AAAA2FBD54",
INIT_20 => X"FEBAA2D5401450051401555D7FC0145F7AEBFFFF08002AA10A2AABFEAAA2FFC0",
INIT_21 => X"D755555517FFEFA280021FF082E974AA5D7BFFE000804000BAAAAAAAB45557FF",
INIT_22 => X"EA8B45005168A10AA8028A10087FD7410557FC21555D51574AAA2FFE8B455D7B",
INIT_23 => X"AE95410AA80000005D003FEAAFFAEBFE00A2803FEBA002A820AA0800174BA5D2",
INIT_24 => X"2AEA8A10000417410A2FFE8BEFF7FFE8B45FFFBC00005D003FF45557FC01FFFF",
INIT_25 => X"00000000000000000000000000000000000000557DF5500003DFEFFF84175EFA",
INIT_26 => X"5F524AFE38B780154BAFFF1D54AF0075D75EFEBAE9554540754717F1F8000000",
INIT_27 => X"50B6AABDE12BEA0AF010B7D1F8F47E00A2DB45AA8A3AFD7B68E2AB78550E1255",
INIT_28 => X"E9257F1E816D557095EAAA2D1401D500002A150038038E285D7F78FD7000B6AB",
INIT_29 => X"5A87AAD178A8002D1D21C5E8257D5C7AA854008700249243A412EBFF5542A43F",
INIT_2A => X"52A82000E3A5D2150AB8F401471EDBC0B680900AAF52B474385D75C502D15754",
INIT_2B => X"FD7E9541242FE920AD082E10A28F6A150012A2F02AFFDF40E85F475451D502D1",
INIT_2C => X"0550E87B7A405B52AAD152BD00151EAFEDB52E3F1EFFFF485A2DA3D5D24BD417",
INIT_2D => X"57F40545850000000000000000000000000000000000000000000005AAF55508",
INIT_2E => X"F7AEAABFF5D2A81151FB8635A02FA69574BAF7D5555AF0D79D55FFA2AC974450",
INIT_2F => X"8D46F6ABE7082AAAAF2FAC77FE00FF16565B2FA9075F4F7B3EBDF50FEAEAAB55",
INIT_30 => X"56803CE3AEB038662E5D81406014D5D51F5E08A394003A908B8410E707EF34A0",
INIT_31 => X"4AF0151555AF58794040077D774FAE8C798A11A0EAEF75F7AA84001A7052C952",
INIT_32 => X"4E1870108B11020AD4AA05542A0A05051023F9A9D57B63BFBF906CB45FABC095",
INIT_33 => X"F5F0DA6BC9525688C1A2A0C06E9FEE5555BE48AB2A2AE0A0F20C43EAC562245B",
INIT_34 => X"000000FF80F55E25C00A0BA7FBED407A97F6F35F498B96BEB12DAAB77558ABD5",
INIT_35 => X"8000000FF8000000FF8000000FF8000000FF8000000FF8000000FF8000000FF8",
INIT_36 => X"00000000000000000000000000FF8000000FF8000000FF8000000FF8000000FF",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000008000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(0),               -- Port A write enable input
DIA(0)   => data_write_a(0),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(0),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(0),               -- Port B write enable input
DIB(0)   => data_write_b(0),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(0),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_1_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"212C001411984004084D000508C53810A03D1450E839B003342114428A000803",
INIT_01 => X"08000010400A0008010600000084005000400002000000000000000000140000",
INIT_02 => X"C084484000002014400205851002007030450E0000A606C8C44CB4C6666C00E0",
INIT_03 => X"CCF7CE0002058001000000800240200001018CA1800001091408463061120118",
INIT_04 => X"082800100000000040000900010000100040000000008411600401C02100000C",
INIT_05 => X"10800202080422000020012200000000810000200000000004020C00200011A0",
INIT_06 => X"56BDBFBC48C315A8660C18305750C008940D8000011000820001000104050004",
INIT_07 => X"8B4344400004000150248912154404C6060A2FE24555013E13060C158AC97F01",
INIT_08 => X"00082080087A000559102400200281000469000008B000000090108000400430",
INIT_09 => X"0000000000001004140545402820020000010010208000008041060008200001",
INIT_0A => X"2102210182004840007845004044020000200080080844200000048088000000",
INIT_0B => X"48800000190191064620646A06468064680646A0646A06468064690321503234",
INIT_0C => X"02008100200800A1100707040101E20BE0B002605C1C110848200C0000000800",
INIT_0D => X"F000A000C0000012187087010AE4B00000000810010040108104100408020401",
INIT_0E => X"F000A000CC4200002F08E03080000010F18058000003C0F000A000C4000003C0",
INIT_0F => X"000000078808C00000023461C0E00000012704000003C0F000A000C4000003C0",
INIT_10 => X"201803000000240218C0044200001E1878060000000AAC00680000001F10E038",
INIT_11 => X"2100B00048230C200009A0001303204800025200040A00D000000202090C281F",
INIT_12 => X"00000002C9000260640900004D0000904618400012900001EC03F00000000039",
INIT_13 => X"80025A0A3C020000002A8400B00007806070308000000961002880204A901C0E",
INIT_14 => X"000801046004308A185000020128000904285C0C0312A0020000000838810028",
INIT_15 => X"0401004010040100401004010040100010410C002000040280100000000008D0",
INIT_16 => X"4010040100401004010040100401004010040100401004010040100401004010",
INIT_17 => X"0100401004010040100401004010040100401004010040100401004010040100",
INIT_18 => X"48D757DF8A9410218E8A56085142020000000000000000004010040100401004",
INIT_19 => X"555555555555555555555555555554514514514514550431A581924924B02651",
INIT_1A => X"4BA5D2E974BA5D2E974BA5D2E974BA5D2EB75BADD6EB75BADD6EB75555555555",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800005D2E974BA5D2E974BA5D2E97",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000607FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"10AAAABFFFFFF803FE10F7D17FEBA55556AAAAAA800000000000000000000000",
INIT_1F => X"EBAFFD555400557BD54BA5D7FFDF45A2FBD75EFA2AE97555F7FBFFF45FFAE800",
INIT_20 => X"ABEFA2D568A005D5157400AA8028AAAF7FBD54AA002A955555D7FE8ABA082EBF",
INIT_21 => X"FDF55AAFBC0010555540010550417555AA8028BEFAAAE97555082A80000AA802",
INIT_22 => X"BD7410550428ABA5D5168ABA552EBDFEF5D7FEAA00AAAABFEAA007BC0145FFFF",
INIT_23 => X"FFEAB55557FFFEBAAAD568B45A2D5575555D7FC2155F7AEA8BEFAAAA954BA557",
INIT_24 => X"D7BD74000804154BA082ABFF55FFD57DF45F7D568ABAF7AABFFFF082ABFFFFFF",
INIT_25 => X"000000000000000000000000000000000000002EBFFEFA280021FF082E974AA5",
INIT_26 => X"5E175EFF57BF8FC2000BEA4BAE97F78A3FE28E3D17DEAA485FE8E02B50000000",
INIT_27 => X"455571E8A2A087BF8EAAEB8E0016D5D75D54BA5D7BFFF7DA2FFD55EFAAA49554",
INIT_28 => X"157428145A00AA8A2FBD7B6DF6AA28550E10405F7A4AFE38EAA0924921C2FD55",
INIT_29 => X"8E971471C7010B7D168F47400A07A28415A001684104155C5B6DF6DBEFBFAA07",
INIT_2A => X"BFBD7B6A0BF492415FC20105D24AAABF1FFBC7010FF8A38FEF557FEAB78B6AAB",
INIT_2B => X"017EBA4A8EB8F6FFD5FE8B7D557495EAAA2D16D1FDBED56A55557A43DE385FD4",
INIT_2C => X"854008700249243A417FFF41542F5D717FE2AAAA56DEBD17FE3DF7FB7FEBFE38",
INIT_2D => X"07DFCA127B8000000000000000000000000000000000000000000002A3D5C7AA",
INIT_2E => X"AAFBD55FFAA8416545A6FB60F47AF2A00010F78028B15F7823FEAAA2D57DFBA0",
INIT_2F => X"22A38C20B2552E975F758516AAAA0869AAAB8A7C19C55550E8574BA557BFFFEF",
INIT_30 => X"55FFEFBCEE5FBAACB10085EE5DE10A2AEBFF55F7BAAA8565DBAC1112FFAC21A0",
INIT_31 => X"BEA097BEAAFAF2863FA00DD574201E7AD1FFF5575841DE08007FC20480028957",
INIT_32 => X"54FF57EFBFA18D4FBFFF40FF809D4000D7FC00FC5D062BBA05ED5034472A02EA",
INIT_33 => X"7DFBFF6963FCAAA2283CF14050062B0A2F7AE8B5D5D51F5E18ABD5EAFFF2AF95",
INIT_34 => X"000000002CB75F7AA84001A7052C95256807DC31AA8114DE55F5BED201FFFED1",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000008000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(0),               -- Port A write enable input
DIA(0)   => data_write_a(1),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(1),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(0),               -- Port B write enable input
DIB(0)   => data_write_b(1),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(1),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_2_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10E44660018259B2843913100062C98004802322D3E030235201006009B2813",
INIT_01 => X"000AC188084900481C8024A542400340404000720885800802000906E4910204",
INIT_02 => X"82040072AC248C31010204880000007401044C0550200000480E0080001300E0",
INIT_03 => X"0080812C130D0A0D1193088802182142494D218220021100001A8020C1004A00",
INIT_04 => X"090D0AD62824A44A428408540D1610020C6E510818923441A4908B0503404201",
INIT_05 => X"5000A004081122242420480A14A99C428908122144244150906124248C002168",
INIT_06 => X"1400088400450000460000001308890094082015800011012D41D518044C1100",
INIT_07 => X"26731111491C1541324C1114BD880004002040204050413F1400100480000201",
INIT_08 => X"02410582881E0C1511D02082AAAB016A2463288549B044605201D10AE11B0020",
INIT_09 => X"E80394280E40158020B591000800481051241A4A404B5035C60904502054E000",
INIT_0A => X"0102C9E12202EA6014D027C418428E220A5500024808922801A0900A84454458",
INIT_0B => X"4600070110C10D04340043400434A043420434A04342043480434102184021A0",
INIT_0C => X"E9CA34328E44CA1401306100A246000402100C088104010AC8005C5681812B04",
INIT_0D => X"0000A0000801487334E34C1A980001550055481204090A4C01351253A728D194",
INIT_0E => X"0000A000013800004000080000000000500000B01480010000A0000150148001",
INIT_0F => X"0000000608000A500409000800000000012001501480010000A00000B0148001",
INIT_10 => X"1000000000002400000001A100004002000000000000A0000360018040001000",
INIT_11 => X"380001C01048000000090298040440000002400008C400022042004080028000",
INIT_12 => X"0000000009530080880000004813802090000000120C94000200000000000001",
INIT_13 => X"4C000100000000000002E0000950002018000000000001580002508010440000",
INIT_14 => X"7120642000000400015020500004221018000082008000000000000820180002",
INIT_15 => X"5094A5294A5294A52942509425094209461468000822241A03835D88482AB001",
INIT_16 => X"09465094A5294A5294A5294250942509425094A5294A5294A529425094250942",
INIT_17 => X"94650946509465294E5294E5294E5094650946509465294E5294E5294E509465",
INIT_18 => X"080271AE180616A38A18FA204452A7F03F03F07E07E07E05294E5294E5294E50",
INIT_19 => X"20820820820820820820820820820820820820820820490C04102CB2CB2EB2C0",
INIT_1A => X"8944A25128944A25128944A25128944A25128944A25128944A25128208208208",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF1F804A25128944A25128944A2512",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000787FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"AAAA843DFFFAAD1554005D7FD74AA00040015500000000000000000000000000",
INIT_1F => X"F45AAAAA8A10A2AE80010A2AA975FF5D003FE10F7D17FEBAF7D5420AA0855420",
INIT_20 => X"FF45A2AA975EFA2FFD7555FFFBFFF45AAFBC20AAF7D1575EF55517DF555D2EBF",
INIT_21 => X"95555552E974105D517DF55AAAAAABEFAAD1575EFAAAE974AA5D51554BA5D7FF",
INIT_22 => X"E82010F7AABFE10FFD542145FFD5554AA555555555557FE8ABA082EBFFFFAAAE",
INIT_23 => X"FBC0010AA802ABEFAAD540000FFD540000AA802AABAF7FFC2010AAAE821EF552",
INIT_24 => X"A8028BEFAAAE821550851420AA002E800AA08042AB45007FC00BAFFD168BEFF7",
INIT_25 => X"000000000000000000000000000000000000002E80010555540010550417555A",
INIT_26 => X"AE95F40002157F470AABE803AE97A2DF55400557FD54AA1D04001C5150000000",
INIT_27 => X"EF55517DFC5552ABDF45B6AEAFFD5F7A482000BEAE905C755003FE28E3D17DEA",
INIT_28 => X"0BA5FD0154BA5D7BFAF7DA2AE955EFAAA495545E3F5EFF57F7FE80082FFDE105",
INIT_29 => X"8AAF082AB8EAAEB8E0016D5D2A924105D5B7FF7DB6AAAABC7BEDB505EFBEA407",
INIT_2A => X"95038AAAEAF1D7410E80000FF8438E00B6DF68FEF4871D24BA495B5556D5571E",
INIT_2B => X"1ED1EFEAF1EFFFDEAD1C5010AA8E2FBD7B6DF47A00EBDB50000A380AAE28E804",
INIT_2C => X"5A001684104155C5B68E2DBEFBFFBC703AE2DF42AAA002A851C214003FF68007",
INIT_2D => X"50002155510000000000000000000000000000000000000000000002087A2841",
INIT_2E => X"55003FEAAAAD57DEBAA2FDDC01051FBD74BAF7802AB05AAFBD5400557BD54AA5",
INIT_2F => X"7AF7FC20B2F7FBC015D58517FF555D2ABDF55F782BEB47AFAD00010F7AA82155",
INIT_30 => X"55FFFFC20FFF3AE544108410174BA557BEABEFAAEBD55FFAA1456547A2D360F4",
INIT_31 => X"0BA547FD75FF58516AAAA0828AAAB4A78016545540400010557BFDFFFF7822A9",
INIT_32 => X"550AAFACAAA122AA8954BAA2AE9D545002A800A8FF862BA00F2F9E8F0050D442",
INIT_33 => X"954505C417FFFF08555555BAAD335B57AB5155400A2AEBFF45FFFB404007FFBD",
INIT_34 => X"00000000061DE08007FC2048002895755FFAEBCFE57BBA57002DF3C4AAAA002E",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000010000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(0),               -- Port A write enable input
DIA(0)   => data_write_a(2),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(2),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(0),               -- Port B write enable input
DIB(0)   => data_write_b(2),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(2),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_3_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"210C44A20020248B08431120001604B8156023104C40771B3430400A02380206",
INIT_01 => X"015A2A4050B009683C0422C992000B61404040028804A0080A000C16A8990A0C",
INIT_02 => X"C0A406500CE0A95011000D1501005274B5041AB330860281CC08008222170060",
INIT_03 => X"AB488054270F08E1289084C8020420E005A48DA16C021100003A46B06900C91A",
INIT_04 => X"848966150DA0A02941A4080C612A104201C689044382FD403C17E491829B259B",
INIT_05 => X"D006620608843116942508120A208D18A5050160C600D4C894600094B49CA068",
INIT_06 => X"12002D9401C70008060408141788E2C094887033080071913209CC8004640100",
INIT_07 => X"221111454874CCC4122C0932155400C2023940284000003E15020525CE805E11",
INIT_08 => X"020103C9984A0AC511102029869D974214EDBA132891000052C1750B48290020",
INIT_09 => X"60808C8A2E41351020004148A289428730A51E5E644C8233A0090E1020208100",
INIT_0A => X"A4000041A600417914506F955D6422000934000A090A94A020229603A414144D",
INIT_0B => X"469100841001000406D04065040650406D0406D04065040670406C8201782032",
INIT_0C => X"6A4AF532A8040AF821042D01F14084030070262810340402C0000CCE4CC12520",
INIT_0D => X"000800000401C333494594532980733302CCC81300094E5C91200257AD2AD795",
INIT_0E => X"00080000051C0000400000000000000800000190148000000800000450148000",
INIT_0F => X"0000010000000B100409000000000004000005101480000008000004F0148000",
INIT_10 => X"0000000002000000000001B00000400000000000000400000168018040000000",
INIT_11 => X"1000034010480000010002D804044000004000812E4400002440014080028000",
INIT_12 => X"0000000100570080880000080015C02090000002000CCC000200000000000040",
INIT_13 => X"1C0001000000000000104000094C002018000000000040100006418010440000",
INIT_14 => X"4128652000004404010E20500004208018800082008000000000010000100006",
INIT_15 => X"5795A5595A5595A5595A5595A5595E1152556D008028341B13924D80C2E67009",
INIT_16 => X"69565795A5595A5595A5595A5595A5595A559525795257952579525795257952",
INIT_17 => X"95256956579525495E5595A5495E5595A5495E5595A569565795256956579525",
INIT_18 => X"7818F18E0C8514298B0C52A0115009AA9556AAD552AAD5556956579525695657",
INIT_19 => X"24924924924924924924924924924820820820820825042C0000249249202A60",
INIT_1A => X"8D46A351A8D46A351A8D46A351A8D46A353A9D4EA753A9D4EA753A9249249249",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF248086A351A8D46A351A8D46A351A",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"EFAAFFD54AAF7D168B45AAAABDF5500002AA1000000000000000000000000000",
INIT_1F => X"F45FFD168AAA0855420AAAA843DFFFAAD1554005D7FD74AAA284001550055421",
INIT_20 => X"55FF5D003FE10F7803FEBAFFD5420AA080400155AAD5554AAF7802AB4500043D",
INIT_21 => X"28B45A2AE82155A2FBFFEBA0800021550855555FFAA84001FFAAAE80010A2AA9",
INIT_22 => X"168ABAFFFBD54BAAAAE97400A2FBC20AAA284175EF55517DF555D2EBFE00AA80",
INIT_23 => X"AA954AA5D7FFFF45AAAA975EF007BD7555FFFBFDF55AAFBD55EF5D2EBFE10085",
INIT_24 => X"AD1575EFAAAE974AA5D00175555D0015410F7AAAAAAA55043DE00FFFFD5555AA",
INIT_25 => X"0000000000000000000000000000000000000004174105D517DF55AAAAAABEFA",
INIT_26 => X"ABC04001C51551471D7AAF1D05D2EBD56DB7DBEAEBFF551C042AA101D0000000",
INIT_27 => X"92EB842FB5508043FF55EBD56ABD75D5B470AABE8A3AFD7A2DF55400557FD54A",
INIT_28 => X"557FD2082000BEAE905C755003FE28E3D17DEAAEBDF40002550F47155AADB504",
INIT_29 => X"DF40552ABDF45B6AEAFFD5F7A48017DAAFFFAE821C0A0717D1C5B575FFB68E82",
INIT_2A => X"C55D7492E90E3808756DA92EBFFD74BAE3AE85480FFFFC00AABE8E105C755517",
INIT_2B => X"43AE10EAF5C5547FF80954AA5D7FFAF7DA2AE905EF0075D5545E3F5EFF57F7D5",
INIT_2C => X"5B7FF7DB6AAAABC7BEDB505EFBEF5C7092FF801756D490A10438EBA4B8E92410",
INIT_2D => X"D0028A00510000000000000000000000000000000000000000000000E124105D",
INIT_2E => X"AAFBD54005D7BD54AAF78002155515157555AAD142040A2D57FFFFFFAEBFF555",
INIT_2F => X"051AE955F7AAFBC0000AF843FF5500003FF55AAFD6AB455157D74BAF7AAA8B45",
INIT_30 => X"FF557BD74EFFBACD41577B8400010F7AA8215555003FEAAAAC53DEB8A2FDDC01",
INIT_31 => X"0BAF7AA8015558517FF555D2ABDF51F782BCB47ABAE801FFAAFBEAA105D2E955",
INIT_32 => X"214FA2D3EAF57AFFDD7555082AA0AAA00557FEA8A2FDD64BAAF8282012AFFEC2",
INIT_33 => X"820AAAB842AA00000028AB0AAFF48547AE04174BA557BEABEFA2AA951FF88554",
INIT_34 => X"000000002A80010557BFDFFFF7822A955FFFFC21FFF3BE40412DE02955FF082A",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000008000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(0),               -- Port A write enable input
DIA(0)   => data_write_a(3),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(3),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(0),               -- Port B write enable input
DIB(0)   => data_write_b(3),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(3),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_4_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A108400020612C80284210081034849800A000303100048B3432C82904204006",
INIT_01 => X"210668000008004C1C20250E12100368403008418984014902030906A8910200",
INIT_02 => X"120404C0024C0600000206100008402404040C00F104008040080080001310E0",
INIT_03 => X"7728805052470B5C1B873C04121D03845D0020CA0822018000080084C1000002",
INIT_04 => X"0B899E43891686690790485D5C3E02000E9892201D306D03A9835C16029AC186",
INIT_05 => X"C001E080005030767434C0003C8A01D6B81C5703C82CDBC000072400089C8120",
INIT_06 => X"1000088100410000460002041300004084080070D00030032009700024641102",
INIT_07 => X"4261950408CCBC2012048310951000000003402A4000143E1008912480000211",
INIT_08 => X"00811007AC0A1EB5131120C79E7D176251E53E80E8B361604041340838452020",
INIT_09 => X"C08360820C0912800035F1801630A8260900180C00C8021C800FEE522020A108",
INIT_0A => X"8400F88C166262E940D00D410D62AD02091704024D0A02882192020DA0544043",
INIT_0B => X"4011078510C90D143142430C243042430C24304243042430C24305121A612186",
INIT_0C => X"C08060101000C00401008800F004140009400E4002A0010240000DC3C080002C",
INIT_0D => X"000800100001C07261C51C42390240F050C3C000950008088130040100018000",
INIT_0E => X"00080010003510004000000000000048010002E0100000000800100220100000",
INIT_0F => X"0000014008001550000800000000000400800280100000000800100360100000",
INIT_10 => X"00000000020000080080009410004000000000000044080000D8008000000000",
INIT_11 => X"000005800008000001040168000040000041000100EC00004002214000008000",
INIT_12 => X"00000041003C000008000008200D00001000000208050C000200000000002040",
INIT_13 => X"17000100000000000090000002C8000008000000000060000004480000400000",
INIT_14 => X"8400C00208004844C00800000000528008000000008000000000010040000000",
INIT_15 => X"0100800004030080000C010000A00D1804404912802A261B53104810DB1E0028",
INIT_16 => X"000C030000200C01000020040300800004030000000C03000000040100802004",
INIT_17 => X"008020040100C010000200800004010040300800000020040100C03000020000",
INIT_18 => X"40C700FC0A000280C68A08A950520E964C3269B2C9864D30000C030040100800",
INIT_19 => X"555555555555555555555555555554514514514514526991A199A28A28981451",
INIT_1A => X"41A0D068341A0D068341A0D068341A0D06A351A8D46A351A8D46A35555555555",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF771F60D068341A0D068341A0D0683",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FF087FFDF5508003FEBA087FD54BAAA841540055000000000000000000000000",
INIT_1F => X"F5500003DF455555421EFAAFFD54AAF7D168B45AAAABDF55A2802AA1000002AB",
INIT_20 => X"DFFFAAD1554005D7FD74AAAA840015500002AABA082E954005500021FF5D2EBF",
INIT_21 => X"68BEF080028BFF0855555455500174BAA2AABDE0055517FF555555420AAAA843",
INIT_22 => X"168ABA0055574BA5555554BA5D0400155AAD1554AAF7802AB4500043DF45FFD1",
INIT_23 => X"0400010A2AA955FF55003FE10F7803FEBAFFD5420BA085168A00007BFDE10085",
INIT_24 => X"855555FFAA84001FFAAFBEAB45002A97545F7D1555EF55043DF5555517DEAA5D",
INIT_25 => X"000000000000000000000000000000000000002A82155A2FBFFEBA0800021550",
INIT_26 => X"5BC042AA101D0A28BC7007FFDF45080A3AEAA007BD2482BE84124285C0000000",
INIT_27 => X"004100021FF492AB8F7D1C0438E381451471D7AAFBD0492EBD56DB7DBEAEBFF5",
INIT_28 => X"FED1C5F470AABE8A3AFD7A2DF55400557FD54AABE84001C5550A28ABA1424974",
INIT_29 => X"FB5508043FF55EBD56ABD75D0428BEF005557545490012482B6A0BAE2849557A",
INIT_2A => X"6DA101475FDE10145F68A921C55504924955524AA140E0717DAADB50492EB842",
INIT_2B => X"43AF6D405F78E3A1C2002000BEAA905C755003FE28E3803DEAAEBDF40002557F",
INIT_2C => X"FFFAE821C0A0717D1C5B575FFB6DF425575D7BEFB55002097555FFD5401EF5D0",
INIT_2D => X"784000AA59000000000000000000000000000000000000000000000208017DAA",
INIT_2E => X"A2D57FFFFF7AEBFF55FF8028A00512EAAB45007FFFF55082EA8AAA087FC2010F",
INIT_2F => X"5512AAAA085D04174100800021FF002EA8BEF5D0428ABA595557555AAFBC2000",
INIT_30 => X"00FF802ABAA04552ABFF597FD74BAF7AAA8B45AAFBD54005D7BD54AAF7800215",
INIT_31 => X"5FFAAFBC0000AF843FF5500003FF55AAFD6AB4551002ABEF0055555550004020",
INIT_32 => X"DEB0A2FD5600051537DE005D557DE005D7BE8AA85555400100879560AA592F95",
INIT_33 => X"17545FFD5421FF5D0428BEF0079FCABA598400010F7AA8215555003FEAAAA843",
INIT_34 => X"0000000004001FFAAFBEAA105D2E955FF557BD75EFFBBCD415521FBFDF450004",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000010000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(0),               -- Port A write enable input
DIA(0)   => data_write_a(4),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(4),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(0),               -- Port B write enable input
DIB(0)   => data_write_b(4),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(4),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_5_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50DB0A0791B1B41694368283C81F9996A091A32152007AB36B20E03C040C002",
INIT_01 => X"880015C49830884C446A40000C34C24841280A00084000C8C212892EEA953231",
INIT_02 => X"408F417400B1D9100002171C1FA20171124E6AA00D8633F8CD09DBFBBB972F7C",
INIT_03 => X"88538F0182058082D800C3314722DC08A34084A100C4D7C99208521063D00148",
INIT_04 => X"F45E41AFAF420996B8411CA282F80A9091224800A2C61490363080C8A4000308",
INIT_05 => X"0EA416069640420901A01505C4410020C6E228DC30532839B043289D9C005031",
INIT_06 => X"13992D9AF8C74E92B7B568D19708C038AFFA89F0B9348C9204C389672407EF12",
INIT_07 => X"6255000016053C18162589725146F442222CE6AF844012BE795224458BA4DE0F",
INIT_08 => X"4F3F00503B4AE104B5347230418190420821006016FC18843630D285FC416CB4",
INIT_09 => X"EEA33E700340902C4424C442B0344724066C56C2248130A2D9C185B24A24832B",
INIT_0A => X"315325008348CC40AB570500204462508135D5AA593E043731E9B18A98440137",
INIT_0B => X"E0CD463C5813804E0258E0358E02D8E03D8E0258E03D8E02D8E03447012C701E",
INIT_0C => X"F8DE3C27CA181E5D710664A5F140C14BD32A2E281992940AFAA15C3FC0836310",
INIT_0D => X"F000BE0FC80020130841840308653FF0313FE92C23FB1EECB367C0F3E378F0BC",
INIT_0E => X"F000BE0FCD806FFFAF0AE83080E2AEB2F0F1E01BE53FE1F000BE0FC41BE53FE1",
INIT_0F => X"0231F0BF9E3F02A7FFD63669C0E008C3CB7F041BE1BFE1F000BE0FC41BE1BFE1",
INIT_10 => X"30180309A0F83FE2B87C7D006FFF9F1A7806013879BAA78FC103FF5F1F12F038",
INIT_11 => X"39E9C1DBF8A30C2098DBE2FF7F2320483136F200A822CBACAB9DDEB7F9BC291F",
INIT_12 => X"004C72BEC95FEF64E4090626DF15B7D1C6184131B7980DFFFC03F00003F01FB9",
INIT_13 => X"1DFFFA0A3C0202B8776AE7A7C9CBFFF060703080E29F1B79E9F6427EFE901C0E",
INIT_14 => X"2B716CA5C56620590350ACD3A7D5B7EFAC6DFC8C0312A0024B83F07F3999E9F2",
INIT_15 => X"F0BCAF3BC2F3BC6F0BCEF2BC2F3BC6DBC67C251104A2261253904580207E1C81",
INIT_16 => X"1BCEF0BC2F3BC2F1BCEF0BC6F2BC2F1BCAF1BC6F2BC6F2BCAF1BC2F3BC6F2BCE",
INIT_17 => X"BCEF0BC2F3BC2F1BCAF1BCAF3BC6F0BCEF0BCEF2BC6F2BCAF1BCAF1BC2F3BCAF",
INIT_18 => X"69CFEF73B6FFE7436DB6FD0831518424965B4D2492CB69AF1BCEF0BC6F2BC6F0",
INIT_19 => X"F7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF3EF9FBFBB9E79E7BEBCB7",
INIT_1A => X"DEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDF7DF7DF7D",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF29FDAF77BBDDEEF77BBDDEEF77BBD",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"AAA2802AA10FFFFFDE0008556AABA5D2ABFFEFFF800000000000000000000000",
INIT_1F => X"ABAF7AAA8BFFAA802ABFF087FFDF5508003FEBA087FD54BA0804154005555574",
INIT_20 => X"54AAF7D168B45AAAABDF55AA802AA1000003FEBA00002AABA5D2EBFEBAAAD16A",
INIT_21 => X"3DE005555575EFA2D142145A2FFE8B45FF80001555D2E955FFFFD5421EFAAFFD",
INIT_22 => X"FC00BA5D5568AAAF7AAAAAAAAA802AABA082E954005500021FF5D2EBFF550000",
INIT_23 => X"D5420AAAA843DFFFAAD1554005D7FD74AAAA840014500517FFEF007BEABFF5D7",
INIT_24 => X"2AABDE0055517FF555504154BAA2FBEAA105D2E97410FFD16AAAA5D2ABDEBAFF",
INIT_25 => X"000000000000000000000000000000000000000028BFF0855555455500174BAA",
INIT_26 => X"21E84124285C51574BAB68A2DA00FFFFFFE38085F6FA92552AB8FEFF78000000",
INIT_27 => X"925D2AB8EBABEDB6AA92F7AAA8BC7B68A28BC70075FDF45080A3AEAA007BD248",
INIT_28 => X"5FFFFD1471D7AAFBD0492EBD56DB7DBEAEBFF55BE842AA105D0A38EBA1C0428A",
INIT_29 => X"21FF492AB8F7D1C0438E38145B575EFA2DB45145B6F5EFB6DF78E05145552A92",
INIT_2A => X"7DFC70875EABC7557FC20AA415F68AAAF7AAAAA82BE8A28A9214249740041000",
INIT_2B => X"B6FABA542ABAE2AF7DF470AABE8A3AFD7A2DF55400557FD54AABE84001C55551",
INIT_2C => X"5557545490012482B6A0BAE2849043AFED1C0E10492B6FFEFA105D2A95410FFD",
INIT_2D => X"D2AAABEFFB8000000000000000000000000000000000000000000000428BEF00",
INIT_2E => X"082EA8AAA087FC20105504000AA5955554BAFFAEBDE10F7FBFDEBA007BFDE005",
INIT_2F => X"0512AA8AAA5D0028A005D2AA8ABAF7FBE8A00FFAEAAB45F3AAAAB4500557FF55",
INIT_30 => X"EFFFAA97545552A821EFFBD557555AAFBC2000A2D57FFFFF7AEBFF55FF8028A0",
INIT_31 => X"A005D04174100800021FF002EA8BEF5D0428ABA597FD55FFA2FFD5555FFD57FF",
INIT_32 => X"54AAF7800015551517DF45005168B55557FC0012087FEAABAF7AAAAA10F3AAAA",
INIT_33 => X"FFE005D2A95410F7FFFFEBA5D2EA8ABAFBFFD74BAF7AAA8B45AAFBD54005D7BD",
INIT_34 => X"00000000002ABEF005555555000402000FF802AAAA04452ABFF592E80010FFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000060000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(0),               -- Port A write enable input
DIA(0)   => data_write_a(5),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(5),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(0),               -- Port B write enable input
DIB(0)   => data_write_b(5),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(5),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_6_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10800B0061A01002840002C030028180004003220200403312301C4389B2082",
INIT_01 => X"060009C838394848188160000C42426041000000090800090210090000510200",
INIT_02 => X"00043040009001100000061000018070002408000000000648080000001210E0",
INIT_03 => X"0000800002054081020080801200A0000300008000201184681A0000410C4800",
INIT_04 => X"0808801040000001401048008100022401400002024024053200020089000100",
INIT_05 => X"0240040408402202002000C200400020A50000A0000010010001260808000520",
INIT_06 => X"44000881064500004600000013088002840C240F5048011200010000440C0146",
INIT_07 => X"0241914041FE83E010040110110003040020402A0000003E1000000488000201",
INIT_08 => X"8001BF002C4A01041B112020200110024029006FE09081002004902000012068",
INIT_09 => X"0083FE38A040100281353150ACB645AEF8C01404448000008011061204200108",
INIT_0A => X"3103AD0413424E4014D627C470462200011504420C0A962A2189002881404060",
INIT_0B => X"46C1060C16C96D15B0425B0425B1425B1425B0C25B0C25B1C25B1512D8212D82",
INIT_0C => X"009000140401100601016600A040220203A004480598010248000D0010420C0C",
INIT_0D => X"0000A01033A00013000000000018800F2400091081100C0090A5008200410020",
INIT_0E => X"0000A0103142000000000000000000455D0018100000000000A0103410000000",
INIT_0F => X"000000466800C200000000000000000001A0F4100000000000A0103410000000",
INIT_10 => X"00000000000024094680014200000000000000000041E8002900000000000000",
INIT_11 => X"F000322000000000000D1A000000000000034D240C2000502000000000000000",
INIT_12 => X"000000403F4000000000000068D24000000000001A60F0000000000000002007",
INIT_13 => X"C0000000000000000087C0003014000000000000000025D00008958000000000",
INIT_14 => X"02000000000814C219500150002800101280000000000000000000086670000C",
INIT_15 => X"8120C82208812048120882208892055A0060011280222413130449010301F051",
INIT_16 => X"3200802008320C82200802048320C82200812048320880200812048220880204",
INIT_17 => X"20C83208812048020883204802048120882204812008220C8220081204822088",
INIT_18 => X"79CFF1FE1E9F52ABEF9EFE8150120EC718638E38E30C71C812088220C8120080",
INIT_19 => X"71C71C71C71C71C71C71C71C71C71C71C71C71C71C736D9DBD9BBEFBEFBEBEF1",
INIT_1A => X"CFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FC71C71C71C",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCF29A7F3F9FCFE7F3F9FCFE7F3F9F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000607FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"EFA2FBD54BA5555554BAAAFBC20BA5D7BEAAAAFF800000000000000000000000",
INIT_1F => X"EBA0855421455555574AAA2802AA10FFFFFDE0008556AABA5D2ABFFEFFF843DF",
INIT_20 => X"DF5508003FEBA087FD54BA000415400550428AAAAA84021FF007BD54BAAAD17D",
INIT_21 => X"A8BFFAAD1554BA002A95555A28417400AAFBE8ABAF7FFD54AAAA802ABFF087FF",
INIT_22 => X"BD5545080417555A2D17FE1000003FEBA00002AABA5D2EBFEBAAAD16AABAF7AA",
INIT_23 => X"D5421EFAAFFD54AAF7D168B45AAAABDF55AA802AA100000001EF087FEAA00FFF",
INIT_24 => X"F80001555D2E955FFFF843DEAAA2803DFEF0855401FF082EA8B555D7FC21FFFF",
INIT_25 => X"0000000000000000000000000000000000000055575EFA2D142145A2FFE8B45F",
INIT_26 => X"2552AB8FEFF78E3DFFFAAFFD04AA415B52492B6F5C20825D7FE8A92FF8000000",
INIT_27 => X"EF147BD2482BED57AE921451421555551574BAB68A2DA00FFFFFFE38085F6FA9",
INIT_28 => X"4BAB68A28BC70075FDF45080A3AEAA007BD24821C04124281C0E2DA82BE8E001",
INIT_29 => X"8EBABEDB6AA92F7AAA8BC7B6D5524AA14209557DA28E15400BEF1EFA92FFFFD2",
INIT_2A => X"071FF0071EDA38F7F1D5555000417545B6D178E281C0A38EBA1C0428A925D2AB",
INIT_2B => X"4A8B555C7FC2147F7D1471D7AAFBD0492EBD56DB7DBEAEBFF55BE842AA105D0E",
INIT_2C => X"DB45145B6F5EFB6DF78E05145552A925FFFF8E3DE82BE8E38FFF0851401C7082",
INIT_2D => X"57FE8A00F38000000000000000000000000000000000000000000005B575EFA2",
INIT_2E => X"F7FBFDEBA007BFDE005D2AAABEFFBAABDFEFAAFBC00BA007BC0000FFD5420005",
INIT_2F => X"A592ABFE00F7AA821FF557FC0010F7D168A105D55421455155554BAFFAEBDE10",
INIT_30 => X"10F7D57DE00FFFBC00AAFBAAAAB4500557FF55082EA8AAA087FC20105504000A",
INIT_31 => X"AAA5D0028A005D2AA8ABAF7FBE8A00FFAEAAB45F3D5400BA5504155EFAAAE954",
INIT_32 => X"FF55FF8028A00512E975FF08557FEAAF7D157545080417545F7D56AAAA592AA8",
INIT_33 => X"AABEF005542155000028B555D7FC2145F3D557555AAFBC2000A2D57FFFFF7AEB",
INIT_34 => X"000000007FD55FFA2FFD5555FFD57FFEFFFAA97545552A821EFFBAABDE00F7AA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000048000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(0),               -- Port A write enable input
DIA(0)   => data_write_a(6),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(6),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(0),               -- Port B write enable input
DIB(0)   => data_write_b(6),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(6),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_7_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10844B00482258A2842112C02450418800002300500030B313300C418992002",
INIT_01 => X"020009C23838684D1C20E0000E11424840000000080000080200000000110204",
INIT_02 => X"000520700CA08910000206101180803081144880010400044808000000122160",
INIT_03 => X"000080040305208000008000328080040304008020303194289A000041484800",
INIT_04 => X"08088000000000010000CA008008060441000000028234493410820191000000",
INIT_05 => X"03500404000022020020044000000C208400408000001000984005949C002928",
INIT_06 => X"54000881044500004680000013008002940C24001A4A010200018920646410C7",
INIT_07 => X"22510040400500011204813015012204002040280000013E1000000488000201",
INIT_08 => X"9001A0602C4A01051B132820208001024069004008908002120851420001226A",
INIT_09 => X"01100020A2401008A20404E08200A05000A4264640800022C8198C4E05200018",
INIT_0A => X"20002000024040400050450440C48A0041140C420B0904208800904286000008",
INIT_0B => X"50822002120D2134800648006480064800648106481064810648193240432404",
INIT_0C => X"284A142288042A5C24202451505E00A621A5220A8091444040188C001B41210A",
INIT_0D => X"00F001F021141A12004104020810B000100000000109064C80010050A3285194",
INIT_0E => X"00F001F027420000400004C3201C514408081C1014800000F001F02810148000",
INIT_0F => X"E00E0E404100E200040900000B0380383480C81014800000F001F02810148000",
INIT_10 => X"4160C0301D07001D0402034200004000019860078641004039000180400002C0",
INIT_11 => X"08103BA0104810C8462416E8040446120C890814600010512000000080028400",
INIT_12 => X"98038D4030DD008088C2419120B740209021908C4846FC000200030F000FE006",
INIT_13 => X"DD000100411C81078884204035DC00201804C3201C60A408100DD58010440130",
INIT_14 => X"412024202211148019064200402A32901A8000B2048902C0807C0E00C448100D",
INIT_15 => X"50942509425194651946519465894619421421102000269243854D8002000250",
INIT_16 => X"19465194E50942509425094E51946519465094A50942509425194E5194651942",
INIT_17 => X"9425094251946539465094250946539465194250942509465194650942509425",
INIT_18 => X"0000000000000000000000080150890820800041041000052942509465194653",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF21E6C000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"AAF7D5575455D557DFEF002AAAB55002E820AAAA800000000000000000000000",
INIT_1F => X"B55007FD74AAAA843DFEFA2FBD54BA5555554BAAAFBC20BA5D7BEAAAAFFFBC00",
INIT_20 => X"AA10FFFFFDE0008556AABA5D2ABFFEFFFAAAAAAAF7D57FFEFF7D555555A2AEAA",
INIT_21 => X"42145552ABDFEFFFAA801EFFFFBFDF550000175555504175450055574AAA2802",
INIT_22 => X"A975EF00003DF55555168A00000428AAAAA84021FF007BD54BAAAD17DEBA0855",
INIT_23 => X"802ABFF087FFDF5508003FEBA087FD54BA000415400557BD74BAFFD140000082",
INIT_24 => X"AFBE8ABAF7FFD54AAAAAEA8ABA55557FEAAA2843FF55A2AEA8B55AAAABDEAAFF",
INIT_25 => X"0000000000000000000000000000000000000051554BA002A95555A28417400A",
INIT_26 => X"25D7FE8A92FFFFC70BAE3D155555415178FD7082EAAB550820870BAAA8000000",
INIT_27 => X"FFEBD55557DBEA4AFB550871D7482AA8E3DFFFAAFFD04AA415B52492B6F5C208",
INIT_28 => X"5550051574BAB68A2DA00FFFFFFE38085F6FA92552AB8FEFF7A0ADABAEBD578F",
INIT_29 => X"2482BED57AE921451421555524BDFD7FFA4801D7F7F5FDF55000E17545410E17",
INIT_2A => X"D2482E3D1450381C20905EF08003AF55415F6DA38080E2DA82BE8E001EF147BD",
INIT_2B => X"AAFB55ABA0BDE02EB8A28BC70075FDF45080A3AEAA007BD24821C04124281C7B",
INIT_2C => X"209557DA28E15400BEF1EFA92FFFFD24BAB6A4A8A82495F78E92AA843DF45BEA",
INIT_2D => X"800174BAA680000000000000000000000000000000000000000000055524AA14",
INIT_2E => X"007BC0000FFD542000557FE8A00F3FFD54BAAAD15754508556AB45002AA8B450",
INIT_2F => X"FFB803DEAAAAD56ABEFAAD5575EFF7803DF45085557410AEAABDFEFAAFBC00BA",
INIT_30 => X"55082E97555002E955550C55554BAFFAEBDE10F7FBFDEBA007BFDE005D2AAABE",
INIT_31 => X"E00F7AA821FF557FC0010F7D168A105D554214551003FF45FF8400145FFD57FF",
INIT_32 => X"20105504000AA597FC2010A2D1554AA5500021EF000028B55087BFDEBA042ABF",
INIT_33 => X"E8A00A2803FF45F7AABDF55AA843FE10AEAAAAB4500557FF55082EA8AAA087FC",
INIT_34 => X"0000000055400BA5504155EFAAAE95410F7D57DE00FFFBC00AAFB8028A00007F",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000007FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(0),               -- Port A write enable input
DIA(0)   => data_write_a(7),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(7),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(0),               -- Port B write enable input
DIB(0)   => data_write_b(7),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(7),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_8_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000B0000040042840002C0000001800000070000000033022000000000086",
INIT_01 => X"000009C21838284D1C2160000E12426840000000180800080200080040510200",
INIT_02 => X"0001004000900110000006100080003000240800014400004808000000122160",
INIT_03 => X"00008000020440810002A0801010A0044300000000200086011A000040404800",
INIT_04 => X"8000801000020401400040408108022029400000124004041200000089000100",
INIT_05 => X"02080424085022020000040200480020850010A0002010010120060800040400",
INIT_06 => X"50000880006500000680000011008006840C200018C1010200018920E0640102",
INIT_07 => X"426000404005000112048130150120240020400A0000013E1000000488000010",
INIT_08 => X"220100402C42010413110020200100024029004000A200002004902200012141",
INIT_09 => X"0000000080400008010410A2940A45240040140440800022C8388E1200A00008",
INIT_0A => X"00420100020048405000070440C0000001140412090000000021002081000048",
INIT_0B => X"0000000800000100011000010000100001000010000100001000010000880008",
INIT_0C => X"001000040001100008012008004020102180800804802000C0080D00100A0008",
INIT_0D => X"0FF0000002200A1200410402080080003000091085100C008124008000400020",
INIT_0E => X"0FF000000140000040F517CF600000000104081010001E0FF00000001010001E",
INIT_0F => X"E000000000804200000809963F1F80000000001010001E0FF00000001010001E",
INIT_10 => X"CFE7C0F00000000000810140000040E587F9E000000008100900008000ED0FC7",
INIT_11 => X"00021040030C73D80000021000585F3600000020240020102000000802419660",
INIT_12 => X"F80000000042000B0BD6C0000010800618E7B000000C000003F80FFF00000000",
INIT_13 => X"800005D5C3FD800000000008180000078A8FCF600000000002028001006AA3F1",
INIT_14 => X"020000000008808219002100100C000041120370DCAD1FC18000000000000202",
INIT_15 => X"8020080200812048120481204812055A04604930A02026934215410102000110",
INIT_16 => X"0200802008020080200802048120481204812048120481204802008020080200",
INIT_17 => X"2008020081204812048120481200802008020080200802048120481204812048",
INIT_18 => X"414A87D78AF42143CEBAC88151120A0000000000000000081204812008020080",
INIT_19 => X"F3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF7E799B1BEB65B65948051",
INIT_1A => X"C3E9F0FA7C3E9F0FA7C3E9F0FA7C3E9F0F87C3E1F0F87C3E1F0F87CF3CF3CF3C",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF1B5DA9F0FA7C3E9F0FA7C3E9F0FA7",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"0000043DF55087BC01EF007FD75FFFF84000AAFF800000000000000000000000",
INIT_1F => X"E10A28028AAAAAFBC00AAF7D5575455D557DFEF002AAAB55002E820AAAA84000",
INIT_20 => X"54BA5555554BAAAFBC20BA5D7BEAAAAFFAA95545552ABFE00087BC00AA082EBF",
INIT_21 => X"D74AAAAD57FF45002A975FF007BE8BFFA2FBFFFFFAAD5400AAFF843DFEFA2FBD",
INIT_22 => X"BE8A00082A97410F7D5555EFAAAAAAAAAF7D57FFEFF7D555555A2AEAAB55007F",
INIT_23 => X"55574AAA2802AA10FFFFFDE0008556AABA5D2ABFFEFFFAA82000555555545AAF",
INIT_24 => X"00017555550417545000015545087BC2010AAD54014500516ABFFA2AABDF4500",
INIT_25 => X"000000000000000000000000000000000000002ABDFEFFFAA801EFFFFBFDF550",
INIT_26 => X"50820870BAAA8407000140038F450075C71FF087BD75D7FF84050BAEB8000000",
INIT_27 => X"10007FC50BA002ABFE00AA8A2AABABEFFC70BAE3D155555415178FD7082EAAB5",
INIT_28 => X"082EB8E3DFFFAAFFD04AA415B52492B6F5C20825D7FE8A92FFA497545552AB8E",
INIT_29 => X"557DBEA4AFB550871D7482AAD17DF451C24955EF0875EFBD7B6F1FFFC7BEDB45",
INIT_2A => X"87000415B5057DAAFBE8A10082092410EBD5505EFB6A0ADABAEBD578FFFEBD55",
INIT_2B => X"B6ABC7B6AABFFED0051574BAB68A2DA00FFFFFFE38085F6FA92552AB8FEFF7AA",
INIT_2C => X"A4801D7F7F5FDF55000E17545410E17555000E17545007BC0000BED14217D005",
INIT_2D => X"784174AAA280000000000000000000000000000000000000000000024BDFD7FF",
INIT_2E => X"08556AB45002AA8B450800174BAA684174105D042AB550055555FF007BD7555F",
INIT_2F => X"0F384175555D2EA8A00087BD74BA082EBDE10AAAEA8ABAF7FFD54BAAAD157545",
INIT_30 => X"55FFD57DF55FFFBD5400A2AABDFEFAAFBC00BA007BC0000FFD542000557FE8A0",
INIT_31 => X"EAAAAD56ABEFAAD5575EFF7803DF45085557410AED17FF455D04155FF00557DF",
INIT_32 => X"DE005D2AAABEFFBAE97410087BC21EFA2FFEAA00000002010A2D5421FFFF803D",
INIT_33 => X"C0010FFD1401EF087FE8B55FFAEBDFEF0855554BAFFAEBDE10F7FBFDEBA007BF",
INIT_34 => X"00000000003FF45FF8400145FFD57FF55082E97555002E955550C2E95555087B",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000020000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(1),               -- Port A write enable input
DIA(0)   => data_write_a(8),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(8),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(1),               -- Port B write enable input
DIB(0)   => data_write_b(8),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(8),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_9_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00018248A2840112C00002C18000002300500030B3132000400812002",
INIT_01 => X"A140098218302849180060000C004240413C0A61590001D90213C90008510204",
INIT_02 => X"102008700CB089100002061031285074810448800104008048080080001210E2",
INIT_03 => X"00008015074608840390A0040040800203140000A00010800408108448020042",
INIT_04 => X"082080400004A00100000100840602020100000002C2344156108201811801C0",
INIT_05 => X"0200048480011502049500280020CC2084000080008010019161249C9C002188",
INIT_06 => X"70000881004500004E01020411D08000940C00001800010200018B20206C0102",
INIT_07 => X"EA70C0040005000312048130150100040020404A0000017E10408104C8000110",
INIT_08 => X"000000402C220104131004202081120050A5104000A204617201D10801002000",
INIT_09 => X"000800002F4924003085E51420A0100400641E4E40800022C8088C1220200908",
INIT_0A => X"20102000024040484028450001648C2229150400080244000401900284000440",
INIT_0B => X"0880110901081110411204112040120411204012041120401204111020090208",
INIT_0C => X"685B34A688841A5C21200101A01A0004009024028004044248404D00104B2100",
INIT_0D => X"0000A01000000213000000000000B0001000010000190E44802002D1A168D0B4",
INIT_0E => X"0000A010014000000000000000000040500008100400000000A0100410040000",
INIT_0F => X"0000004608004200040000000000000001A004100080000000A0100410008000",
INIT_10 => X"00000000000024080000014000000000000000000040A0000900010000000000",
INIT_11 => X"300013E010000000000D00F804000000000340000C0000102000000080000000",
INIT_12 => X"00000040091F0000800000006807C000800000001A0CFC000000000000002001",
INIT_13 => X"DD000000000000000082C00019DC002000000000000021500006D58010000000",
INIT_14 => X"03206420000000C019502050000C32901A800080000000000000000860100006",
INIT_15 => X"D1B46D1B46D0B42D0B42D0B42D8B424342342832002A24921082158802001011",
INIT_16 => X"0B42D0B42D0B42D0B42D0B46D1B46D1B46D1B46D1B46D1B46D1B46D1B46D1B46",
INIT_17 => X"B42D0B42D1B46D1B46D1B46D1B46D1B46D1B46D1B46D1B42D0B42D0B42D0B42D",
INIT_18 => X"89999E91BCD1512B871C4A0100000000000000000000000D0B42D0B42D0B42D0",
INIT_19 => X"A28A28A28A28A28A28A28A28A28A29A69A69A69A69A51C200807249041202AE6",
INIT_1A => X"8349A4D068341A0D269341A0D269341A0D068341A0D068341A0D068A28A28A28",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF2DA921A0D269341A0D068349A4D06",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"45A280154BA5555401EFFFD5421EFA2FFFFF555D000000000000000000000000",
INIT_1F => X"5EF00557DF555D040000000043DF55087BC01EF007FD75FFFF84000AAFFD57DF",
INIT_20 => X"75455D557DFEF002AAAB55002E820AAAA843DFEF00517DEBA007BFDFEFFFD157",
INIT_21 => X"28AAAAAAABDF45F7803FFEF555568AAAF7802AA00FFFBD7555087BC00AAF7D55",
INIT_22 => X"BD54BA550417400085155555082A95545552ABFE00087BC00AA082EBFE10A280",
INIT_23 => X"043DFEFA2FBD54BA5555554BAAAFBC20BA5D7BEAAAAFFFBC00AA552E95545087",
INIT_24 => X"2FBFFFFFAAD5400AAFF8402000A2FFFDF555D7BE8BFF5D51575EFA280175555D",
INIT_25 => X"00000000000000000000000000000000000000557FF45002A975FF007BE8BFFA",
INIT_26 => X"7FF84050BAEBDF78F45B68010482415B471C7E3DF451EFBEFBFAF45490000000",
INIT_27 => X"82007FFAFEFE3DB505EF1C5B7AF45490407000140038F450075C71FF087BD75D",
INIT_28 => X"5451C7FC70BAE3D155555415178FD7082EAAB550820870BAAA8438FFF00517DE",
INIT_29 => X"50BA002ABFE00AA8A2AABABEAEB8F45F78A3DFD741516DAAAE38E2DA28EBFFD5",
INIT_2A => X"C20BA5D2E905550071D54825D0A1543808515756D1C2497545552AB8E10007FC",
INIT_2B => X"5505FFBE801256D490E3DFFFAAFFD04AA415B52492B6F5C20825D7FE8A92FFFF",
INIT_2C => X"24955EF0875EFBD7B6F1FFFC7BEDB45082EB8002000AAFFFDF6D417FEABEF5D5",
INIT_2D => X"7FBE8B5500000000000000000000000000000000000000000000000517DF451C",
INIT_2E => X"0055555FF007BD7555F784174AAA2FBEAB45F78402010007BD5545AAFFD55EFF",
INIT_2F => X"AA68028BEF00517FE10007BE8BFFAAFFC01FF557FE8B550004174105D042AB55",
INIT_30 => X"AAAAAEBFEAAAAFFD5545557FD54BAAAD15754508556AB45002AA8B450800174B",
INIT_31 => X"5555D2EA8A00087BD74BA082EBDE10AAAEA8ABAF7AAAAB45F7AEBFF4508557FE",
INIT_32 => X"2000557FE8A00F3FFC00BA552E80145005557400552A954BA0051575EF550417",
INIT_33 => X"FDFFF007FE8BFF5551401EFF784021FF002ABDFEFAAFBC00BA007BC0000FFD54",
INIT_34 => X"00000000517FF455D04155FF00557DF55FFD57DF55FFFBD5400A28400010A2FB",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000040000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(1),               -- Port A write enable input
DIA(0)   => data_write_a(9),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(9),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(1),               -- Port B write enable input
DIB(0)   => data_write_b(9),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(9),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_10_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00018248A2840112C00002C18000202300500030B3132000400992006",
INIT_01 => X"A140098218302849180060000C00424040000000080000080200090008510204",
INIT_02 => X"102100400C8001100000061000A8503401044880010400004808000000122160",
INIT_03 => X"000080150746088401908000100080020304000020201080001A108448404842",
INIT_04 => X"800080400004A001000040008406020201000000020004401000000180180080",
INIT_05 => X"02000484800133020495040800208C20A4000080000010000001249010042008",
INIT_06 => X"50000881004500004681020411808000940C20001800010200018920206C0102",
INIT_07 => X"024084044005000112048130150120040020400A0000013E10408104C8000010",
INIT_08 => X"000100402C020105131100200000124250A51040088084614001110801012000",
INIT_09 => X"00080082CD09240820800000000000040000180840800022C8088C1220200108",
INIT_0A => X"841201000200484910000F050560262229140402080200A00402000484140400",
INIT_0B => X"0010118900080010000200102001020000200002001020010200001000010008",
INIT_0C => X"408120900404004821202001F05E00040180260A8080044240004C0010800228",
INIT_0D => X"0000A01000000813004104020800800030000800010008088124020102008100",
INIT_0E => X"0000A010014000004000000000000040500008101480000000A0100410148000",
INIT_0F => X"0000004608004200040900000000000001A004101480000000A0100410148000",
INIT_10 => X"00000000000024080000014000004000000000000040A0000900018040000000",
INIT_11 => X"3800100010480000000D00000404400000034000282000102000000080028000",
INIT_12 => X"00000040090000808800000068000020900000001A0000000200000000002001",
INIT_13 => X"80000100000000000082E0001000002018000000000021580000800010440000",
INIT_14 => X"00004000000004C0195000500008000000000082008000000000000860180000",
INIT_15 => X"0100401004010040100401004090055804404110802A24921317580802001011",
INIT_16 => X"0000000000000000000000040100401004010040100401004010040100401004",
INIT_17 => X"0040100400000000000000000000000000000000000000000000000000000000",
INIT_18 => X"215281FC1A72E2486AAA40A85052020000000000000000001004010040100401",
INIT_19 => X"51451451451451451451451451451451451451451452AA83330A8A28A29EA8D1",
INIT_1A => X"5CA6532994CA6532B95CAE572994CA6532994CA6532994CA6532994514514514",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF31CE2E572994CA6532994CAE572B9",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"10AAFBE8AAAA2D540000F7D57DF55A2AABFFEF08000000000000000000000000",
INIT_1F => X"F45FFFBC2010AAD57DF45A280154BA5555401EFFFD5421EFA2FFFFF555D003FE",
INIT_20 => X"DF55087BC01EF007FD75FFFF84000AAFF8002155AAFFE8B45AAD540000087FFD",
INIT_21 => X"7DF555D517FEBA082A801EFF7FBD5400FFD568B555D00155EF08040000000043",
INIT_22 => X"BFDE00A2FBC0145005168A10AA843DFEF00517DEBA007BFDFEFFFD1575EF0055",
INIT_23 => X"7BC00AAF7D5575455D557DFEF002AAAB55002E820AAAA803FEBA082AAAAAAF7F",
INIT_24 => X"7802AA00FFFBD7555082E82155FFAEAAB55AAD568B455D00154BAFFFBD75EF5D",
INIT_25 => X"000000000000000000000000000000000000002ABDF45F7803FFEF555568AAAF",
INIT_26 => X"FBEFBFAF4549003DE10BEF5EDAAAAAD547038EBD57DF7DA2AEB8FC7000000000",
INIT_27 => X"6DAADF470280075FFF45E3F1C7038A2DF78F45B68010482415B471C7E3DF451E",
INIT_28 => X"5C7000407000140038F450075C71FF087BD75D7FF84050BAEB8002155BEF5EDB",
INIT_29 => X"AFEFE3DB505EF1C5B7AF45495B7DEAA0824851EFEBFBD2410EBD168B7D410A17",
INIT_2A => X"38EAA0824A8AAAEBF5FAE28AAF1C2155005F68A10A28438FFF00517DE82007FF",
INIT_2B => X"4104AAF7F1D75EF557FC70BAE3D155555415178FD7082EAAB550820870BAAA80",
INIT_2C => X"8A3DFD741516DAAAE38E2DA28EBFFD55451C2087155EBA4A8B7DAADF68B7D410",
INIT_2D => X"2AEAAB55000000000000000000000000000000000000000000000002EB8F45F7",
INIT_2E => X"007BD5545AAFFD55EFF7FBE8B5500043FE00F7D17FEBAA2D5574BAAAD17DFEFA",
INIT_2F => X"AA28002155FFD17FFFFA2FBD74BA00557FF45A2D5554AAA2FBEAB45F78402010",
INIT_30 => X"00AAD16ABFF002A975450004174105D042AB550055555FF007BD7555F784174A",
INIT_31 => X"BEF00517FE10007BE8BFFAAFFC01FF557FE8B55007FFDEAA0004175FFA2FBC20",
INIT_32 => X"8B450800174BAA68428AAA08042AABAAAD56AABAAAD140155087FEAA10A28028",
INIT_33 => X"2ABEFAAFBE8BFF0004020AAFFD5555EF557FD54BAAAD15754508556AB45002AA",
INIT_34 => X"000000002AAAB45F7AEBFF4508557FEAAAAAEBFEAAAAFFD5545550015555A284",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000047FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(1),               -- Port A write enable input
DIA(0)   => data_write_a(10),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(10),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(1),               -- Port B write enable input
DIB(0)   => data_write_b(10),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(10),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_11_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10180B05A0010402840602C2D001019000000300000000330A20080EC180002",
INIT_01 => X"AB400984B830084C1820E0000C36424840000000080000088200000802112220",
INIT_02 => X"102A68440080011000000618062AD03502640800010410424908136019920868",
INIT_03 => X"001282118644C88481908001106088022300000080F4925CDC9A10844A9A4842",
INIT_04 => X"401280480004A1011000418084460002E12000000200040010000040A8000000",
INIT_05 => X"0FC8048484011502059511488020802084400888001110000000050000005400",
INIT_06 => X"1011088AE24500001631024511C08004A70AA40008B90D0200018B60A0650D45",
INIT_07 => X"020011005405000910040150110041040024400D800002BE18408104C9205908",
INIT_08 => X"89390040280241041D175820000001020061004004800567403512A801014C46",
INIT_09 => X"050800E20D09A424C5840400808000040680180840800022D8288E946CA00833",
INIT_0A => X"85002000024040410A000D0504408C32E915D9C208050084840201A099100400",
INIT_0B => X"B01011934A005101431CA821CA831CA821CA831CA831CA821CA83165410E5410",
INIT_0C => X"00010080028000010402214850444091019B02080885200042A9CC001000003A",
INIT_0D => X"5A5018C5A0A00812004104020808B00030000808024008008325820000000000",
INIT_0E => X"5A5018C5AB0062C38A4DB680A0D8241500D5761B011986695014A96E1A811986",
INIT_0F => X"42056A289A1BB2078A922DA2A8B180A2600AAE1A811986695014A96E1B011986",
INIT_10 => X"05AA429189B60AC43C6C7F0272C3841DB528802CAB18468F4101621B1BAC8455",
INIT_11 => X"C003104289A668B8CAB270106338317A3D94392020224ACDE215883078681B5C",
INIT_12 => X"804B020A06020C67061BC785938085134CD551BCA1C90006C0C2958502861120",
INIT_13 => X"80819A5539D503336D61056ABA006282806CA64090B89E015AAA880E48382EB8",
INIT_14 => X"40000000E808989003066E03513E41470126C6284B2D20410AB4503089C00A82",
INIT_15 => X"0000000000000000000000000000041800400110200026124202500802000800",
INIT_16 => X"1004010040100401004010000000000000000000000000000000000000000000",
INIT_17 => X"0040100401004010040100401004010040100401004010040100401004010040",
INIT_18 => X"C110083018162148420840280050800000000000000000001004010040100401",
INIT_19 => X"000000000000000000000000000001041041041041003882928E0000000AA0C4",
INIT_1A => X"0000000000008040000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3E0FC000000000000020100000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"EFAA842ABEFA280155EFFFFBC01EF08554000055000000000000000000000000",
INIT_1F => X"F4508514000000003FE10AAFBE8AAAA2D540000F7D57DF55A2AABFFEF0804155",
INIT_20 => X"54BA5555401EFFFD5421EFA2FFFFF555D51575FFA2FFD75FF550015400FFFBFF",
INIT_21 => X"C2010AAD568AAAAAD142145FF80155EF0051555FF0804155FFF7D57DF45A2801",
INIT_22 => X"01540008514215555003DFFFA28002155AAFFE8B45AAD540000087FFDF45FFFB",
INIT_23 => X"040000000043DF55087BC01EF007FD75FFFF84000AAFF802ABFFA2AABFE10080",
INIT_24 => X"FD568B555D00155EF085168B45085142010FFAE800AA5D7BFDF45F7FFEAA0000",
INIT_25 => X"00000000000000000000000000000000000000517FEBA082A801EFF7FBD5400F",
INIT_26 => X"DA2AEB8FC70000175EFB6802DBC7BE8A155EFE3FBC71FF145B42038550000000",
INIT_27 => X"EF550E15400E3F1FFF7D085B420381C003DE10BEF5EDAAAAAD547038EBD57DF7",
INIT_28 => X"5C7F7DF78F45B68010482415B471C7E3DF451EFBEFBFAF45495F575FFBEF5D05",
INIT_29 => X"70280075FFF45E3F1C7038A2DB68ABAB6D145145FF84155D7085B555C7140410",
INIT_2A => X"28BEFBEA4BDE28140A1543800514515549003FFC7BE8002155BEF5EDB6DAADF4",
INIT_2B => X"FFFF7DE3F1EFA10140407000140038F450075C71FF087BD75D7FF84050BAEB84",
INIT_2C => X"24851EFEBFBD2410EBD168B7D410A175C7005B6DB55145140000FFAE85082417",
INIT_2D => X"57BC20AA5D0000000000000000000000000000000000000000000005B7DEAA08",
INIT_2E => X"A2D5574BAAAD17DFEFA2AEAAB550004175FFF7803DF45FFAE955EFAAFBD55EF5",
INIT_2F => X"5007FD75FFF7D5401EF5D2E97410AAD17DFEF007FC20AA5D043FE00F7D17FEBA",
INIT_30 => X"55007FD5545550400145FFFBEAB45F78402010007BD5545AAFFD55EFF7FBE8B5",
INIT_31 => X"155FFD17FFFFA2FBD74BA00557FF45A2D5554AAA2FBEAAAAFFD555545FF80155",
INIT_32 => X"7555F784174AAA2842ABEFFF803DEAA5D2E974AA00515754500003FF55FF8002",
INIT_33 => X"40000FFAE97410007BFFFFFA2D57FE105D04174105D042AB550055555FF007BD",
INIT_34 => X"000000007FFDEAA0004175FFA2FBC2000AAD16ABFF002A97545007FFFF455555",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000040000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(1),               -- Port A write enable input
DIA(0)   => data_write_a(11),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(11),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(1),               -- Port B write enable input
DIB(0)   => data_write_b(11),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(11),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_12_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50080B01BC002006940202C0DE041196A83183000000023322287E0FC000006",
INIT_01 => X"0E000C068000E04D40238000001702484000000008000008820009280A553231",
INIT_02 => X"400B71440C8001100000171C0283813013766A800586235ECC09C8423B962966",
INIT_03 => X"CC618E048306E082000081000040900003548421A080025EDF08421042DC0108",
INIT_04 => X"00028020000000812000012080080000E100001002000448100000C1BC18008C",
INIT_05 => X"0FF8060610000402010015E100004C2084800090000310000000079010007C19",
INIT_06 => X"33992D98DEC74A003EA468D01510C03E8F580C800A3F018200418927E0668645",
INIT_07 => X"0204000406050013142409121142F746222EE2498000007E111204058B84C50C",
INIT_08 => X"E826A0602902A10491165C200000820018A5104010C01086003C13E000004EDF",
INIT_09 => X"023000000000000867000000000000040000600060801022C9F88D244FA40133",
INIT_0A => X"00100000820040482B28050001600010C13499F01B334015980001E09F000000",
INIT_0B => X"B80460124F16F06BC20CBC30CBC20CBC20CBC30CBC20CBC20CBC3065E1865E10",
INIT_0C => X"00000000029D204B7C0382FD0100F3F9F80FA0200E0BF40063F99C0010000012",
INIT_0D => X"93900F6EE230301208008001007A80001100002002801000A042000000000000",
INIT_0E => X"93900F6EEC421392C96B1237E0D8BD9629F97E0B348EDAC3900F6EFA0B158EDA",
INIT_0F => X"622DBC31D73F6006A5891533EF9500EAE64BCA0B158EDAC3900F6EFA0B348EDA",
INIT_10 => X"C2B083798D341B10DEFE14400392C74CAEAD412EDD2B4FCFF812A383430C669E",
INIT_11 => X"49FAB442994B3238D4E2FB104636652E19B8BA30C022DAD8C100CA39E8CEBE66",
INIT_12 => X"30469392526208C6CC95C33717D88532966471A9C5DD00B12728D5360234D62A",
INIT_13 => X"828C4999AF580395542D27CDBA0020F0FABAC800DA550C29F36A8A2554E48A64",
INIT_14 => X"40000000873FB80B8A00EF03F56CC12B416A51B60585A5C28895962502E9F36A",
INIT_15 => X"0000000000000000000000000000008000000410802A26924010000002000EE0",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"28C1111026C152A121960A884042020000000000000000000000000000000000",
INIT_19 => X"2082082082082082082082082082092492492492492400200005A8A28A200A37",
INIT_1A => X"964B2592C964B2592C964B2592C964B2590C86432190C86432190C8208208208",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF400FEB2592C964B2592C964B2592C",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FF00042ABEFFF8400010082EAABFF55002ABEF08000000000000000000000000",
INIT_1F => X"BEFFFFBD54000004155EFAA842ABEFA280155EFFFFBC01EF0855400005555421",
INIT_20 => X"8AAAA2D540000F7D57DF55A2AABFFEF08556AA10000028AAAFFD15541000002A",
INIT_21 => X"40000005168AAA087BFFFFF5D04001FF00041554555557FE005D003FE10AAFBE",
INIT_22 => X"1555FF082AA8B55F7AEA8BEF5551575FFA2FFD75FF550015400FFFBFFF450851",
INIT_23 => X"D57DF45A280154BA5555401EFFFD5421EFA2FFFFF555D0000145082E955FF085",
INIT_24 => X"051555FF0804155FFF7842AA100000020BAAA801541055042ABEFFFFBD5410AA",
INIT_25 => X"000000000000000000000000000000000000005568AAAAAD142145FF80155EF0",
INIT_26 => X"F145B42038555F401D71C0A2DBC7EB80000280824ADBD7490E28BEF080000000",
INIT_27 => X"82FFDB5243800002FBD7EBFBD24101C00175EFB6802DBC7BE8A155EFE3FBC71F",
INIT_28 => X"E1041003DE10BEF5EDAAAAAD547038EBD57DF7DA2AEB8FC7005F6AA381C0A2DA",
INIT_29 => X"5400E3F1FFF7D085B420381C5B6AA82147FF8FEF410E001FF000E17555555B7A",
INIT_2A => X"0017D142E905EF1451525C7082AADB45F7AEA8BEF555F575FFBEF5D05EF550E1",
INIT_2B => X"02FBEFEBFBD2410AADF78F45B68010482415B471C7E3DF451EFBEFBFAF454900",
INIT_2C => X"D145145FF84155D7085B555C71404105C7F7842FA381C0A00082AA8A10410410",
INIT_2D => X"02AA8BEF000000000000000000000000000000000000000000000005B68ABAB6",
INIT_2E => X"FFAE955EFAAFBD55EF557BC20AA5D7BC01555D2EBFF55A284000AA08003FF550",
INIT_2F => X"5007BE8AAA5D2EBDE00FFFFC00AA08003FF55A2FBC00105D04175FFF7803DF45",
INIT_30 => X"FF082A97555557FE8A0000043FE00F7D17FEBAA2D5574BAAAD17DFEFA2AEAAB5",
INIT_31 => X"5FFF7D5401EF5D2E97410AAD17DFEF007FC20AA5D7BE8A005D7FEABFF002E821",
INIT_32 => X"55EFF7FBE8B550004001FF5D2A801EF5D5142145082EBFF55F7AAAABEF5D7FD7",
INIT_33 => X"82010A2AA8000008043FFFFA2FBC2010A2FBEAB45F78402010007BD5545AAFFD",
INIT_34 => X"000000007BEAAAAFFD555545FF8015555007FD5545550400145FF843DEAA552A",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000007FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(1),               -- Port A write enable input
DIA(0)   => data_write_a(12),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(12),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(1),               -- Port B write enable input
DIB(0)   => data_write_b(12),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(12),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_13_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10110A0441812402840402822007818000E00700000000330A3000000008042",
INIT_01 => X"A1400986B830E84D182260000C1042484001000008220008A20019080A510200",
INIT_02 => X"10A108600C9141100000C6180CA85035010E4880010431004908135980122D60",
INIT_03 => X"0013881507460886C190832175809C02030400002020124C441A108468424842",
INIT_04 => X"203080680204A0113801D600864E0C96C12000008244244052200201801802C0",
INIT_05 => X"030004849601110204950409C0208C2084E0009C0000100120A00C9918002098",
INIT_06 => X"10000882804544921681428591908000AF28A8002BC00D020003896020658FC4",
INIT_07 => X"CA20400450050009100501501102E0042020448D0000023E10408144C800D800",
INIT_08 => X"1D2B00402B220104B53100200001020218A5104016CC1C616401910801010100",
INIT_09 => X"050800404D49A42EB08000000000000406481C8C408000A2D8088D1820200B00",
INIT_0A => X"0010000002004048AA08050401604462E9144002090740148441200484000500",
INIT_0B => X"000A112100000000010000000001000000000000001000000000000000800000",
INIT_0C => X"509528954404144C200425010040000001B020081094040072005C0030864208",
INIT_0D => X"1C10B3831034081200000000000430003000206822F20CA8826AC2A14250A128",
INIT_0E => X"1C10B383110218CB0E54C2EA404A4F03D404A41AA5B7344C10B383081BA4B734",
INIT_0F => X"8001CE3E20A5B284ED1132909C72885A2B2C381BA4B7344C10B383081AA5B734",
INIT_10 => X"AC3CC0C0B8182597A801610218CB0C3548B3A008E730A01AB113A5524E6ACA67",
INIT_11 => X"A151EC5952E44128CA194517354C180A3C066430202021252991C22C99731014",
INIT_12 => X"1804C8A0ADA2E6A983014780CA28B2A5C8825194332B018A444AEA2701288A15",
INIT_13 => X"02D09852745F80112C428562EE0353635232D50048A411C158BB0A7910142C77",
INIT_14 => X"4240480068001C9B9150A0000297046E4023F8BE8E3E1E0109472C3EB50158BB",
INIT_15 => X"A1284A1284A1284A1284A1284A12851A84284110406A26924302590806000110",
INIT_16 => X"1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284",
INIT_17 => X"284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A",
INIT_18 => X"7DDFE7EFBEFFE7D3EFBEFC48A0550000000000000000000A1284A1284A1284A1",
INIT_19 => X"D75D75D75D75D75D75D75D75D75D75D75D75D75D75D7EFBFBFBBAAAAAABEFDF7",
INIT_1A => X"5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5D75D75D75",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000FEFD7EBF5FAFD7EBF5FAFD7EBF",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"AA5D043FFFFAAAABDEAA557BFDE00FFD140155F7800000000000000000000000",
INIT_1F => X"400AAD540155A2D5421FF00042ABEFFF8400010082EAABFF55002ABEF08556AA",
INIT_20 => X"ABEFA280155EFFFFBC01EF08554000055043DEBAF7843FFFFF7AABDF55A2AA97",
INIT_21 => X"D5400005568A1055043DEBAAAFFE8B45557FD7410552EAAABAAA84155EFAA842",
INIT_22 => X"FE8ABAAA8428A00087BD7555FFD56AA10000028AAAFFD15541000002ABEFFFFB",
INIT_23 => X"803FE10AAFBE8AAAA2D540000F7D57DF55A2AABFFEF085557545FFD17DEBAA2F",
INIT_24 => X"0041554555557FE005D0000155557BEAABA5D2ABDF450851420AA5D7FD5555A2",
INIT_25 => X"000000000000000000000000000000000000005168AAA087BFFFFF5D04001FF0",
INIT_26 => X"7490E28BEF08516DA82410A3FFD7AAA4B8E824971F8E38E3DF45155EB8000000",
INIT_27 => X"D7EBA4BDF45AAAA90410BEDF45155A2DF401D71C0A2DBC7EB80000280824ADBD",
INIT_28 => X"A82B680175EFB6802DBC7BE8A155EFE3FBC71FF145B42038550E38E92EB803FF",
INIT_29 => X"243800002FBD7EBFBD24101C556FA38490A3FE92BEFFEAB45417FD24385D2AAF",
INIT_2A => X"5056DE3D17FE92BEF1EFA92AA8428A10007FD557DFFDF6AA381C0A2DA82FFDB5",
INIT_2B => X"B400925D7FD557DA2803DE10BEF5EDAAAAAD547038EBD57DF7DA2AEB8FC70051",
INIT_2C => X"7FF8FEF410E001FF000E17555555B7AE10410E00155497FEFABA4120B8F55085",
INIT_2D => X"2FBD7545AA8000000000000000000000000000000000000000000005B6AA8214",
INIT_2E => X"A284000AA08003FF55002AA8BEF00517FE00082EBDF45AA8428A10085568ABAA",
INIT_2F => X"A5D2EA8A00A2803DF45AA843DF55AAAE82000F7FBD5545AAFBC01555D2EBFF55",
INIT_30 => X"55087FC00BA552ABFE10F784175FFF7803DF45FFAE955EFAAFBD55EF557BC20A",
INIT_31 => X"AAA5D2EBDE00FFFFC00AA08003FF55A2FBC00105D517FEAA082EBFE10F7FFE8B",
INIT_32 => X"DFEFA2AEAAB550051401FFA2D57FE10F7D57DE00AA842AA00007FD75FFF7FBE8",
INIT_33 => X"FDEAA08042AB45087FC0010557FD55FFAA843FE00F7D17FEBAA2D5574BAAAD17",
INIT_34 => X"000000007BE8A005D7FEABFF002E821FF082A97555557FE8A00002E82155007B",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000067FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(1),               -- Port A write enable input
DIA(0)   => data_write_a(13),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(13),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(1),               -- Port B write enable input
DIB(0)   => data_write_b(13),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(13),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_14_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10020A000180000284008280000281800000030000000033022000000580002",
INIT_01 => X"A14009821830284D186860000C30C24840000000084000084200090008510200",
INIT_02 => X"102100600C9001100000061020A8503401044880010400204908012018122F64",
INIT_03 => X"00008015074608840190800010008002030400002074F401209A108448404842",
INIT_04 => X"000080400004A00100004000840E000201000000024024401200020180180080",
INIT_05 => X"0A000484800111020495040800208C2084000080000010010020049818002008",
INIT_06 => X"1000088020450402B6A1420511C080008468A80008000D0200018B202067AF10",
INIT_07 => X"422000044005000910040110510260040024400C800000BE3850A144C924080E",
INIT_08 => X"000B004028020104111100200001020210A51040008004616001910801010000",
INIT_09 => X"000800004D492408208000000000000406401C0C40800022C8088DB420200900",
INIT_0A => X"0010000002004048000005040160042229140002090200000401000484000400",
INIT_0B => X"0000110100000000010000100000000000000100000000000000100000000000",
INIT_0C => X"409120940404104C2000210100400000011020080084040040005C0010820208",
INIT_0D => X"E0E0A0000190081200000000000000003000000000100C088020028102408120",
INIT_0E => X"E0E0A0000B02740421A0E5D1A024002050805210040000B0E0A0000210040000",
INIT_0F => X"E01200860008920106460D4501CB000111300210008000B0E0A0000210008000",
INIT_10 => X"0ABBC00905C33C6000400F02740412C0715C40110080A4006110510C14D18178",
INIT_11 => X"20000041DB011CC000090012565306500002411420220080220C0093C3892324",
INIT_12 => X"5809240C09024A4AE0CA00004800839682398000120800658992F3C700C30181",
INIT_13 => X"002B46867DBC002A830280000800F7B7A0B1E240240A8340000200067EAA8CB6",
INIT_14 => X"42004005800004801150A00341244000845C7DB0D0200900422ACA4B28000002",
INIT_15 => X"8120481204812048120481204812051A04204110002A26924302590802000000",
INIT_16 => X"1204812048120481204812048120481204812048120481204812048120481204",
INIT_17 => X"2048120481204812048120481204812048120481204812048120481204812048",
INIT_18 => X"69CB91FE1EF7D3ABEFBECA080050000000000000000000081204812048120481",
INIT_19 => X"F3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF7EFBBBBBF9E79E7BEAAF3",
INIT_1A => X"CFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCF3CF3CF3C",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FF007F3F9FCFE7F3F9FCFE7F3F9F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"45AAD157400007BEAAAAAAAE955555D5568A105D000000000000000000000000",
INIT_1F => X"0AAF784020AAF7D56AAAA5D043FFFFAAAABDEAA557BFDE00FFD140155F7D17DF",
INIT_20 => X"ABEFFF8400010082EAABFF55002ABEF085155400FFD1420100055574AAA2AA80",
INIT_21 => X"40155A28028B550051574005D7FFFE105D7BD7545A284020BA0055421FF00042",
INIT_22 => X"1421FF5D7FFDEBA085168B45FF843DEBAF7843FFFFF7AABDF55A2AA97400AAD5",
INIT_23 => X"04155EFAA842ABEFA280155EFFFFBC01EF08554000055002AB455D5142010085",
INIT_24 => X"57FD7410552EAAABAAA8017400AAD140000002EBFFEFA2AAA8BEFF780021FF55",
INIT_25 => X"000000000000000000000000000000000000005568A1055043DEBAAAFFE8B455",
INIT_26 => X"8E3DF45155EBD17FF6DAADB504001C71EDA82AAA0955455D556DA00490000000",
INIT_27 => X"101C55554AAAAA480082FF84000BAEBD16DA82410A3FFD7AAA4B8E824971F8E3",
INIT_28 => X"092085F401D71C0A2DBC7EB80000280824ADBD7490E28BEF085157428FFDB420",
INIT_29 => X"DF45AAAA90410BEDF45155A28E2AB7D0051504005D71F8E004975D556DB68405",
INIT_2A => X"28B6D5D51420101C5B401EF417BFAEAA08516AB45E38E38E92EB803FFD7EBA4B",
INIT_2B => X"EAFBC7EB80071FF5500175EFB6802DBC7BE8A155EFE3FBC71FF145B420385500",
INIT_2C => X"0A3FE92BEFFEAB45417FD24385D2AAFA82B68015400AADB40000082EBFFC7A2A",
INIT_2D => X"5557FE1000000000000000000000000000000000000000000000000556FA3849",
INIT_2E => X"AA8428A10085568ABAA2FBD7545AAD17DFFFAAFFC200055557DE00A280155455",
INIT_2F => X"F0051554AAFFFFC00105D55554BAA28400000F784020BAAAD17FE00082EBDF45",
INIT_30 => X"000051575FFF78415410087BC01555D2EBFF55A284000AA08003FF55002AA8BE",
INIT_31 => X"A00A2803DF45AA843DF55AAAE82000F7FBD5545AAAEAABFF0051400105D5568A",
INIT_32 => X"55EF557BC20AA5D042ABFF555142000557FC01EF007FEAABA00556AB55A2AEA8",
INIT_33 => X"C0010082EBDF55A2AABDF45A284175FF5D04175FFF7803DF45FFAE955EFAAFBD",
INIT_34 => X"00000000517FEAA082EBFE10F7FFE8B55087FC00BA552ABFE10F78415400A2FB",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000007FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(1),               -- Port A write enable input
DIA(0)   => data_write_a(14),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(14),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(1),               -- Port B write enable input
DIB(0)   => data_write_b(14),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(14),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_15_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000A000000000284000280000001800020030000000033022000000180002",
INIT_01 => X"A140098018300848180060000C00426040000000080000080200000000110200",
INIT_02 => X"1020004000801110000006100028503400040800010430004808000180120278",
INIT_03 => X"00008011064408840190800000228002A3000000000010000008108448000042",
INIT_04 => X"701280400004A991000000A28406000211000000220004941000000880000000",
INIT_05 => X"02000484800155020495000800218020C4002880005310000000040000000001",
INIT_06 => X"10000880004540000711224491C08000850A880008000D020001892020656300",
INIT_07 => X"8A04000016050009140501505100000420204008000000BE70408104C8000000",
INIT_08 => X"001F004028026104111002200000000200210040008004614001100801010000",
INIT_09 => X"000800000D09240000800000000000040600180840800022C8088C1020200000",
INIT_0A => X"0000000002004040000105000040042229140002080000000400000080000400",
INIT_0B => X"0000110100000000010000100001000010000000000000000000100000800008",
INIT_0C => X"0001008000000000000025000040000001300008009400006200580010000000",
INIT_0D => X"0000000002300012000000000004200030000000000008008020020000000000",
INIT_0E => X"0000000001000000400000000000000000000010108000000000000010108000",
INIT_0F => X"0000000000000200000900000000000000000010140000000000000010140000",
INIT_10 => X"0140000000000000000001000000400000000000000000000100008040000000",
INIT_11 => X"0000004000480000000000100004400000000030002000406000000000068409",
INIT_12 => X"8000000000020080080000000000802010000000000800000201000800000000",
INIT_13 => X"00000100000000000000000008000000184400A0000000000002000000441108",
INIT_14 => X"4000000000000000010620000004000000000242038B82800000000000000002",
INIT_15 => X"0000000000000000000000000000041800000110000024130202500802000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000080050000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"000804154AA5D00001EFF78428AAA007BC2145F7800000000000000000000000",
INIT_1F => X"0AA007FC2000F7D17DF45AAD157400007BEAAAAAAAE955555D5568A105D7FC00",
INIT_20 => X"FFFFAAAABDEAA557BFDE00FFD140155F7FBD74AAAAD17DF45F7D1421EF005540",
INIT_21 => X"020AAF7FFFDF45FF84000BA552ABDFEF08517DF55A2FBEAB555D556AAAA5D043",
INIT_22 => X"FEAB45F7843FF45082A801FF005155400FFD1420100055574AAA2AA800AAF784",
INIT_23 => X"D5421FF00042ABEFFF8400010082EAABFF55002ABEF087BE8ABA555168B55AAF",
INIT_24 => X"D7BD7545A284020BA007FFFE10A284000AA0055401550055574005D2E800AAA2",
INIT_25 => X"000000000000000000000000000000000000000028B550051574005D7FFFE105",
INIT_26 => X"55D556DA004971C7038140012482550E021C7EB8028A821C7BC516DFF8000000",
INIT_27 => X"45E3DF471C70851400BA0071C5028FFD17FF6DAADB504001C71EDA82AAA09554",
INIT_28 => X"B555D516DA82410A3FFD7AAA4B8E824971F8E38E3DF45155EBF1D5492BED17FF",
INIT_29 => X"54AAAAA480082FF84000BAEBF1FFF7DEB8000092552ABFFEF08517DF6DB6FBE8",
INIT_2A => X"EFA8241516DB55A2FFEAB6DEB843DF551C20801C71C5157428FFDB420101C555",
INIT_2B => X"550428412A85082BEDF401D71C0A2DBC7EB80000280824ADBD7490E28BEF087F",
INIT_2C => X"51504005D71F8E004975D556DB68405092087FF8E00BE8A02082005F47145085",
INIT_2D => X"57BD75EFF78000000000000000000000000000000000000000000000E2AB7D00",
INIT_2E => X"55557DE00A2801554555557FE100055554BA5504000105D2A80145AA842AA005",
INIT_2F => X"5AAD557410F7D57DF55AAFBD55450055420BA0055574BAF7D17DFFFAAFFC2000",
INIT_30 => X"FF08517FFFFF7FBEAB455D517FE00082EBDF45AA8428A10085568ABAA2FBD754",
INIT_31 => X"4AAFFFFC00105D55554BAA28400000F784020BAAAD57FFEFA28402010552ABDF",
INIT_32 => X"FF55002AA8BEF007FFDE1000557DF45AAFBE8BEFA2803FF45550400155555155",
INIT_33 => X"80000087BD55450855400BA002A95400F7FBC01555D2EBFF55A284000AA08003",
INIT_34 => X"000000002EAABFF0051400105D5568A000051575FFF78415410087FEAA10F7AE",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000060000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(1),               -- Port A write enable input
DIA(0)   => data_write_a(15),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(15),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(1),               -- Port B write enable input
DIB(0)   => data_write_b(15),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(15),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_16_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"DA22C618B1000482B688B186588884862A400438255FC38381441205BA803003",
INIT_01 => X"264AC80028404C211203A952A90341080B173340412000E1005D628000820484",
INIT_02 => X"400034C206C405000001A48202084004003008255040826EE008B440200E2042",
INIT_03 => X"2916704900606AC82B49CC56DF8CC1E50E4800202115005760010010000C0400",
INIT_04 => X"052DCA856DC7504B82BF6614C86D2B7F85AAD17F4B100000B88148C4804A428A",
INIT_05 => X"373CB02A00C0502F301180141A42A5720E0F43C17A8479580001AC20000000E2",
INIT_06 => X"303E2094282B85242C85001038D5710E8410D5959BC4800015001219D0550077",
INIT_07 => X"880100000159954501280B0080146F7112D949A0015018220540000382805001",
INIT_08 => X"30015452880C8D90409A05B2CB2CA400200209E5601044A24000000462A60018",
INIT_09 => X"452D54000C0907000330000000000096480050000685400005FC014743E0DC92",
INIT_0A => X"00014808A02004200E540480212000A448C0080024AEA00C9688000000000005",
INIT_0B => X"000D58460018F6D3D84400044000440004400044000440004400042000220002",
INIT_0C => X"0001004010A8812831605DA0000A054052E40000817680220040025699200002",
INIT_0D => X"AAADA0C343F1AC1B01040A002024895514554485D00000012400240000000000",
INIT_0E => X"AAADA0CC421CA003B694B68018FAAA708E2CB5320018CAC99BA0A3B9320018CA",
INIT_0F => X"B1443A1891E4A928C29020E6A8524CE7A3EE59320018CAC99BA0ACB9320018CA",
INIT_10 => X"04B2A5A40B1E6644AF0F021EA003AC24352AB2449A3FF2FA04E5E09B128834AD",
INIT_11 => X"60ED838E890B703C6260D8E3A21275714C902375B801324301AB0067622E5E54",
INIT_12 => X"064F70DBDB1C74424E91E1C194C71D1216F50A8C241815FEB6A9158863F638FB",
INIT_13 => X"45FDF9D364DBD9435A6D45C9E81BED555E4C15F11133D171727A2550EE2F1BA0",
INIT_14 => X"08150013F162119014204373517700ACCC59432A2B2D001F803471A9A960E572",
INIT_15 => X"000000000000000000000000000000880002054000229088542210206B2AB015",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"2A898D21B4C98389ED146C080000000000000000000000000000000000000000",
INIT_19 => X"A29A29A29A29A29A29A29A29A29A28A28A28A28A28A53CBF0F0D3CF3CF0AB1A2",
INIT_1A => X"8F47A3D1E8F4FA7D3E9F4FA7D3E9F4FA7D3E8F4FA3D3E8F4FA3D3E9A29A29A29",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000FA7D3E9F4FA7D1E8F47A3D1E",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFF7FBE8B45AAD568BFFFFAA975FF00003FE0055000000000000000000000000",
INIT_1F => X"0005D2A95410FFFFC00000804154AA5D00001EFF78428AAA007BC2145F7843FF",
INIT_20 => X"7400007BEAAAAAAAE955555D5568A105D2E974BAF7FBEAB45FFFFC00BAF78002",
INIT_21 => X"C2000F78000010552E800AA002E821FFA2AAAAA00000417555FFD17DF45AAD15",
INIT_22 => X"43FEBA5D55575FFF7AABFE00557BD74AAAAD17DF45F7D1421EF0055400AA007F",
INIT_23 => X"D56AAAA5D043FFFFAAAABDEAA557BFDE00FFD140155F7AABDF55F7AE820AA080",
INIT_24 => X"8517DF55A2FBEAB555D04154BAA2FBE8B55FFFFD55FF557FC2000FF8015410FF",
INIT_25 => X"000000000000000000000000000000000000007FFDF45FF84000BA552ABDFEF0",
INIT_26 => X"21C7BC516DFF8438FC7E3F1EAB55B6DF6DBFFF7AA955C71C043FE10490000000",
INIT_27 => X"55FFF1C70BAF78A000005D2097438FFF1C7038140012482550E021C7EB8028A8",
INIT_28 => X"57DEBD17FF6DAADB504001C71EDA82AAA0955455D556DA00492490492F7FBE8B",
INIT_29 => X"71C70851400BA0071C5028FF84020285D2085092002A801FFB6AAA8A10080E17",
INIT_2A => X"BAF6DE3AA8709208043FEBA555B555FFE3AABFE005D71D5492BED17FF45E3DF4",
INIT_2B => X"BC0028E38412428EBD16DA82410A3FFD7AAA4B8E824971F8E38E3DF45155EBA4",
INIT_2C => X"8000092552ABFFEF08517DF6DB6FBE8B555D04124BAB6FBE8B45E3FBD55D7557",
INIT_2D => X"5003DE000000000000000000000000000000000000000000000000071FFF7DEB",
INIT_2E => X"5D2A80145AA842AA00557BD75EFF78428B55AAD168B55F7FFFDFEFFFAA955555",
INIT_2F => X"0000000010F7FBEAB45FFD1554AAFFAE820105500154AAF7D5554BA550400010",
INIT_30 => X"EFF7AEA8A10002E955FFA2D17DFFFAAFFC200055557DE00A2801554555557FE1",
INIT_31 => X"410F7D57DF55AAFBD55450055420BA0055574BAF784000BA5D0017410082E801",
INIT_32 => X"8ABAA2FBD7545AA802ABEFA2AA9541000003DEBA557BD75EFA2AEBDE105D5557",
INIT_33 => X"EAB45AAFFD55555D7FC20AAA280000AAAAD17FE00082EBDF45AA8428A1008556",
INIT_34 => X"00000000557FFEFA28402010552ABDFFF08517FFFFF7FBEAB455D04020AAFFFB",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000020000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(2),               -- Port A write enable input
DIA(0)   => data_write_a(16),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(16),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(2),               -- Port B write enable input
DIB(0)   => data_write_b(16),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(16),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_17_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"5284CE4FB7BD2C8994A13392DBD02E14006B82AC7E800D44D3DD2FD5F9B961C0",
INIT_01 => X"F9BA301F7E03FC6793F2199B39FC233C11D93AE6F3BB92B32091DBC339B24542",
INIT_02 => X"1D5FC0C08F040404446965C0607FB8A217C400C33A908078551BD04222186338",
INIT_03 => X"A14124C28DFD960832C90446DF8400A5055C25295B695FF97E1B5AC757F06D6B",
INIT_04 => X"04A106866DA3D02A01FB660C08A4AB7F840EDB6F48100DFC8081081D78AC7402",
INIT_05 => X"51E072F0C0C58D9C125EBFC00A46CF0388054100F680E0CE0107B8D040DAFCDA",
INIT_06 => X"019A4D00786B048112C58B16307F15DE8408B233661C10BBA5DAAFA9DDA1194D",
INIT_07 => X"8E00001660700CE170284A00891C7C03D29DE26814515835902AC089A2801540",
INIT_08 => X"C009F3A1B0120A1C51DFF881861CBE0305A12A0321810217C01D34EDC98FFA1C",
INIT_09 => X"747E6610052CDEE97FF1F9F63E3EF790380078002CE976AB6BF769769E4D437D",
INIT_0A => X"00185C44B91BC1740B7605040BE0018CFC7429F326B9D045FF8000E9AB415606",
INIT_0B => X"3A28FC1AAF5CF6F3D3EF3D3EF3D3EF3D3EF3D3EF3D3EF3D3EF3D3EF9E9F79E9E",
INIT_0C => X"0000020012E9E10A31EB5FF9296A67F5B4FFBD2FAD7FE653C3FBFF33E10C001B",
INIT_0D => X"333EA16031F2BD47BDA2CA5D8164FCCFE833C5C3D00018006C68170000000000",
INIT_0E => X"333EA160391BEFF2C32FB695F919110D5ECE542A6FEEB2533EA160782A6FEEB2",
INIT_0F => X"D18C0D06638A207CFDE1F7DDAD76D5282400F82A6FEEB2533EA160782A6FEEB2",
INIT_10 => X"E6E43E59AFE4A59B57679D19EFF2C7573FAD5A86840354D1706FFFA3EF6E24B6",
INIT_11 => X"F7D7A0ABD6DAAAB96529382B74E4E1FE4ACA4D77FAAB77CE3AF3EE78F58DB737",
INIT_12 => X"2D1281017F056E9C9C3FC95949C157ADB55572CA52606DFED6CA55334C04C04F",
INIT_13 => X"59FDEB974F486905001FDF5FA0D719F9956EAA1A184045D5D7A870D2F5A5D752",
INIT_14 => X"60158015177F916A039EF41FDB34A91F432EA58949D5B5C85F97871876F7D7E8",
INIT_15 => X"000000000000000000000000000004DC200005E705B7B3D9FC22F00BE419FB55",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"06013DB9880A5D22E229F3030018000000000000000000000000000000000000",
INIT_19 => X"D35D74D35D74D34D35D74D35D74D34D34D34D34D34D0D30D0D303AEBAE886E40",
INIT_1A => X"51A8D46A351A0D068341A0D068341A0D068341A8D468341A8D46834D35D74D34",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000008D46A351A8D46A351A8D46A3",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFF7FBFDF55A28402000F7D56ABFF55000000000000000000000000",
INIT_1F => X"A00F7843FEBA55043FFFFF7FBE8B45AAD568BFFFFAA975FF00003FE0055043FF",
INIT_20 => X"54AA5D00001EFF78428AAA007BC2145F7D568B45000002010552EBDF45A28028",
INIT_21 => X"95410FFAE800105D2A95410002A95410AAAEBFF55AAFFC00BAF7FFC000008041",
INIT_22 => X"57DE00F7AE800AAAAAABDFEF5D2E974BAF7FBEAB45FFFFC00BAF780020005D2A",
INIT_23 => X"517DF45AAD157400007BEAAAAAAAE955555D5568A105D7FFFFEFA2D568BFFFFD",
INIT_24 => X"2AAAAA00000417555FF8028B55082A974105D003FF55F7802AAAAAAD168AAA5D",
INIT_25 => X"000000000000000000000000000000000000000000010552E800AA002E821FFA",
INIT_26 => X"71C043FE10490A3FFFFFFFFFDFEFE3F5FAF45AA8000038F7DB6FBD7490000000",
INIT_27 => X"384124BFF7DB68A28A38F7803DE82490438FC7E3F1EAB55B6DF6DBFFF7AA955C",
INIT_28 => X"0BAFFF1C7038140012482550E021C7EB8028A821C7BC516DFFDF68B551C0E050",
INIT_29 => X"70BAF78A000005D2097438FFAA85000492495428082E95400AAA0BDF7DB6F5C7",
INIT_2A => X"FAFFFB6D56FBFFEBDB78E38F7AA800BAB6AEBDFD75D2490492F7FBE8B55FFF1C",
INIT_2B => X"028AAAB6D16FA8249517FF6DAADB504001C71EDA82AAA0955455D556DA00497F",
INIT_2C => X"2085092002A801FFB6AAA8A10080E1757DEB8A2DB5514249243841003FF6DEB8",
INIT_2D => X"7FFFDF550000000000000000000000000000000000000000000000004020285D",
INIT_2E => X"F7FFFDFEFFFAA9555555003DE00002ABFFEFF7FBFDFFFAAD168B55AA80000BAF",
INIT_2F => X"FF7FBEAB45552E954BA08003DFFFFFAAA8AAAF7843FE10000428B55AAD168B55",
INIT_30 => X"10AA843FFFFF7D5554BAF7D5554BA5504000105D2A80145AA842AA00557BD75E",
INIT_31 => X"010F7FBEAB45FFD1554AAFFAE820105500154AAF7AE974000800154AA002E954",
INIT_32 => X"554555557FE10007FEABEFFFD57FFEFAAFFE8ABAFFAA820BAF7AEBFF55550000",
INIT_33 => X"020AA08003DFFFA28028AAAF7D17DE0000517DFFFAAFFC200055557DE00A2801",
INIT_34 => X"0000000004000BA5D0017410082E801EFF7AEA8A10002E955FFA2AABFF455500",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000067FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(2),               -- Port A write enable input
DIA(0)   => data_write_a(17),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(17),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(2),               -- Port B write enable input
DIB(0)   => data_write_b(17),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(17),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_18_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"69844019080000A21A611406840014122A641074155FC28A2024001001801003",
INIT_01 => X"01067920034004180005E9E3C90360C0041C0181002001602025800008440084",
INIT_02 => X"40AC3CAA22D605200000856E2481902400344A20F802C22054001000021E2379",
INIT_03 => X"A95308ECD3207AC81D91C4002004C08A06008080BA868007E58040102B0E0100",
INIT_04 => X"044CC183800CA00780808004C8DB841405A80A100B586200FAC24AE4805242CA",
INIT_05 => X"771C10000000000B1135883C08A115320E0401C0200038394230070A19000020",
INIT_06 => X"3001499C602A8A003E800A042D8132A00098408F79E3901218050018024110D6",
INIT_07 => X"5029401000C983E60004010030400353C05806800104004E0000042E52800E20",
INIT_08 => X"0000117088080990419005B0C309402030060860E01004A828408800440405E3",
INIT_09 => X"6B8186185C42900693A002004040001E1950850C848601008708114A2030B480",
INIT_0A => X"100180A8062026000DC425C0301311324AA237108857220BA089420440000030",
INIT_0B => X"C44703657083080C2800C2000C2000C2000C2000C2000C2000C2000610006100",
INIT_0C => X"C1B0609C05013065CC042004040808084001E000108010230400800FD9B286C4",
INIT_0D => X"CCC15F9CBA45505640000A402019003F140FC2060014250B9080008306C18360",
INIT_0E => X"CCC15F9FB1962FCB69E08AAAEAEBCDDF7C728582081483ACC15F9C3982081483",
INIT_0F => X"EBF1CFFF7670ACC3811A28AB57523CDFEBFBF982081483ACC15F9F3982081483",
INIT_10 => X"C9002BF05800D875E63CC9962FCB52CAA02FE3F8E7F5E3AC3620805298B15A3F",
INIT_11 => X"F1B72A8A800B7546DB9F1CA320037F01BD67DC4041D4CF03138DD865103EFEEA",
INIT_12 => X"81CCFAFDBF9464006FD037AEFAE5150016EA8DB7BFE25208E8F46A228BF8A757",
INIT_13 => X"641256EC844B8AF92FD7CEDC24A9E181A8A29509EAAE7FD3B749471C48F8A459",
INIT_14 => X"0297D086E00036D2440E0880AAD62BEFF5778802A3AF8E8FB0440CE78773B709",
INIT_15 => X"8360D8360D8360D8360D8360D83609220D20D00000080C0601400B402307E480",
INIT_16 => X"360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D",
INIT_17 => X"60D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8",
INIT_18 => X"D9D701DC2E784601EFBE2C00000000000000000000000008360D8360D8360D83",
INIT_19 => X"5155555545145145155555545145145145145145145220B22A0B820820965177",
INIT_1A => X"44A25128944A25128944A25128944A25128944AA552A954A2512895554514514",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000025128944A25128944A251289",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFEFF7AE954BA5D04174AA00000000000000000000000000",
INIT_1F => X"145AA801741000043FFFFFFFFFFFFFF7FBFDF55A28402000F7D56ABFF55043FF",
INIT_20 => X"8B45AAD568BFFFFAA975FF00003FE0055043FFFFFFFFFDFEFA2D56AB45AA8400",
INIT_21 => X"3FEBA55557FFEFA2D168B55AAFBFFFFFFF80021EF0855421EF00043FFFFF7FBE",
INIT_22 => X"A82155F7AEBFEBAFFD56AA00A2D568B45000002010552EBDF45A28028A00F784",
INIT_23 => X"FFC00000804154AA5D00001EFF78428AAA007BC2145F7D5400000004020AA5D2",
INIT_24 => X"AAEBFF55AAFFC00BAF7AE80010082E954BA0004174AAAA8428B45082ABFEBAA2",
INIT_25 => X"000000000000000000000000000000000000002E800105D2A95410002A95410A",
INIT_26 => X"8F7DB6FBD7490E3FFFFFFFFFFFFFFFFBFDFEFFFAE954AA550415492140000000",
INIT_27 => X"D7AAD16FB6DBE8E00155BE8015410140A3FFFFFFFFFDFEFE3F5FAF45AA800003",
INIT_28 => X"1C7140438FC7E3F1EAB55B6DF6DBFFF7AA955C71C043FE1049043FFEFE3F1F8F",
INIT_29 => X"FF7DB68A28A38F7803DE82495B78FC7AAD56FB6DBEF1FAFD7E384001EF145B47",
INIT_2A => X"420381C0A02082492A85155E3A4BDE92FFD56FA28B6DF68B551C0E050384124B",
INIT_2B => X"E28B7D1420BDEAAA2F1C7038140012482550E021C7EB8028A821C7BC516DFFD1",
INIT_2C => X"2495428082E95400AAA0BDF7DB6F5C70BAFFAE870280024904BA1400174AABE8",
INIT_2D => X"50415410550000000000000000000000000000000000000000000002A8500049",
INIT_2E => X"AAD168B55AA80000BAF7FFFDF55002ABFFFFFFFFFFFEFF7FBFDFFFF7AA974BA5",
INIT_2F => X"000043DFEFA2D56AB45AAD57DFEFF7AA82155F78015400552ABFFEFF7FBFDFFF",
INIT_30 => X"55A280021EF557FD7555550428B55AAD168B55F7FFFDFEFFFAA9555555003DE0",
INIT_31 => X"B45552E954BA08003DFFFFFAAA8AAAF7843FE10007FEAB55A2D17FFEFFFD568B",
INIT_32 => X"AA00557BD75EFF7D1400AA5D2A82000002A95545A2843FE00F7D17FEAAF7FBEA",
INIT_33 => X"020AA5D04154BAF7AEA8BEF55003DEAAA2D5554BA5504000105D2A80145AA842",
INIT_34 => X"000000002E974000800154AA002E95410AA843FFFFF7D5554BAF7AE974BA0004",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000020000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(2),               -- Port A write enable input
DIA(0)   => data_write_a(18),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(18),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(2),               -- Port B write enable input
DIB(0)   => data_write_b(18),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(18),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_19_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"042200000000000041088001001AA00000000000000000000000500802000003",
INIT_01 => X"074018000024000000000404000000000A22000800000800004A200000000001",
INIT_02 => X"0000048002C405000000000006A84000000000200893C246A20000000020031A",
INIT_03 => X"020A9639044012C80001C4000004C08006000000001025000000000000000000",
INIT_04 => X"0400C0800000000380800004C8000000058800000B1000009880480480024200",
INIT_05 => X"420410000000000B10804004080001320E0401C0200038080000000000000000",
INIT_06 => X"2002409006F00A8428050A000280493104004500480090080A01120220140020",
INIT_07 => X"0000000000418026090240923240002190400000000000C0054A912054004021",
INIT_08 => X"0000115080000990000000B0C308000000000860200160000000000038380000",
INIT_09 => X"8000F80001012590001000000000001618000000020280008180810200000000",
INIT_0A => X"0000000000000000000000000000000100008000110000000000000000000017",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000840007600000000000000000800259000000",
INIT_0D => X"0008A0034078104B41A41000000000031400C002000000000000000000000000",
INIT_0E => X"0008A0004263C0343EDD414004042228DC0D385598035D0008A003B05598035D",
INIT_0F => X"040231068187C39F5A4F985C008902041124505598035D0008A000B05598035D",
INIT_10 => X"1BFBD406451B02000E033263C0343CB740500401180DE053A98F6ECC739D8140",
INIT_11 => X"420851546B2400000040D8549B5800000010227848D4303807FC8CC5508AEAED",
INIT_12 => X"52210402120A936B0000000004C2A8D6480000000018A700FCF980CC300318A2",
INIT_13 => X"B1427ED430B41402D025082359700181C21140E40511802208D6B30C48F8A8A4",
INIT_14 => X"9C000018440021011821B35254E99AF9E9410006362A2B6424287B08286208D6",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000023006000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"7747E18E0218CC18E88324000000000000000000000000000000000000000000",
INIT_19 => X"34C30C30C30C30D34C30C30C30C30C30C30C30C30C3504118982A69A6980E411",
INIT_1A => X"C26130984C26130984C26130984C261309A4D26130984C26130984C30C30C30D",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000130984C26130984C26130984",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAA954BA5500020BA5D000000000000000000000000",
INIT_1F => X"4BA5D517FFFF08043FFFFFFFFFFFFFFFFFFFFEFF7AE954BA5D04174AA007BFFF",
INIT_20 => X"FFFFF7FBFDF55A28402000F7D56ABFF557BFFFFFFFFFFFFFFFFFBFDFEFFFAA97",
INIT_21 => X"17410007BFFFFFFFFFFFFEFF7D16AB45AA8002000F7D5575455D043FFFFFFFFF",
INIT_22 => X"568B55F7AE955FFAA840201008043FFFFFFFFFDFEFA2D56AB45AA8400145AA80",
INIT_23 => X"043FFFFF7FBE8B45AAD568BFFFFAA975FF00003FE00557BFFFFFFFFBFDF45AAD",
INIT_24 => X"F80021EF0855421EF002ABFFEFF7D168B55AAD17FFEFF7AE975FF00557FFFF5D",
INIT_25 => X"00000000000000000000000000000000000000557FFEFA2D168B55AAFBFFFFFF",
INIT_26 => X"A5504154921471FFFFFFFFFFFFFFFFFFFFFFFF7AA954BA550000082550000000",
INIT_27 => X"EFF7FBFAFD7E3A4954BA555B7AFC7080E3FFFFFFFFFFFFFFFFBFDFEFFFAE954A",
INIT_28 => X"545550A3FFFFFFFFFDFEFE3F5FAF45AA8000038F7DB6FBD74975FFFFFFFFFFFF",
INIT_29 => X"FB6DBE8E00155BE8015410147FFFFFFF7FBF8FC7EBD568B55A28000000FFDF52",
INIT_2A => X"FDFC7E3F1FAF55A2DB6FB7DF7AE955C7BE800000008043FFEFE3F1F8FD7AAD16",
INIT_2B => X"0955FF145B7AFC7410438FC7E3F1EAB55B6DF6DBFFF7AA955C71C043FE10497B",
INIT_2C => X"D56FB6DBEF1FAFD7E384001EF145B471C71424B8FC7E3D56AB6DB6DF7AFC7EBA",
INIT_2D => X"50002000550000000000000000000000000000000000000000000005B78FC7AA",
INIT_2E => X"F7FBFDFFFF7AA974BA55041541055517FFFFFFFFFFFFFFFFFFFFEFF7AA974AA5",
INIT_2F => X"500517FFFFFFFBFDFEFFFFFEAB45AA80154AA557BEAB45002ABFFFFFFFFFFFEF",
INIT_30 => X"55A28002000F7FFC2155552ABFFEFF7FBFDFFFAAD168B55AA80000BAF7FFFDF5",
INIT_31 => X"FEFA2D56AB45AAD57DFEFF7AA82155F78015400557BFDFEFF7FBEAB55A2D56AB",
INIT_32 => X"555555003DE00007FFDF45AAD568B45AAFBFFFFFFFAA95545F7840201000043D",
INIT_33 => X"6ABFFFFFBEAB45A280155EF557FE8B55000428B55AAD168B55F7FFFDFEFFFAA9",
INIT_34 => X"000000007FEAB55A2D17FFEFFFD568B55A280021EF557FD755555042AB55AAD1",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000040000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(2),               -- Port A write enable input
DIA(0)   => data_write_a(19),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(19),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(2),               -- Port B write enable input
DIB(0)   => data_write_b(19),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(19),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_20_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000003",
INIT_01 => X"A65FF80000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000048002CC070000000000000000000000002FF86100200000000220002362",
INIT_03 => X"00000000000203D80025DC18004DC3D01E000000000000000000000000000000",
INIT_04 => X"07E5DF808071026F87C4191DD8005080679800000F300002998058068002C000",
INIT_05 => X"C205F23A2100557F70000004390021F61E1E87C3FD0CFBF80880072042000044",
INIT_06 => X"1209244C2000100006800000020010000008407FC800B0000000100600040000",
INIT_07 => X"8802000009FFBFE51886018002040020000800000554003E0000000002800000",
INIT_08 => X"30801F5780259FB0000000F7DF78020004011FEFE00000000020031502000083",
INIT_09 => X"00000000001000000000000000000056F8000001000000040000040141800802",
INIT_0A => X"0000000000000008000800000000000000000000000000000010010014800000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"00010240001721214E000004000000080000008000001000040080FFDB000000",
INIT_0D => X"0000000F3008001E00000000001803FF14FFC006000000008010200000000000",
INIT_0E => X"0000000F3040200000020000000026A70C0008020000200000000F3002000020",
INIT_0F => X"000030B86000400080000200000000004A58F0020000200000000F3002000020",
INIT_10 => X"0000000002183E61E6000040200001000000000019B140000800800000020000",
INIT_11 => X"C00010080000000000525801000000000014AC08000000508001030A0A400100",
INIT_12 => X"000002BC360020000000000292C0100000000000A56000090100000000001F86",
INIT_13 => X"8010000000000000574500001001060600000000001716800000803102020000",
INIT_14 => X"00000000000040040040002000080506049CDF70C08040100000706707600000",
INIT_15 => X"00000000000000000000000000802040200200604040000000000024FB7FE008",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"060070400020112240209A408004000000000000000000000000000000000000",
INIT_19 => X"65965965965965965965965965965861861861861860D30424343CF3CF340E00",
INIT_1A => X"90C86432190C86432190C86432190C86432190C86432190C8643219659659659",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000086432190C86432190C864321",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974AA55040201008000000000000000000000000",
INIT_1F => X"4AA550002000007BFFFFFFFFFFFFFFFFFFFFFFFFFAA954BA5500020BA5D7FFFF",
INIT_20 => X"FFFFFFFFFFFEFF7AE954BA5D04174AA00003FFFFFFFFFFFFFFFFFFFFFFF7AA97",
INIT_21 => X"7FFFF087FFFFFFFFFFFFFFFFFFFFDFEFFFAE974AA5D003FE005D043FFFFFFFFF",
INIT_22 => X"BFDFFFAA84000105D556AB55557BFFFFFFFFFFFFFFFFFBFDFEFFFAA974BA5D51",
INIT_23 => X"043FFFFFFFFFFFFFF7FBFDF55A28402000F7D56ABFF55003FFFFFFFFFFFFFF7F",
INIT_24 => X"A8002000F7D5575455D2EBFFFFFFFFFFFEFF7FBEAB55A28000010F7D16ABEF08",
INIT_25 => X"000000000000000000000000000000000000007BFFFFFFFFFFFFEFF7D16AB45A",
INIT_26 => X"A550000082557FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550400028000000000",
INIT_27 => X"FFFFFFFDFEFF7AE974BA5500050380071FFFFFFFFFFFFFFFFFFFFFFFF7AA954B",
INIT_28 => X"E285D0E3FFFFFFFFFFFFFFFFBFDFEFFFAE954AA55041549214043FFFFFFFFFFF",
INIT_29 => X"AFD7E3A4954BA555B7AFC70871FFFFFFFFFFFFFFF7FBFDFFFFFAA974BA550038",
INIT_2A => X"3FFFFFFFFFDFEFF7F1FAFC7A28002028555F6FB7D5D75FFFFFFFFFFFFEFF7FBF",
INIT_2B => X"402010FFDB6ABEF140A3FFFFFFFFFDFEFE3F5FAF45AA8000038F7DB6FBD7490E",
INIT_2C => X"FBF8FC7EBD568B55A28000000FFDF525455524BFFFFFFFBFDFC7E3F5E8B45A28",
INIT_2D => X"504000BA080000000000000000000000000000000000000000000007FFFFFFF7",
INIT_2E => X"FFFFFFFEFF7AA974AA550002000557FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5",
INIT_2F => X"055043FFFFFFFFFFFFFF7FBFDFEFFFAE954BA5500174AA08517FFFFFFFFFFFFF",
INIT_30 => X"EFF7AE974AA550028AAA5D2ABFFFFFFFFFFFEFF7FBFDFFFF7AA974BA55041541",
INIT_31 => X"FFFFFFBFDFEFFFFFEAB45AA80154AA557BEAB4500557FFFFFFFFFDFEFF7FFFFF",
INIT_32 => X"00BAF7FFFDF55002EBFFFFF7FBFDFEFFFD568B55A284020BA557FFFFFF5D517F",
INIT_33 => X"FFF55A2D16AB45AA8402000F7FBEABEF5D2ABFFEFF7FBFDFFFAAD168B55AA800",
INIT_34 => X"000000007BFDFEFF7FBEAB55A2D56AB55A28002000F7FFC215555043DFEFF7FB",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000007FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(2),               -- Port A write enable input
DIA(0)   => data_write_a(20),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(20),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(2),               -- Port B write enable input
DIB(0)   => data_write_b(20),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(20),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_21_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"4A302428B824900A128C090A5C1800261500213C005FE812D10420054085A202",
INIT_01 => X"081FFE3440B609703B0427F801A40B8115BC4F655300340288A40D30040E4DD8",
INIT_02 => X"04CA478082CC1740002019824E0203100640303FF8C0B31061096E21A1840814",
INIT_03 => X"230CA7A4810083F80095DE00102DC3823EA821094EC68248923200013290C800",
INIT_04 => X"07CFFFC04904AA7F8780409DF84A0202879800000F3000029980780EA2C3C002",
INIT_05 => X"DE87F0280000407FF900D914382091FE1E1C0FC3E01EFFF8000480200008D062",
INIT_06 => X"010E2182002BC107A03448808F0D7C002822987FC830F40134CC74D002016612",
INIT_07 => X"0401000011FBFFE00520000200422033025C4209104500000012004C004D8C0B",
INIT_08 => X"00EF1F5FA0041FF080AC70FFDF78220010841EFFE7116E144071268DFD3E4C24",
INIT_09 => X"FC8BFE18008083B4443151462A28C6DFF80010002605302248088950484550A3",
INIT_0A => X"10018C241102068006C620C03882019480E631A0855E924E2598038938404037",
INIT_0B => X"A641165448C80C103648A3648A3648A3648A3648A3648A3648A366451B2451B2",
INIT_0C => X"011100841200D001000624000100C002804A08221890004806A310FFDF000454",
INIT_0D => X"5004D8158809C86065941840B1014FFF56FFC0281280080180B2948004400220",
INIT_0E => X"5004D815810D42E04A08A80098C02450025360694101816002D41A4068C10181",
INIT_0F => X"134160C8125B0B271802242880A04482418A0068C101816002D41A4069410181",
INIT_10 => X"10080E05C0B06AA8B12CFD0D42E0441A300012682960828F05C96A001B029010",
INIT_11 => X"00010362A8A20826A88660D86B202049F115100920C54E8EA256ECF078BA081C",
INIT_12 => X"064802C0081B0D64040936443306C55144104F30A8801406D002900062803201",
INIT_13 => X"4581BA0038005A706680012280506A8010602011819E290048A2118EC8140C08",
INIT_14 => X"CC158092C044600466208CC5091011C322A4C40A0300600C0A80509F41800880",
INIT_15 => X"80200802008020080200802008020412002001000000381C02004000FBFFF80D",
INIT_16 => X"0200802008020080200802008020080200802008020080200802008020080200",
INIT_17 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_18 => X"FDDFEFFFBEFFE7C7BFBEFC000000000000000000000000080200802008020080",
INIT_19 => X"F7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7FFBFBFFF9E79E7FFFDF3",
INIT_1A => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFDFEFF7FBFDFEFF7FBFDF7DF7DF7D",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00001FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D000200008000000000000000000000000",
INIT_1F => X"4AA5D00020AA5D7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550402010087FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAA954BA5500020BA5D7FFFFFFFFFFFFFFFFFFFFFFFFFFAE95",
INIT_21 => X"0200000003FFFFFFFFFFFFFFFFFFFFFFF7AA974BA5D0402000557BFFFFFFFFFF",
INIT_22 => X"FFFFEFF7AE974BA5D00174BA00003FFFFFFFFFFFFFFFFFFFFFFF7AA974AA5500",
INIT_23 => X"043FFFFFFFFFFFFFFFFFFFFEFF7AE954BA5D04174AA00003FFFFFFFFFFFFFFFF",
INIT_24 => X"FAE974AA5D003FE005D2EBFFFFFFFFFFFFFFFFFFDFEFF7AE954AA5500174BA5D",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFDFEFF",
INIT_26 => X"A550400028007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0000010000000000",
INIT_27 => X"FFFFFFFFFFFFFAA954BA5D00000BA557FFFFFFFFFFFFFFFFFFFFFFFFFFAE974A",
INIT_28 => X"0005571FFFFFFFFFFFFFFFFFFFFFFFF7AA954BA550000082557BFFFFFFFFFFFF",
INIT_29 => X"DFEFF7AE974BA55000503800003FFFFFFFFFFFFFFFFFFFFEFF7AA974AA5D0405",
INIT_2A => X"3FFFFFFFFFFFFFFFFFFDFEFF7AE954BA5D00154AA00043FFFFFFFFFFFFFFFFFF",
INIT_2B => X"A974BA5D00104925D0E3FFFFFFFFFFFFFFFFBFDFEFFFAE954AA550415492140E",
INIT_2C => X"FFFFFFFF7FBFDFFFFFAA974BA550038E285D2ABFFFFFFFFFFFFFFFFBFDFEFFFA",
INIT_2D => X"D00000100000000000000000000000000000000000000000000000071FFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE954AA5504000BA087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0557BFFFFFFFFFFFFFFFFFFFFFFFF7AA954BA5D00000BA5D7FFFFFFFFFFFFFFF",
INIT_30 => X"EFF7AE954AA5D041740055517FFFFFFFFFFFFFFFFFFFFEFF7AA974AA55000200",
INIT_31 => X"FFFFFFFFFFFFF7FBFDFEFFFAE954BA5500174AA08043FFFFFFFFFFFFFFFFBFDF",
INIT_32 => X"74BA550415410552ABFFFFFFFFFFFFFF7FBFDFFFFFAA974AA5D00174BA08043F",
INIT_33 => X"FDFEFF7FBFFFFFF7AE954BA5D0000010552ABFFFFFFFFFFFEFF7FBFDFFFF7AA9",
INIT_34 => X"00000000557FFFFFFFFFDFEFF7FFFFFEFF7AE974AA550028AAA5D2EBFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(2),               -- Port A write enable input
DIA(0)   => data_write_a(21),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(21),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(2),               -- Port B write enable input
DIB(0)   => data_write_b(21),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(21),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_22_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"5290F4CDE914905A14A43D33F488243E17122300F55FEB189B343A1140548380",
INIT_01 => X"A94007B259F6A975386262000C344BA9573C6FF57B18A5FB0ABFCD3C2C5F4F0C",
INIT_02 => X"D56B4302AC01005111011BD506AA5205274056900596A539584E2E6DFE4B2418",
INIT_03 => X"9AC0FCBD854688207C90007A1000047A00E588632CA213C8903AD6B55AD0EB5A",
INIT_04 => X"30002047A6FCA110086C402022F2124A8022492580040440002021C922D9109B",
INIT_05 => X"14A206B6838151008D95DD1847811C08002380041F1104002205AC4140DAD060",
INIT_06 => X"1727FF2EB9EF113A10BD32F44289D1F840C1710010344DB9A808FDFF3DE03130",
INIT_07 => X"050700154A00401D00495A06A8D464C5F6B54AA8551040818F4C997AC80CBE05",
INIT_08 => X"0141008801018040E48D50080002B00A0C00801014541E9504703680017F6CB4",
INIT_09 => X"02680000010937986481514E2A29CE010708C0804C6A033F7FCFF9426A41F1AB",
INIT_0A => X"00500001840000C80B410014088040F4A944B1AA313C004554002381B8000500",
INIT_0B => X"A004D1594832824A070AA070AA070AA070AA070AA070AA070AA0725503855038",
INIT_0C => X"501428054278142151262CA50343854E506A2C6898B2950AA6A35B0004284058",
INIT_0D => X"90078E1F840A2B0114020104022460002200050F60E220A06880D2A14050A028",
INIT_0E => X"90078E1F891C239F8908003099C1ACF06273612B3482C0C0078E1F412B1582C0",
INIT_0F => X"1BA1B0FD16770236A4091621C08055C2C0DB012B1582C0C0078E1F412B3482C0",
INIT_10 => X"00101F09C030AB28B03C111C239F870828041BA859F213AFC14AA38043006018",
INIT_11 => X"10E8822A984B0025B0DE6089462660095337B08AA600CA88B143AB11880C2806",
INIT_12 => X"055412D4481128C4CC012A66F304553096004B61BD8068B92400D0004E303689",
INIT_13 => X"589C48082C006A9057CA4385809520F07830001AC2173B00E162563454C40804",
INIT_14 => X"00460848952220592745AC11A544B1BF006850840180A00E1C81900C4190E160",
INIT_15 => X"22088220882208822088220882208CD888088D940D2A3A9D5002001300800C8C",
INIT_16 => X"0080200882208822088220882208822088220882208822088220882208822088",
INIT_17 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_18 => X"FBDFD1FE3EFBD7BBEFBEFA0A245120000000007FFFFFFFF20080200802008020",
INIT_19 => X"F3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF7FFBFAFBBBEFBEFBEFBF7",
INIT_1A => X"CFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCF3CF3CF3C",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000007F3F9FCFE7F3F9FCFE7F3F9F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040000000000000000000000000000000",
INIT_1F => X"4BA550000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0002000087FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974AA550402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"020AA5D7FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5D00000AA007FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAA954BA5504000AA557FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5D00",
INIT_23 => X"7BFFFFFFFFFFFFFFFFFFFFFFFFFAA954BA5500020BA5D7FFFFFFFFFFFFFFFFFF",
INIT_24 => X"7AA974BA5D040200055517FFFFFFFFFFFFFFFFFFFFFFFFAA954BA5500000BA5D",
INIT_25 => X"00000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000080000000",
INIT_27 => X"FFFFFFFFFFFFFAE974AA550002010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"0BA087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550400028007FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAA954BA5D00000BA557FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5D0002",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAA954BA5504020AA5D7BFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"A974AA5D00070925D71FFFFFFFFFFFFFFFFFFFFFFFF7AA954BA5500000825571",
INIT_2C => X"FFFFFFFFFFFFFFEFF7AA974AA5D040500055517FFFFFFFFFFFFFFFFFFFFFFF7A",
INIT_2D => X"D040200008000000000000000000000000000000000000000000000003FFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"A087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550002000087FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAA954AA5D00020AA007FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5504000B",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFF7AA954BA5D00000BA5D7BFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"74AA55000200055517FFFFFFFFFFFFFFFFFFFFEFF7AA974BA5504020BA557BFF",
INIT_33 => X"FFFFFFFFFFDFEFF7AE974AA5D00154105D517FFFFFFFFFFFFFFFFFFFFEFF7AA9",
INIT_34 => X"00000000043FFFFFFFFFFFFFFFFBFDFEFF7AE954AA5D041740055557FFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000007FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(2),               -- Port A write enable input
DIA(0)   => data_write_a(22),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(22),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(2),               -- Port B write enable input
DIB(0)   => data_write_b(22),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(22),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_23_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"EF20906D902424807BC8241BC81801B97D38AD3C0800103362A6741C80A12A02",
INIT_01 => X"001FFF8409F089003B4422000D80C80106804A7951C5B9D1C828043EA28838F9",
INIT_02 => X"028406A002DC176444683862400003111001303FFC00F240D50146013B300500",
INIT_03 => X"0006C90C010203F80005DC00C52FC380BEAC25886C02034800200200A1008008",
INIT_04 => X"17DFFF8049000BFF878314BFF8488890979800002F702002BB807A068403C280",
INIT_05 => X"DA07F0000000007FF020C814380011FE5E1C2FC3E05FFFF90020000808900010",
INIT_06 => X"10004C9690A8CA008024685184097E81E872C8FFE900FC31348EFDF03BE15E22",
INIT_07 => X"402000001FFBFFFD00080200B8140011F0D8C108155542018D1A302193E94004",
INIT_08 => X"41BE1F5F80003FF0002023FFDF79000000000EFFE309606020008005FC000000",
INIT_09 => X"FC83FE1840C0902400300000000000DFFD4004040C4D32BF7C0EE860003CE680",
INIT_0A => X"10018C24110A860006C620C0312241C482B20420CC56924E2199000C00415037",
INIT_0B => X"4669070510C90C14304043040430404304043040430404304043040218202182",
INIT_0C => X"008000105400C00400100000A018000801000C024000004A940000FFDF820604",
INIT_0D => X"100152100801C17E61841950B1C10FFF57FFC02812F00429DC92C40002000100",
INIT_0E => X"10015210088528E00E02C8200A430A424202A1CAF13F214001521001CBF03F21",
INIT_0F => X"01C1C044006D0C94FB94320880603C420B8001CBF03F214001521001CAF13F21",
INIT_10 => X"30182800A018D9CA8000648528E00D12480202C86040902AC60BACDF0E02D020",
INIT_11 => X"0445C19960A00026880C006739000009B00300010AF5052419D1964419028014",
INIT_12 => X"01844068880CE72000013600600332C140004D101808458A5602E00089202911",
INIT_13 => X"41D0B9023402085020825132C8CB5B4040301009408021144CB042F880100C06",
INIT_14 => X"8E17C0D240406519400500840A9524EE38A1F80E02120018390320F050144CB2",
INIT_15 => X"01004010040100401004010040100100040040000000000001000900FBFFE000",
INIT_16 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_17 => X"0040100401004010040100401004010040100401004010040100401004010040",
INIT_18 => X"0000000000000000000000000000000000000000000000001004010040100401",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000000000000000000000000",
INIT_1F => X"4BA5D0400010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000007FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974BA5D0002000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"00010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA550002000007FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAE974AA550400000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5500",
INIT_23 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550402010087FFFFFFFFFFFFFFFFFF",
INIT_24 => X"FAE954AA5D00000AA007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA55040200008",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010000000000",
INIT_27 => X"FFFFFFFFFFFFFAE974BA5D0400010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0000010007FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAE974AA550002010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA550002",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550400010087FFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"E954AA5D0402038007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550400028007F",
INIT_2C => X"FFFFFFFFFFFFFFFFFFAE954AA5D00020BA087FFFFFFFFFFFFFFFFFFFFFFFFFFA",
INIT_2D => X"D0402010000000000000000000000000000000000000000000000007FFFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000087FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAE974BA550002010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D000001",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFFFAE974AA550002000087FFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"54AA5504000BA087FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA550400010007FFF",
INIT_33 => X"FFFFFFFFFFFFFFFFAA954AA5D04000AA087FFFFFFFFFFFFFFFFFFFFFFFFFFAE9",
INIT_34 => X"000000007BFFFFFFFFFFFFFFFFFFFFFFFFFAA954AA5D00020AA007BFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000007FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(2),               -- Port A write enable input
DIA(0)   => data_write_a(23),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(23),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(2),               -- Port B write enable input
DIB(0)   => data_write_b(23),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(23),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_24_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100600007FFF000080108004000800020000840041000080808",
INIT_02 => X"0000068002CC07400000090C080002000000103FF811F150231000520ABE4404",
INIT_03 => X"210A0600000203F80005DC00000DC3801EA000000745C4010220000000008000",
INIT_04 => X"07C5FF804900026F8780001DF8000000079800000F300002998078068003C080",
INIT_05 => X"C207F0000000007FF0000004380001FE1E1C07C3E00CFFF80000000000000000",
INIT_06 => X"0002648240F20035A0102000BD0000002802C87FC800FCAA035400001B918600",
INIT_07 => X"0000000001FBFFEC4D2B4AD0B8129063B2CC0000100042018408142F16C01848",
INIT_08 => X"008E1F5F80001FF0000000FFDF78000000000EFFE001600000000005FC000000",
INIT_09 => X"E883FE180000000000300000000000DFFD0000002A80D500000671000004A000",
INIT_0A => X"10018C0411020600048620C030020502000200000400920A2198000800404037",
INIT_0B => X"0641060400C00C00304003040030400304003040030400304003040018200182",
INIT_0C => X"000000001000C00000000000000240058000000000000000000000FFDF000404",
INIT_0D => X"E00880104809C1666594584031010FFF56FFC000104000000010440000000000",
INIT_0E => X"E0088010492064206100E81084200048C0804012500021B00880108012500021",
INIT_0F => X"04100144800803419043064900C0020501840012500021B00880108012500021",
INIT_10 => X"1018140F02C0000809408D206420530270040410004C840041A0D80054109038",
INIT_11 => X"110002C9E8010C00010480B35A0300400041020902F60002260D65B361BAA104",
INIT_12 => X"0228204300166B4060080008240593D0021800020818B06D9802F00030C02060",
INIT_13 => X"143B62023C00142800B04400095DFF90203020042108603100061516EE800C06",
INIT_14 => X"DC1180C7804400044029208301040214AE4C7C02000040206602C10B48110006",
INIT_15 => X"00000000000000000000000000000000000000000000000000000000FBFFE000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"DD5EDCF9822659B6888332000000000000000000000000000000000000000000",
INIT_19 => X"F3CF3CF3CF3CF3DF7DF7DF7DF7DF7DF3DF3DF3DF3DF4D30C2432AEBAEBFE5A15",
INIT_1A => X"C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783DF7DF7DF7C",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000F0783C1E0F0783C1E0F0783",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201008000000000000000000000000",
INIT_1F => X"4BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974BA5D0400000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"00010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000007FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAE974BA5D0000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_23 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0002000087FFFFFFFFFFFFFFFFFF",
INIT_24 => X"FAE974BA550002000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D000200000",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010080000000",
INIT_27 => X"FFFFFFFFFFFFFAE974BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000087FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAE974BA5D0400010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0000010007FFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"E974BA550002000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0000010007F",
INIT_2C => X"FFFFFFFFFFFFFFFFFFAE974BA550002000007FFFFFFFFFFFFFFFFFFFFFFFFFFA",
INIT_2D => X"D0402010080000000000000000000000000000000000000000000007FFFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAE974BA5D0400000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040200",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000087FFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"74BA5D0000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0000010087FFF",
INIT_33 => X"FFFFFFFFFFFFFFFFAE974BA550000010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE9",
INIT_34 => X"000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA550002010087FFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(3),               -- Port A write enable input
DIA(0)   => data_write_a(24),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(24),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(3),               -- Port B write enable input
DIB(0)   => data_write_b(24),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(24),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_25_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100200002000000080100004000000020000800041000080808",
INIT_02 => X"0000068002CC474000000800000002000000103FFCE302008000000880844A04",
INIT_03 => X"00000040700803FC0105DE00020DC3801EA00000040000000020000000008000",
INIT_04 => X"47C5FFC04904026F8780081DFC040000079C92484F30499299837C168003E400",
INIT_05 => X"C207F0382004407FF0000004382281FF1E1C07C3E00CFFFC090004B05000200A",
INIT_06 => X"1009015C4000000020000000390C10002802C87FC800F8000000000019810600",
INIT_07 => X"0501000001FBFFFD480A0280A816002010800001000054018408102000000002",
INIT_08 => X"0C8E1F5FA21C9FF8004000FFDF7C062031863EFFF75D78004001010DFC000020",
INIT_09 => X"E883FE180C00000000300000000000DFFF00180800000000000660100000A000",
INIT_0A => X"1001DCCC31222730A49620C030020100000200000400921A21D8000804404037",
INIT_0B => X"0641062400C00C00304003040030400304003040030400304003040018200182",
INIT_0C => X"C11160845004D04820000000000000000000000000000000940000FFDF000404",
INIT_0D => X"000800000801C0786184185031810FFF56FFC02812E0182000F2C48304418220",
INIT_0E => X"0008000000002020000008000000000800800002400001000800000002400001",
INIT_0F => X"0000010000000000900000080000000400000002400001000800000002400001",
INIT_10 => X"1000000002002000004000002020000200000000000404000000880000001000",
INIT_11 => X"010000082000000001000001080000000040000100C600800001040000040009",
INIT_12 => X"0000000100002100000000080000104000000002000000081001000000000040",
INIT_13 => X"0010200000000000001004000001080000400080000040010000001080001008",
INIT_14 => X"8C11808200400000400000C20000000420000000030280000000010000010000",
INIT_15 => X"82208822088220882208822088A20C52082081A30080000002005008FBFFF001",
INIT_16 => X"2208822088220882208822088220882208822088220882208822088220882208",
INIT_17 => X"2088220882208822088220882208822088220882208822088220882208822088",
INIT_18 => X"29432D518B45265D82BB4101000005FFFFFFFFFFFFFFFFF82208822088220882",
INIT_19 => X"24924924924924820820820820820820924820924824000A6242B4D34D7F7451",
INIT_1A => X"AC562B158AC562B158AC562B158AC562B1188C46231188C46231189249249249",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000162B158AC562B158AC562B158",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000000000000000000000000",
INIT_1F => X"4BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"02000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAE974BA5D0402000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_23 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000007FFFFFFFFFFFFFFFFFF",
INIT_24 => X"FAE974BA5D0400000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040000008",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010000000000",
INIT_27 => X"FFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAE974BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000007FFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"E974BA5D0400000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000087F",
INIT_2C => X"FFFFFFFFFFFFFFFFFFAE974BA5D0400000007FFFFFFFFFFFFFFFFFFFFFFFFFFA",
INIT_2D => X"D0402010000000000000000000000000000000000000000000000007FFFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"74BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000007FFF",
INIT_33 => X"FFFFFFFFFFFFFFFFAE974BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE9",
INIT_34 => X"000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000007FFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000007FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(3),               -- Port A write enable input
DIA(0)   => data_write_a(25),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(25),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(3),               -- Port B write enable input
DIB(0)   => data_write_b(25),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(25),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_26_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"E9264EAB20190CA3BA4997AA9002AE9C001006B0778015CFA17E0811039879C7",
INIT_01 => X"F1FFF9BB1F773C7F9BB07DFFFDD863FC5FFF3FEFFBBF9FFB22FFFBC7B9F30686",
INIT_02 => X"9B3184F8AFDEAF300029E4E300FC78A6258548EFFA71C00172082400003A2161",
INIT_03 => X"0084F0FF7FFF1FDD3FEFDCDE981DC3FF5F0D294A7B2B18A0001B9CE6CC606E73",
INIT_04 => X"0FC5DFD7EDFFD66F87FE605DDDBFF3690F9EDB7F5F7AFF639BD7DE37C2FEF591",
INIT_05 => X"F205F0F8E9D199FF76DFEE1C3FCC3FF7BE1FD7C3FFACFBFFDFF7B4FEFFDAA10E",
INIT_06 => X"042648C40179912406C1830639AFBEC14489737FDC00B13BB79DFDB83BF4112A",
INIT_07 => X"763A844769FFBFE4398E4390BB9C28B1D0F049080414583F9468D1AEFC000060",
INIT_08 => X"02C05FD7BC471FBD13D981F7DF7D7E6171AF3FEFE8A3E679FAC1FD1FFFBEB000",
INIT_09 => X"F8CFFE38FF7F6BD928F1ABB47476B5FEF9F59F5FCEEDE73FEE0EFC53B079F5CC",
INIT_0A => X"315BDDCC3B336F7C548667D47B7737AF3FD62601EDC2B66A67B9D60FE4C4427F",
INIT_0B => X"06E19F4DA0E80E903DE3035E3035E3035E3035E3035E3035E3035E981AF181AE",
INIT_0C => X"EBFBF7FEBD66DBFCA3F87501AE7B080607307DCFE1D4077B4D026FFFFBFFAFCD",
INIT_0D => X"0007E010084BCD7FF1B61B5C33813FFFFCFFC7D7D51D6F5FDCB935D7AFEBD7F5",
INIT_0E => X"0007E01001BD8020500008001F010040520201F45EC0010007E01001F45EC001",
INIT_0F => X"1DC0004600400F781429C0080000770001A001F45EC0010007E01001F45EC001",
INIT_10 => X"10003C064000E408010081BD8020600200001EC00040B02007EC09A0E0001000",
INIT_11 => X"360403E434588007200D00F88C84C081C203404B3BFD0402346235408402C080",
INIT_12 => X"07B00040091F1190982038406807C868B1000E401A08FE0012040000FC002001",
INIT_13 => X"7D00212000007C400082D81009FC08281D00001F010021560406758091454000",
INIT_14 => X"FFBFF5FA1040076065F730FC08043A903A80008320C0403C3400008860160406",
INIT_15 => X"D7F5FD7F5FD7F5FD7F5FD7F5FDFF7F7F7F77F9F761FFBFDFFDE5BFFFFF7FF005",
INIT_16 => X"7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5F",
INIT_17 => X"F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD",
INIT_18 => X"B79E923C2CD990AA7F0DDB6B910C8DFFFFFFFFFFFFFFFFFD7F5FD7F5FD7F5FD7",
INIT_19 => X"30C30C30C30C30C30C30C30C30C30C30D34D34C30C35F7AA9ABF0E38E3A8EB62",
INIT_1A => X"C26130984C26130984C26130984C26130984C26130984C26130984C30C30C30C",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000130984C26130984C26130984",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000000000000000000000000",
INIT_1F => X"4BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"02010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_23 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFF",
INIT_24 => X"FAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010000000000",
INIT_27 => X"FFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"E974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007F",
INIT_2C => X"FFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFA",
INIT_2D => X"D0402010000000000000000000000000000000000000000000000007FFFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"74BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFF",
INIT_33 => X"FFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE9",
INIT_34 => X"000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(3),               -- Port A write enable input
DIA(0)   => data_write_a(26),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(26),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(3),               -- Port B write enable input
DIB(0)   => data_write_b(26),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(26),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_27_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"00080A40000A41248002029000050A088000008242A0004404480002000A1155",
INIT_01 => X"F1FFF1C11F781C129C107DFFFE0860941E81258CA2B71C2220EC1B86E1A00002",
INIT_02 => X"183080988B2EAE00002BE001117C78C6848140CFFA0000800042008000011081",
INIT_03 => X"000000FF7CF91F1D3DEF3CDA881D23FB5C0C21085B0B0820001318C60C204C63",
INIT_04 => X"8FC51FD7EDFDD66E47EE205D1DB7F1490E5EDB7D5CBADB2385D79C3643D4E580",
INIT_05 => X"E001F0C0C991BBFC76DFEA1A3F8C3BC7391F9723FF2CE3FCD6D13096B79C8106",
INIT_06 => X"40000001000000084041830600A40C415004637FC4003021259CFDB01BF80028",
INIT_07 => X"3158954761FA3FE402088220AC1108001080400A400041018468D1A060000050",
INIT_08 => X"02005F0784411E390A4881C7BEFC5F6171CE2F8FE823E778DAC16C1FFBBC9000",
INIT_09 => X"F0C7FEBABF3F6BD108F40E04C0C084F0F8B58B5B8849673F6C0E7A01B00914C4",
INIT_0A => X"B51BFDCC39732F3554866AD57C37BEAF1C152201A4C0B6EA63AAD60B60D4427F",
INIT_0B => X"06F18FC5A0E00F0038D1030D1030D1030D1030D1030D1030D1030F0818688186",
INIT_0C => X"AB6AD7EAB962CBD8A3A83101F47E08040510768EA0C406630D0226FFE375ADE5",
INIT_0D => X"000760000843C561E5C55C42B9011FFF48FFCC57550D63564D1D2556ADAB56D5",
INIT_0E => X"0007600004BD8020100008001F010000130201E44A40010007600005E44A4001",
INIT_0F => X"1DC0000208400D781020C00800007700002005E44A40010007600005E44A4001",
INIT_10 => X"10003C064000C400018080BD8020200200001EC00000382006EC0820A0001000",
INIT_11 => X"3E0403A424108007200102E888808081C20040431BC504021462354004004080",
INIT_12 => X"07B00000015D1110102038400817484821000E400204FE0010040000FC000000",
INIT_13 => X"7D00202000007C400000F81001FC08080500001F0100005E0404758081014000",
INIT_14 => X"8DBBB5FA10400360649310FC08003A903A8000012040403C34000080201E0404",
INIT_15 => X"56D5B56D5B56D5B56D5B56D5B56D7E3D7B57B1C4E17F0944B8D596EEFC7FF001",
INIT_16 => X"6D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B",
INIT_17 => X"D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B5",
INIT_18 => X"2D0200903950C080420948E2D10E8FFFFFFFFFFFFFFFFFF56D5B56D5B56D5B56",
INIT_19 => X"00000000000000000000000000000104000000000004000E5E420000002921C4",
INIT_1A => X"28140A05028140A05028140A05028140A0100804020100804020100000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000140A05028140A05028140A050",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000000000000000000000000",
INIT_1F => X"4BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_23 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFF",
INIT_24 => X"FAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201008",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010000000000",
INIT_27 => X"FFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"E974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087F",
INIT_2C => X"FFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFA",
INIT_2D => X"D0402010000000000000000000000000000000000000000000000007FFFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"74BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFF",
INIT_33 => X"FFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE9",
INIT_34 => X"000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000007FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(3),               -- Port A write enable input
DIA(0)   => data_write_a(27),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(27),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(3),               -- Port B write enable input
DIB(0)   => data_write_b(27),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(27),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_28_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"02200AA400180030808802A900002A08001280A08A801044104A1000001818C3",
INIT_01 => X"50A00011460214428114180000882214413D0A71592A01D92213D28005210202",
INIT_02 => X"8A54800A210200111100C2110054289220810440030404010844000444410001",
INIT_03 => X"1080010208B51400007800000A000001000108C21008092000018C6295200631",
INIT_04 => X"0008000000017000000028000001610300000010000802202040012040040011",
INIT_05 => X"2000044440048880026A22000026A20000000000000000004994140203000064",
INIT_06 => X"1400922401041008004891224228810080010200040001020800000004000008",
INIT_07 => X"150B001328000001404010040084088404200020455514000224489028492201",
INIT_08 => X"00414000201800004080A0000002480B04008100011000088800081002C19020",
INIT_09 => X"000400001036584108415B4A6A694A0000100101C08200000001000190200044",
INIT_0A => X"004800210C19808400500010009110091500020B408820000200400040811600",
INIT_0B => X"40000800B00100040D8140581405814058140581405814058140580A02C0A02C",
INIT_0C => X"00200248010201008298150006210802043058C46054032981002D00201C8081",
INIT_0D => X"0000A00000400600841041108280300008000140000401028008330000800040",
INIT_0E => X"0000A000000080001000000000000000500000040A40000000A00000040A4000",
INIT_0F => X"00000006000000080020C00000000000012000040A40000000A00000040A4000",
INIT_10 => X"00000000000024000000000080002000000000000000A00000040020A0000000",
INIT_11 => X"2200000404108000000900008080808000024040152000000020000004004080",
INIT_12 => X"0000000009001010102000004800080821000000120002000004000000000001",
INIT_13 => X"2000002000000000000288000020000805000000000001420000200001014000",
INIT_14 => X"408010000000022000D610280000080000000001204000000000000820020000",
INIT_15 => X"00401004010040100401004010042024210218734CD52150A840827504000000",
INIT_16 => X"0401004010040100401004010040100401004010040100401004010040100401",
INIT_17 => X"4010040100401004010040100401004010040100401004010040100401004010",
INIT_18 => X"05822140048D2E57B1348141845C200000000000000000000401004010040100",
INIT_19 => X"04104104104104104104104104104104104104104101A6A0A0EB1861863BC422",
INIT_1A => X"2C160B0582C160B0582C160B0582C160B0180C06030180C06030181041041041",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000160B0582C160B0582C160B058",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000000000000000000000000",
INIT_1F => X"4BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_23 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFF",
INIT_24 => X"FAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010000000000",
INIT_27 => X"FFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"E974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007F",
INIT_2C => X"FFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFA",
INIT_2D => X"D0402010000000000000000000000000000000000000000000000007FFFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"74BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFF",
INIT_33 => X"FFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE9",
INIT_34 => X"000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000007FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(3),               -- Port A write enable input
DIA(0)   => data_write_a(28),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(28),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(3),               -- Port B write enable input
DIB(0)   => data_write_b(28),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(28),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_29_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"79964E4BA01DACAB9E659792D00AAE160002829C7FDFEFCEE97C2815039D70C3",
INIT_01 => X"50BFF9AB0775343F9AB01DF80D5821FC0FFF3FEFD1AF9FF1207FFBC7B9720586",
INIT_02 => X"0D15846807D207200021C4E200D428A2018408600271C000720A0000003A2161",
INIT_03 => X"0000B0027BBF17C43E6DC05E1A0DC07D1F0000803B2819A00019084345606421",
INIT_04 => X"07CDC047A4FB526F807C681DC4B97369078249370F482E62BA414627C2FE3000",
INIT_05 => X"F204007861C088FF0EFF260407C427F19E03C7C01F8CF80749B390EA4BCA202C",
INIT_06 => X"000248C00079800406C081023B233E804488527FDC008019968D74982C94110A",
INIT_07 => X"5229000221FF8000398641903B082831D05000200000083F942850AEB4000221",
INIT_08 => X"00805FD0180E1F8C1111A0F041056A0100A11FE000916249A800B915FE82B020",
INIT_09 => X"F80C000055FF7C492840AAB45456B55E015015058665A31DA603A4539058F54C",
INIT_0A => X"000850400A11414C005005000B51158936D20601A98A204006114005C4800217",
INIT_0B => X"40201948B029029409A3401A3401A3401A3401A3401A3401A3401A9A00D1A00C",
INIT_0C => X"40B1225C1506512C83E85500AC3A080406305587A154023141006DFFF89E82C9",
INIT_0D => X"0000A01008480D3EB4A24A0C910037FFFC0007C7C0140D0B50A8218102C08160",
INIT_0E => X"0000A010010080005000000000000040520000141EC0000000A01000141EC000",
INIT_0F => X"00000046000002080429C0000000000001A000141EC0000000A01000141EC000",
INIT_10 => X"00000000000024080100010080006000000000000040B000010401A0E0000000",
INIT_11 => X"3600004414588000000D00108484C080000340483B590000202000008402C080",
INIT_12 => X"00000040090210909820000068008828B10000001A0802000204000000002001",
INIT_13 => X"20000120000000000082D800082000281D000000000021560002200011454000",
INIT_14 => X"B29450580000066021F6303C000408000000008320C000000000000860160002",
INIT_15 => X"816058160581605816058160589625662522506344FF9FCFFF62EB6DFF001004",
INIT_16 => X"1605816058160581605816058160581605816058160581605816058160581605",
INIT_17 => X"6058160581605816058160581605816058160581605816058160581605816058",
INIT_18 => X"F2DDCFFFBEFFCF07FFBFFD41800C05FFFFFFFFFFFFFFFFF81605816058160581",
INIT_19 => X"7DF7DF7DF7DF7DF7DF7DF7DF7DF7DD75D75D75D75D77FFBF3F7DFFFFFFD779F3",
INIT_1A => X"FEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDF7DF7DF7DF",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00001F7FBFDFEFF7FBFDFEFF7FBFD",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000000000000000000000000",
INIT_1F => X"4BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_23 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFF",
INIT_24 => X"FAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010000000000",
INIT_27 => X"FFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"E974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007F",
INIT_2C => X"FFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFA",
INIT_2D => X"D0402010000000000000000000000000000000000000000000000007FFFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"74BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFF",
INIT_33 => X"FFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE9",
INIT_34 => X"000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(3),               -- Port A write enable input
DIA(0)   => data_write_a(29),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(29),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(3),               -- Port B write enable input
DIB(0)   => data_write_b(29),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(29),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_30_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"FFDFF3FC3EFFF7FFFFBFFA000000000000000000000000000000000000000000",
INIT_19 => X"F3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF5F7AEBEBFBEFBEFFEFFF7",
INIT_1A => X"CFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCF3CF3CF3C",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000007F3F9FCFE7F3F9FCFE7F3F9F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000000000000000000000000",
INIT_1F => X"4BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_23 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFF",
INIT_24 => X"FAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010000000000",
INIT_27 => X"FFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"E974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007F",
INIT_2C => X"FFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFA",
INIT_2D => X"D0402010000000000000000000000000000000000000000000000007FFFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"74BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFF",
INIT_33 => X"FFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE9",
INIT_34 => X"000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(3),               -- Port A write enable input
DIA(0)   => data_write_a(30),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(30),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(3),               -- Port B write enable input
DIB(0)   => data_write_b(30),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(30),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_31_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"129000008004A00804A40000400800020000000C005FEA005800200400050100",
INIT_01 => X"A15FF18019700810180065FFFC0040801E80258CA2951C2200EC0906A0804140",
INIT_02 => X"146000808A0C060444692000402850040400408FF80000000010000000004000",
INIT_03 => X"000000FD74480B1C3D951C5A800D03FA1C0C21084B0300000012108518004842",
INIT_04 => X"07C51FC7EDFCA26E07EE001D1CB6904A061EDB6D4C30490281831C1602D0E480",
INIT_05 => X"C001F0808181117C7C95C8183FA099C7181F8703FF0CE3FC0201209010988002",
INIT_06 => X"00000000000000010001020400840C41C000617FC0003021259CFDB01BF00020",
INIT_07 => X"0000000441FA3FE400080200A810000010804008100040018448912040000040",
INIT_08 => X"00011F0780011E38004801C79E7C162231862E8FE00166704041240DF93D0000",
INIT_09 => X"F0C3FE180D89279000B00000000000D0F80088080849673F6C0E780020091480",
INIT_0A => X"1011DCCC31222730048620C4382204A608142002A440924A6188020920404437",
INIT_0B => X"0661874500E00E00304003040030400304003040030400304003060018200182",
INIT_0C => X"810040801060C04821202001A05A00040100240A80800442040202FFC3200444",
INIT_0D => X"000740000803C0616184184031010FFF40FFC407500020004C10060204010200",
INIT_0E => X"0007400000BD0020000008001F010000020201E04000010007400001E0400001",
INIT_0F => X"1DC0000000400D701000000800007700000001E04000010007400001E0400001",
INIT_10 => X"10003C064000C000010080BD0020000200001EC00000102006E8080000001000",
INIT_11 => X"140403A020000007200000E808000001C200000308C504021442354000000000",
INIT_12 => X"07B00000001D0100000038400007404000000E400000FC0010000000FC000000",
INIT_13 => X"5D00200000007C400000501001DC08000000001F010000140404558080000000",
INIT_14 => X"8C1380DA10400140640100D4080032903A8000000000403C3400008000140404",
INIT_15 => X"02008020080200802008020080200C1808008184012A08041202500AF87FF001",
INIT_16 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_17 => X"0080200802008020080200802008020080200802008020080200802008020080",
INIT_18 => X"000000000000000000000002001005FFFFFFFFFFFFFFFFF02008020080200802",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000000000000000000000000",
INIT_1F => X"4BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_23 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFF",
INIT_24 => X"FAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010000000000",
INIT_27 => X"FFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"E974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007F",
INIT_2C => X"FFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFA",
INIT_2D => X"D0402010000000000000000000000000000000000000000000000007FFFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"74BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFF",
INIT_33 => X"FFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE9",
INIT_34 => X"000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(3),               -- Port A write enable input
DIA(0)   => data_write_a(31),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(31),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(3),               -- Port B write enable input
DIB(0)   => data_write_b(31),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(31),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_0_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"ED39BA795990D275FB4A6E96ACC4731DEA4598B0AFB54867F6EE4618C3749807",
INIT_01 => X"58A0047D8607944AC7DA180001ECA2444042106208408208C20022E9173734B3",
INIT_02 => X"8B1E49562021F8051500147A0E162923024F28000415F5787B09FBF999BB1EFC",
INIT_03 => X"1013BF028A959403C06A23A147723C01E140088280C4CF6996088862C7922221",
INIT_04 => X"781A003802015D9078011DE20340699198600000B08694916434804825241311",
INIT_05 => X"2CA000587E10C880036A3103C00F2000E1E0383C00730002B4409845E4425171",
INIT_06 => X"179B48CFF95DCF9EF730E1C3BB731138AF7B888025340C0888430047040FEE18",
INIT_07 => X"AF155113160400185F87C1F05707D415E664A6E7C5551EBE783060CEB164833F",
INIT_08 => X"4D7E40002B7AE005FDB47600208229010C6101001EFE198C96B0528202C0DCB4",
INIT_09 => X"062400608234D864444081048A80CC00062D42D30222108091C107A1DA040267",
INIT_0A => X"204A21008E514844EB5145000255DA599581D3A9583C24351240B58298011308",
INIT_0B => X"E08C4830F81380CE0F89E07A9E0789E07A9E0789E07A9E0789E070CF0184F038",
INIT_0C => X"3A4E9D63EA180EB150CA1CA45C254D4AF4AA414568729139F2A12C0000016110",
INIT_0D => X"F0009E0FC048211E9C11C31F82E4A000890022B827EB52F52347F174E93A749D",
INIT_0E => X"F0009E0FCC42EFDFBF0AE03080E2AEB2E0F1F80FA97FE0F0009E0FC40FA97FE0",
INIT_0F => X"0231F0BD9E3FC08FEBD6F661C0E008C3CB5F040FAB3FE0F0009E0FC40FAB3FE0",
INIT_10 => X"20180309A0F83BE2B87C7C42EFDFBF187806013879BA878FE807F65FBF12E038",
INIT_11 => X"0BE9F01FC8B38C2098DAE007F323A0C83136B248831ACBFC8BBDCAB779BC699F",
INIT_12 => X"004C72BEC800FE7464290626D7003F9947184131B59003FFEC07F00003F01FB9",
INIT_13 => X"A0FFDA2A3C0202B8776A2FA7F023F7D065703080E29F1B2BE9F8A27E6E915C0E",
INIT_14 => X"016C2D25E52630BB1AE49C2BA7F98D6F846DFC0C2352A0024B83F07F198BE9F8",
INIT_15 => X"749D2749D2749D2749D2749D2749F285F25D2C500815A5522CB5A4B400000CD4",
INIT_16 => X"49D2749D2749D2749D2749D2749D2749D2749D2749D2749D2749D2749D2749D2",
INIT_17 => X"9D2749D2749D2749D2749D2749D2749D2749D2749D2749D2749D2749D2749D27",
INIT_18 => X"31C136AD8E9B562BA39E2600654BA800000000000000000749D2749D2749D274",
INIT_19 => X"4104104104104104104104104104104104104104104104109C83B8E38E2ABE71",
INIT_1A => X"0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0410410410",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000007C3E1F0F87C3E1F0F87C3E1F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000187FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"BAF7FFD55EF007FD75EFFFAE97555557BD75EF5D000000000000000000000000",
INIT_1F => X"000AA843FE00AAFBE8B45AA803DFEFA28428B455D0017410A28428AAAA2FBD54",
INIT_20 => X"FEBAA2D5401450051401555D7FC0145F7AEBFFFF08002AA10A2AABFEAAA2FFC0",
INIT_21 => X"D755555517FFEFA280021FF082E974AA5D7BFFE000804000BAAAAAAAB45557FF",
INIT_22 => X"EA8B45005168A10AA8028A10087FD7410557FC21555D51574AAA2FFE8B455D7B",
INIT_23 => X"AE95410AA80000005D003FEAAFFAEBFE00A2803FEBA002A820AA0800174BA5D2",
INIT_24 => X"2AEA8A10000417410A2FFE8BEFF7FFE8B45FFFBC00005D003FF45557FC01FFFF",
INIT_25 => X"00000000000000000000000000000000000000557DF5500003DFEFFF84175EFA",
INIT_26 => X"5F524AFE38B780154BAFFF1D54AF0075D75EFEBAE9554540754717F1F8000000",
INIT_27 => X"50B6AABDE12BEA0AF010B7D1F8F47E00A2DB45AA8A3AFD7B68E2AB78550E1255",
INIT_28 => X"E9257F1E816D557095EAAA2D1401D500002A150038038E285D7F78FD7000B6AB",
INIT_29 => X"5A87AAD178A8002D1D21C5E8257D5C7AA854008700249243A412EBFF5542A43F",
INIT_2A => X"52A82000E3A5D2150AB8F401471EDBC0B680900AAF52B474385D75C502D15754",
INIT_2B => X"FD7E9541242FE920AD082E10A28F6A150012A2F02AFFDF40E85F475451D502D1",
INIT_2C => X"0550E87B7A405B52AAD152BD00151EAFEDB52E3F1EFFFF485A2DA3D5D24BD417",
INIT_2D => X"57F40545850000000000000000000000000000000000000000000005AAF55508",
INIT_2E => X"F7AEAABFF5D2A81151FB8635A02FA69574BAF7D5555AF0D79D55FFA2AC974450",
INIT_2F => X"8D46F6ABE7082AAAAF2FAC77FE00FF16565B2FA9075F4F7B3EBDF50FEAEAAB55",
INIT_30 => X"56803CE3AEB038662E5D81406014D5D51F5E08A394003A908B8410E707EF34A0",
INIT_31 => X"4AF0151555AF58794040077D774FAE8C798A11A0EAEF75F7AA84001A7052C952",
INIT_32 => X"4E1870108B11020AD4AA05542A0A05051023F9A9D57B63BFBF906CB45FABC095",
INIT_33 => X"F5F0DA6BC9525688C1A2A0C06E9FEE5555BE48AB2A2AE0A0F20C43EAC562245B",
INIT_34 => X"000000FF80F55E25C00A0BA7FBED407A97F6F35F498B96BEB12DAAB77558ABD5",
INIT_35 => X"8000000FF8000000FF8000000FF8000000FF8000000FF8000000FF8000000FF8",
INIT_36 => X"00000000000000000000000000FF8000000FF8000000FF8000000FF8000000FF",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000008000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(0),               -- Port A write enable input
DIA(0)   => data_write_a(0),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(0),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(0),               -- Port B write enable input
DIB(0)   => data_write_b(0),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(0),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_1_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"212C001411984004084D000508C53810A03D1450E839B003342114428A000803",
INIT_01 => X"08000010400A0008010600000084005000400002000000000000000000140000",
INIT_02 => X"C084484000002014400205851002007030450E0000A606C8C44CB4C6666C00E0",
INIT_03 => X"CCF7CE0002058001000000800240200001018CA1800001091408463061120118",
INIT_04 => X"082800100000000040000900010000100040000000008411600401C02100000C",
INIT_05 => X"10800202080422000020012200000000810000200000000004020C00200011A0",
INIT_06 => X"56BDBFBC48C315A8660C18305750C008940D8000011000820001000104050004",
INIT_07 => X"8B4344400004000150248912154404C6060A2FE24555013E13060C158AC97F01",
INIT_08 => X"00082080087A000559102400200281000469000008B000000090108000400430",
INIT_09 => X"0000000000001004140545402820020000010010208000008041060008200001",
INIT_0A => X"2102210182004840007845004044020000200080080844200000048088000000",
INIT_0B => X"48800000190191064620646A06468064680646A0646A06468064690321503234",
INIT_0C => X"02008100200800A1100707040101E20BE0B002605C1C110848200C0000000800",
INIT_0D => X"F000A000C0000012187087010AE4B00000000810010040108104100408020401",
INIT_0E => X"F000A000CC4200002F08E03080000010F18058000003C0F000A000C4000003C0",
INIT_0F => X"000000078808C00000023461C0E00000012704000003C0F000A000C4000003C0",
INIT_10 => X"201803000000240218C0044200001E1878060000000AAC00680000001F10E038",
INIT_11 => X"2100B00048230C200009A0001303204800025200040A00D000000202090C281F",
INIT_12 => X"00000002C9000260640900004D0000904618400012900001EC03F00000000039",
INIT_13 => X"80025A0A3C020000002A8400B00007806070308000000961002880204A901C0E",
INIT_14 => X"000801046004308A185000020128000904285C0C0312A0020000000838810028",
INIT_15 => X"0401004010040100401004010040100010410C002000040280100000000008D0",
INIT_16 => X"4010040100401004010040100401004010040100401004010040100401004010",
INIT_17 => X"0100401004010040100401004010040100401004010040100401004010040100",
INIT_18 => X"48D757DF8A9410218E8A56085142020000000000000000004010040100401004",
INIT_19 => X"555555555555555555555555555554514514514514550431A581924924B02651",
INIT_1A => X"4BA5D2E974BA5D2E974BA5D2E974BA5D2EB75BADD6EB75BADD6EB75555555555",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800005D2E974BA5D2E974BA5D2E97",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000607FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"10AAAABFFFFFF803FE10F7D17FEBA55556AAAAAA800000000000000000000000",
INIT_1F => X"EBAFFD555400557BD54BA5D7FFDF45A2FBD75EFA2AE97555F7FBFFF45FFAE800",
INIT_20 => X"ABEFA2D568A005D5157400AA8028AAAF7FBD54AA002A955555D7FE8ABA082EBF",
INIT_21 => X"FDF55AAFBC0010555540010550417555AA8028BEFAAAE97555082A80000AA802",
INIT_22 => X"BD7410550428ABA5D5168ABA552EBDFEF5D7FEAA00AAAABFEAA007BC0145FFFF",
INIT_23 => X"FFEAB55557FFFEBAAAD568B45A2D5575555D7FC2155F7AEA8BEFAAAA954BA557",
INIT_24 => X"D7BD74000804154BA082ABFF55FFD57DF45F7D568ABAF7AABFFFF082ABFFFFFF",
INIT_25 => X"000000000000000000000000000000000000002EBFFEFA280021FF082E974AA5",
INIT_26 => X"5E175EFF57BF8FC2000BEA4BAE97F78A3FE28E3D17DEAA485FE8E02B50000000",
INIT_27 => X"455571E8A2A087BF8EAAEB8E0016D5D75D54BA5D7BFFF7DA2FFD55EFAAA49554",
INIT_28 => X"157428145A00AA8A2FBD7B6DF6AA28550E10405F7A4AFE38EAA0924921C2FD55",
INIT_29 => X"8E971471C7010B7D168F47400A07A28415A001684104155C5B6DF6DBEFBFAA07",
INIT_2A => X"BFBD7B6A0BF492415FC20105D24AAABF1FFBC7010FF8A38FEF557FEAB78B6AAB",
INIT_2B => X"017EBA4A8EB8F6FFD5FE8B7D557495EAAA2D16D1FDBED56A55557A43DE385FD4",
INIT_2C => X"854008700249243A417FFF41542F5D717FE2AAAA56DEBD17FE3DF7FB7FEBFE38",
INIT_2D => X"07DFCA127B8000000000000000000000000000000000000000000002A3D5C7AA",
INIT_2E => X"AAFBD55FFAA8416545A6FB60F47AF2A00010F78028B15F7823FEAAA2D57DFBA0",
INIT_2F => X"22A38C20B2552E975F758516AAAA0869AAAB8A7C19C55550E8574BA557BFFFEF",
INIT_30 => X"55FFEFBCEE5FBAACB10085EE5DE10A2AEBFF55F7BAAA8565DBAC1112FFAC21A0",
INIT_31 => X"BEA097BEAAFAF2863FA00DD574201E7AD1FFF5575841DE08007FC20480028957",
INIT_32 => X"54FF57EFBFA18D4FBFFF40FF809D4000D7FC00FC5D062BBA05ED5034472A02EA",
INIT_33 => X"7DFBFF6963FCAAA2283CF14050062B0A2F7AE8B5D5D51F5E18ABD5EAFFF2AF95",
INIT_34 => X"000000002CB75F7AA84001A7052C95256807DC31AA8114DE55F5BED201FFFED1",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000008000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(0),               -- Port A write enable input
DIA(0)   => data_write_a(1),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(1),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(0),               -- Port B write enable input
DIB(0)   => data_write_b(1),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(1),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_2_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10E44660018259B2843913100062C98004802322D3E030235201006009B2813",
INIT_01 => X"000AC188084900481C8024A542400340404000720885800802000906E4910204",
INIT_02 => X"82040072AC248C31010204880000007401044C0550200000480E0080001300E0",
INIT_03 => X"0080812C130D0A0D1193088802182142494D218220021100001A8020C1004A00",
INIT_04 => X"090D0AD62824A44A428408540D1610020C6E510818923441A4908B0503404201",
INIT_05 => X"5000A004081122242420480A14A99C428908122144244150906124248C002168",
INIT_06 => X"1400088400450000460000001308890094082015800011012D41D518044C1100",
INIT_07 => X"26731111491C1541324C1114BD880004002040204050413F1400100480000201",
INIT_08 => X"02410582881E0C1511D02082AAAB016A2463288549B044605201D10AE11B0020",
INIT_09 => X"E80394280E40158020B591000800481051241A4A404B5035C60904502054E000",
INIT_0A => X"0102C9E12202EA6014D027C418428E220A5500024808922801A0900A84454458",
INIT_0B => X"4600070110C10D04340043400434A043420434A04342043480434102184021A0",
INIT_0C => X"E9CA34328E44CA1401306100A246000402100C088104010AC8005C5681812B04",
INIT_0D => X"0000A0000801487334E34C1A980001550055481204090A4C01351253A728D194",
INIT_0E => X"0000A000013800004000080000000000500000B01480010000A0000150148001",
INIT_0F => X"0000000608000A500409000800000000012001501480010000A00000B0148001",
INIT_10 => X"1000000000002400000001A100004002000000000000A0000360018040001000",
INIT_11 => X"380001C01048000000090298040440000002400008C400022042004080028000",
INIT_12 => X"0000000009530080880000004813802090000000120C94000200000000000001",
INIT_13 => X"4C000100000000000002E0000950002018000000000001580002508010440000",
INIT_14 => X"7120642000000400015020500004221018000082008000000000000820180002",
INIT_15 => X"5094A5294A5294A52942509425094209461468000822241A03835D88482AB001",
INIT_16 => X"09465094A5294A5294A5294250942509425094A5294A5294A529425094250942",
INIT_17 => X"94650946509465294E5294E5294E5094650946509465294E5294E5294E509465",
INIT_18 => X"080271AE180616A38A18FA204452A7F03F03F07E07E07E05294E5294E5294E50",
INIT_19 => X"20820820820820820820820820820820820820820820490C04102CB2CB2EB2C0",
INIT_1A => X"8944A25128944A25128944A25128944A25128944A25128944A25128208208208",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF1F804A25128944A25128944A2512",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000787FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"AAAA843DFFFAAD1554005D7FD74AA00040015500000000000000000000000000",
INIT_1F => X"F45AAAAA8A10A2AE80010A2AA975FF5D003FE10F7D17FEBAF7D5420AA0855420",
INIT_20 => X"FF45A2AA975EFA2FFD7555FFFBFFF45AAFBC20AAF7D1575EF55517DF555D2EBF",
INIT_21 => X"95555552E974105D517DF55AAAAAABEFAAD1575EFAAAE974AA5D51554BA5D7FF",
INIT_22 => X"E82010F7AABFE10FFD542145FFD5554AA555555555557FE8ABA082EBFFFFAAAE",
INIT_23 => X"FBC0010AA802ABEFAAD540000FFD540000AA802AABAF7FFC2010AAAE821EF552",
INIT_24 => X"A8028BEFAAAE821550851420AA002E800AA08042AB45007FC00BAFFD168BEFF7",
INIT_25 => X"000000000000000000000000000000000000002E80010555540010550417555A",
INIT_26 => X"AE95F40002157F470AABE803AE97A2DF55400557FD54AA1D04001C5150000000",
INIT_27 => X"EF55517DFC5552ABDF45B6AEAFFD5F7A482000BEAE905C755003FE28E3D17DEA",
INIT_28 => X"0BA5FD0154BA5D7BFAF7DA2AE955EFAAA495545E3F5EFF57F7FE80082FFDE105",
INIT_29 => X"8AAF082AB8EAAEB8E0016D5D2A924105D5B7FF7DB6AAAABC7BEDB505EFBEA407",
INIT_2A => X"95038AAAEAF1D7410E80000FF8438E00B6DF68FEF4871D24BA495B5556D5571E",
INIT_2B => X"1ED1EFEAF1EFFFDEAD1C5010AA8E2FBD7B6DF47A00EBDB50000A380AAE28E804",
INIT_2C => X"5A001684104155C5B68E2DBEFBFFBC703AE2DF42AAA002A851C214003FF68007",
INIT_2D => X"50002155510000000000000000000000000000000000000000000002087A2841",
INIT_2E => X"55003FEAAAAD57DEBAA2FDDC01051FBD74BAF7802AB05AAFBD5400557BD54AA5",
INIT_2F => X"7AF7FC20B2F7FBC015D58517FF555D2ABDF55F782BEB47AFAD00010F7AA82155",
INIT_30 => X"55FFFFC20FFF3AE544108410174BA557BEABEFAAEBD55FFAA1456547A2D360F4",
INIT_31 => X"0BA547FD75FF58516AAAA0828AAAB4A78016545540400010557BFDFFFF7822A9",
INIT_32 => X"550AAFACAAA122AA8954BAA2AE9D545002A800A8FF862BA00F2F9E8F0050D442",
INIT_33 => X"954505C417FFFF08555555BAAD335B57AB5155400A2AEBFF45FFFB404007FFBD",
INIT_34 => X"00000000061DE08007FC2048002895755FFAEBCFE57BBA57002DF3C4AAAA002E",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000010000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(0),               -- Port A write enable input
DIA(0)   => data_write_a(2),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(2),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(0),               -- Port B write enable input
DIB(0)   => data_write_b(2),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(2),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_3_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"210C44A20020248B08431120001604B8156023104C40771B3430400A02380206",
INIT_01 => X"015A2A4050B009683C0422C992000B61404040028804A0080A000C16A8990A0C",
INIT_02 => X"C0A406500CE0A95011000D1501005274B5041AB330860281CC08008222170060",
INIT_03 => X"AB488054270F08E1289084C8020420E005A48DA16C021100003A46B06900C91A",
INIT_04 => X"848966150DA0A02941A4080C612A104201C689044382FD403C17E491829B259B",
INIT_05 => X"D006620608843116942508120A208D18A5050160C600D4C894600094B49CA068",
INIT_06 => X"12002D9401C70008060408141788E2C094887033080071913209CC8004640100",
INIT_07 => X"221111454874CCC4122C0932155400C2023940284000003E15020525CE805E11",
INIT_08 => X"020103C9984A0AC511102029869D974214EDBA132891000052C1750B48290020",
INIT_09 => X"60808C8A2E41351020004148A289428730A51E5E644C8233A0090E1020208100",
INIT_0A => X"A4000041A600417914506F955D6422000934000A090A94A020229603A414144D",
INIT_0B => X"469100841001000406D04065040650406D0406D04065040670406C8201782032",
INIT_0C => X"6A4AF532A8040AF821042D01F14084030070262810340402C0000CCE4CC12520",
INIT_0D => X"000800000401C333494594532980733302CCC81300094E5C91200257AD2AD795",
INIT_0E => X"00080000051C0000400000000000000800000190148000000800000450148000",
INIT_0F => X"0000010000000B100409000000000004000005101480000008000004F0148000",
INIT_10 => X"0000000002000000000001B00000400000000000000400000168018040000000",
INIT_11 => X"1000034010480000010002D804044000004000812E4400002440014080028000",
INIT_12 => X"0000000100570080880000080015C02090000002000CCC000200000000000040",
INIT_13 => X"1C0001000000000000104000094C002018000000000040100006418010440000",
INIT_14 => X"4128652000004404010E20500004208018800082008000000000010000100006",
INIT_15 => X"5795A5595A5595A5595A5595A5595E1152556D008028341B13924D80C2E67009",
INIT_16 => X"69565795A5595A5595A5595A5595A5595A559525795257952579525795257952",
INIT_17 => X"95256956579525495E5595A5495E5595A5495E5595A569565795256956579525",
INIT_18 => X"7818F18E0C8514298B0C52A0115009AA9556AAD552AAD5556956579525695657",
INIT_19 => X"24924924924924924924924924924820820820820825042C0000249249202A60",
INIT_1A => X"8D46A351A8D46A351A8D46A351A8D46A353A9D4EA753A9D4EA753A9249249249",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF248086A351A8D46A351A8D46A351A",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"EFAAFFD54AAF7D168B45AAAABDF5500002AA1000000000000000000000000000",
INIT_1F => X"F45FFD168AAA0855420AAAA843DFFFAAD1554005D7FD74AAA284001550055421",
INIT_20 => X"55FF5D003FE10F7803FEBAFFD5420AA080400155AAD5554AAF7802AB4500043D",
INIT_21 => X"28B45A2AE82155A2FBFFEBA0800021550855555FFAA84001FFAAAE80010A2AA9",
INIT_22 => X"168ABAFFFBD54BAAAAE97400A2FBC20AAA284175EF55517DF555D2EBFE00AA80",
INIT_23 => X"AA954AA5D7FFFF45AAAA975EF007BD7555FFFBFDF55AAFBD55EF5D2EBFE10085",
INIT_24 => X"AD1575EFAAAE974AA5D00175555D0015410F7AAAAAAA55043DE00FFFFD5555AA",
INIT_25 => X"0000000000000000000000000000000000000004174105D517DF55AAAAAABEFA",
INIT_26 => X"ABC04001C51551471D7AAF1D05D2EBD56DB7DBEAEBFF551C042AA101D0000000",
INIT_27 => X"92EB842FB5508043FF55EBD56ABD75D5B470AABE8A3AFD7A2DF55400557FD54A",
INIT_28 => X"557FD2082000BEAE905C755003FE28E3D17DEAAEBDF40002550F47155AADB504",
INIT_29 => X"DF40552ABDF45B6AEAFFD5F7A48017DAAFFFAE821C0A0717D1C5B575FFB68E82",
INIT_2A => X"C55D7492E90E3808756DA92EBFFD74BAE3AE85480FFFFC00AABE8E105C755517",
INIT_2B => X"43AE10EAF5C5547FF80954AA5D7FFAF7DA2AE905EF0075D5545E3F5EFF57F7D5",
INIT_2C => X"5B7FF7DB6AAAABC7BEDB505EFBEF5C7092FF801756D490A10438EBA4B8E92410",
INIT_2D => X"D0028A00510000000000000000000000000000000000000000000000E124105D",
INIT_2E => X"AAFBD54005D7BD54AAF78002155515157555AAD142040A2D57FFFFFFAEBFF555",
INIT_2F => X"051AE955F7AAFBC0000AF843FF5500003FF55AAFD6AB455157D74BAF7AAA8B45",
INIT_30 => X"FF557BD74EFFBACD41577B8400010F7AA8215555003FEAAAAC53DEB8A2FDDC01",
INIT_31 => X"0BAF7AA8015558517FF555D2ABDF51F782BCB47ABAE801FFAAFBEAA105D2E955",
INIT_32 => X"214FA2D3EAF57AFFDD7555082AA0AAA00557FEA8A2FDD64BAAF8282012AFFEC2",
INIT_33 => X"820AAAB842AA00000028AB0AAFF48547AE04174BA557BEABEFA2AA951FF88554",
INIT_34 => X"000000002A80010557BFDFFFF7822A955FFFFC21FFF3BE40412DE02955FF082A",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000008000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(0),               -- Port A write enable input
DIA(0)   => data_write_a(3),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(3),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(0),               -- Port B write enable input
DIB(0)   => data_write_b(3),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(3),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_4_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A108400020612C80284210081034849800A000303100048B3432C82904204006",
INIT_01 => X"210668000008004C1C20250E12100368403008418984014902030906A8910200",
INIT_02 => X"120404C0024C0600000206100008402404040C00F104008040080080001310E0",
INIT_03 => X"7728805052470B5C1B873C04121D03845D0020CA0822018000080084C1000002",
INIT_04 => X"0B899E43891686690790485D5C3E02000E9892201D306D03A9835C16029AC186",
INIT_05 => X"C001E080005030767434C0003C8A01D6B81C5703C82CDBC000072400089C8120",
INIT_06 => X"1000088100410000460002041300004084080070D00030032009700024641102",
INIT_07 => X"4261950408CCBC2012048310951000000003402A4000143E1008912480000211",
INIT_08 => X"00811007AC0A1EB5131120C79E7D176251E53E80E8B361604041340838452020",
INIT_09 => X"C08360820C0912800035F1801630A8260900180C00C8021C800FEE522020A108",
INIT_0A => X"8400F88C166262E940D00D410D62AD02091704024D0A02882192020DA0544043",
INIT_0B => X"4011078510C90D143142430C243042430C24304243042430C24305121A612186",
INIT_0C => X"C08060101000C00401008800F004140009400E4002A0010240000DC3C080002C",
INIT_0D => X"000800100001C07261C51C42390240F050C3C000950008088130040100018000",
INIT_0E => X"00080010003510004000000000000048010002E0100000000800100220100000",
INIT_0F => X"0000014008001550000800000000000400800280100000000800100360100000",
INIT_10 => X"00000000020000080080009410004000000000000044080000D8008000000000",
INIT_11 => X"000005800008000001040168000040000041000100EC00004002214000008000",
INIT_12 => X"00000041003C000008000008200D00001000000208050C000200000000002040",
INIT_13 => X"17000100000000000090000002C8000008000000000060000004480000400000",
INIT_14 => X"8400C00208004844C00800000000528008000000008000000000010040000000",
INIT_15 => X"0100800004030080000C010000A00D1804404912802A261B53104810DB1E0028",
INIT_16 => X"000C030000200C01000020040300800004030000000C03000000040100802004",
INIT_17 => X"008020040100C010000200800004010040300800000020040100C03000020000",
INIT_18 => X"40C700FC0A000280C68A08A950520E964C3269B2C9864D30000C030040100800",
INIT_19 => X"555555555555555555555555555554514514514514526991A199A28A28981451",
INIT_1A => X"41A0D068341A0D068341A0D068341A0D06A351A8D46A351A8D46A35555555555",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF771F60D068341A0D068341A0D0683",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FF087FFDF5508003FEBA087FD54BAAA841540055000000000000000000000000",
INIT_1F => X"F5500003DF455555421EFAAFFD54AAF7D168B45AAAABDF55A2802AA1000002AB",
INIT_20 => X"DFFFAAD1554005D7FD74AAAA840015500002AABA082E954005500021FF5D2EBF",
INIT_21 => X"68BEF080028BFF0855555455500174BAA2AABDE0055517FF555555420AAAA843",
INIT_22 => X"168ABA0055574BA5555554BA5D0400155AAD1554AAF7802AB4500043DF45FFD1",
INIT_23 => X"0400010A2AA955FF55003FE10F7803FEBAFFD5420BA085168A00007BFDE10085",
INIT_24 => X"855555FFAA84001FFAAFBEAB45002A97545F7D1555EF55043DF5555517DEAA5D",
INIT_25 => X"000000000000000000000000000000000000002A82155A2FBFFEBA0800021550",
INIT_26 => X"5BC042AA101D0A28BC7007FFDF45080A3AEAA007BD2482BE84124285C0000000",
INIT_27 => X"004100021FF492AB8F7D1C0438E381451471D7AAFBD0492EBD56DB7DBEAEBFF5",
INIT_28 => X"FED1C5F470AABE8A3AFD7A2DF55400557FD54AABE84001C5550A28ABA1424974",
INIT_29 => X"FB5508043FF55EBD56ABD75D0428BEF005557545490012482B6A0BAE2849557A",
INIT_2A => X"6DA101475FDE10145F68A921C55504924955524AA140E0717DAADB50492EB842",
INIT_2B => X"43AF6D405F78E3A1C2002000BEAA905C755003FE28E3803DEAAEBDF40002557F",
INIT_2C => X"FFFAE821C0A0717D1C5B575FFB6DF425575D7BEFB55002097555FFD5401EF5D0",
INIT_2D => X"784000AA59000000000000000000000000000000000000000000000208017DAA",
INIT_2E => X"A2D57FFFFF7AEBFF55FF8028A00512EAAB45007FFFF55082EA8AAA087FC2010F",
INIT_2F => X"5512AAAA085D04174100800021FF002EA8BEF5D0428ABA595557555AAFBC2000",
INIT_30 => X"00FF802ABAA04552ABFF597FD74BAF7AAA8B45AAFBD54005D7BD54AAF7800215",
INIT_31 => X"5FFAAFBC0000AF843FF5500003FF55AAFD6AB4551002ABEF0055555550004020",
INIT_32 => X"DEB0A2FD5600051537DE005D557DE005D7BE8AA85555400100879560AA592F95",
INIT_33 => X"17545FFD5421FF5D0428BEF0079FCABA598400010F7AA8215555003FEAAAA843",
INIT_34 => X"0000000004001FFAAFBEAA105D2E955FF557BD75EFFBBCD415521FBFDF450004",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000010000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(0),               -- Port A write enable input
DIA(0)   => data_write_a(4),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(4),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(0),               -- Port B write enable input
DIB(0)   => data_write_b(4),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(4),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_5_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50DB0A0791B1B41694368283C81F9996A091A32152007AB36B20E03C040C002",
INIT_01 => X"880015C49830884C446A40000C34C24841280A00084000C8C212892EEA953231",
INIT_02 => X"408F417400B1D9100002171C1FA20171124E6AA00D8633F8CD09DBFBBB972F7C",
INIT_03 => X"88538F0182058082D800C3314722DC08A34084A100C4D7C99208521063D00148",
INIT_04 => X"F45E41AFAF420996B8411CA282F80A9091224800A2C61490363080C8A4000308",
INIT_05 => X"0EA416069640420901A01505C4410020C6E228DC30532839B043289D9C005031",
INIT_06 => X"13992D9AF8C74E92B7B568D19708C038AFFA89F0B9348C9204C389672407EF12",
INIT_07 => X"6255000016053C18162589725146F442222CE6AF844012BE795224458BA4DE0F",
INIT_08 => X"4F3F00503B4AE104B5347230418190420821006016FC18843630D285FC416CB4",
INIT_09 => X"EEA33E700340902C4424C442B0344724066C56C2248130A2D9C185B24A24832B",
INIT_0A => X"315325008348CC40AB570500204462508135D5AA593E043731E9B18A98440137",
INIT_0B => X"E0CD463C5813804E0258E0358E02D8E03D8E0258E03D8E02D8E03447012C701E",
INIT_0C => X"F8DE3C27CA181E5D710664A5F140C14BD32A2E281992940AFAA15C3FC0836310",
INIT_0D => X"F000BE0FC80020130841840308653FF0313FE92C23FB1EECB367C0F3E378F0BC",
INIT_0E => X"F000BE0FCD806FFFAF0AE83080E2AEB2F0F1E01BE53FE1F000BE0FC41BE53FE1",
INIT_0F => X"0231F0BF9E3F02A7FFD63669C0E008C3CB7F041BE1BFE1F000BE0FC41BE1BFE1",
INIT_10 => X"30180309A0F83FE2B87C7D006FFF9F1A7806013879BAA78FC103FF5F1F12F038",
INIT_11 => X"39E9C1DBF8A30C2098DBE2FF7F2320483136F200A822CBACAB9DDEB7F9BC291F",
INIT_12 => X"004C72BEC95FEF64E4090626DF15B7D1C6184131B7980DFFFC03F00003F01FB9",
INIT_13 => X"1DFFFA0A3C0202B8776AE7A7C9CBFFF060703080E29F1B79E9F6427EFE901C0E",
INIT_14 => X"2B716CA5C56620590350ACD3A7D5B7EFAC6DFC8C0312A0024B83F07F3999E9F2",
INIT_15 => X"F0BCAF3BC2F3BC6F0BCEF2BC2F3BC6DBC67C251104A2261253904580207E1C81",
INIT_16 => X"1BCEF0BC2F3BC2F1BCEF0BC6F2BC2F1BCAF1BC6F2BC6F2BCAF1BC2F3BC6F2BCE",
INIT_17 => X"BCEF0BC2F3BC2F1BCAF1BCAF3BC6F0BCEF0BCEF2BC6F2BCAF1BCAF1BC2F3BCAF",
INIT_18 => X"69CFEF73B6FFE7436DB6FD0831518424965B4D2492CB69AF1BCEF0BC6F2BC6F0",
INIT_19 => X"F7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF3EF9FBFBB9E79E7BEBCB7",
INIT_1A => X"DEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDF7DF7DF7D",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF29FDAF77BBDDEEF77BBDDEEF77BBD",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"AAA2802AA10FFFFFDE0008556AABA5D2ABFFEFFF800000000000000000000000",
INIT_1F => X"ABAF7AAA8BFFAA802ABFF087FFDF5508003FEBA087FD54BA0804154005555574",
INIT_20 => X"54AAF7D168B45AAAABDF55AA802AA1000003FEBA00002AABA5D2EBFEBAAAD16A",
INIT_21 => X"3DE005555575EFA2D142145A2FFE8B45FF80001555D2E955FFFFD5421EFAAFFD",
INIT_22 => X"FC00BA5D5568AAAF7AAAAAAAAA802AABA082E954005500021FF5D2EBFF550000",
INIT_23 => X"D5420AAAA843DFFFAAD1554005D7FD74AAAA840014500517FFEF007BEABFF5D7",
INIT_24 => X"2AABDE0055517FF555504154BAA2FBEAA105D2E97410FFD16AAAA5D2ABDEBAFF",
INIT_25 => X"000000000000000000000000000000000000000028BFF0855555455500174BAA",
INIT_26 => X"21E84124285C51574BAB68A2DA00FFFFFFE38085F6FA92552AB8FEFF78000000",
INIT_27 => X"925D2AB8EBABEDB6AA92F7AAA8BC7B68A28BC70075FDF45080A3AEAA007BD248",
INIT_28 => X"5FFFFD1471D7AAFBD0492EBD56DB7DBEAEBFF55BE842AA105D0A38EBA1C0428A",
INIT_29 => X"21FF492AB8F7D1C0438E38145B575EFA2DB45145B6F5EFB6DF78E05145552A92",
INIT_2A => X"7DFC70875EABC7557FC20AA415F68AAAF7AAAAA82BE8A28A9214249740041000",
INIT_2B => X"B6FABA542ABAE2AF7DF470AABE8A3AFD7A2DF55400557FD54AABE84001C55551",
INIT_2C => X"5557545490012482B6A0BAE2849043AFED1C0E10492B6FFEFA105D2A95410FFD",
INIT_2D => X"D2AAABEFFB8000000000000000000000000000000000000000000000428BEF00",
INIT_2E => X"082EA8AAA087FC20105504000AA5955554BAFFAEBDE10F7FBFDEBA007BFDE005",
INIT_2F => X"0512AA8AAA5D0028A005D2AA8ABAF7FBE8A00FFAEAAB45F3AAAAB4500557FF55",
INIT_30 => X"EFFFAA97545552A821EFFBD557555AAFBC2000A2D57FFFFF7AEBFF55FF8028A0",
INIT_31 => X"A005D04174100800021FF002EA8BEF5D0428ABA597FD55FFA2FFD5555FFD57FF",
INIT_32 => X"54AAF7800015551517DF45005168B55557FC0012087FEAABAF7AAAAA10F3AAAA",
INIT_33 => X"FFE005D2A95410F7FFFFEBA5D2EA8ABAFBFFD74BAF7AAA8B45AAFBD54005D7BD",
INIT_34 => X"00000000002ABEF005555555000402000FF802AAAA04452ABFF592E80010FFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000060000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(0),               -- Port A write enable input
DIA(0)   => data_write_a(5),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(5),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(0),               -- Port B write enable input
DIB(0)   => data_write_b(5),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(5),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_6_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10800B0061A01002840002C030028180004003220200403312301C4389B2082",
INIT_01 => X"060009C838394848188160000C42426041000000090800090210090000510200",
INIT_02 => X"00043040009001100000061000018070002408000000000648080000001210E0",
INIT_03 => X"0000800002054081020080801200A0000300008000201184681A0000410C4800",
INIT_04 => X"0808801040000001401048008100022401400002024024053200020089000100",
INIT_05 => X"0240040408402202002000C200400020A50000A0000010010001260808000520",
INIT_06 => X"44000881064500004600000013088002840C240F5048011200010000440C0146",
INIT_07 => X"0241914041FE83E010040110110003040020402A0000003E1000000488000201",
INIT_08 => X"8001BF002C4A01041B112020200110024029006FE09081002004902000012068",
INIT_09 => X"0083FE38A040100281353150ACB645AEF8C01404448000008011061204200108",
INIT_0A => X"3103AD0413424E4014D627C470462200011504420C0A962A2189002881404060",
INIT_0B => X"46C1060C16C96D15B0425B0425B1425B1425B0C25B0C25B1C25B1512D8212D82",
INIT_0C => X"009000140401100601016600A040220203A004480598010248000D0010420C0C",
INIT_0D => X"0000A01033A00013000000000018800F2400091081100C0090A5008200410020",
INIT_0E => X"0000A0103142000000000000000000455D0018100000000000A0103410000000",
INIT_0F => X"000000466800C200000000000000000001A0F4100000000000A0103410000000",
INIT_10 => X"00000000000024094680014200000000000000000041E8002900000000000000",
INIT_11 => X"F000322000000000000D1A000000000000034D240C2000502000000000000000",
INIT_12 => X"000000403F4000000000000068D24000000000001A60F0000000000000002007",
INIT_13 => X"C0000000000000000087C0003014000000000000000025D00008958000000000",
INIT_14 => X"02000000000814C219500150002800101280000000000000000000086670000C",
INIT_15 => X"8120C82208812048120882208892055A0060011280222413130449010301F051",
INIT_16 => X"3200802008320C82200802048320C82200812048320880200812048220880204",
INIT_17 => X"20C83208812048020883204802048120882204812008220C8220081204822088",
INIT_18 => X"79CFF1FE1E9F52ABEF9EFE8150120EC718638E38E30C71C812088220C8120080",
INIT_19 => X"71C71C71C71C71C71C71C71C71C71C71C71C71C71C736D9DBD9BBEFBEFBEBEF1",
INIT_1A => X"CFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FC71C71C71C",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCF29A7F3F9FCFE7F3F9FCFE7F3F9F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000607FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"EFA2FBD54BA5555554BAAAFBC20BA5D7BEAAAAFF800000000000000000000000",
INIT_1F => X"EBA0855421455555574AAA2802AA10FFFFFDE0008556AABA5D2ABFFEFFF843DF",
INIT_20 => X"DF5508003FEBA087FD54BA000415400550428AAAAA84021FF007BD54BAAAD17D",
INIT_21 => X"A8BFFAAD1554BA002A95555A28417400AAFBE8ABAF7FFD54AAAA802ABFF087FF",
INIT_22 => X"BD5545080417555A2D17FE1000003FEBA00002AABA5D2EBFEBAAAD16AABAF7AA",
INIT_23 => X"D5421EFAAFFD54AAF7D168B45AAAABDF55AA802AA100000001EF087FEAA00FFF",
INIT_24 => X"F80001555D2E955FFFF843DEAAA2803DFEF0855401FF082EA8B555D7FC21FFFF",
INIT_25 => X"0000000000000000000000000000000000000055575EFA2D142145A2FFE8B45F",
INIT_26 => X"2552AB8FEFF78E3DFFFAAFFD04AA415B52492B6F5C20825D7FE8A92FF8000000",
INIT_27 => X"EF147BD2482BED57AE921451421555551574BAB68A2DA00FFFFFFE38085F6FA9",
INIT_28 => X"4BAB68A28BC70075FDF45080A3AEAA007BD24821C04124281C0E2DA82BE8E001",
INIT_29 => X"8EBABEDB6AA92F7AAA8BC7B6D5524AA14209557DA28E15400BEF1EFA92FFFFD2",
INIT_2A => X"071FF0071EDA38F7F1D5555000417545B6D178E281C0A38EBA1C0428A925D2AB",
INIT_2B => X"4A8B555C7FC2147F7D1471D7AAFBD0492EBD56DB7DBEAEBFF55BE842AA105D0E",
INIT_2C => X"DB45145B6F5EFB6DF78E05145552A925FFFF8E3DE82BE8E38FFF0851401C7082",
INIT_2D => X"57FE8A00F38000000000000000000000000000000000000000000005B575EFA2",
INIT_2E => X"F7FBFDEBA007BFDE005D2AAABEFFBAABDFEFAAFBC00BA007BC0000FFD5420005",
INIT_2F => X"A592ABFE00F7AA821FF557FC0010F7D168A105D55421455155554BAFFAEBDE10",
INIT_30 => X"10F7D57DE00FFFBC00AAFBAAAAB4500557FF55082EA8AAA087FC20105504000A",
INIT_31 => X"AAA5D0028A005D2AA8ABAF7FBE8A00FFAEAAB45F3D5400BA5504155EFAAAE954",
INIT_32 => X"FF55FF8028A00512E975FF08557FEAAF7D157545080417545F7D56AAAA592AA8",
INIT_33 => X"AABEF005542155000028B555D7FC2145F3D557555AAFBC2000A2D57FFFFF7AEB",
INIT_34 => X"000000007FD55FFA2FFD5555FFD57FFEFFFAA97545552A821EFFBAABDE00F7AA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000048000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(0),               -- Port A write enable input
DIA(0)   => data_write_a(6),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(6),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(0),               -- Port B write enable input
DIB(0)   => data_write_b(6),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(6),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_7_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10844B00482258A2842112C02450418800002300500030B313300C418992002",
INIT_01 => X"020009C23838684D1C20E0000E11424840000000080000080200000000110204",
INIT_02 => X"000520700CA08910000206101180803081144880010400044808000000122160",
INIT_03 => X"000080040305208000008000328080040304008020303194289A000041484800",
INIT_04 => X"08088000000000010000CA008008060441000000028234493410820191000000",
INIT_05 => X"03500404000022020020044000000C208400408000001000984005949C002928",
INIT_06 => X"54000881044500004680000013008002940C24001A4A010200018920646410C7",
INIT_07 => X"22510040400500011204813015012204002040280000013E1000000488000201",
INIT_08 => X"9001A0602C4A01051B132820208001024069004008908002120851420001226A",
INIT_09 => X"01100020A2401008A20404E08200A05000A4264640800022C8198C4E05200018",
INIT_0A => X"20002000024040400050450440C48A0041140C420B0904208800904286000008",
INIT_0B => X"50822002120D2134800648006480064800648106481064810648193240432404",
INIT_0C => X"284A142288042A5C24202451505E00A621A5220A8091444040188C001B41210A",
INIT_0D => X"00F001F021141A12004104020810B000100000000109064C80010050A3285194",
INIT_0E => X"00F001F027420000400004C3201C514408081C1014800000F001F02810148000",
INIT_0F => X"E00E0E404100E200040900000B0380383480C81014800000F001F02810148000",
INIT_10 => X"4160C0301D07001D0402034200004000019860078641004039000180400002C0",
INIT_11 => X"08103BA0104810C8462416E8040446120C890814600010512000000080028400",
INIT_12 => X"98038D4030DD008088C2419120B740209021908C4846FC000200030F000FE006",
INIT_13 => X"DD000100411C81078884204035DC00201804C3201C60A408100DD58010440130",
INIT_14 => X"412024202211148019064200402A32901A8000B2048902C0807C0E00C448100D",
INIT_15 => X"50942509425194651946519465894619421421102000269243854D8002000250",
INIT_16 => X"19465194E50942509425094E51946519465094A50942509425194E5194651942",
INIT_17 => X"9425094251946539465094250946539465194250942509465194650942509425",
INIT_18 => X"0000000000000000000000080150890820800041041000052942509465194653",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF21E6C000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"AAF7D5575455D557DFEF002AAAB55002E820AAAA800000000000000000000000",
INIT_1F => X"B55007FD74AAAA843DFEFA2FBD54BA5555554BAAAFBC20BA5D7BEAAAAFFFBC00",
INIT_20 => X"AA10FFFFFDE0008556AABA5D2ABFFEFFFAAAAAAAF7D57FFEFF7D555555A2AEAA",
INIT_21 => X"42145552ABDFEFFFAA801EFFFFBFDF550000175555504175450055574AAA2802",
INIT_22 => X"A975EF00003DF55555168A00000428AAAAA84021FF007BD54BAAAD17DEBA0855",
INIT_23 => X"802ABFF087FFDF5508003FEBA087FD54BA000415400557BD74BAFFD140000082",
INIT_24 => X"AFBE8ABAF7FFD54AAAAAEA8ABA55557FEAAA2843FF55A2AEA8B55AAAABDEAAFF",
INIT_25 => X"0000000000000000000000000000000000000051554BA002A95555A28417400A",
INIT_26 => X"25D7FE8A92FFFFC70BAE3D155555415178FD7082EAAB550820870BAAA8000000",
INIT_27 => X"FFEBD55557DBEA4AFB550871D7482AA8E3DFFFAAFFD04AA415B52492B6F5C208",
INIT_28 => X"5550051574BAB68A2DA00FFFFFFE38085F6FA92552AB8FEFF7A0ADABAEBD578F",
INIT_29 => X"2482BED57AE921451421555524BDFD7FFA4801D7F7F5FDF55000E17545410E17",
INIT_2A => X"D2482E3D1450381C20905EF08003AF55415F6DA38080E2DA82BE8E001EF147BD",
INIT_2B => X"AAFB55ABA0BDE02EB8A28BC70075FDF45080A3AEAA007BD24821C04124281C7B",
INIT_2C => X"209557DA28E15400BEF1EFA92FFFFD24BAB6A4A8A82495F78E92AA843DF45BEA",
INIT_2D => X"800174BAA680000000000000000000000000000000000000000000055524AA14",
INIT_2E => X"007BC0000FFD542000557FE8A00F3FFD54BAAAD15754508556AB45002AA8B450",
INIT_2F => X"FFB803DEAAAAD56ABEFAAD5575EFF7803DF45085557410AEAABDFEFAAFBC00BA",
INIT_30 => X"55082E97555002E955550C55554BAFFAEBDE10F7FBFDEBA007BFDE005D2AAABE",
INIT_31 => X"E00F7AA821FF557FC0010F7D168A105D554214551003FF45FF8400145FFD57FF",
INIT_32 => X"20105504000AA597FC2010A2D1554AA5500021EF000028B55087BFDEBA042ABF",
INIT_33 => X"E8A00A2803FF45F7AABDF55AA843FE10AEAAAAB4500557FF55082EA8AAA087FC",
INIT_34 => X"0000000055400BA5504155EFAAAE95410F7D57DE00FFFBC00AAFB8028A00007F",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000007FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(0),               -- Port A write enable input
DIA(0)   => data_write_a(7),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(7),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(0),               -- Port B write enable input
DIB(0)   => data_write_b(7),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(7),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_8_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000B0000040042840002C0000001800000070000000033022000000000086",
INIT_01 => X"000009C21838284D1C2160000E12426840000000180800080200080040510200",
INIT_02 => X"0001004000900110000006100080003000240800014400004808000000122160",
INIT_03 => X"00008000020440810002A0801010A0044300000000200086011A000040404800",
INIT_04 => X"8000801000020401400040408108022029400000124004041200000089000100",
INIT_05 => X"02080424085022020000040200480020850010A0002010010120060800040400",
INIT_06 => X"50000880006500000680000011008006840C200018C1010200018920E0640102",
INIT_07 => X"426000404005000112048130150120240020400A0000013E1000000488000010",
INIT_08 => X"220100402C42010413110020200100024029004000A200002004902200012141",
INIT_09 => X"0000000080400008010410A2940A45240040140440800022C8388E1200A00008",
INIT_0A => X"00420100020048405000070440C0000001140412090000000021002081000048",
INIT_0B => X"0000000800000100011000010000100001000010000100001000010000880008",
INIT_0C => X"001000040001100008012008004020102180800804802000C0080D00100A0008",
INIT_0D => X"0FF0000002200A1200410402080080003000091085100C008124008000400020",
INIT_0E => X"0FF000000140000040F517CF600000000104081010001E0FF00000001010001E",
INIT_0F => X"E000000000804200000809963F1F80000000001010001E0FF00000001010001E",
INIT_10 => X"CFE7C0F00000000000810140000040E587F9E000000008100900008000ED0FC7",
INIT_11 => X"00021040030C73D80000021000585F3600000020240020102000000802419660",
INIT_12 => X"F80000000042000B0BD6C0000010800618E7B000000C000003F80FFF00000000",
INIT_13 => X"800005D5C3FD800000000008180000078A8FCF600000000002028001006AA3F1",
INIT_14 => X"020000000008808219002100100C000041120370DCAD1FC18000000000000202",
INIT_15 => X"8020080200812048120481204812055A04604930A02026934215410102000110",
INIT_16 => X"0200802008020080200802048120481204812048120481204802008020080200",
INIT_17 => X"2008020081204812048120481200802008020080200802048120481204812048",
INIT_18 => X"414A87D78AF42143CEBAC88151120A0000000000000000081204812008020080",
INIT_19 => X"F3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF7E799B1BEB65B65948051",
INIT_1A => X"C3E9F0FA7C3E9F0FA7C3E9F0FA7C3E9F0F87C3E1F0F87C3E1F0F87CF3CF3CF3C",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF1B5DA9F0FA7C3E9F0FA7C3E9F0FA7",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"0000043DF55087BC01EF007FD75FFFF84000AAFF800000000000000000000000",
INIT_1F => X"E10A28028AAAAAFBC00AAF7D5575455D557DFEF002AAAB55002E820AAAA84000",
INIT_20 => X"54BA5555554BAAAFBC20BA5D7BEAAAAFFAA95545552ABFE00087BC00AA082EBF",
INIT_21 => X"D74AAAAD57FF45002A975FF007BE8BFFA2FBFFFFFAAD5400AAFF843DFEFA2FBD",
INIT_22 => X"BE8A00082A97410F7D5555EFAAAAAAAAAF7D57FFEFF7D555555A2AEAAB55007F",
INIT_23 => X"55574AAA2802AA10FFFFFDE0008556AABA5D2ABFFEFFFAA82000555555545AAF",
INIT_24 => X"00017555550417545000015545087BC2010AAD54014500516ABFFA2AABDF4500",
INIT_25 => X"000000000000000000000000000000000000002ABDFEFFFAA801EFFFFBFDF550",
INIT_26 => X"50820870BAAA8407000140038F450075C71FF087BD75D7FF84050BAEB8000000",
INIT_27 => X"10007FC50BA002ABFE00AA8A2AABABEFFC70BAE3D155555415178FD7082EAAB5",
INIT_28 => X"082EB8E3DFFFAAFFD04AA415B52492B6F5C20825D7FE8A92FFA497545552AB8E",
INIT_29 => X"557DBEA4AFB550871D7482AAD17DF451C24955EF0875EFBD7B6F1FFFC7BEDB45",
INIT_2A => X"87000415B5057DAAFBE8A10082092410EBD5505EFB6A0ADABAEBD578FFFEBD55",
INIT_2B => X"B6ABC7B6AABFFED0051574BAB68A2DA00FFFFFFE38085F6FA92552AB8FEFF7AA",
INIT_2C => X"A4801D7F7F5FDF55000E17545410E17555000E17545007BC0000BED14217D005",
INIT_2D => X"784174AAA280000000000000000000000000000000000000000000024BDFD7FF",
INIT_2E => X"08556AB45002AA8B450800174BAA684174105D042AB550055555FF007BD7555F",
INIT_2F => X"0F384175555D2EA8A00087BD74BA082EBDE10AAAEA8ABAF7FFD54BAAAD157545",
INIT_30 => X"55FFD57DF55FFFBD5400A2AABDFEFAAFBC00BA007BC0000FFD542000557FE8A0",
INIT_31 => X"EAAAAD56ABEFAAD5575EFF7803DF45085557410AED17FF455D04155FF00557DF",
INIT_32 => X"DE005D2AAABEFFBAE97410087BC21EFA2FFEAA00000002010A2D5421FFFF803D",
INIT_33 => X"C0010FFD1401EF087FE8B55FFAEBDFEF0855554BAFFAEBDE10F7FBFDEBA007BF",
INIT_34 => X"00000000003FF45FF8400145FFD57FF55082E97555002E955550C2E95555087B",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000020000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(1),               -- Port A write enable input
DIA(0)   => data_write_a(8),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(8),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(1),               -- Port B write enable input
DIB(0)   => data_write_b(8),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(8),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_9_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00018248A2840112C00002C18000002300500030B3132000400812002",
INIT_01 => X"A140098218302849180060000C004240413C0A61590001D90213C90008510204",
INIT_02 => X"102008700CB089100002061031285074810448800104008048080080001210E2",
INIT_03 => X"00008015074608840390A0040040800203140000A00010800408108448020042",
INIT_04 => X"082080400004A00100000100840602020100000002C2344156108201811801C0",
INIT_05 => X"0200048480011502049500280020CC2084000080008010019161249C9C002188",
INIT_06 => X"70000881004500004E01020411D08000940C00001800010200018B20206C0102",
INIT_07 => X"EA70C0040005000312048130150100040020404A0000017E10408104C8000110",
INIT_08 => X"000000402C220104131004202081120050A5104000A204617201D10801002000",
INIT_09 => X"000800002F4924003085E51420A0100400641E4E40800022C8088C1220200908",
INIT_0A => X"20102000024040484028450001648C2229150400080244000401900284000440",
INIT_0B => X"0880110901081110411204112040120411204012041120401204111020090208",
INIT_0C => X"685B34A688841A5C21200101A01A0004009024028004044248404D00104B2100",
INIT_0D => X"0000A01000000213000000000000B0001000010000190E44802002D1A168D0B4",
INIT_0E => X"0000A010014000000000000000000040500008100400000000A0100410040000",
INIT_0F => X"0000004608004200040000000000000001A004100080000000A0100410008000",
INIT_10 => X"00000000000024080000014000000000000000000040A0000900010000000000",
INIT_11 => X"300013E010000000000D00F804000000000340000C0000102000000080000000",
INIT_12 => X"00000040091F0000800000006807C000800000001A0CFC000000000000002001",
INIT_13 => X"DD000000000000000082C00019DC002000000000000021500006D58010000000",
INIT_14 => X"03206420000000C019502050000C32901A800080000000000000000860100006",
INIT_15 => X"D1B46D1B46D0B42D0B42D0B42D8B424342342832002A24921082158802001011",
INIT_16 => X"0B42D0B42D0B42D0B42D0B46D1B46D1B46D1B46D1B46D1B46D1B46D1B46D1B46",
INIT_17 => X"B42D0B42D1B46D1B46D1B46D1B46D1B46D1B46D1B46D1B42D0B42D0B42D0B42D",
INIT_18 => X"89999E91BCD1512B871C4A0100000000000000000000000D0B42D0B42D0B42D0",
INIT_19 => X"A28A28A28A28A28A28A28A28A28A29A69A69A69A69A51C200807249041202AE6",
INIT_1A => X"8349A4D068341A0D269341A0D269341A0D068341A0D068341A0D068A28A28A28",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF2DA921A0D269341A0D068349A4D06",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"45A280154BA5555401EFFFD5421EFA2FFFFF555D000000000000000000000000",
INIT_1F => X"5EF00557DF555D040000000043DF55087BC01EF007FD75FFFF84000AAFFD57DF",
INIT_20 => X"75455D557DFEF002AAAB55002E820AAAA843DFEF00517DEBA007BFDFEFFFD157",
INIT_21 => X"28AAAAAAABDF45F7803FFEF555568AAAF7802AA00FFFBD7555087BC00AAF7D55",
INIT_22 => X"BD54BA550417400085155555082A95545552ABFE00087BC00AA082EBFE10A280",
INIT_23 => X"043DFEFA2FBD54BA5555554BAAAFBC20BA5D7BEAAAAFFFBC00AA552E95545087",
INIT_24 => X"2FBFFFFFAAD5400AAFF8402000A2FFFDF555D7BE8BFF5D51575EFA280175555D",
INIT_25 => X"00000000000000000000000000000000000000557FF45002A975FF007BE8BFFA",
INIT_26 => X"7FF84050BAEBDF78F45B68010482415B471C7E3DF451EFBEFBFAF45490000000",
INIT_27 => X"82007FFAFEFE3DB505EF1C5B7AF45490407000140038F450075C71FF087BD75D",
INIT_28 => X"5451C7FC70BAE3D155555415178FD7082EAAB550820870BAAA8438FFF00517DE",
INIT_29 => X"50BA002ABFE00AA8A2AABABEAEB8F45F78A3DFD741516DAAAE38E2DA28EBFFD5",
INIT_2A => X"C20BA5D2E905550071D54825D0A1543808515756D1C2497545552AB8E10007FC",
INIT_2B => X"5505FFBE801256D490E3DFFFAAFFD04AA415B52492B6F5C20825D7FE8A92FFFF",
INIT_2C => X"24955EF0875EFBD7B6F1FFFC7BEDB45082EB8002000AAFFFDF6D417FEABEF5D5",
INIT_2D => X"7FBE8B5500000000000000000000000000000000000000000000000517DF451C",
INIT_2E => X"0055555FF007BD7555F784174AAA2FBEAB45F78402010007BD5545AAFFD55EFF",
INIT_2F => X"AA68028BEF00517FE10007BE8BFFAAFFC01FF557FE8B550004174105D042AB55",
INIT_30 => X"AAAAAEBFEAAAAFFD5545557FD54BAAAD15754508556AB45002AA8B450800174B",
INIT_31 => X"5555D2EA8A00087BD74BA082EBDE10AAAEA8ABAF7AAAAB45F7AEBFF4508557FE",
INIT_32 => X"2000557FE8A00F3FFC00BA552E80145005557400552A954BA0051575EF550417",
INIT_33 => X"FDFFF007FE8BFF5551401EFF784021FF002ABDFEFAAFBC00BA007BC0000FFD54",
INIT_34 => X"00000000517FF455D04155FF00557DF55FFD57DF55FFFBD5400A28400010A2FB",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000040000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(1),               -- Port A write enable input
DIA(0)   => data_write_a(9),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(9),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(1),               -- Port B write enable input
DIB(0)   => data_write_b(9),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(9),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_10_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00018248A2840112C00002C18000202300500030B3132000400992006",
INIT_01 => X"A140098218302849180060000C00424040000000080000080200090008510204",
INIT_02 => X"102100400C8001100000061000A8503401044880010400004808000000122160",
INIT_03 => X"000080150746088401908000100080020304000020201080001A108448404842",
INIT_04 => X"800080400004A001000040008406020201000000020004401000000180180080",
INIT_05 => X"02000484800133020495040800208C20A4000080000010000001249010042008",
INIT_06 => X"50000881004500004681020411808000940C20001800010200018920206C0102",
INIT_07 => X"024084044005000112048130150120040020400A0000013E10408104C8000010",
INIT_08 => X"000100402C020105131100200000124250A51040088084614001110801012000",
INIT_09 => X"00080082CD09240820800000000000040000180840800022C8088C1220200108",
INIT_0A => X"841201000200484910000F050560262229140402080200A00402000484140400",
INIT_0B => X"0010118900080010000200102001020000200002001020010200001000010008",
INIT_0C => X"408120900404004821202001F05E00040180260A8080044240004C0010800228",
INIT_0D => X"0000A01000000813004104020800800030000800010008088124020102008100",
INIT_0E => X"0000A010014000004000000000000040500008101480000000A0100410148000",
INIT_0F => X"0000004608004200040900000000000001A004101480000000A0100410148000",
INIT_10 => X"00000000000024080000014000004000000000000040A0000900018040000000",
INIT_11 => X"3800100010480000000D00000404400000034000282000102000000080028000",
INIT_12 => X"00000040090000808800000068000020900000001A0000000200000000002001",
INIT_13 => X"80000100000000000082E0001000002018000000000021580000800010440000",
INIT_14 => X"00004000000004C0195000500008000000000082008000000000000860180000",
INIT_15 => X"0100401004010040100401004090055804404110802A24921317580802001011",
INIT_16 => X"0000000000000000000000040100401004010040100401004010040100401004",
INIT_17 => X"0040100400000000000000000000000000000000000000000000000000000000",
INIT_18 => X"215281FC1A72E2486AAA40A85052020000000000000000001004010040100401",
INIT_19 => X"51451451451451451451451451451451451451451452AA83330A8A28A29EA8D1",
INIT_1A => X"5CA6532994CA6532B95CAE572994CA6532994CA6532994CA6532994514514514",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF31CE2E572994CA6532994CAE572B9",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"10AAFBE8AAAA2D540000F7D57DF55A2AABFFEF08000000000000000000000000",
INIT_1F => X"F45FFFBC2010AAD57DF45A280154BA5555401EFFFD5421EFA2FFFFF555D003FE",
INIT_20 => X"DF55087BC01EF007FD75FFFF84000AAFF8002155AAFFE8B45AAD540000087FFD",
INIT_21 => X"7DF555D517FEBA082A801EFF7FBD5400FFD568B555D00155EF08040000000043",
INIT_22 => X"BFDE00A2FBC0145005168A10AA843DFEF00517DEBA007BFDFEFFFD1575EF0055",
INIT_23 => X"7BC00AAF7D5575455D557DFEF002AAAB55002E820AAAA803FEBA082AAAAAAF7F",
INIT_24 => X"7802AA00FFFBD7555082E82155FFAEAAB55AAD568B455D00154BAFFFBD75EF5D",
INIT_25 => X"000000000000000000000000000000000000002ABDF45F7803FFEF555568AAAF",
INIT_26 => X"FBEFBFAF4549003DE10BEF5EDAAAAAD547038EBD57DF7DA2AEB8FC7000000000",
INIT_27 => X"6DAADF470280075FFF45E3F1C7038A2DF78F45B68010482415B471C7E3DF451E",
INIT_28 => X"5C7000407000140038F450075C71FF087BD75D7FF84050BAEB8002155BEF5EDB",
INIT_29 => X"AFEFE3DB505EF1C5B7AF45495B7DEAA0824851EFEBFBD2410EBD168B7D410A17",
INIT_2A => X"38EAA0824A8AAAEBF5FAE28AAF1C2155005F68A10A28438FFF00517DE82007FF",
INIT_2B => X"4104AAF7F1D75EF557FC70BAE3D155555415178FD7082EAAB550820870BAAA80",
INIT_2C => X"8A3DFD741516DAAAE38E2DA28EBFFD55451C2087155EBA4A8B7DAADF68B7D410",
INIT_2D => X"2AEAAB55000000000000000000000000000000000000000000000002EB8F45F7",
INIT_2E => X"007BD5545AAFFD55EFF7FBE8B5500043FE00F7D17FEBAA2D5574BAAAD17DFEFA",
INIT_2F => X"AA28002155FFD17FFFFA2FBD74BA00557FF45A2D5554AAA2FBEAB45F78402010",
INIT_30 => X"00AAD16ABFF002A975450004174105D042AB550055555FF007BD7555F784174A",
INIT_31 => X"BEF00517FE10007BE8BFFAAFFC01FF557FE8B55007FFDEAA0004175FFA2FBC20",
INIT_32 => X"8B450800174BAA68428AAA08042AABAAAD56AABAAAD140155087FEAA10A28028",
INIT_33 => X"2ABEFAAFBE8BFF0004020AAFFD5555EF557FD54BAAAD15754508556AB45002AA",
INIT_34 => X"000000002AAAB45F7AEBFF4508557FEAAAAAEBFEAAAAFFD5545550015555A284",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000047FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(1),               -- Port A write enable input
DIA(0)   => data_write_a(10),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(10),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(1),               -- Port B write enable input
DIB(0)   => data_write_b(10),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(10),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_11_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10180B05A0010402840602C2D001019000000300000000330A20080EC180002",
INIT_01 => X"AB400984B830084C1820E0000C36424840000000080000088200000802112220",
INIT_02 => X"102A68440080011000000618062AD03502640800010410424908136019920868",
INIT_03 => X"001282118644C88481908001106088022300000080F4925CDC9A10844A9A4842",
INIT_04 => X"401280480004A1011000418084460002E12000000200040010000040A8000000",
INIT_05 => X"0FC8048484011502059511488020802084400888001110000000050000005400",
INIT_06 => X"1011088AE24500001631024511C08004A70AA40008B90D0200018B60A0650D45",
INIT_07 => X"020011005405000910040150110041040024400D800002BE18408104C9205908",
INIT_08 => X"89390040280241041D175820000001020061004004800567403512A801014C46",
INIT_09 => X"050800E20D09A424C5840400808000040680180840800022D8288E946CA00833",
INIT_0A => X"85002000024040410A000D0504408C32E915D9C208050084840201A099100400",
INIT_0B => X"B01011934A005101431CA821CA831CA821CA831CA831CA821CA83165410E5410",
INIT_0C => X"00010080028000010402214850444091019B02080885200042A9CC001000003A",
INIT_0D => X"5A5018C5A0A00812004104020808B00030000808024008008325820000000000",
INIT_0E => X"5A5018C5AB0062C38A4DB680A0D8241500D5761B011986695014A96E1A811986",
INIT_0F => X"42056A289A1BB2078A922DA2A8B180A2600AAE1A811986695014A96E1B011986",
INIT_10 => X"05AA429189B60AC43C6C7F0272C3841DB528802CAB18468F4101621B1BAC8455",
INIT_11 => X"C003104289A668B8CAB270106338317A3D94392020224ACDE215883078681B5C",
INIT_12 => X"804B020A06020C67061BC785938085134CD551BCA1C90006C0C2958502861120",
INIT_13 => X"80819A5539D503336D61056ABA006282806CA64090B89E015AAA880E48382EB8",
INIT_14 => X"40000000E808989003066E03513E41470126C6284B2D20410AB4503089C00A82",
INIT_15 => X"0000000000000000000000000000041800400110200026124202500802000800",
INIT_16 => X"1004010040100401004010000000000000000000000000000000000000000000",
INIT_17 => X"0040100401004010040100401004010040100401004010040100401004010040",
INIT_18 => X"C110083018162148420840280050800000000000000000001004010040100401",
INIT_19 => X"000000000000000000000000000001041041041041003882928E0000000AA0C4",
INIT_1A => X"0000000000008040000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3E0FC000000000000020100000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"EFAA842ABEFA280155EFFFFBC01EF08554000055000000000000000000000000",
INIT_1F => X"F4508514000000003FE10AAFBE8AAAA2D540000F7D57DF55A2AABFFEF0804155",
INIT_20 => X"54BA5555401EFFFD5421EFA2FFFFF555D51575FFA2FFD75FF550015400FFFBFF",
INIT_21 => X"C2010AAD568AAAAAD142145FF80155EF0051555FF0804155FFF7D57DF45A2801",
INIT_22 => X"01540008514215555003DFFFA28002155AAFFE8B45AAD540000087FFDF45FFFB",
INIT_23 => X"040000000043DF55087BC01EF007FD75FFFF84000AAFF802ABFFA2AABFE10080",
INIT_24 => X"FD568B555D00155EF085168B45085142010FFAE800AA5D7BFDF45F7FFEAA0000",
INIT_25 => X"00000000000000000000000000000000000000517FEBA082A801EFF7FBD5400F",
INIT_26 => X"DA2AEB8FC70000175EFB6802DBC7BE8A155EFE3FBC71FF145B42038550000000",
INIT_27 => X"EF550E15400E3F1FFF7D085B420381C003DE10BEF5EDAAAAAD547038EBD57DF7",
INIT_28 => X"5C7F7DF78F45B68010482415B471C7E3DF451EFBEFBFAF45495F575FFBEF5D05",
INIT_29 => X"70280075FFF45E3F1C7038A2DB68ABAB6D145145FF84155D7085B555C7140410",
INIT_2A => X"28BEFBEA4BDE28140A1543800514515549003FFC7BE8002155BEF5EDB6DAADF4",
INIT_2B => X"FFFF7DE3F1EFA10140407000140038F450075C71FF087BD75D7FF84050BAEB84",
INIT_2C => X"24851EFEBFBD2410EBD168B7D410A175C7005B6DB55145140000FFAE85082417",
INIT_2D => X"57BC20AA5D0000000000000000000000000000000000000000000005B7DEAA08",
INIT_2E => X"A2D5574BAAAD17DFEFA2AEAAB550004175FFF7803DF45FFAE955EFAAFBD55EF5",
INIT_2F => X"5007FD75FFF7D5401EF5D2E97410AAD17DFEF007FC20AA5D043FE00F7D17FEBA",
INIT_30 => X"55007FD5545550400145FFFBEAB45F78402010007BD5545AAFFD55EFF7FBE8B5",
INIT_31 => X"155FFD17FFFFA2FBD74BA00557FF45A2D5554AAA2FBEAAAAFFD555545FF80155",
INIT_32 => X"7555F784174AAA2842ABEFFF803DEAA5D2E974AA00515754500003FF55FF8002",
INIT_33 => X"40000FFAE97410007BFFFFFA2D57FE105D04174105D042AB550055555FF007BD",
INIT_34 => X"000000007FFDEAA0004175FFA2FBC2000AAD16ABFF002A97545007FFFF455555",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000040000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(1),               -- Port A write enable input
DIA(0)   => data_write_a(11),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(11),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(1),               -- Port B write enable input
DIB(0)   => data_write_b(11),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(11),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_12_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50080B01BC002006940202C0DE041196A83183000000023322287E0FC000006",
INIT_01 => X"0E000C068000E04D40238000001702484000000008000008820009280A553231",
INIT_02 => X"400B71440C8001100000171C0283813013766A800586235ECC09C8423B962966",
INIT_03 => X"CC618E048306E082000081000040900003548421A080025EDF08421042DC0108",
INIT_04 => X"00028020000000812000012080080000E100001002000448100000C1BC18008C",
INIT_05 => X"0FF8060610000402010015E100004C2084800090000310000000079010007C19",
INIT_06 => X"33992D98DEC74A003EA468D01510C03E8F580C800A3F018200418927E0668645",
INIT_07 => X"0204000406050013142409121142F746222EE2498000007E111204058B84C50C",
INIT_08 => X"E826A0602902A10491165C200000820018A5104010C01086003C13E000004EDF",
INIT_09 => X"023000000000000867000000000000040000600060801022C9F88D244FA40133",
INIT_0A => X"00100000820040482B28050001600010C13499F01B334015980001E09F000000",
INIT_0B => X"B80460124F16F06BC20CBC30CBC20CBC20CBC30CBC20CBC20CBC3065E1865E10",
INIT_0C => X"00000000029D204B7C0382FD0100F3F9F80FA0200E0BF40063F99C0010000012",
INIT_0D => X"93900F6EE230301208008001007A80001100002002801000A042000000000000",
INIT_0E => X"93900F6EEC421392C96B1237E0D8BD9629F97E0B348EDAC3900F6EFA0B158EDA",
INIT_0F => X"622DBC31D73F6006A5891533EF9500EAE64BCA0B158EDAC3900F6EFA0B348EDA",
INIT_10 => X"C2B083798D341B10DEFE14400392C74CAEAD412EDD2B4FCFF812A383430C669E",
INIT_11 => X"49FAB442994B3238D4E2FB104636652E19B8BA30C022DAD8C100CA39E8CEBE66",
INIT_12 => X"30469392526208C6CC95C33717D88532966471A9C5DD00B12728D5360234D62A",
INIT_13 => X"828C4999AF580395542D27CDBA0020F0FABAC800DA550C29F36A8A2554E48A64",
INIT_14 => X"40000000873FB80B8A00EF03F56CC12B416A51B60585A5C28895962502E9F36A",
INIT_15 => X"0000000000000000000000000000008000000410802A26924010000002000EE0",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"28C1111026C152A121960A884042020000000000000000000000000000000000",
INIT_19 => X"2082082082082082082082082082092492492492492400200005A8A28A200A37",
INIT_1A => X"964B2592C964B2592C964B2592C964B2590C86432190C86432190C8208208208",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF400FEB2592C964B2592C964B2592C",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FF00042ABEFFF8400010082EAABFF55002ABEF08000000000000000000000000",
INIT_1F => X"BEFFFFBD54000004155EFAA842ABEFA280155EFFFFBC01EF0855400005555421",
INIT_20 => X"8AAAA2D540000F7D57DF55A2AABFFEF08556AA10000028AAAFFD15541000002A",
INIT_21 => X"40000005168AAA087BFFFFF5D04001FF00041554555557FE005D003FE10AAFBE",
INIT_22 => X"1555FF082AA8B55F7AEA8BEF5551575FFA2FFD75FF550015400FFFBFFF450851",
INIT_23 => X"D57DF45A280154BA5555401EFFFD5421EFA2FFFFF555D0000145082E955FF085",
INIT_24 => X"051555FF0804155FFF7842AA100000020BAAA801541055042ABEFFFFBD5410AA",
INIT_25 => X"000000000000000000000000000000000000005568AAAAAD142145FF80155EF0",
INIT_26 => X"F145B42038555F401D71C0A2DBC7EB80000280824ADBD7490E28BEF080000000",
INIT_27 => X"82FFDB5243800002FBD7EBFBD24101C00175EFB6802DBC7BE8A155EFE3FBC71F",
INIT_28 => X"E1041003DE10BEF5EDAAAAAD547038EBD57DF7DA2AEB8FC7005F6AA381C0A2DA",
INIT_29 => X"5400E3F1FFF7D085B420381C5B6AA82147FF8FEF410E001FF000E17555555B7A",
INIT_2A => X"0017D142E905EF1451525C7082AADB45F7AEA8BEF555F575FFBEF5D05EF550E1",
INIT_2B => X"02FBEFEBFBD2410AADF78F45B68010482415B471C7E3DF451EFBEFBFAF454900",
INIT_2C => X"D145145FF84155D7085B555C71404105C7F7842FA381C0A00082AA8A10410410",
INIT_2D => X"02AA8BEF000000000000000000000000000000000000000000000005B68ABAB6",
INIT_2E => X"FFAE955EFAAFBD55EF557BC20AA5D7BC01555D2EBFF55A284000AA08003FF550",
INIT_2F => X"5007BE8AAA5D2EBDE00FFFFC00AA08003FF55A2FBC00105D04175FFF7803DF45",
INIT_30 => X"FF082A97555557FE8A0000043FE00F7D17FEBAA2D5574BAAAD17DFEFA2AEAAB5",
INIT_31 => X"5FFF7D5401EF5D2E97410AAD17DFEF007FC20AA5D7BE8A005D7FEABFF002E821",
INIT_32 => X"55EFF7FBE8B550004001FF5D2A801EF5D5142145082EBFF55F7AAAABEF5D7FD7",
INIT_33 => X"82010A2AA8000008043FFFFA2FBC2010A2FBEAB45F78402010007BD5545AAFFD",
INIT_34 => X"000000007BEAAAAFFD555545FF8015555007FD5545550400145FF843DEAA552A",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000007FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(1),               -- Port A write enable input
DIA(0)   => data_write_a(12),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(12),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(1),               -- Port B write enable input
DIB(0)   => data_write_b(12),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(12),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_13_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10110A0441812402840402822007818000E00700000000330A3000000008042",
INIT_01 => X"A1400986B830E84D182260000C1042484001000008220008A20019080A510200",
INIT_02 => X"10A108600C9141100000C6180CA85035010E4880010431004908135980122D60",
INIT_03 => X"0013881507460886C190832175809C02030400002020124C441A108468424842",
INIT_04 => X"203080680204A0113801D600864E0C96C12000008244244052200201801802C0",
INIT_05 => X"030004849601110204950409C0208C2084E0009C0000100120A00C9918002098",
INIT_06 => X"10000882804544921681428591908000AF28A8002BC00D020003896020658FC4",
INIT_07 => X"CA20400450050009100501501102E0042020448D0000023E10408144C800D800",
INIT_08 => X"1D2B00402B220104B53100200001020218A5104016CC1C616401910801010100",
INIT_09 => X"050800404D49A42EB08000000000000406481C8C408000A2D8088D1820200B00",
INIT_0A => X"0010000002004048AA08050401604462E9144002090740148441200484000500",
INIT_0B => X"000A112100000000010000000001000000000000001000000000000000800000",
INIT_0C => X"509528954404144C200425010040000001B020081094040072005C0030864208",
INIT_0D => X"1C10B3831034081200000000000430003000206822F20CA8826AC2A14250A128",
INIT_0E => X"1C10B383110218CB0E54C2EA404A4F03D404A41AA5B7344C10B383081BA4B734",
INIT_0F => X"8001CE3E20A5B284ED1132909C72885A2B2C381BA4B7344C10B383081AA5B734",
INIT_10 => X"AC3CC0C0B8182597A801610218CB0C3548B3A008E730A01AB113A5524E6ACA67",
INIT_11 => X"A151EC5952E44128CA194517354C180A3C066430202021252991C22C99731014",
INIT_12 => X"1804C8A0ADA2E6A983014780CA28B2A5C8825194332B018A444AEA2701288A15",
INIT_13 => X"02D09852745F80112C428562EE0353635232D50048A411C158BB0A7910142C77",
INIT_14 => X"4240480068001C9B9150A0000297046E4023F8BE8E3E1E0109472C3EB50158BB",
INIT_15 => X"A1284A1284A1284A1284A1284A12851A84284110406A26924302590806000110",
INIT_16 => X"1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284",
INIT_17 => X"284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A",
INIT_18 => X"7DDFE7EFBEFFE7D3EFBEFC48A0550000000000000000000A1284A1284A1284A1",
INIT_19 => X"D75D75D75D75D75D75D75D75D75D75D75D75D75D75D7EFBFBFBBAAAAAABEFDF7",
INIT_1A => X"5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5D75D75D75",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000FEFD7EBF5FAFD7EBF5FAFD7EBF",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"AA5D043FFFFAAAABDEAA557BFDE00FFD140155F7800000000000000000000000",
INIT_1F => X"400AAD540155A2D5421FF00042ABEFFF8400010082EAABFF55002ABEF08556AA",
INIT_20 => X"ABEFA280155EFFFFBC01EF08554000055043DEBAF7843FFFFF7AABDF55A2AA97",
INIT_21 => X"D5400005568A1055043DEBAAAFFE8B45557FD7410552EAAABAAA84155EFAA842",
INIT_22 => X"FE8ABAAA8428A00087BD7555FFD56AA10000028AAAFFD15541000002ABEFFFFB",
INIT_23 => X"803FE10AAFBE8AAAA2D540000F7D57DF55A2AABFFEF085557545FFD17DEBAA2F",
INIT_24 => X"0041554555557FE005D0000155557BEAABA5D2ABDF450851420AA5D7FD5555A2",
INIT_25 => X"000000000000000000000000000000000000005168AAA087BFFFFF5D04001FF0",
INIT_26 => X"7490E28BEF08516DA82410A3FFD7AAA4B8E824971F8E38E3DF45155EB8000000",
INIT_27 => X"D7EBA4BDF45AAAA90410BEDF45155A2DF401D71C0A2DBC7EB80000280824ADBD",
INIT_28 => X"A82B680175EFB6802DBC7BE8A155EFE3FBC71FF145B42038550E38E92EB803FF",
INIT_29 => X"243800002FBD7EBFBD24101C556FA38490A3FE92BEFFEAB45417FD24385D2AAF",
INIT_2A => X"5056DE3D17FE92BEF1EFA92AA8428A10007FD557DFFDF6AA381C0A2DA82FFDB5",
INIT_2B => X"B400925D7FD557DA2803DE10BEF5EDAAAAAD547038EBD57DF7DA2AEB8FC70051",
INIT_2C => X"7FF8FEF410E001FF000E17555555B7AE10410E00155497FEFABA4120B8F55085",
INIT_2D => X"2FBD7545AA8000000000000000000000000000000000000000000005B6AA8214",
INIT_2E => X"A284000AA08003FF55002AA8BEF00517FE00082EBDF45AA8428A10085568ABAA",
INIT_2F => X"A5D2EA8A00A2803DF45AA843DF55AAAE82000F7FBD5545AAFBC01555D2EBFF55",
INIT_30 => X"55087FC00BA552ABFE10F784175FFF7803DF45FFAE955EFAAFBD55EF557BC20A",
INIT_31 => X"AAA5D2EBDE00FFFFC00AA08003FF55A2FBC00105D517FEAA082EBFE10F7FFE8B",
INIT_32 => X"DFEFA2AEAAB550051401FFA2D57FE10F7D57DE00AA842AA00007FD75FFF7FBE8",
INIT_33 => X"FDEAA08042AB45087FC0010557FD55FFAA843FE00F7D17FEBAA2D5574BAAAD17",
INIT_34 => X"000000007BE8A005D7FEABFF002E821FF082A97555557FE8A00002E82155007B",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000067FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(1),               -- Port A write enable input
DIA(0)   => data_write_a(13),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(13),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(1),               -- Port B write enable input
DIB(0)   => data_write_b(13),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(13),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_14_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10020A000180000284008280000281800000030000000033022000000580002",
INIT_01 => X"A14009821830284D186860000C30C24840000000084000084200090008510200",
INIT_02 => X"102100600C9001100000061020A8503401044880010400204908012018122F64",
INIT_03 => X"00008015074608840190800010008002030400002074F401209A108448404842",
INIT_04 => X"000080400004A00100004000840E000201000000024024401200020180180080",
INIT_05 => X"0A000484800111020495040800208C2084000080000010010020049818002008",
INIT_06 => X"1000088020450402B6A1420511C080008468A80008000D0200018B202067AF10",
INIT_07 => X"422000044005000910040110510260040024400C800000BE3850A144C924080E",
INIT_08 => X"000B004028020104111100200001020210A51040008004616001910801010000",
INIT_09 => X"000800004D492408208000000000000406401C0C40800022C8088DB420200900",
INIT_0A => X"0010000002004048000005040160042229140002090200000401000484000400",
INIT_0B => X"0000110100000000010000100000000000000100000000000000100000000000",
INIT_0C => X"409120940404104C2000210100400000011020080084040040005C0010820208",
INIT_0D => X"E0E0A0000190081200000000000000003000000000100C088020028102408120",
INIT_0E => X"E0E0A0000B02740421A0E5D1A024002050805210040000B0E0A0000210040000",
INIT_0F => X"E01200860008920106460D4501CB000111300210008000B0E0A0000210008000",
INIT_10 => X"0ABBC00905C33C6000400F02740412C0715C40110080A4006110510C14D18178",
INIT_11 => X"20000041DB011CC000090012565306500002411420220080220C0093C3892324",
INIT_12 => X"5809240C09024A4AE0CA00004800839682398000120800658992F3C700C30181",
INIT_13 => X"002B46867DBC002A830280000800F7B7A0B1E240240A8340000200067EAA8CB6",
INIT_14 => X"42004005800004801150A00341244000845C7DB0D0200900422ACA4B28000002",
INIT_15 => X"8120481204812048120481204812051A04204110002A26924302590802000000",
INIT_16 => X"1204812048120481204812048120481204812048120481204812048120481204",
INIT_17 => X"2048120481204812048120481204812048120481204812048120481204812048",
INIT_18 => X"69CB91FE1EF7D3ABEFBECA080050000000000000000000081204812048120481",
INIT_19 => X"F3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF7EFBBBBBF9E79E7BEAAF3",
INIT_1A => X"CFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCF3CF3CF3C",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FF007F3F9FCFE7F3F9FCFE7F3F9F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"45AAD157400007BEAAAAAAAE955555D5568A105D000000000000000000000000",
INIT_1F => X"0AAF784020AAF7D56AAAA5D043FFFFAAAABDEAA557BFDE00FFD140155F7D17DF",
INIT_20 => X"ABEFFF8400010082EAABFF55002ABEF085155400FFD1420100055574AAA2AA80",
INIT_21 => X"40155A28028B550051574005D7FFFE105D7BD7545A284020BA0055421FF00042",
INIT_22 => X"1421FF5D7FFDEBA085168B45FF843DEBAF7843FFFFF7AABDF55A2AA97400AAD5",
INIT_23 => X"04155EFAA842ABEFA280155EFFFFBC01EF08554000055002AB455D5142010085",
INIT_24 => X"57FD7410552EAAABAAA8017400AAD140000002EBFFEFA2AAA8BEFF780021FF55",
INIT_25 => X"000000000000000000000000000000000000005568A1055043DEBAAAFFE8B455",
INIT_26 => X"8E3DF45155EBD17FF6DAADB504001C71EDA82AAA0955455D556DA00490000000",
INIT_27 => X"101C55554AAAAA480082FF84000BAEBD16DA82410A3FFD7AAA4B8E824971F8E3",
INIT_28 => X"092085F401D71C0A2DBC7EB80000280824ADBD7490E28BEF085157428FFDB420",
INIT_29 => X"DF45AAAA90410BEDF45155A28E2AB7D0051504005D71F8E004975D556DB68405",
INIT_2A => X"28B6D5D51420101C5B401EF417BFAEAA08516AB45E38E38E92EB803FFD7EBA4B",
INIT_2B => X"EAFBC7EB80071FF5500175EFB6802DBC7BE8A155EFE3FBC71FF145B420385500",
INIT_2C => X"0A3FE92BEFFEAB45417FD24385D2AAFA82B68015400AADB40000082EBFFC7A2A",
INIT_2D => X"5557FE1000000000000000000000000000000000000000000000000556FA3849",
INIT_2E => X"AA8428A10085568ABAA2FBD7545AAD17DFFFAAFFC200055557DE00A280155455",
INIT_2F => X"F0051554AAFFFFC00105D55554BAA28400000F784020BAAAD17FE00082EBDF45",
INIT_30 => X"000051575FFF78415410087BC01555D2EBFF55A284000AA08003FF55002AA8BE",
INIT_31 => X"A00A2803DF45AA843DF55AAAE82000F7FBD5545AAAEAABFF0051400105D5568A",
INIT_32 => X"55EF557BC20AA5D042ABFF555142000557FC01EF007FEAABA00556AB55A2AEA8",
INIT_33 => X"C0010082EBDF55A2AABDF45A284175FF5D04175FFF7803DF45FFAE955EFAAFBD",
INIT_34 => X"00000000517FEAA082EBFE10F7FFE8B55087FC00BA552ABFE10F78415400A2FB",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000007FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(1),               -- Port A write enable input
DIA(0)   => data_write_a(14),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(14),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(1),               -- Port B write enable input
DIB(0)   => data_write_b(14),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(14),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_15_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000A000000000284000280000001800020030000000033022000000180002",
INIT_01 => X"A140098018300848180060000C00426040000000080000080200000000110200",
INIT_02 => X"1020004000801110000006100028503400040800010430004808000180120278",
INIT_03 => X"00008011064408840190800000228002A3000000000010000008108448000042",
INIT_04 => X"701280400004A991000000A28406000211000000220004941000000880000000",
INIT_05 => X"02000484800155020495000800218020C4002880005310000000040000000001",
INIT_06 => X"10000880004540000711224491C08000850A880008000D020001892020656300",
INIT_07 => X"8A04000016050009140501505100000420204008000000BE70408104C8000000",
INIT_08 => X"001F004028026104111002200000000200210040008004614001100801010000",
INIT_09 => X"000800000D09240000800000000000040600180840800022C8088C1020200000",
INIT_0A => X"0000000002004040000105000040042229140002080000000400000080000400",
INIT_0B => X"0000110100000000010000100001000010000000000000000000100000800008",
INIT_0C => X"0001008000000000000025000040000001300008009400006200580010000000",
INIT_0D => X"0000000002300012000000000004200030000000000008008020020000000000",
INIT_0E => X"0000000001000000400000000000000000000010108000000000000010108000",
INIT_0F => X"0000000000000200000900000000000000000010140000000000000010140000",
INIT_10 => X"0140000000000000000001000000400000000000000000000100008040000000",
INIT_11 => X"0000004000480000000000100004400000000030002000406000000000068409",
INIT_12 => X"8000000000020080080000000000802010000000000800000201000800000000",
INIT_13 => X"00000100000000000000000008000000184400A0000000000002000000441108",
INIT_14 => X"4000000000000000010620000004000000000242038B82800000000000000002",
INIT_15 => X"0000000000000000000000000000041800000110000024130202500802000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000080050000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"000804154AA5D00001EFF78428AAA007BC2145F7800000000000000000000000",
INIT_1F => X"0AA007FC2000F7D17DF45AAD157400007BEAAAAAAAE955555D5568A105D7FC00",
INIT_20 => X"FFFFAAAABDEAA557BFDE00FFD140155F7FBD74AAAAD17DF45F7D1421EF005540",
INIT_21 => X"020AAF7FFFDF45FF84000BA552ABDFEF08517DF55A2FBEAB555D556AAAA5D043",
INIT_22 => X"FEAB45F7843FF45082A801FF005155400FFD1420100055574AAA2AA800AAF784",
INIT_23 => X"D5421FF00042ABEFFF8400010082EAABFF55002ABEF087BE8ABA555168B55AAF",
INIT_24 => X"D7BD7545A284020BA007FFFE10A284000AA0055401550055574005D2E800AAA2",
INIT_25 => X"000000000000000000000000000000000000000028B550051574005D7FFFE105",
INIT_26 => X"55D556DA004971C7038140012482550E021C7EB8028A821C7BC516DFF8000000",
INIT_27 => X"45E3DF471C70851400BA0071C5028FFD17FF6DAADB504001C71EDA82AAA09554",
INIT_28 => X"B555D516DA82410A3FFD7AAA4B8E824971F8E38E3DF45155EBF1D5492BED17FF",
INIT_29 => X"54AAAAA480082FF84000BAEBF1FFF7DEB8000092552ABFFEF08517DF6DB6FBE8",
INIT_2A => X"EFA8241516DB55A2FFEAB6DEB843DF551C20801C71C5157428FFDB420101C555",
INIT_2B => X"550428412A85082BEDF401D71C0A2DBC7EB80000280824ADBD7490E28BEF087F",
INIT_2C => X"51504005D71F8E004975D556DB68405092087FF8E00BE8A02082005F47145085",
INIT_2D => X"57BD75EFF78000000000000000000000000000000000000000000000E2AB7D00",
INIT_2E => X"55557DE00A2801554555557FE100055554BA5504000105D2A80145AA842AA005",
INIT_2F => X"5AAD557410F7D57DF55AAFBD55450055420BA0055574BAF7D17DFFFAAFFC2000",
INIT_30 => X"FF08517FFFFF7FBEAB455D517FE00082EBDF45AA8428A10085568ABAA2FBD754",
INIT_31 => X"4AAFFFFC00105D55554BAA28400000F784020BAAAD57FFEFA28402010552ABDF",
INIT_32 => X"FF55002AA8BEF007FFDE1000557DF45AAFBE8BEFA2803FF45550400155555155",
INIT_33 => X"80000087BD55450855400BA002A95400F7FBC01555D2EBFF55A284000AA08003",
INIT_34 => X"000000002EAABFF0051400105D5568A000051575FFF78415410087FEAA10F7AE",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000060000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(1),               -- Port A write enable input
DIA(0)   => data_write_a(15),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(15),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(1),               -- Port B write enable input
DIB(0)   => data_write_b(15),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(15),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_16_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"DA22C618B1000482B688B186588884862A400438255FC38381441205BA803003",
INIT_01 => X"264AC80028404C211203A952A90341080B173340412000E1005D628000820484",
INIT_02 => X"400034C206C405000001A48202084004003008255040826EE008B440200E2042",
INIT_03 => X"2916704900606AC82B49CC56DF8CC1E50E4800202115005760010010000C0400",
INIT_04 => X"052DCA856DC7504B82BF6614C86D2B7F85AAD17F4B100000B88148C4804A428A",
INIT_05 => X"373CB02A00C0502F301180141A42A5720E0F43C17A8479580001AC20000000E2",
INIT_06 => X"303E2094282B85242C85001038D5710E8410D5959BC4800015001219D0550077",
INIT_07 => X"880100000159954501280B0080146F7112D949A0015018220540000382805001",
INIT_08 => X"30015452880C8D90409A05B2CB2CA400200209E5601044A24000000462A60018",
INIT_09 => X"452D54000C0907000330000000000096480050000685400005FC014743E0DC92",
INIT_0A => X"00014808A02004200E540480212000A448C0080024AEA00C9688000000000005",
INIT_0B => X"000D58460018F6D3D84400044000440004400044000440004400042000220002",
INIT_0C => X"0001004010A8812831605DA0000A054052E40000817680220040025699200002",
INIT_0D => X"AAADA0C343F1AC1B01040A002024895514554485D00000012400240000000000",
INIT_0E => X"AAADA0CC421CA003B694B68018FAAA708E2CB5320018CAC99BA0A3B9320018CA",
INIT_0F => X"B1443A1891E4A928C29020E6A8524CE7A3EE59320018CAC99BA0ACB9320018CA",
INIT_10 => X"04B2A5A40B1E6644AF0F021EA003AC24352AB2449A3FF2FA04E5E09B128834AD",
INIT_11 => X"60ED838E890B703C6260D8E3A21275714C902375B801324301AB0067622E5E54",
INIT_12 => X"064F70DBDB1C74424E91E1C194C71D1216F50A8C241815FEB6A9158863F638FB",
INIT_13 => X"45FDF9D364DBD9435A6D45C9E81BED555E4C15F11133D171727A2550EE2F1BA0",
INIT_14 => X"08150013F162119014204373517700ACCC59432A2B2D001F803471A9A960E572",
INIT_15 => X"000000000000000000000000000000880002054000229088542210206B2AB015",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"2A898D21B4C98389ED146C080000000000000000000000000000000000000000",
INIT_19 => X"A29A29A29A29A29A29A29A29A29A28A28A28A28A28A53CBF0F0D3CF3CF0AB1A2",
INIT_1A => X"8F47A3D1E8F4FA7D3E9F4FA7D3E9F4FA7D3E8F4FA3D3E8F4FA3D3E9A29A29A29",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000FA7D3E9F4FA7D1E8F47A3D1E",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFF7FBE8B45AAD568BFFFFAA975FF00003FE0055000000000000000000000000",
INIT_1F => X"0005D2A95410FFFFC00000804154AA5D00001EFF78428AAA007BC2145F7843FF",
INIT_20 => X"7400007BEAAAAAAAE955555D5568A105D2E974BAF7FBEAB45FFFFC00BAF78002",
INIT_21 => X"C2000F78000010552E800AA002E821FFA2AAAAA00000417555FFD17DF45AAD15",
INIT_22 => X"43FEBA5D55575FFF7AABFE00557BD74AAAAD17DF45F7D1421EF0055400AA007F",
INIT_23 => X"D56AAAA5D043FFFFAAAABDEAA557BFDE00FFD140155F7AABDF55F7AE820AA080",
INIT_24 => X"8517DF55A2FBEAB555D04154BAA2FBE8B55FFFFD55FF557FC2000FF8015410FF",
INIT_25 => X"000000000000000000000000000000000000007FFDF45FF84000BA552ABDFEF0",
INIT_26 => X"21C7BC516DFF8438FC7E3F1EAB55B6DF6DBFFF7AA955C71C043FE10490000000",
INIT_27 => X"55FFF1C70BAF78A000005D2097438FFF1C7038140012482550E021C7EB8028A8",
INIT_28 => X"57DEBD17FF6DAADB504001C71EDA82AAA0955455D556DA00492490492F7FBE8B",
INIT_29 => X"71C70851400BA0071C5028FF84020285D2085092002A801FFB6AAA8A10080E17",
INIT_2A => X"BAF6DE3AA8709208043FEBA555B555FFE3AABFE005D71D5492BED17FF45E3DF4",
INIT_2B => X"BC0028E38412428EBD16DA82410A3FFD7AAA4B8E824971F8E38E3DF45155EBA4",
INIT_2C => X"8000092552ABFFEF08517DF6DB6FBE8B555D04124BAB6FBE8B45E3FBD55D7557",
INIT_2D => X"5003DE000000000000000000000000000000000000000000000000071FFF7DEB",
INIT_2E => X"5D2A80145AA842AA00557BD75EFF78428B55AAD168B55F7FFFDFEFFFAA955555",
INIT_2F => X"0000000010F7FBEAB45FFD1554AAFFAE820105500154AAF7D5554BA550400010",
INIT_30 => X"EFF7AEA8A10002E955FFA2D17DFFFAAFFC200055557DE00A2801554555557FE1",
INIT_31 => X"410F7D57DF55AAFBD55450055420BA0055574BAF784000BA5D0017410082E801",
INIT_32 => X"8ABAA2FBD7545AA802ABEFA2AA9541000003DEBA557BD75EFA2AEBDE105D5557",
INIT_33 => X"EAB45AAFFD55555D7FC20AAA280000AAAAD17FE00082EBDF45AA8428A1008556",
INIT_34 => X"00000000557FFEFA28402010552ABDFFF08517FFFFF7FBEAB455D04020AAFFFB",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000020000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(2),               -- Port A write enable input
DIA(0)   => data_write_a(16),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(16),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(2),               -- Port B write enable input
DIB(0)   => data_write_b(16),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(16),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_17_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"5284CE4FB7BD2C8994A13392DBD02E14006B82AC7E800D44D3DD2FD5F9B961C0",
INIT_01 => X"F9BA301F7E03FC6793F2199B39FC233C11D93AE6F3BB92B32091DBC339B24542",
INIT_02 => X"1D5FC0C08F040404446965C0607FB8A217C400C33A908078551BD04222186338",
INIT_03 => X"A14124C28DFD960832C90446DF8400A5055C25295B695FF97E1B5AC757F06D6B",
INIT_04 => X"04A106866DA3D02A01FB660C08A4AB7F840EDB6F48100DFC8081081D78AC7402",
INIT_05 => X"51E072F0C0C58D9C125EBFC00A46CF0388054100F680E0CE0107B8D040DAFCDA",
INIT_06 => X"019A4D00786B048112C58B16307F15DE8408B233661C10BBA5DAAFA9DDA1194D",
INIT_07 => X"8E00001660700CE170284A00891C7C03D29DE26814515835902AC089A2801540",
INIT_08 => X"C009F3A1B0120A1C51DFF881861CBE0305A12A0321810217C01D34EDC98FFA1C",
INIT_09 => X"747E6610052CDEE97FF1F9F63E3EF790380078002CE976AB6BF769769E4D437D",
INIT_0A => X"00185C44B91BC1740B7605040BE0018CFC7429F326B9D045FF8000E9AB415606",
INIT_0B => X"3A28FC1AAF5CF6F3D3EF3D3EF3D3EF3D3EF3D3EF3D3EF3D3EF3D3EF9E9F79E9E",
INIT_0C => X"0000020012E9E10A31EB5FF9296A67F5B4FFBD2FAD7FE653C3FBFF33E10C001B",
INIT_0D => X"333EA16031F2BD47BDA2CA5D8164FCCFE833C5C3D00018006C68170000000000",
INIT_0E => X"333EA160391BEFF2C32FB695F919110D5ECE542A6FEEB2533EA160782A6FEEB2",
INIT_0F => X"D18C0D06638A207CFDE1F7DDAD76D5282400F82A6FEEB2533EA160782A6FEEB2",
INIT_10 => X"E6E43E59AFE4A59B57679D19EFF2C7573FAD5A86840354D1706FFFA3EF6E24B6",
INIT_11 => X"F7D7A0ABD6DAAAB96529382B74E4E1FE4ACA4D77FAAB77CE3AF3EE78F58DB737",
INIT_12 => X"2D1281017F056E9C9C3FC95949C157ADB55572CA52606DFED6CA55334C04C04F",
INIT_13 => X"59FDEB974F486905001FDF5FA0D719F9956EAA1A184045D5D7A870D2F5A5D752",
INIT_14 => X"60158015177F916A039EF41FDB34A91F432EA58949D5B5C85F97871876F7D7E8",
INIT_15 => X"000000000000000000000000000004DC200005E705B7B3D9FC22F00BE419FB55",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"06013DB9880A5D22E229F3030018000000000000000000000000000000000000",
INIT_19 => X"D35D74D35D74D34D35D74D35D74D34D34D34D34D34D0D30D0D303AEBAE886E40",
INIT_1A => X"51A8D46A351A0D068341A0D068341A0D068341A8D468341A8D46834D35D74D34",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000008D46A351A8D46A351A8D46A3",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFF7FBFDF55A28402000F7D56ABFF55000000000000000000000000",
INIT_1F => X"A00F7843FEBA55043FFFFF7FBE8B45AAD568BFFFFAA975FF00003FE0055043FF",
INIT_20 => X"54AA5D00001EFF78428AAA007BC2145F7D568B45000002010552EBDF45A28028",
INIT_21 => X"95410FFAE800105D2A95410002A95410AAAEBFF55AAFFC00BAF7FFC000008041",
INIT_22 => X"57DE00F7AE800AAAAAABDFEF5D2E974BAF7FBEAB45FFFFC00BAF780020005D2A",
INIT_23 => X"517DF45AAD157400007BEAAAAAAAE955555D5568A105D7FFFFEFA2D568BFFFFD",
INIT_24 => X"2AAAAA00000417555FF8028B55082A974105D003FF55F7802AAAAAAD168AAA5D",
INIT_25 => X"000000000000000000000000000000000000000000010552E800AA002E821FFA",
INIT_26 => X"71C043FE10490A3FFFFFFFFFDFEFE3F5FAF45AA8000038F7DB6FBD7490000000",
INIT_27 => X"384124BFF7DB68A28A38F7803DE82490438FC7E3F1EAB55B6DF6DBFFF7AA955C",
INIT_28 => X"0BAFFF1C7038140012482550E021C7EB8028A821C7BC516DFFDF68B551C0E050",
INIT_29 => X"70BAF78A000005D2097438FFAA85000492495428082E95400AAA0BDF7DB6F5C7",
INIT_2A => X"FAFFFB6D56FBFFEBDB78E38F7AA800BAB6AEBDFD75D2490492F7FBE8B55FFF1C",
INIT_2B => X"028AAAB6D16FA8249517FF6DAADB504001C71EDA82AAA0955455D556DA00497F",
INIT_2C => X"2085092002A801FFB6AAA8A10080E1757DEB8A2DB5514249243841003FF6DEB8",
INIT_2D => X"7FFFDF550000000000000000000000000000000000000000000000004020285D",
INIT_2E => X"F7FFFDFEFFFAA9555555003DE00002ABFFEFF7FBFDFFFAAD168B55AA80000BAF",
INIT_2F => X"FF7FBEAB45552E954BA08003DFFFFFAAA8AAAF7843FE10000428B55AAD168B55",
INIT_30 => X"10AA843FFFFF7D5554BAF7D5554BA5504000105D2A80145AA842AA00557BD75E",
INIT_31 => X"010F7FBEAB45FFD1554AAFFAE820105500154AAF7AE974000800154AA002E954",
INIT_32 => X"554555557FE10007FEABEFFFD57FFEFAAFFE8ABAFFAA820BAF7AEBFF55550000",
INIT_33 => X"020AA08003DFFFA28028AAAF7D17DE0000517DFFFAAFFC200055557DE00A2801",
INIT_34 => X"0000000004000BA5D0017410082E801EFF7AEA8A10002E955FFA2AABFF455500",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000067FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(2),               -- Port A write enable input
DIA(0)   => data_write_a(17),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(17),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(2),               -- Port B write enable input
DIB(0)   => data_write_b(17),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(17),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_18_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"69844019080000A21A611406840014122A641074155FC28A2024001001801003",
INIT_01 => X"01067920034004180005E9E3C90360C0041C0181002001602025800008440084",
INIT_02 => X"40AC3CAA22D605200000856E2481902400344A20F802C22054001000021E2379",
INIT_03 => X"A95308ECD3207AC81D91C4002004C08A06008080BA868007E58040102B0E0100",
INIT_04 => X"044CC183800CA00780808004C8DB841405A80A100B586200FAC24AE4805242CA",
INIT_05 => X"771C10000000000B1135883C08A115320E0401C0200038394230070A19000020",
INIT_06 => X"3001499C602A8A003E800A042D8132A00098408F79E3901218050018024110D6",
INIT_07 => X"5029401000C983E60004010030400353C05806800104004E0000042E52800E20",
INIT_08 => X"0000117088080990419005B0C309402030060860E01004A828408800440405E3",
INIT_09 => X"6B8186185C42900693A002004040001E1950850C848601008708114A2030B480",
INIT_0A => X"100180A8062026000DC425C0301311324AA237108857220BA089420440000030",
INIT_0B => X"C44703657083080C2800C2000C2000C2000C2000C2000C2000C2000610006100",
INIT_0C => X"C1B0609C05013065CC042004040808084001E000108010230400800FD9B286C4",
INIT_0D => X"CCC15F9CBA45505640000A402019003F140FC2060014250B9080008306C18360",
INIT_0E => X"CCC15F9FB1962FCB69E08AAAEAEBCDDF7C728582081483ACC15F9C3982081483",
INIT_0F => X"EBF1CFFF7670ACC3811A28AB57523CDFEBFBF982081483ACC15F9F3982081483",
INIT_10 => X"C9002BF05800D875E63CC9962FCB52CAA02FE3F8E7F5E3AC3620805298B15A3F",
INIT_11 => X"F1B72A8A800B7546DB9F1CA320037F01BD67DC4041D4CF03138DD865103EFEEA",
INIT_12 => X"81CCFAFDBF9464006FD037AEFAE5150016EA8DB7BFE25208E8F46A228BF8A757",
INIT_13 => X"641256EC844B8AF92FD7CEDC24A9E181A8A29509EAAE7FD3B749471C48F8A459",
INIT_14 => X"0297D086E00036D2440E0880AAD62BEFF5778802A3AF8E8FB0440CE78773B709",
INIT_15 => X"8360D8360D8360D8360D8360D83609220D20D00000080C0601400B402307E480",
INIT_16 => X"360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D",
INIT_17 => X"60D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8",
INIT_18 => X"D9D701DC2E784601EFBE2C00000000000000000000000008360D8360D8360D83",
INIT_19 => X"5155555545145145155555545145145145145145145220B22A0B820820965177",
INIT_1A => X"44A25128944A25128944A25128944A25128944AA552A954A2512895554514514",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000025128944A25128944A251289",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFEFF7AE954BA5D04174AA00000000000000000000000000",
INIT_1F => X"145AA801741000043FFFFFFFFFFFFFF7FBFDF55A28402000F7D56ABFF55043FF",
INIT_20 => X"8B45AAD568BFFFFAA975FF00003FE0055043FFFFFFFFFDFEFA2D56AB45AA8400",
INIT_21 => X"3FEBA55557FFEFA2D168B55AAFBFFFFFFF80021EF0855421EF00043FFFFF7FBE",
INIT_22 => X"A82155F7AEBFEBAFFD56AA00A2D568B45000002010552EBDF45A28028A00F784",
INIT_23 => X"FFC00000804154AA5D00001EFF78428AAA007BC2145F7D5400000004020AA5D2",
INIT_24 => X"AAEBFF55AAFFC00BAF7AE80010082E954BA0004174AAAA8428B45082ABFEBAA2",
INIT_25 => X"000000000000000000000000000000000000002E800105D2A95410002A95410A",
INIT_26 => X"8F7DB6FBD7490E3FFFFFFFFFFFFFFFFBFDFEFFFAE954AA550415492140000000",
INIT_27 => X"D7AAD16FB6DBE8E00155BE8015410140A3FFFFFFFFFDFEFE3F5FAF45AA800003",
INIT_28 => X"1C7140438FC7E3F1EAB55B6DF6DBFFF7AA955C71C043FE1049043FFEFE3F1F8F",
INIT_29 => X"FF7DB68A28A38F7803DE82495B78FC7AAD56FB6DBEF1FAFD7E384001EF145B47",
INIT_2A => X"420381C0A02082492A85155E3A4BDE92FFD56FA28B6DF68B551C0E050384124B",
INIT_2B => X"E28B7D1420BDEAAA2F1C7038140012482550E021C7EB8028A821C7BC516DFFD1",
INIT_2C => X"2495428082E95400AAA0BDF7DB6F5C70BAFFAE870280024904BA1400174AABE8",
INIT_2D => X"50415410550000000000000000000000000000000000000000000002A8500049",
INIT_2E => X"AAD168B55AA80000BAF7FFFDF55002ABFFFFFFFFFFFEFF7FBFDFFFF7AA974BA5",
INIT_2F => X"000043DFEFA2D56AB45AAD57DFEFF7AA82155F78015400552ABFFEFF7FBFDFFF",
INIT_30 => X"55A280021EF557FD7555550428B55AAD168B55F7FFFDFEFFFAA9555555003DE0",
INIT_31 => X"B45552E954BA08003DFFFFFAAA8AAAF7843FE10007FEAB55A2D17FFEFFFD568B",
INIT_32 => X"AA00557BD75EFF7D1400AA5D2A82000002A95545A2843FE00F7D17FEAAF7FBEA",
INIT_33 => X"020AA5D04154BAF7AEA8BEF55003DEAAA2D5554BA5504000105D2A80145AA842",
INIT_34 => X"000000002E974000800154AA002E95410AA843FFFFF7D5554BAF7AE974BA0004",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000020000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(2),               -- Port A write enable input
DIA(0)   => data_write_a(18),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(18),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(2),               -- Port B write enable input
DIB(0)   => data_write_b(18),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(18),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_19_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"042200000000000041088001001AA00000000000000000000000500802000003",
INIT_01 => X"074018000024000000000404000000000A22000800000800004A200000000001",
INIT_02 => X"0000048002C405000000000006A84000000000200893C246A20000000020031A",
INIT_03 => X"020A9639044012C80001C4000004C08006000000001025000000000000000000",
INIT_04 => X"0400C0800000000380800004C8000000058800000B1000009880480480024200",
INIT_05 => X"420410000000000B10804004080001320E0401C0200038080000000000000000",
INIT_06 => X"2002409006F00A8428050A000280493104004500480090080A01120220140020",
INIT_07 => X"0000000000418026090240923240002190400000000000C0054A912054004021",
INIT_08 => X"0000115080000990000000B0C308000000000860200160000000000038380000",
INIT_09 => X"8000F80001012590001000000000001618000000020280008180810200000000",
INIT_0A => X"0000000000000000000000000000000100008000110000000000000000000017",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000840007600000000000000000800259000000",
INIT_0D => X"0008A0034078104B41A41000000000031400C002000000000000000000000000",
INIT_0E => X"0008A0004263C0343EDD414004042228DC0D385598035D0008A003B05598035D",
INIT_0F => X"040231068187C39F5A4F985C008902041124505598035D0008A000B05598035D",
INIT_10 => X"1BFBD406451B02000E033263C0343CB740500401180DE053A98F6ECC739D8140",
INIT_11 => X"420851546B2400000040D8549B5800000010227848D4303807FC8CC5508AEAED",
INIT_12 => X"52210402120A936B0000000004C2A8D6480000000018A700FCF980CC300318A2",
INIT_13 => X"B1427ED430B41402D025082359700181C21140E40511802208D6B30C48F8A8A4",
INIT_14 => X"9C000018440021011821B35254E99AF9E9410006362A2B6424287B08286208D6",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000023006000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"7747E18E0218CC18E88324000000000000000000000000000000000000000000",
INIT_19 => X"34C30C30C30C30D34C30C30C30C30C30C30C30C30C3504118982A69A6980E411",
INIT_1A => X"C26130984C26130984C26130984C261309A4D26130984C26130984C30C30C30D",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000130984C26130984C26130984",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAA954BA5500020BA5D000000000000000000000000",
INIT_1F => X"4BA5D517FFFF08043FFFFFFFFFFFFFFFFFFFFEFF7AE954BA5D04174AA007BFFF",
INIT_20 => X"FFFFF7FBFDF55A28402000F7D56ABFF557BFFFFFFFFFFFFFFFFFBFDFEFFFAA97",
INIT_21 => X"17410007BFFFFFFFFFFFFEFF7D16AB45AA8002000F7D5575455D043FFFFFFFFF",
INIT_22 => X"568B55F7AE955FFAA840201008043FFFFFFFFFDFEFA2D56AB45AA8400145AA80",
INIT_23 => X"043FFFFF7FBE8B45AAD568BFFFFAA975FF00003FE00557BFFFFFFFFBFDF45AAD",
INIT_24 => X"F80021EF0855421EF002ABFFEFF7D168B55AAD17FFEFF7AE975FF00557FFFF5D",
INIT_25 => X"00000000000000000000000000000000000000557FFEFA2D168B55AAFBFFFFFF",
INIT_26 => X"A5504154921471FFFFFFFFFFFFFFFFFFFFFFFF7AA954BA550000082550000000",
INIT_27 => X"EFF7FBFAFD7E3A4954BA555B7AFC7080E3FFFFFFFFFFFFFFFFBFDFEFFFAE954A",
INIT_28 => X"545550A3FFFFFFFFFDFEFE3F5FAF45AA8000038F7DB6FBD74975FFFFFFFFFFFF",
INIT_29 => X"FB6DBE8E00155BE8015410147FFFFFFF7FBF8FC7EBD568B55A28000000FFDF52",
INIT_2A => X"FDFC7E3F1FAF55A2DB6FB7DF7AE955C7BE800000008043FFEFE3F1F8FD7AAD16",
INIT_2B => X"0955FF145B7AFC7410438FC7E3F1EAB55B6DF6DBFFF7AA955C71C043FE10497B",
INIT_2C => X"D56FB6DBEF1FAFD7E384001EF145B471C71424B8FC7E3D56AB6DB6DF7AFC7EBA",
INIT_2D => X"50002000550000000000000000000000000000000000000000000005B78FC7AA",
INIT_2E => X"F7FBFDFFFF7AA974BA55041541055517FFFFFFFFFFFFFFFFFFFFEFF7AA974AA5",
INIT_2F => X"500517FFFFFFFBFDFEFFFFFEAB45AA80154AA557BEAB45002ABFFFFFFFFFFFEF",
INIT_30 => X"55A28002000F7FFC2155552ABFFEFF7FBFDFFFAAD168B55AA80000BAF7FFFDF5",
INIT_31 => X"FEFA2D56AB45AAD57DFEFF7AA82155F78015400557BFDFEFF7FBEAB55A2D56AB",
INIT_32 => X"555555003DE00007FFDF45AAD568B45AAFBFFFFFFFAA95545F7840201000043D",
INIT_33 => X"6ABFFFFFBEAB45A280155EF557FE8B55000428B55AAD168B55F7FFFDFEFFFAA9",
INIT_34 => X"000000007FEAB55A2D17FFEFFFD568B55A280021EF557FD755555042AB55AAD1",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000040000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(2),               -- Port A write enable input
DIA(0)   => data_write_a(19),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(19),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(2),               -- Port B write enable input
DIB(0)   => data_write_b(19),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(19),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_20_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000003",
INIT_01 => X"A65FF80000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000048002CC070000000000000000000000002FF86100200000000220002362",
INIT_03 => X"00000000000203D80025DC18004DC3D01E000000000000000000000000000000",
INIT_04 => X"07E5DF808071026F87C4191DD8005080679800000F300002998058068002C000",
INIT_05 => X"C205F23A2100557F70000004390021F61E1E87C3FD0CFBF80880072042000044",
INIT_06 => X"1209244C2000100006800000020010000008407FC800B0000000100600040000",
INIT_07 => X"8802000009FFBFE51886018002040020000800000554003E0000000002800000",
INIT_08 => X"30801F5780259FB0000000F7DF78020004011FEFE00000000020031502000083",
INIT_09 => X"00000000001000000000000000000056F8000001000000040000040141800802",
INIT_0A => X"0000000000000008000800000000000000000000000000000010010014800000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"00010240001721214E000004000000080000008000001000040080FFDB000000",
INIT_0D => X"0000000F3008001E00000000001803FF14FFC006000000008010200000000000",
INIT_0E => X"0000000F3040200000020000000026A70C0008020000200000000F3002000020",
INIT_0F => X"000030B86000400080000200000000004A58F0020000200000000F3002000020",
INIT_10 => X"0000000002183E61E6000040200001000000000019B140000800800000020000",
INIT_11 => X"C00010080000000000525801000000000014AC08000000508001030A0A400100",
INIT_12 => X"000002BC360020000000000292C0100000000000A56000090100000000001F86",
INIT_13 => X"8010000000000000574500001001060600000000001716800000803102020000",
INIT_14 => X"00000000000040040040002000080506049CDF70C08040100000706707600000",
INIT_15 => X"00000000000000000000000000802040200200604040000000000024FB7FE008",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"060070400020112240209A408004000000000000000000000000000000000000",
INIT_19 => X"65965965965965965965965965965861861861861860D30424343CF3CF340E00",
INIT_1A => X"90C86432190C86432190C86432190C86432190C86432190C8643219659659659",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000086432190C86432190C864321",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974AA55040201008000000000000000000000000",
INIT_1F => X"4AA550002000007BFFFFFFFFFFFFFFFFFFFFFFFFFAA954BA5500020BA5D7FFFF",
INIT_20 => X"FFFFFFFFFFFEFF7AE954BA5D04174AA00003FFFFFFFFFFFFFFFFFFFFFFF7AA97",
INIT_21 => X"7FFFF087FFFFFFFFFFFFFFFFFFFFDFEFFFAE974AA5D003FE005D043FFFFFFFFF",
INIT_22 => X"BFDFFFAA84000105D556AB55557BFFFFFFFFFFFFFFFFFBFDFEFFFAA974BA5D51",
INIT_23 => X"043FFFFFFFFFFFFFF7FBFDF55A28402000F7D56ABFF55003FFFFFFFFFFFFFF7F",
INIT_24 => X"A8002000F7D5575455D2EBFFFFFFFFFFFEFF7FBEAB55A28000010F7D16ABEF08",
INIT_25 => X"000000000000000000000000000000000000007BFFFFFFFFFFFFEFF7D16AB45A",
INIT_26 => X"A550000082557FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550400028000000000",
INIT_27 => X"FFFFFFFDFEFF7AE974BA5500050380071FFFFFFFFFFFFFFFFFFFFFFFF7AA954B",
INIT_28 => X"E285D0E3FFFFFFFFFFFFFFFFBFDFEFFFAE954AA55041549214043FFFFFFFFFFF",
INIT_29 => X"AFD7E3A4954BA555B7AFC70871FFFFFFFFFFFFFFF7FBFDFFFFFAA974BA550038",
INIT_2A => X"3FFFFFFFFFDFEFF7F1FAFC7A28002028555F6FB7D5D75FFFFFFFFFFFFEFF7FBF",
INIT_2B => X"402010FFDB6ABEF140A3FFFFFFFFFDFEFE3F5FAF45AA8000038F7DB6FBD7490E",
INIT_2C => X"FBF8FC7EBD568B55A28000000FFDF525455524BFFFFFFFBFDFC7E3F5E8B45A28",
INIT_2D => X"504000BA080000000000000000000000000000000000000000000007FFFFFFF7",
INIT_2E => X"FFFFFFFEFF7AA974AA550002000557FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5",
INIT_2F => X"055043FFFFFFFFFFFFFF7FBFDFEFFFAE954BA5500174AA08517FFFFFFFFFFFFF",
INIT_30 => X"EFF7AE974AA550028AAA5D2ABFFFFFFFFFFFEFF7FBFDFFFF7AA974BA55041541",
INIT_31 => X"FFFFFFBFDFEFFFFFEAB45AA80154AA557BEAB4500557FFFFFFFFFDFEFF7FFFFF",
INIT_32 => X"00BAF7FFFDF55002EBFFFFF7FBFDFEFFFD568B55A284020BA557FFFFFF5D517F",
INIT_33 => X"FFF55A2D16AB45AA8402000F7FBEABEF5D2ABFFEFF7FBFDFFFAAD168B55AA800",
INIT_34 => X"000000007BFDFEFF7FBEAB55A2D56AB55A28002000F7FFC215555043DFEFF7FB",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000007FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(2),               -- Port A write enable input
DIA(0)   => data_write_a(20),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(20),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(2),               -- Port B write enable input
DIB(0)   => data_write_b(20),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(20),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_21_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"4A302428B824900A128C090A5C1800261500213C005FE812D10420054085A202",
INIT_01 => X"081FFE3440B609703B0427F801A40B8115BC4F655300340288A40D30040E4DD8",
INIT_02 => X"04CA478082CC1740002019824E0203100640303FF8C0B31061096E21A1840814",
INIT_03 => X"230CA7A4810083F80095DE00102DC3823EA821094EC68248923200013290C800",
INIT_04 => X"07CFFFC04904AA7F8780409DF84A0202879800000F3000029980780EA2C3C002",
INIT_05 => X"DE87F0280000407FF900D914382091FE1E1C0FC3E01EFFF8000480200008D062",
INIT_06 => X"010E2182002BC107A03448808F0D7C002822987FC830F40134CC74D002016612",
INIT_07 => X"0401000011FBFFE00520000200422033025C4209104500000012004C004D8C0B",
INIT_08 => X"00EF1F5FA0041FF080AC70FFDF78220010841EFFE7116E144071268DFD3E4C24",
INIT_09 => X"FC8BFE18008083B4443151462A28C6DFF80010002605302248088950484550A3",
INIT_0A => X"10018C241102068006C620C03882019480E631A0855E924E2598038938404037",
INIT_0B => X"A641165448C80C103648A3648A3648A3648A3648A3648A3648A366451B2451B2",
INIT_0C => X"011100841200D001000624000100C002804A08221890004806A310FFDF000454",
INIT_0D => X"5004D8158809C86065941840B1014FFF56FFC0281280080180B2948004400220",
INIT_0E => X"5004D815810D42E04A08A80098C02450025360694101816002D41A4068C10181",
INIT_0F => X"134160C8125B0B271802242880A04482418A0068C101816002D41A4069410181",
INIT_10 => X"10080E05C0B06AA8B12CFD0D42E0441A300012682960828F05C96A001B029010",
INIT_11 => X"00010362A8A20826A88660D86B202049F115100920C54E8EA256ECF078BA081C",
INIT_12 => X"064802C0081B0D64040936443306C55144104F30A8801406D002900062803201",
INIT_13 => X"4581BA0038005A706680012280506A8010602011819E290048A2118EC8140C08",
INIT_14 => X"CC158092C044600466208CC5091011C322A4C40A0300600C0A80509F41800880",
INIT_15 => X"80200802008020080200802008020412002001000000381C02004000FBFFF80D",
INIT_16 => X"0200802008020080200802008020080200802008020080200802008020080200",
INIT_17 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_18 => X"FDDFEFFFBEFFE7C7BFBEFC000000000000000000000000080200802008020080",
INIT_19 => X"F7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7FFBFBFFF9E79E7FFFDF3",
INIT_1A => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFDFEFF7FBFDFEFF7FBFDF7DF7DF7D",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00001FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D000200008000000000000000000000000",
INIT_1F => X"4AA5D00020AA5D7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550402010087FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAA954BA5500020BA5D7FFFFFFFFFFFFFFFFFFFFFFFFFFAE95",
INIT_21 => X"0200000003FFFFFFFFFFFFFFFFFFFFFFF7AA974BA5D0402000557BFFFFFFFFFF",
INIT_22 => X"FFFFEFF7AE974BA5D00174BA00003FFFFFFFFFFFFFFFFFFFFFFF7AA974AA5500",
INIT_23 => X"043FFFFFFFFFFFFFFFFFFFFEFF7AE954BA5D04174AA00003FFFFFFFFFFFFFFFF",
INIT_24 => X"FAE974AA5D003FE005D2EBFFFFFFFFFFFFFFFFFFDFEFF7AE954AA5500174BA5D",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFDFEFF",
INIT_26 => X"A550400028007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0000010000000000",
INIT_27 => X"FFFFFFFFFFFFFAA954BA5D00000BA557FFFFFFFFFFFFFFFFFFFFFFFFFFAE974A",
INIT_28 => X"0005571FFFFFFFFFFFFFFFFFFFFFFFF7AA954BA550000082557BFFFFFFFFFFFF",
INIT_29 => X"DFEFF7AE974BA55000503800003FFFFFFFFFFFFFFFFFFFFEFF7AA974AA5D0405",
INIT_2A => X"3FFFFFFFFFFFFFFFFFFDFEFF7AE954BA5D00154AA00043FFFFFFFFFFFFFFFFFF",
INIT_2B => X"A974BA5D00104925D0E3FFFFFFFFFFFFFFFFBFDFEFFFAE954AA550415492140E",
INIT_2C => X"FFFFFFFF7FBFDFFFFFAA974BA550038E285D2ABFFFFFFFFFFFFFFFFBFDFEFFFA",
INIT_2D => X"D00000100000000000000000000000000000000000000000000000071FFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE954AA5504000BA087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0557BFFFFFFFFFFFFFFFFFFFFFFFF7AA954BA5D00000BA5D7FFFFFFFFFFFFFFF",
INIT_30 => X"EFF7AE954AA5D041740055517FFFFFFFFFFFFFFFFFFFFEFF7AA974AA55000200",
INIT_31 => X"FFFFFFFFFFFFF7FBFDFEFFFAE954BA5500174AA08043FFFFFFFFFFFFFFFFBFDF",
INIT_32 => X"74BA550415410552ABFFFFFFFFFFFFFF7FBFDFFFFFAA974AA5D00174BA08043F",
INIT_33 => X"FDFEFF7FBFFFFFF7AE954BA5D0000010552ABFFFFFFFFFFFEFF7FBFDFFFF7AA9",
INIT_34 => X"00000000557FFFFFFFFFDFEFF7FFFFFEFF7AE974AA550028AAA5D2EBFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(2),               -- Port A write enable input
DIA(0)   => data_write_a(21),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(21),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(2),               -- Port B write enable input
DIB(0)   => data_write_b(21),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(21),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_22_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"5290F4CDE914905A14A43D33F488243E17122300F55FEB189B343A1140548380",
INIT_01 => X"A94007B259F6A975386262000C344BA9573C6FF57B18A5FB0ABFCD3C2C5F4F0C",
INIT_02 => X"D56B4302AC01005111011BD506AA5205274056900596A539584E2E6DFE4B2418",
INIT_03 => X"9AC0FCBD854688207C90007A1000047A00E588632CA213C8903AD6B55AD0EB5A",
INIT_04 => X"30002047A6FCA110086C402022F2124A8022492580040440002021C922D9109B",
INIT_05 => X"14A206B6838151008D95DD1847811C08002380041F1104002205AC4140DAD060",
INIT_06 => X"1727FF2EB9EF113A10BD32F44289D1F840C1710010344DB9A808FDFF3DE03130",
INIT_07 => X"050700154A00401D00495A06A8D464C5F6B54AA8551040818F4C997AC80CBE05",
INIT_08 => X"0141008801018040E48D50080002B00A0C00801014541E9504703680017F6CB4",
INIT_09 => X"02680000010937986481514E2A29CE010708C0804C6A033F7FCFF9426A41F1AB",
INIT_0A => X"00500001840000C80B410014088040F4A944B1AA313C004554002381B8000500",
INIT_0B => X"A004D1594832824A070AA070AA070AA070AA070AA070AA070AA0725503855038",
INIT_0C => X"501428054278142151262CA50343854E506A2C6898B2950AA6A35B0004284058",
INIT_0D => X"90078E1F840A2B0114020104022460002200050F60E220A06880D2A14050A028",
INIT_0E => X"90078E1F891C239F8908003099C1ACF06273612B3482C0C0078E1F412B1582C0",
INIT_0F => X"1BA1B0FD16770236A4091621C08055C2C0DB012B1582C0C0078E1F412B3482C0",
INIT_10 => X"00101F09C030AB28B03C111C239F870828041BA859F213AFC14AA38043006018",
INIT_11 => X"10E8822A984B0025B0DE6089462660095337B08AA600CA88B143AB11880C2806",
INIT_12 => X"055412D4481128C4CC012A66F304553096004B61BD8068B92400D0004E303689",
INIT_13 => X"589C48082C006A9057CA4385809520F07830001AC2173B00E162563454C40804",
INIT_14 => X"00460848952220592745AC11A544B1BF006850840180A00E1C81900C4190E160",
INIT_15 => X"22088220882208822088220882208CD888088D940D2A3A9D5002001300800C8C",
INIT_16 => X"0080200882208822088220882208822088220882208822088220882208822088",
INIT_17 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_18 => X"FBDFD1FE3EFBD7BBEFBEFA0A245120000000007FFFFFFFF20080200802008020",
INIT_19 => X"F3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF7FFBFAFBBBEFBEFBEFBF7",
INIT_1A => X"CFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCF3CF3CF3C",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000007F3F9FCFE7F3F9FCFE7F3F9F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040000000000000000000000000000000",
INIT_1F => X"4BA550000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0002000087FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974AA550402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"020AA5D7FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5D00000AA007FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAA954BA5504000AA557FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5D00",
INIT_23 => X"7BFFFFFFFFFFFFFFFFFFFFFFFFFAA954BA5500020BA5D7FFFFFFFFFFFFFFFFFF",
INIT_24 => X"7AA974BA5D040200055517FFFFFFFFFFFFFFFFFFFFFFFFAA954BA5500000BA5D",
INIT_25 => X"00000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000080000000",
INIT_27 => X"FFFFFFFFFFFFFAE974AA550002010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"0BA087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550400028007FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAA954BA5D00000BA557FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5D0002",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAA954BA5504020AA5D7BFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"A974AA5D00070925D71FFFFFFFFFFFFFFFFFFFFFFFF7AA954BA5500000825571",
INIT_2C => X"FFFFFFFFFFFFFFEFF7AA974AA5D040500055517FFFFFFFFFFFFFFFFFFFFFFF7A",
INIT_2D => X"D040200008000000000000000000000000000000000000000000000003FFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"A087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550002000087FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAA954AA5D00020AA007FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5504000B",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFF7AA954BA5D00000BA5D7BFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"74AA55000200055517FFFFFFFFFFFFFFFFFFFFEFF7AA974BA5504020BA557BFF",
INIT_33 => X"FFFFFFFFFFDFEFF7AE974AA5D00154105D517FFFFFFFFFFFFFFFFFFFFEFF7AA9",
INIT_34 => X"00000000043FFFFFFFFFFFFFFFFBFDFEFF7AE954AA5D041740055557FFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000007FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(2),               -- Port A write enable input
DIA(0)   => data_write_a(22),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(22),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(2),               -- Port B write enable input
DIB(0)   => data_write_b(22),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(22),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_23_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"EF20906D902424807BC8241BC81801B97D38AD3C0800103362A6741C80A12A02",
INIT_01 => X"001FFF8409F089003B4422000D80C80106804A7951C5B9D1C828043EA28838F9",
INIT_02 => X"028406A002DC176444683862400003111001303FFC00F240D50146013B300500",
INIT_03 => X"0006C90C010203F80005DC00C52FC380BEAC25886C02034800200200A1008008",
INIT_04 => X"17DFFF8049000BFF878314BFF8488890979800002F702002BB807A068403C280",
INIT_05 => X"DA07F0000000007FF020C814380011FE5E1C2FC3E05FFFF90020000808900010",
INIT_06 => X"10004C9690A8CA008024685184097E81E872C8FFE900FC31348EFDF03BE15E22",
INIT_07 => X"402000001FFBFFFD00080200B8140011F0D8C108155542018D1A302193E94004",
INIT_08 => X"41BE1F5F80003FF0002023FFDF79000000000EFFE309606020008005FC000000",
INIT_09 => X"FC83FE1840C0902400300000000000DFFD4004040C4D32BF7C0EE860003CE680",
INIT_0A => X"10018C24110A860006C620C0312241C482B20420CC56924E2199000C00415037",
INIT_0B => X"4669070510C90C14304043040430404304043040430404304043040218202182",
INIT_0C => X"008000105400C00400100000A018000801000C024000004A940000FFDF820604",
INIT_0D => X"100152100801C17E61841950B1C10FFF57FFC02812F00429DC92C40002000100",
INIT_0E => X"10015210088528E00E02C8200A430A424202A1CAF13F214001521001CBF03F21",
INIT_0F => X"01C1C044006D0C94FB94320880603C420B8001CBF03F214001521001CAF13F21",
INIT_10 => X"30182800A018D9CA8000648528E00D12480202C86040902AC60BACDF0E02D020",
INIT_11 => X"0445C19960A00026880C006739000009B00300010AF5052419D1964419028014",
INIT_12 => X"01844068880CE72000013600600332C140004D101808458A5602E00089202911",
INIT_13 => X"41D0B9023402085020825132C8CB5B4040301009408021144CB042F880100C06",
INIT_14 => X"8E17C0D240406519400500840A9524EE38A1F80E02120018390320F050144CB2",
INIT_15 => X"01004010040100401004010040100100040040000000000001000900FBFFE000",
INIT_16 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_17 => X"0040100401004010040100401004010040100401004010040100401004010040",
INIT_18 => X"0000000000000000000000000000000000000000000000001004010040100401",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000000000000000000000000",
INIT_1F => X"4BA5D0400010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000007FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974BA5D0002000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"00010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA550002000007FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAE974AA550400000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5500",
INIT_23 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550402010087FFFFFFFFFFFFFFFFFF",
INIT_24 => X"FAE954AA5D00000AA007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA55040200008",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010000000000",
INIT_27 => X"FFFFFFFFFFFFFAE974BA5D0400010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0000010007FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAE974AA550002010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA550002",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550400010087FFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"E954AA5D0402038007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550400028007F",
INIT_2C => X"FFFFFFFFFFFFFFFFFFAE954AA5D00020BA087FFFFFFFFFFFFFFFFFFFFFFFFFFA",
INIT_2D => X"D0402010000000000000000000000000000000000000000000000007FFFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000087FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAE974BA550002010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D000001",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFFFAE974AA550002000087FFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"54AA5504000BA087FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA550400010007FFF",
INIT_33 => X"FFFFFFFFFFFFFFFFAA954AA5D04000AA087FFFFFFFFFFFFFFFFFFFFFFFFFFAE9",
INIT_34 => X"000000007BFFFFFFFFFFFFFFFFFFFFFFFFFAA954AA5D00020AA007BFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000007FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(2),               -- Port A write enable input
DIA(0)   => data_write_a(23),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(23),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(2),               -- Port B write enable input
DIB(0)   => data_write_b(23),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(23),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_24_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100600007FFF000080108004000800020000840041000080808",
INIT_02 => X"0000068002CC07400000090C080002000000103FF811F150231000520ABE4404",
INIT_03 => X"210A0600000203F80005DC00000DC3801EA000000745C4010220000000008000",
INIT_04 => X"07C5FF804900026F8780001DF8000000079800000F300002998078068003C080",
INIT_05 => X"C207F0000000007FF0000004380001FE1E1C07C3E00CFFF80000000000000000",
INIT_06 => X"0002648240F20035A0102000BD0000002802C87FC800FCAA035400001B918600",
INIT_07 => X"0000000001FBFFEC4D2B4AD0B8129063B2CC0000100042018408142F16C01848",
INIT_08 => X"008E1F5F80001FF0000000FFDF78000000000EFFE001600000000005FC000000",
INIT_09 => X"E883FE180000000000300000000000DFFD0000002A80D500000671000004A000",
INIT_0A => X"10018C0411020600048620C030020502000200000400920A2198000800404037",
INIT_0B => X"0641060400C00C00304003040030400304003040030400304003040018200182",
INIT_0C => X"000000001000C00000000000000240058000000000000000000000FFDF000404",
INIT_0D => X"E00880104809C1666594584031010FFF56FFC000104000000010440000000000",
INIT_0E => X"E0088010492064206100E81084200048C0804012500021B00880108012500021",
INIT_0F => X"04100144800803419043064900C0020501840012500021B00880108012500021",
INIT_10 => X"1018140F02C0000809408D206420530270040410004C840041A0D80054109038",
INIT_11 => X"110002C9E8010C00010480B35A0300400041020902F60002260D65B361BAA104",
INIT_12 => X"0228204300166B4060080008240593D0021800020818B06D9802F00030C02060",
INIT_13 => X"143B62023C00142800B04400095DFF90203020042108603100061516EE800C06",
INIT_14 => X"DC1180C7804400044029208301040214AE4C7C02000040206602C10B48110006",
INIT_15 => X"00000000000000000000000000000000000000000000000000000000FBFFE000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"DD5EDCF9822659B6888332000000000000000000000000000000000000000000",
INIT_19 => X"F3CF3CF3CF3CF3DF7DF7DF7DF7DF7DF3DF3DF3DF3DF4D30C2432AEBAEBFE5A15",
INIT_1A => X"C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783DF7DF7DF7C",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000F0783C1E0F0783C1E0F0783",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201008000000000000000000000000",
INIT_1F => X"4BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974BA5D0400000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"00010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000007FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAE974BA5D0000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_23 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0002000087FFFFFFFFFFFFFFFFFF",
INIT_24 => X"FAE974BA550002000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D000200000",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010080000000",
INIT_27 => X"FFFFFFFFFFFFFAE974BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000087FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAE974BA5D0400010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0000010007FFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"E974BA550002000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0000010007F",
INIT_2C => X"FFFFFFFFFFFFFFFFFFAE974BA550002000007FFFFFFFFFFFFFFFFFFFFFFFFFFA",
INIT_2D => X"D0402010080000000000000000000000000000000000000000000007FFFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAE974BA5D0400000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040200",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000087FFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"74BA5D0000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0000010087FFF",
INIT_33 => X"FFFFFFFFFFFFFFFFAE974BA550000010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE9",
INIT_34 => X"000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA550002010087FFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(3),               -- Port A write enable input
DIA(0)   => data_write_a(24),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(24),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(3),               -- Port B write enable input
DIB(0)   => data_write_b(24),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(24),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_25_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100200002000000080100004000000020000800041000080808",
INIT_02 => X"0000068002CC474000000800000002000000103FFCE302008000000880844A04",
INIT_03 => X"00000040700803FC0105DE00020DC3801EA00000040000000020000000008000",
INIT_04 => X"47C5FFC04904026F8780081DFC040000079C92484F30499299837C168003E400",
INIT_05 => X"C207F0382004407FF0000004382281FF1E1C07C3E00CFFFC090004B05000200A",
INIT_06 => X"1009015C4000000020000000390C10002802C87FC800F8000000000019810600",
INIT_07 => X"0501000001FBFFFD480A0280A816002010800001000054018408102000000002",
INIT_08 => X"0C8E1F5FA21C9FF8004000FFDF7C062031863EFFF75D78004001010DFC000020",
INIT_09 => X"E883FE180C00000000300000000000DFFF00180800000000000660100000A000",
INIT_0A => X"1001DCCC31222730A49620C030020100000200000400921A21D8000804404037",
INIT_0B => X"0641062400C00C00304003040030400304003040030400304003040018200182",
INIT_0C => X"C11160845004D04820000000000000000000000000000000940000FFDF000404",
INIT_0D => X"000800000801C0786184185031810FFF56FFC02812E0182000F2C48304418220",
INIT_0E => X"0008000000002020000008000000000800800002400001000800000002400001",
INIT_0F => X"0000010000000000900000080000000400000002400001000800000002400001",
INIT_10 => X"1000000002002000004000002020000200000000000404000000880000001000",
INIT_11 => X"010000082000000001000001080000000040000100C600800001040000040009",
INIT_12 => X"0000000100002100000000080000104000000002000000081001000000000040",
INIT_13 => X"0010200000000000001004000001080000400080000040010000001080001008",
INIT_14 => X"8C11808200400000400000C20000000420000000030280000000010000010000",
INIT_15 => X"82208822088220882208822088A20C52082081A30080000002005008FBFFF001",
INIT_16 => X"2208822088220882208822088220882208822088220882208822088220882208",
INIT_17 => X"2088220882208822088220882208822088220882208822088220882208822088",
INIT_18 => X"29432D518B45265D82BB4101000005FFFFFFFFFFFFFFFFF82208822088220882",
INIT_19 => X"24924924924924820820820820820820924820924824000A6242B4D34D7F7451",
INIT_1A => X"AC562B158AC562B158AC562B158AC562B1188C46231188C46231189249249249",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000162B158AC562B158AC562B158",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000000000000000000000000",
INIT_1F => X"4BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"02000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAE974BA5D0402000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_23 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000007FFFFFFFFFFFFFFFFFF",
INIT_24 => X"FAE974BA5D0400000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040000008",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010000000000",
INIT_27 => X"FFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAE974BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000007FFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"E974BA5D0400000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000087F",
INIT_2C => X"FFFFFFFFFFFFFFFFFFAE974BA5D0400000007FFFFFFFFFFFFFFFFFFFFFFFFFFA",
INIT_2D => X"D0402010000000000000000000000000000000000000000000000007FFFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"74BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000007FFF",
INIT_33 => X"FFFFFFFFFFFFFFFFAE974BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE9",
INIT_34 => X"000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000007FFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000007FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(3),               -- Port A write enable input
DIA(0)   => data_write_a(25),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(25),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(3),               -- Port B write enable input
DIB(0)   => data_write_b(25),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(25),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_26_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"E9264EAB20190CA3BA4997AA9002AE9C001006B0778015CFA17E0811039879C7",
INIT_01 => X"F1FFF9BB1F773C7F9BB07DFFFDD863FC5FFF3FEFFBBF9FFB22FFFBC7B9F30686",
INIT_02 => X"9B3184F8AFDEAF300029E4E300FC78A6258548EFFA71C00172082400003A2161",
INIT_03 => X"0084F0FF7FFF1FDD3FEFDCDE981DC3FF5F0D294A7B2B18A0001B9CE6CC606E73",
INIT_04 => X"0FC5DFD7EDFFD66F87FE605DDDBFF3690F9EDB7F5F7AFF639BD7DE37C2FEF591",
INIT_05 => X"F205F0F8E9D199FF76DFEE1C3FCC3FF7BE1FD7C3FFACFBFFDFF7B4FEFFDAA10E",
INIT_06 => X"042648C40179912406C1830639AFBEC14489737FDC00B13BB79DFDB83BF4112A",
INIT_07 => X"763A844769FFBFE4398E4390BB9C28B1D0F049080414583F9468D1AEFC000060",
INIT_08 => X"02C05FD7BC471FBD13D981F7DF7D7E6171AF3FEFE8A3E679FAC1FD1FFFBEB000",
INIT_09 => X"F8CFFE38FF7F6BD928F1ABB47476B5FEF9F59F5FCEEDE73FEE0EFC53B079F5CC",
INIT_0A => X"315BDDCC3B336F7C548667D47B7737AF3FD62601EDC2B66A67B9D60FE4C4427F",
INIT_0B => X"06E19F4DA0E80E903DE3035E3035E3035E3035E3035E3035E3035E981AF181AE",
INIT_0C => X"EBFBF7FEBD66DBFCA3F87501AE7B080607307DCFE1D4077B4D026FFFFBFFAFCD",
INIT_0D => X"0007E010084BCD7FF1B61B5C33813FFFFCFFC7D7D51D6F5FDCB935D7AFEBD7F5",
INIT_0E => X"0007E01001BD8020500008001F010040520201F45EC0010007E01001F45EC001",
INIT_0F => X"1DC0004600400F781429C0080000770001A001F45EC0010007E01001F45EC001",
INIT_10 => X"10003C064000E408010081BD8020600200001EC00040B02007EC09A0E0001000",
INIT_11 => X"360403E434588007200D00F88C84C081C203404B3BFD0402346235408402C080",
INIT_12 => X"07B00040091F1190982038406807C868B1000E401A08FE0012040000FC002001",
INIT_13 => X"7D00212000007C400082D81009FC08281D00001F010021560406758091454000",
INIT_14 => X"FFBFF5FA1040076065F730FC08043A903A80008320C0403C3400008860160406",
INIT_15 => X"D7F5FD7F5FD7F5FD7F5FD7F5FDFF7F7F7F77F9F761FFBFDFFDE5BFFFFF7FF005",
INIT_16 => X"7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5F",
INIT_17 => X"F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD",
INIT_18 => X"B79E923C2CD990AA7F0DDB6B910C8DFFFFFFFFFFFFFFFFFD7F5FD7F5FD7F5FD7",
INIT_19 => X"30C30C30C30C30C30C30C30C30C30C30D34D34C30C35F7AA9ABF0E38E3A8EB62",
INIT_1A => X"C26130984C26130984C26130984C26130984C26130984C26130984C30C30C30C",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000130984C26130984C26130984",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000000000000000000000000",
INIT_1F => X"4BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"02010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_23 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFF",
INIT_24 => X"FAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010000000000",
INIT_27 => X"FFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"E974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007F",
INIT_2C => X"FFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFA",
INIT_2D => X"D0402010000000000000000000000000000000000000000000000007FFFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"74BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFF",
INIT_33 => X"FFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE9",
INIT_34 => X"000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(3),               -- Port A write enable input
DIA(0)   => data_write_a(26),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(26),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(3),               -- Port B write enable input
DIB(0)   => data_write_b(26),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(26),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_27_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"00080A40000A41248002029000050A088000008242A0004404480002000A1155",
INIT_01 => X"F1FFF1C11F781C129C107DFFFE0860941E81258CA2B71C2220EC1B86E1A00002",
INIT_02 => X"183080988B2EAE00002BE001117C78C6848140CFFA0000800042008000011081",
INIT_03 => X"000000FF7CF91F1D3DEF3CDA881D23FB5C0C21085B0B0820001318C60C204C63",
INIT_04 => X"8FC51FD7EDFDD66E47EE205D1DB7F1490E5EDB7D5CBADB2385D79C3643D4E580",
INIT_05 => X"E001F0C0C991BBFC76DFEA1A3F8C3BC7391F9723FF2CE3FCD6D13096B79C8106",
INIT_06 => X"40000001000000084041830600A40C415004637FC4003021259CFDB01BF80028",
INIT_07 => X"3158954761FA3FE402088220AC1108001080400A400041018468D1A060000050",
INIT_08 => X"02005F0784411E390A4881C7BEFC5F6171CE2F8FE823E778DAC16C1FFBBC9000",
INIT_09 => X"F0C7FEBABF3F6BD108F40E04C0C084F0F8B58B5B8849673F6C0E7A01B00914C4",
INIT_0A => X"B51BFDCC39732F3554866AD57C37BEAF1C152201A4C0B6EA63AAD60B60D4427F",
INIT_0B => X"06F18FC5A0E00F0038D1030D1030D1030D1030D1030D1030D1030F0818688186",
INIT_0C => X"AB6AD7EAB962CBD8A3A83101F47E08040510768EA0C406630D0226FFE375ADE5",
INIT_0D => X"000760000843C561E5C55C42B9011FFF48FFCC57550D63564D1D2556ADAB56D5",
INIT_0E => X"0007600004BD8020100008001F010000130201E44A40010007600005E44A4001",
INIT_0F => X"1DC0000208400D781020C00800007700002005E44A40010007600005E44A4001",
INIT_10 => X"10003C064000C400018080BD8020200200001EC00000382006EC0820A0001000",
INIT_11 => X"3E0403A424108007200102E888808081C20040431BC504021462354004004080",
INIT_12 => X"07B00000015D1110102038400817484821000E400204FE0010040000FC000000",
INIT_13 => X"7D00202000007C400000F81001FC08080500001F0100005E0404758081014000",
INIT_14 => X"8DBBB5FA10400360649310FC08003A903A8000012040403C34000080201E0404",
INIT_15 => X"56D5B56D5B56D5B56D5B56D5B56D7E3D7B57B1C4E17F0944B8D596EEFC7FF001",
INIT_16 => X"6D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B",
INIT_17 => X"D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B5",
INIT_18 => X"2D0200903950C080420948E2D10E8FFFFFFFFFFFFFFFFFF56D5B56D5B56D5B56",
INIT_19 => X"00000000000000000000000000000104000000000004000E5E420000002921C4",
INIT_1A => X"28140A05028140A05028140A05028140A0100804020100804020100000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000140A05028140A05028140A050",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000000000000000000000000",
INIT_1F => X"4BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_23 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFF",
INIT_24 => X"FAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201008",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010000000000",
INIT_27 => X"FFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"E974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087F",
INIT_2C => X"FFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFA",
INIT_2D => X"D0402010000000000000000000000000000000000000000000000007FFFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"74BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFF",
INIT_33 => X"FFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE9",
INIT_34 => X"000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000007FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(3),               -- Port A write enable input
DIA(0)   => data_write_a(27),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(27),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(3),               -- Port B write enable input
DIB(0)   => data_write_b(27),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(27),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_28_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"02200AA400180030808802A900002A08001280A08A801044104A1000001818C3",
INIT_01 => X"50A00011460214428114180000882214413D0A71592A01D92213D28005210202",
INIT_02 => X"8A54800A210200111100C2110054289220810440030404010844000444410001",
INIT_03 => X"1080010208B51400007800000A000001000108C21008092000018C6295200631",
INIT_04 => X"0008000000017000000028000001610300000010000802202040012040040011",
INIT_05 => X"2000044440048880026A22000026A20000000000000000004994140203000064",
INIT_06 => X"1400922401041008004891224228810080010200040001020800000004000008",
INIT_07 => X"150B001328000001404010040084088404200020455514000224489028492201",
INIT_08 => X"00414000201800004080A0000002480B04008100011000088800081002C19020",
INIT_09 => X"000400001036584108415B4A6A694A0000100101C08200000001000190200044",
INIT_0A => X"004800210C19808400500010009110091500020B408820000200400040811600",
INIT_0B => X"40000800B00100040D8140581405814058140581405814058140580A02C0A02C",
INIT_0C => X"00200248010201008298150006210802043058C46054032981002D00201C8081",
INIT_0D => X"0000A00000400600841041108280300008000140000401028008330000800040",
INIT_0E => X"0000A000000080001000000000000000500000040A40000000A00000040A4000",
INIT_0F => X"00000006000000080020C00000000000012000040A40000000A00000040A4000",
INIT_10 => X"00000000000024000000000080002000000000000000A00000040020A0000000",
INIT_11 => X"2200000404108000000900008080808000024040152000000020000004004080",
INIT_12 => X"0000000009001010102000004800080821000000120002000004000000000001",
INIT_13 => X"2000002000000000000288000020000805000000000001420000200001014000",
INIT_14 => X"408010000000022000D610280000080000000001204000000000000820020000",
INIT_15 => X"00401004010040100401004010042024210218734CD52150A840827504000000",
INIT_16 => X"0401004010040100401004010040100401004010040100401004010040100401",
INIT_17 => X"4010040100401004010040100401004010040100401004010040100401004010",
INIT_18 => X"05822140048D2E57B1348141845C200000000000000000000401004010040100",
INIT_19 => X"04104104104104104104104104104104104104104101A6A0A0EB1861863BC422",
INIT_1A => X"2C160B0582C160B0582C160B0582C160B0180C06030180C06030181041041041",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000160B0582C160B0582C160B058",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000000000000000000000000",
INIT_1F => X"4BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_23 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFF",
INIT_24 => X"FAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010000000000",
INIT_27 => X"FFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"E974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007F",
INIT_2C => X"FFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFA",
INIT_2D => X"D0402010000000000000000000000000000000000000000000000007FFFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"74BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFF",
INIT_33 => X"FFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE9",
INIT_34 => X"000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000007FFFFFFFF8000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(3),               -- Port A write enable input
DIA(0)   => data_write_a(28),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(28),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(3),               -- Port B write enable input
DIB(0)   => data_write_b(28),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(28),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_29_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"79964E4BA01DACAB9E659792D00AAE160002829C7FDFEFCEE97C2815039D70C3",
INIT_01 => X"50BFF9AB0775343F9AB01DF80D5821FC0FFF3FEFD1AF9FF1207FFBC7B9720586",
INIT_02 => X"0D15846807D207200021C4E200D428A2018408600271C000720A0000003A2161",
INIT_03 => X"0000B0027BBF17C43E6DC05E1A0DC07D1F0000803B2819A00019084345606421",
INIT_04 => X"07CDC047A4FB526F807C681DC4B97369078249370F482E62BA414627C2FE3000",
INIT_05 => X"F204007861C088FF0EFF260407C427F19E03C7C01F8CF80749B390EA4BCA202C",
INIT_06 => X"000248C00079800406C081023B233E804488527FDC008019968D74982C94110A",
INIT_07 => X"5229000221FF8000398641903B082831D05000200000083F942850AEB4000221",
INIT_08 => X"00805FD0180E1F8C1111A0F041056A0100A11FE000916249A800B915FE82B020",
INIT_09 => X"F80C000055FF7C492840AAB45456B55E015015058665A31DA603A4539058F54C",
INIT_0A => X"000850400A11414C005005000B51158936D20601A98A204006114005C4800217",
INIT_0B => X"40201948B029029409A3401A3401A3401A3401A3401A3401A3401A9A00D1A00C",
INIT_0C => X"40B1225C1506512C83E85500AC3A080406305587A154023141006DFFF89E82C9",
INIT_0D => X"0000A01008480D3EB4A24A0C910037FFFC0007C7C0140D0B50A8218102C08160",
INIT_0E => X"0000A010010080005000000000000040520000141EC0000000A01000141EC000",
INIT_0F => X"00000046000002080429C0000000000001A000141EC0000000A01000141EC000",
INIT_10 => X"00000000000024080100010080006000000000000040B000010401A0E0000000",
INIT_11 => X"3600004414588000000D00108484C080000340483B590000202000008402C080",
INIT_12 => X"00000040090210909820000068008828B10000001A0802000204000000002001",
INIT_13 => X"20000120000000000082D800082000281D000000000021560002200011454000",
INIT_14 => X"B29450580000066021F6303C000408000000008320C000000000000860160002",
INIT_15 => X"816058160581605816058160589625662522506344FF9FCFFF62EB6DFF001004",
INIT_16 => X"1605816058160581605816058160581605816058160581605816058160581605",
INIT_17 => X"6058160581605816058160581605816058160581605816058160581605816058",
INIT_18 => X"F2DDCFFFBEFFCF07FFBFFD41800C05FFFFFFFFFFFFFFFFF81605816058160581",
INIT_19 => X"7DF7DF7DF7DF7DF7DF7DF7DF7DF7DD75D75D75D75D77FFBF3F7DFFFFFFD779F3",
INIT_1A => X"FEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDF7DF7DF7DF",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00001F7FBFDFEFF7FBFDFEFF7FBFD",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000000000000000000000000",
INIT_1F => X"4BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_23 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFF",
INIT_24 => X"FAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010000000000",
INIT_27 => X"FFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"E974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007F",
INIT_2C => X"FFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFA",
INIT_2D => X"D0402010000000000000000000000000000000000000000000000007FFFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"74BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFF",
INIT_33 => X"FFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE9",
INIT_34 => X"000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(3),               -- Port A write enable input
DIA(0)   => data_write_a(29),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(29),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(3),               -- Port B write enable input
DIB(0)   => data_write_b(29),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(29),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_30_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"FFDFF3FC3EFFF7FFFFBFFA000000000000000000000000000000000000000000",
INIT_19 => X"F3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF5F7AEBEBFBEFBEFFEFFF7",
INIT_1A => X"CFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCF3CF3CF3C",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000007F3F9FCFE7F3F9FCFE7F3F9F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000000000000000000000000",
INIT_1F => X"4BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_23 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFF",
INIT_24 => X"FAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010000000000",
INIT_27 => X"FFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"E974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007F",
INIT_2C => X"FFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFA",
INIT_2D => X"D0402010000000000000000000000000000000000000000000000007FFFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"74BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFF",
INIT_33 => X"FFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE9",
INIT_34 => X"000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(3),               -- Port A write enable input
DIA(0)   => data_write_a(30),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(30),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(3),               -- Port B write enable input
DIB(0)   => data_write_b(30),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(30),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_31_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"129000008004A00804A40000400800020000000C005FEA005800200400050100",
INIT_01 => X"A15FF18019700810180065FFFC0040801E80258CA2951C2200EC0906A0804140",
INIT_02 => X"146000808A0C060444692000402850040400408FF80000000010000000004000",
INIT_03 => X"000000FD74480B1C3D951C5A800D03FA1C0C21084B0300000012108518004842",
INIT_04 => X"07C51FC7EDFCA26E07EE001D1CB6904A061EDB6D4C30490281831C1602D0E480",
INIT_05 => X"C001F0808181117C7C95C8183FA099C7181F8703FF0CE3FC0201209010988002",
INIT_06 => X"00000000000000010001020400840C41C000617FC0003021259CFDB01BF00020",
INIT_07 => X"0000000441FA3FE400080200A810000010804008100040018448912040000040",
INIT_08 => X"00011F0780011E38004801C79E7C162231862E8FE00166704041240DF93D0000",
INIT_09 => X"F0C3FE180D89279000B00000000000D0F80088080849673F6C0E780020091480",
INIT_0A => X"1011DCCC31222730048620C4382204A608142002A440924A6188020920404437",
INIT_0B => X"0661874500E00E00304003040030400304003040030400304003060018200182",
INIT_0C => X"810040801060C04821202001A05A00040100240A80800442040202FFC3200444",
INIT_0D => X"000740000803C0616184184031010FFF40FFC407500020004C10060204010200",
INIT_0E => X"0007400000BD0020000008001F010000020201E04000010007400001E0400001",
INIT_0F => X"1DC0000000400D701000000800007700000001E04000010007400001E0400001",
INIT_10 => X"10003C064000C000010080BD0020000200001EC00000102006E8080000001000",
INIT_11 => X"140403A020000007200000E808000001C200000308C504021442354000000000",
INIT_12 => X"07B00000001D0100000038400007404000000E400000FC0010000000FC000000",
INIT_13 => X"5D00200000007C400000501001DC08000000001F010000140404558080000000",
INIT_14 => X"8C1380DA10400140640100D4080032903A8000000000403C3400008000140404",
INIT_15 => X"02008020080200802008020080200C1808008184012A08041202500AF87FF001",
INIT_16 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_17 => X"0080200802008020080200802008020080200802008020080200802008020080",
INIT_18 => X"000000000000000000000002001005FFFFFFFFFFFFFFFFF02008020080200802",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"000000000000000000000007FFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000000000000000000000000",
INIT_1F => X"4BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_20 => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_21 => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_22 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_23 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFF",
INIT_24 => X"FAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000",
INIT_25 => X"000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"A5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010000000000",
INIT_27 => X"FFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974B",
INIT_28 => X"010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFF",
INIT_29 => X"FFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402",
INIT_2A => X"FFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFF",
INIT_2B => X"E974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007F",
INIT_2C => X"FFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFA",
INIT_2D => X"D0402010000000000000000000000000000000000000000000000007FFFFFFFF",
INIT_2E => X"FFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5",
INIT_2F => X"0007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFF",
INIT_30 => X"FFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201",
INIT_31 => X"FFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFF",
INIT_32 => X"74BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFF",
INIT_33 => X"FFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE9",
INIT_34 => X"000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(3),               -- Port A write enable input
DIA(0)   => data_write_a(31),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(31),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(3),               -- Port B write enable input
DIB(0)   => data_write_b(31),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(31),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


end;