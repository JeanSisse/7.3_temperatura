library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_misc.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library UNISIM;
use UNISIM.vcomponents.all;

entity ram_master is
	port(clk             : in  std_logic;
        address_a       : in  std_logic_vector(31 downto 2);
        enable_a        : in  std_logic;
        wbe_a           : in  std_logic_vector(3 downto 0);
        data_write_a    : in  std_logic_vector(31 downto 0);
        data_read_a     : out std_logic_vector(31 downto 0);

        address_b       : in  std_logic_vector(31 downto 2);
        enable_b        : in  std_logic;
        wbe_b           : in  std_logic_vector(3 downto 0);
        data_write_b    : in  std_logic_vector(31 downto 0);
        data_read_b     : out std_logic_vector(31 downto 0));
end; --entity ram     

architecture ram_master of ram_master is
signal enable_a_lo       : std_logic;
signal wbe_a_lo          : std_logic_vector(3 downto 0);
signal data_write_a_lo   : std_logic_vector(31 downto 0);
signal data_read_a_lo    : std_logic_vector(31 downto 0);
signal enable_b_lo       : std_logic;
signal wbe_b_lo          : std_logic_vector(3 downto 0);
signal data_read_b_lo    : std_logic_vector(31 downto 0);
signal enable_a_hi       : std_logic;
signal wbe_a_hi          : std_logic_vector(3 downto 0);
signal data_read_a_hi   : std_logic_vector(31 downto 0);
signal enable_b_hi       : std_logic;
signal wbe_b_hi          : std_logic_vector(3 downto 0);
signal data_read_b_hi    : std_logic_vector(31 downto 0);
signal address_a_reg     : std_logic_vector(31 downto 2);
signal address_b_reg     : std_logic_vector(31 downto 2);
signal enable_a_lo_256       : std_logic;
signal wbe_a_lo_256          : std_logic_vector(3 downto 0);
signal data_write_a_lo_256   : std_logic_vector(31 downto 0);
signal data_read_a_lo_256    : std_logic_vector(31 downto 0);
signal enable_b_lo_256       : std_logic;
signal wbe_b_lo_256          : std_logic_vector(3 downto 0);
signal data_read_b_lo_256    : std_logic_vector(31 downto 0);
signal enable_a_hi_256       : std_logic;
signal wbe_a_hi_256          : std_logic_vector(3 downto 0);
signal data_read_a_hi_256   : std_logic_vector(31 downto 0);
signal enable_b_hi_256       : std_logic;
signal wbe_b_hi_256          : std_logic_vector(3 downto 0);
signal data_read_b_hi_256    : std_logic_vector(31 downto 0);
begin
process(clk)
begin
if rising_edge(clk) then
	address_a_reg <= address_a;
	address_b_reg <= address_b;
	end if;
end process;
data_read_a <= data_read_a_lo when (address_a_reg < x"0001000"&"00") else
data_read_a_hi when ((address_a_reg >= x"0001000"&"00") and (address_a_reg < x"0002000"&"00")) else 
data_read_a_lo_256 when ((address_a_reg >= x"0002000"&"00") and (address_a_reg < x"0003000"&"00")) else 
data_read_a_hi_256 when ((address_a_reg >= x"0003000"&"00") and (address_a_reg < x"0004000"&"00"));
data_read_b <= data_read_b_lo when (address_b_reg < x"0001000"&"00") else
data_read_b_hi when ((address_b_reg >= x"0001000"&"00") and (address_b_reg < x"0002000"&"00")) else
data_read_b_lo_256 when ((address_b_reg >= x"0002000"&"00") and (address_a_reg < x"0003000"&"00")) else 
data_read_b_hi_256 when ((address_b_reg >= x"0003000"&"00") and (address_b_reg< x"0004000"&"00"));
enable_a_lo <= enable_a when (address_a < x"0001000"&"00") else '0';
enable_b_lo <= enable_b when (address_b < x"0001000"&"00") else '0';
enable_a_hi <= enable_a when ((address_a >= x"0001000"&"00") and (address_a < x"0002000"&"00")) else '0';
enable_b_hi <= enable_b when ((address_b >= x"0001000"&"00") and (address_b < x"0002000"&"00")) else '0';
enable_a_lo_256 <= enable_a when ((address_a >= x"0002000"&"00") and (address_a < x"0003000"&"00")) else '0';
enable_b_lo_256 <= enable_b when ((address_b >= x"0002000"&"00") and (address_b < x"0003000"&"00")) else '0';
enable_a_hi_256 <= enable_a when ((address_a >= x"0003000"&"00") and (address_a < x"0004000"&"00")) else '0';
enable_b_hi_256 <= enable_b when ((address_b >= x"0003000"&"00") and (address_b < x"0004000"&"00")) else '0';
wbe_a_lo <= wbe_a when  enable_a_lo='1' else x"0";
wbe_a_hi <= wbe_a when  enable_a_hi='1' else x"0";
wbe_b_lo <= wbe_b when  enable_b_lo='1' else x"0";
wbe_b_hi <= wbe_b when  enable_b_hi='1' else x"0";
wbe_a_lo_256 <= wbe_a when  enable_a_lo_256='1' else x"0";
wbe_a_hi_256 <= wbe_a when  enable_a_hi_256='1' else x"0";
wbe_b_lo_256 <= wbe_b when  enable_b_lo_256='1' else x"0";
wbe_b_hi_256 <= wbe_b when  enable_b_hi_256='1' else x"0";



ram_bit_0_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"ED39BA795990D275FB4A6E96ACC4731DEA4598B0AFB54867F6EE4618C3749807",
INIT_01 => X"58A0047D8607944AC7DA180001ECA2544042106208408208C20022E9173734B3",
INIT_02 => X"9F775E7CB273E6CCA7DAAF00001000000478020113C9C38E09FB7CCCDD9F203E",
INIT_03 => X"441406267B4CB04443163C91110C58F24A31000B8028A810A3D0F8B169A01006",
INIT_04 => X"0005802424830120024121209088809DF81454ACA01E03501D0A3B91E00F0A00",
INIT_05 => X"E0F001CC00012034C20B0232838F80D001C0100AEC83C008EF101A034C8CC300",
INIT_06 => X"908A0D058584A45164BE6E58A000000583F08459A2000DA8C40F003C80030780",
INIT_07 => X"E6CCAFDC3870EEEEC44E2BDFE220094D03022210C011C103FB860B28000007C9",
INIT_08 => X"080032BF07C7C1FC3F87253D96C45557ABFF070C19D62C9065EAF36919FCB273",
INIT_09 => X"DB0009EF68EC0000045082984202002DB93119096025040581B9691E8A88262C",
INIT_0A => X"8014546E000344A0488111084048E082D0ED020133A6BF200005F60820B88206",
INIT_0B => X"28000947E16656074EA560F08054490B01280A26900C4800814069B0C8888008",
INIT_0C => X"03DCF03CCF03DCF03CCF03DCF03CCF038E780C6781C008500804708A42255A88",
INIT_0D => X"7095352BD2A90515A1CA44E7EA84B00001010012008700624187C09C0E707CCF",
INIT_0E => X"0B92800224008AE09F8942C48D1BC49120489024481225058860128543287291",
INIT_0F => X"038ABACB83C7E03EA5FF83C002783F103EA5FF83C002783F0120847A70470C7E",
INIT_10 => X"0380230F2D7C103EACFF83C002783F103EACFF83C002783F310BBF7EFC2B80C2",
INIT_11 => X"BF7EFC61E01804E1E6EA1E3FA01FD97EFC4B80E008C7C2F678FF023FAF5BD987",
INIT_12 => X"CC8E8320C4DAC9220C6B2FF22EF72ADDE6F1A67C80600C2683E0EF8AE1F1F10B",
INIT_13 => X"5C00FE651C6104C6D6400FFFB01FC0000FC07EE42FA7C07F22CE3082636B801F",
INIT_14 => X"C08FDF4195C0C2038A7C6CAFA7E289F9BA4570380131CAFB2003F9D190A4189B",
INIT_15 => X"9FE635BE11B7F0308D4A80092E0FC1FC662FA7E283FF68A8F0080AE1DDA8BE9F",
INIT_16 => X"12058312C1241140A056954AB0D680D000003350013024179498C2EC6B9270AE",
INIT_17 => X"2048120481204812048120481204812048120481204812048120481204812048",
INIT_18 => X"0481204812048120481204812048120481204812048120481204812048120481",
INIT_19 => X"2859400000000000000000120481204812048120481204812048120481204812",
INIT_1A => X"082218821390771C71C557C449F3898E09B56C74DAB16787E0760E5D1CF13043",
INIT_1B => X"7C3E1F0F87C3E082082082082082082082082082082082082082082082082082",
INIT_1C => X"87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F8",
INIT_1D => X"D7BD7400000000000000000000000000000000000000000000061007FE00000F",
INIT_1E => X"A2D1574005D0428A10A2AAA8BEF552EBDFFF557BC01FF5D7BFFEBA5D55555EF5",
INIT_1F => X"AFFFFC2000AA8428AAAFFAAA8BFF00002AA10FF802ABEFA2D16AA00F7FBE8A10",
INIT_20 => X"EFFF8002010002EAAAAAAAD1555FFFFAEA8B550051401450055575FF00517DEB",
INIT_21 => X"5FF0855575455D2AA8BFFA2D1575EF5D5555545FFFBE8A00087FC20BA5D2A975",
INIT_22 => X"8A00FFAE800AA082A820005D2E974BAA2D140145A2842AA00A284021FF5D0415",
INIT_23 => X"7FFEF000017400FFD1555FF007FFFEBA55042AA00000017400FFAABFEBAFF802",
INIT_24 => X"000155F7D540000F7FBFFE105D7BE8ABAA284000105D0428BFFA2FBFDFFFA2D1",
INIT_25 => X"7BFAEBA5551501D51C5FC7E00000000000000000000000000000000000000000",
INIT_26 => X"6D16AA28EBF5EDA38AADE1543849557D492BF8E2DE00552EBFFC7552BC01D75D",
INIT_27 => X"A85400E00E38A175FDE3F5C002DAAD42DAAAF784AFA82BC042DF47E3D1F8028B",
INIT_28 => X"50021C0092490E904BAFFD550A90FFA495FC7A05B555C257AAA8B45007540000",
INIT_29 => X"02402ABD4AD1D0E175D7140B455D516A1EAB45E2A000B4748717A095F571EAA1",
INIT_2A => X"4A8BC0ABFF7D03A17D1D5147540B454AA080038E9748542AE3D0051C7B6F02DA",
INIT_2B => X"D4B8FC7BFFFD2168B68F57492F505FF5FA550490BFA482B420B8428A3DA85400",
INIT_2C => X"0000000000000000000016ABD554201543A1EDE9016D4AAB454AF400547ABFB6",
INIT_2D => X"EBDF55556BC35E7557FE8AB25D11415FD0151614000000000000000000000000",
INIT_2E => X"6CBEA41D7D3DECFAF7D43FABAAAD57DEBAAAFFD74AA04547EE18D680BE9A55D2",
INIT_2F => X"78228E5000EA422E10439C1FBCD282351BDAAF9C20AAAABCBEB1DFF803FC5959",
INIT_30 => X"284683ABBDD7DEAA100069C14B25495A00F38EBAC0E198B9760501805357547D",
INIT_31 => X"8FE6A755ED8EFEFE41B2D17EAF02552BC0545556BD61E501001DF5DD3EBA31E6",
INIT_32 => X"F922ACA8AB8283C8310FAB1588916D3861C0422C44082B52A81550A828141440",
INIT_33 => X"DBCD7D262E5AFAC4B6AADDD562AF57D7C369AF25495A23068A8301BA7FB95556",
INIT_34 => X"FE0000003FE0000003FE0000003FE0000003FE03D5789700282E9FEFB501EA5F",
INIT_35 => X"3FE0000003FE0000003FE0000003FE0000003FE0000003FE0000003FE0000003",
INIT_36 => X"00000000000000000000000000000000000000000000000000000003FE000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000020",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(0),        -- Port A data input
DOA(0)   => data_read_a_lo(0),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(0),        -- Port B data input
DOB(0)   => data_read_b_lo(0),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_1_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"212C001411984004084D000508C53810A03D1450E839B003342114428A000807",
INIT_01 => X"08000010400A0008010600000084004000400002000000000000000000140000",
INIT_02 => X"484DEBA0111800C004400D000000000028800001CC404E6008B4933336880010",
INIT_03 => X"650C00000848A0423183089008C604224200000100A200002C280810098C0001",
INIT_04 => X"00000004208B00200E010800006667BE7000102C00080000040012010000080C",
INIT_05 => X"0080000000002020600100208D04414000800000000200004800080000800200",
INIT_06 => X"0000CB008084001C481040080000006050402008080000800488000000020400",
INIT_07 => X"00C00843060C19E2300221036000004400208000400041034001042000000101",
INIT_08 => X"08000290248CC84E0801318000C45555087C60C182B1592FE26AD7B7F7A01118",
INIT_09 => X"D8000AA220480040050080085200001161020001202100008008611687A28000",
INIT_0A => X"2640440000000080081040000040208300041000008004104006840000B80004",
INIT_0B => X"78051112A80000840200202112800001010828008000000105400020082800A8",
INIT_0C => X"2358323483234832358323583234832340190AC191A52801000C1002020883C2",
INIT_0D => X"4417882F82C00181707044212080300001002102010244800400C80C80323183",
INIT_0E => X"0B92C000000000400001004200004010200810040802040080200284401C1C11",
INIT_0F => X"00000043C2016000000F03C00280030000000F03C00280030000004860C60C0C",
INIT_10 => X"03800000049C0000000F03C00280030000000F03C002800321080000BC2380C2",
INIT_11 => X"00007861E0180000002A9001A00000007C4380E00000001E002300000008D187",
INIT_12 => X"4C0C81200009480010280340000008082430A07C80600C000000900861001108",
INIT_13 => X"34400241186100004A500007B00FC000000000E4A402C001208C308000268800",
INIT_14 => X"C0001E0181C0C200000025A400A200812A4070380000000B2500098190240001",
INIT_15 => X"04A0002410A170300C4A800800000020E22400A200096828F008000000AA9002",
INIT_16 => X"0200820040041002000010080014000000002340002004118010C22861400008",
INIT_17 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_18 => X"0080200802008020080200802008020080200802008020080200802008020080",
INIT_19 => X"0A04000000000000000000020080200802008020080200802008020080200802",
INIT_1A => X"8AB2048634B03249249604C061028A46BABEFC54A08170062002340C7452B500",
INIT_1B => X"DD6EB75BADD6EAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA8A28A28A28A2",
INIT_1C => X"A5D2E974BA5D2E974BA5D2E974BA5D2E974BA5D2E974BA5D2E974BA5D6EB75BA",
INIT_1D => X"AAAAAA00000000000000000000000000000000000000000000181FFFFF00000B",
INIT_1E => X"5D7BE8ABA5D557DFEFFFD17FEBA00042AAAAFFFFFFE00FF843DF45FFAE95555A",
INIT_1F => X"F552A800AA5555575FFA2AE820BAFFAEBFF555500155EF552E975FFF7D168BEF",
INIT_20 => X"00A2FBEAABA5D55420AA00002AA00AAFBE8B55A280175455D002AA00A2AABDFE",
INIT_21 => X"5FFAA802AAAAFFAA801EF00517FFFFF7D56ABEF0004155550004154105D556AA",
INIT_22 => X"75FF08557DEBAA2FBEAAAA552E955EF5D0415410A2AE97545A2AE954BAF7FBD7",
INIT_23 => X"7DF55A2AEBDEAAFFFFC20AAFFFFFFFFFAAD5555FFFFAEAAB55A2D168B555D555",
INIT_24 => X"0000BAFFFBE8A00087FC20BA5D2A975EF5D0002010552E820AAFFD57FF55F7D1",
INIT_25 => X"8A38F45F7AA9217FA380AD400000000000000000000000000000000000000000",
INIT_26 => X"52E975EFFFDF68BFF557BEAA925551785D7BFD5EFE3F08002FA92EBA5FDE28FF",
INIT_27 => X"41017DE92BF8E3AA824924870BF5551555C7A28A821EFE3AABAE38005B575D75",
INIT_28 => X"8005A1041055716DB7DB6FBEFEA81C55D0A0516802AA28BEF5EDB7DAA8A15438",
INIT_29 => X"EF1C043FE28E3FBD55FFAADE2DAAAE3A5C51C71C042DF45A3D1D00281E8A1056",
INIT_2A => X"B45B47F6FB55A95555E90F78E17F52FEF5EDA82FD249057F080417492AAAFC7F",
INIT_2B => X"8AAAA95B7AF45FF8F7DFEDFFAFF8E005FAE92A3AE3DBFF57FA2DF555D257AAA8",
INIT_2C => X"000000000000000000000A8F571EAA150021C0092490E905FFFD0550BD75C5FF",
INIT_2D => X"43DE00A2C57DE08FFAAA8B55F7EE801F7F2849EE000000000000000000000000",
INIT_2E => X"AE29F067155543A15D2E955EFFFFBEABEF557FEAA10595169BED83D1EBCA8000",
INIT_2F => X"FD57DEEAAA15976EB0444BFEB086808A8E3082C954BA5D7DD6145AAAA821A6AA",
INIT_30 => X"FFD55D6107782001FF0812000A255D57FFBEF3B97EEAB2C40217B9778428ABAF",
INIT_31 => X"F003F17418AEE817B540D11CA80BAAFA825EFAABEBCA18FE803755D08079EB47",
INIT_32 => X"EBA2D757547D7862AF57ABFFCABE5553FD5FBEFE86353EFFFD03FE027500035F",
INIT_33 => X"1F70C6AA04537957D6FB4807FFFB45F7EFFDA58FF2AA88A0F3C5014018AC28BD",
INIT_34 => X"00000000000000000000000000000000000000B2DD7DEAA100069C14B25495A0",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000020",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(1),        -- Port A data input
DOA(0)   => data_read_a_lo(1),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(1),        -- Port B data input
DOB(0)   => data_read_b_lo(1),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_2_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10E44660018259B2843913100062C98004802322D3E030235201006009B2812",
INIT_01 => X"8005A188084900481C8024A542400340404000720885800802000906E4910204",
INIT_02 => X"5C010802020408040C640850AA055254090541A111240A104A0000000908B510",
INIT_03 => X"0C1101108800004481060A001204102802156020218808002440850008C80550",
INIT_04 => X"8840C08022050400482812C21C0804040968987810688899444090C10A124A69",
INIT_05 => X"4885109105400029210000010340086856B141212252142242A068A080106372",
INIT_06 => X"0082006020044004C240108005540A400440880000908281302852A6710AA420",
INIT_07 => X"08040860400008C022402502100AA00004404B5075460111044014002AAA2100",
INIT_08 => X"382A885244145048C860214020040505487C0800049000004220000110820204",
INIT_09 => X"88582833A24105145404D4694E710A832488C000002205C23600408C872A2A12",
INIT_0A => X"A211100D0828800A022025A81AE3048228002A7080012082C15C859D5073D520",
INIT_0B => X"3E00659A308809540009202A5820068019108A88B1D007285082002B10416820",
INIT_0C => X"1A0021A5021A1021A5021A1021A4021A0010C2010D010887470912171342A683",
INIT_0D => X"89180010084038220410042B2000715A0400200080623400380886086021A002",
INIT_0E => X"40000554015500481000300000C4480810000002040000000913000004C18402",
INIT_0F => X"00000001440002C052000400028000154052000400028000200501CCD28D206A",
INIT_10 => X"00000000048015405200040002800012C05200040002800014E0000100002000",
INIT_11 => X"00010008000000000002A0000D80060100004000000000180000294010240020",
INIT_12 => X"1011000000090000A310000881080102000A0000400000000000900002000684",
INIT_13 => X"204E008240000000483250000800000000000004E00007004120000000240A60",
INIT_14 => X"254000806000000000000560000942004110000000000000254C020220000001",
INIT_15 => X"00108840600002080200000000000020806000093000040000000000000B8000",
INIT_16 => X"008022200100000020A89068084D402120AAC005C00000000000000005408140",
INIT_17 => X"0802008020080601806018060180200802008020080601806018060180200802",
INIT_18 => X"8040080000800008000180401804018040080000800008060180601806018020",
INIT_19 => X"A2852F81F81F83F03F03F0018040180401804008000080000800018040180401",
INIT_1A => X"04609D21808205965965D64CC5B60040138D70C030B54284722B291C50C7D100",
INIT_1B => X"4A25128944A25041041041041041041041041041041041041041041041041041",
INIT_1C => X"44A25128944A25128944A25128944A25128944A25128944A25128944A2512894",
INIT_1D => X"055400000000000000000000000000000000000000000000001E1007FFE3F009",
INIT_1E => X"FF843DF45FFAEBDF55082A82155082AAAA10F7FFEAB455500175FF5D2A800100",
INIT_1F => X"F082ABDF455D7BD5545F7D5574BAFFD16AAAAA28428ABA000428AAA5D7FD7400",
INIT_20 => X"455D7BEAABA5D2A97545552E975FFFFD168AAA5D7BE8BFF5D557FFEFFFD16ABE",
INIT_21 => X"5555555555FFA2AE820BAFFFFEAABA5555554BA5D0417545F7D56AAAAAAFBEAB",
INIT_22 => X"AA00AAAEBDFFF08042AABA087BD54BA08043DEAAFF843FF5508517FF55552A95",
INIT_23 => X"82010AAD1401FF002EBFF45A2FBFDFEF00042AA00AAFBEAB5500003FF5500002",
INIT_24 => X"0000BA0004155550004154105D556AA00A2FBEAABA085542145082A800BA002A",
INIT_25 => X"00155FF552A87410007145400000000000000000000000000000000000000000",
INIT_26 => X"8002FABA4171D5400FF8A38F45F7AABA57D0000855FD1C2AAFA00EBA5E8B7D55",
INIT_27 => X"555178FD7BFD5FDFFA0020BFF78417BD5545F7F1554AAF7D16DABABFF57DE920",
INIT_28 => X"DFFDF6DAAAAAF1EFB6D417BEFA901C2E97F40552E975EFEBDF68ABA557BEAA92",
INIT_29 => X"7DA3FBD21C7492E9256D555B555C7A2ABC20AAE3AABAE38005B574AA49041756",
INIT_2A => X"B7D1E803AF6D400028E02AB8A3A012540E2AABABC75D043A00003FE10E3802DB",
INIT_2B => X"8B7D0AAA800AA147085000FFDA001C7B47BFABC7BFFF7AB4714042AA38BEF5ED",
INIT_2C => X"000000000000000000000821E8A10568005A1041055716DA38B6FBEFFEF1C0EB",
INIT_2D => X"EBDE00AAC16ABEF5500155EF552A954000855544000000000000000000000000",
INIT_2E => X"D57DE0AFAD1EBEB400043DEAA085555400FFAAAAB55F7AEA8BF77004147EF5D2",
INIT_2F => X"AFBEABAF557FEA8515951E8B4D83D1EBDFF082CBDFEF005756145FFD5574AAF7",
INIT_30 => X"5951550100004155EFF7FFFDE08AA557FFFF083FFCEB95104210405D2E955EFA",
INIT_31 => X"A002A3FE18AE803CBE7A3C014351082E951FF5D7FD6145AAAA820A2AAAD29E00",
INIT_32 => X"45550028ABAFFD17FFED01001FFEF5542ABEB2AA848AAA2552EA8ABA7551400A",
INIT_33 => X"EBAF3F95EEE95C00B7CF12AAA800BA551417105FFFFC21555556EAB4CD6D5EAD",
INIT_34 => X"00000000000000000000000000000000000000187782001FF0812000A255D57F",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000040",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(2),        -- Port A data input
DOA(0)   => data_read_a_lo(2),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(2),        -- Port B data input
DOB(0)   => data_read_b_lo(2),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_3_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"210C00A20020000108430020001600B815602110494074133520400E02B92206",
INIT_01 => X"A00C9BC048800168240442C99E004B61404040028804A0080A000D16A0990A08",
INIT_02 => X"4809A902031800444445089866E331352180D468B8200E600C0081110B80ACD0",
INIT_03 => X"6D0A60100C000142B1A30A040AC68428320006010A80881068A80D401C846330",
INIT_04 => X"482218076809C03B24841CD92CDD5A440209127847294C042640102107102D04",
INIT_05 => X"0583180353202129000104E40B04644B32A86D24014A0D204063297092000E34",
INIT_06 => X"0120D000808040181B5000A014CC662814442808805A52C03068280004629414",
INIT_07 => X"00444841428409C038B02523041994001C644C82732001190000B400E6640901",
INIT_08 => X"E8E64010248C4A5AA040308000440005487C285284B1D00BC22AC005B2820318",
INIT_09 => X"A8D588362040534C3B0E80A9DB742641620AC281826816925040408483008A10",
INIT_0A => X"040450A1439800840C32264119D004860110104004010001E732C0DF80F3B174",
INIT_0B => X"7C8575909088A4D010202422520090840B4028209AC1111954DA902230010002",
INIT_0C => X"032920329203692036920329203392036C900BC9019528100A0D30024BC8A283",
INIT_0D => X"446A101C05C0088A42D001032000333931001902010234888C68804808A03692",
INIT_0E => X"8601CCCC8B33004C0001004240140018380818040A0706009000028000903401",
INIT_0F => X"00000120000006000000000020004011000000000020004010072CC92416414C",
INIT_10 => X"0000001002001400000000002000401380000000002000401070000000000000",
INIT_11 => X"00000000000000000110000001A0000000000000000005002000244000000000",
INIT_12 => X"00000000010402049910000011000500000000000000000008000020000002C0",
INIT_13 => X"805500000000000820133000000000000000810000000C000000000004100B20",
INIT_14 => X"0530000000000000000180000011060000000000000001040154000000000020",
INIT_15 => X"0000820062000000000000000000040100000010700000000000000002400000",
INIT_16 => X"0680C2A05104100280A8D06C004044230B998021002004000001011000380000",
INIT_17 => X"280C0280C0280803808038080380803808038080380C0280C0280C0280C0280C",
INIT_18 => X"00C0280E0200C0280E030080380A030080380A030080380C0280C0280C0280C0",
INIT_19 => X"8A145D54AAB556AA9556AA830080380A030080380A030080380A0200C0280E02",
INIT_1A => X"04A20E858000049249240540430303C0C78C706428A141046016224C58629502",
INIT_1B => X"EA753A9D4EA75249249249249249249249249249249249249249041041041041",
INIT_1C => X"46A351A8D46A351A8D46A351A8D46A351A8D46A351A8D46A351A8D46A753A9D4",
INIT_1D => X"A8400000000000000000000000000000000000000000000000001007FEB6FECD",
INIT_1E => X"5500175FF5D2AA8A10005540155087BEABFF552ABDF45A2D16AAAAF7D540000A",
INIT_1F => X"000556AB55552ABDE00AAD140010F7D17FF45A2AA82155082AAAA10F7FFEAB45",
INIT_20 => X"55557FEAA10007FEAABA000428AAA557FD7400FF843DE00FFAEBFF55082A8201",
INIT_21 => X"A105D7BD5545F7D5574BAFF802AA00A2D168ABA085568BEFFFAE820000855421",
INIT_22 => X"FFEFF7D56ABEF557BD74BAFF8402145A2AEBFFEF552EAAABA5D0028BEF082AA8",
INIT_23 => X"3DEAAAAAA95410F7803FFFF55556AAAA552A975FFFFD16AAAA5D7BC01EF5D557",
INIT_24 => X"0000105D0417545F7D56AAAAAAFBEAB455D7BEAABA5D2A974005D55574005504",
INIT_25 => X"DF6FABAFFD547010AA8407400000000000000000000000000000000000000000",
INIT_26 => X"C2AAFA28EBF5E8B7D5500155FF552AAF0100071455451C75EABC74174BAF55B6",
INIT_27 => X"F7AABAF7D00009543D1C556AB6D4124BAE10BED542010FFD57AF55AAF5D756D1",
INIT_28 => X"FEBA0870281C5F4716D5D7FEDA3A0955FF48208002FABA4171D5400FF8A38F45",
INIT_29 => X"BA15203FFFF002AAFA384171D5545F7D0154AAF7D16DABABFF57DE92005F6ABF",
INIT_2A => X"ABA417BC01D7555178FD7BFD5FDF571575D24BA438E021D5B6A4BAFFF5D2EB8E",
INIT_2B => X"FE005D5B52428410E3AE92E3A490410EB843ABD71551FFE02552A975FFEBDF68",
INIT_2C => X"0000000000000000000003849041756DFFDF6DAAAAAF1EFB6D417BEFBD71C24B",
INIT_2D => X"56AB45081028B55FFFFFFEBAFFD557400A280144000000000000000000000000",
INIT_2E => X"D56ABF5AAD15455F5D2EBDEAAA2D16ABEF5500175EF552ABDE000855545455D5",
INIT_2F => X"85555400FFAAAAB14F7AE28BF77004146BA557DEABEF00002BE10FFD540000FF",
INIT_30 => X"F2D1EAEBA007FEABEFAA84174BA557FD55EF5D3BFEEB35055DEE1000043DEAA0",
INIT_31 => X"5FFAA28BF7592EABE0A0804ABFFB082EBDEAA005556145FFD5574AAF7D47DE0A",
INIT_32 => X"105D2E955EFAAFBE8AAA547FE21550853E8B4FABD5EBFF75D55420AA82AA8015",
INIT_33 => X"FFF087FFCEF90104B780A557FC20AA082AAAE10AA8000000A2AC2ABFD2151EB8",
INIT_34 => X"00000000000000000000000000000000000000AA0004155EFF7FFFDE08AA557F",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000020",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(3),        -- Port A data input
DOA(0)   => data_read_a_lo(3),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(3),        -- Port B data input
DOB(0)   => data_read_b_lo(3),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_4_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10804002061080A284201081034809800A00230350007833422C82904204006",
INIT_01 => X"204398001038084C0420050E12100368403008418984014902030906A0910204",
INIT_02 => X"480108A000000000446118E01E80F00A41043118680402000800000009882390",
INIT_03 => X"065140108C0000400026480000009120270072E03000000030808840888100F0",
INIT_04 => X"9100EB826A155C1AF0B81C160033B9440222BA281AE0D8B8E02010E81C22E821",
INIT_05 => X"5C0F20B36F08010924C084C501441C4CF21C48B133483C8042EAE1E0101074C4",
INIT_06 => X"010290102005118043508020543C1E480002820085D9C0C70000F2AA375A6071",
INIT_07 => X"00000860008008D200102502000786000C00C8025C00091B0400B00061F84020",
INIT_08 => X"991E02100C84C0480020010000004404087C8010009800004022800110000000",
INIT_09 => X"B83D6A2620418F7CF8084082425D01D123C2C040816A00708840408483000011",
INIT_0A => X"BB1B585C1304E002000064010E4007F7210010500400400800F0CC249C1401C1",
INIT_0B => X"7A04331814080458100134201A2086441B50A088078106C14540906D004068A0",
INIT_0C => X"186921829218692182921829218692182090D3490C352296CC60B11357088682",
INIT_0D => X"411050002500A9200A8014010001370F03080980912204883C28864860A18A92",
INIT_0E => X"C40903C1430F20025040102200441A040906008300418050501341208002A005",
INIT_0F => X"0000012004000BC01200000020004008C012000000200040000721CD86146108",
INIT_10 => X"0000001002000A40120000002000400DC01200000020004004D4400000000000",
INIT_11 => X"40000000000000000110200007600401000000000000050020005D4010040000",
INIT_12 => X"1010000001040004A3B000018008850200080000000000000800002002000650",
INIT_13 => X"80360082000000082034300000000000000081004000170041000000041005E0",
INIT_14 => X"2B200080400000000001804000192000401000000000010400F8020200000020",
INIT_15 => X"00114A00200002080000000000000401004000085C0000000000000002410000",
INIT_16 => X"459040281181004A8088986D045C24436C7840A6180300082001211304208140",
INIT_17 => X"1106409004110240904411024090040106419004010640900411064090440102",
INIT_18 => X"9024010041104409024190240104411004190240906411024190440102419004",
INIT_19 => X"021074B261934D964C3269C09064110040104409064190240104401004190640",
INIT_1A => X"8A74C1323433345145130282E6228A063807E05000143842130115063450454A",
INIT_1B => X"8D46A351A8D46AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA8A28A28A28A2",
INIT_1C => X"A0D068341A0D068341A0D068341A0D068341A0D068341A0D068341A0D46A351A",
INIT_1D => X"50015400000000000000000000000000000000000000000000001007FEA73FC1",
INIT_1E => X"A2D16AAAAF7D568A00AA8400000AAFFC21FFF7D542000FFAE821FF552EAAA105",
INIT_1F => X"0AAAE820BA550015400087FD74BAFFD540000F7D155555087BEABFF552ABDF45",
INIT_20 => X"AAF78015545FFD555555082AAAA10F7FFEAB455500175FF5D2AAAA1000554000",
INIT_21 => X"B45552ABDE00AAD140010F7D17FF45A2FBC2000A2FFC21555551554005D2EA8A",
INIT_22 => X"FF55082E82145A280001EFF78402145A2AE801555D2E95555552E9741000556A",
INIT_23 => X"7DF45557BD5410F7D555545F7AA97410000428AAA557FD5400FF843DE00FFAEB",
INIT_24 => X"0000AA085568BEFFFAE82000085542155557FEAA10007FEABEFAAD1400AA5D51",
INIT_25 => X"AA801EF4920AFA10490A17000000000000000000000000000000000000000000",
INIT_26 => X"C75EABEF4124BAF55B6DF6FABAFFD56F010AA8407428A2F1C01FFF7D142028EB",
INIT_27 => X"552AAFA10007155428A2AE850925D0010400087FD24AAE3DF47010E38E051451",
INIT_28 => X"55D51524004920ADA82EB8A12555EBFB4717D1C2AAFA28EBF5E8B7D5500155FF",
INIT_29 => X"55492A850381C5F6AB6D4124BAE10BED542010FFD57AF55AAF5D7410A2FBC015",
INIT_2A => X"400FF8A38E00F7AABAF7D0000955FDB684051D7F7840517DA2A4871554124925",
INIT_2B => X"75EFBED5400825D557FF55007BD7410EBDB5017DE38E8708008002FAAA4171D5",
INIT_2C => X"00000000000000000000082005F6ABFFEBA0870281C5F4716D5D7FEDB7D0955D",
INIT_2D => X"1401FFFFD5420BAA2AA821FF08043DE10002A964000000000000000000000000",
INIT_2E => X"FBD7410A2AE965555D556ABEF080028B55FFFFFDEBAFFD57FE00A280144BAAAD",
INIT_2F => X"2D16ABEF5500175EF552ABDE000855544AAAA82174105D0402000087FC00BAA2",
INIT_30 => X"AAD154400AAFBC015555554001008003FE00AAEA81154AAFFD65FF5D2EBDEAAA",
INIT_31 => X"FA2AA155550004021E5582A964BE557FEABEF00002BE10FFD540000FFD56ABF5",
INIT_32 => X"1000043DEAA085555400FFAAAAA10F7AC28BF558001454DF78017555F780175E",
INIT_33 => X"5EF5D7BFEEF35055487EFF7D1400105D517FF55087FD7410A2FBC01E7F2AE966",
INIT_34 => X"0000000000000000000000000000000000000010007FEABEFAA84174BA557FD5",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000040",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(4),        -- Port A data input
DOA(0)   => data_read_a_lo(4),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(4),        -- Port B data input
DOB(0)   => data_read_b_lo(4),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_5_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50DB4A0791B1B4B694369283C81F9996A091832102004AB37B20E07C0C1E006",
INIT_01 => X"285FBC448000804C446A00000034824841280A00084000C8C212892EE2953235",
INIT_02 => X"C809AD5CB118E640A4D118FC011FF0002080000082C8C66609DB7DDDCB1F2036",
INIT_03 => X"250907263A4C90D210A35C82484285720B20648A88800000B8E0F850A8C4500E",
INIT_04 => X"4005122126899100064D20001044429C78243A2C0436C887198AB916E0551A24",
INIT_05 => X"A370C14CA0E900004048002389CFE2F20F7D7A314CB5C20AE51437E044948912",
INIT_06 => X"90184D150505A1D84B7E2A285401412870B20A51842404C44437118630839B88",
INIT_07 => X"E640A94D1AB469D6300E2FFFAA7F8A4D23248130E259C903FBC403A9601A62E8",
INIT_08 => X"0A7E3016250D49CA3F83108186400000EBFD235488B9749BC1AAF325B35CB118",
INIT_09 => X"9B020B7E6AE46082032004904200C03DBC3BCA4860270BFA829968040B0800AC",
INIT_0A => X"22181A2B9203642840124098516CE0C3D825124111A79F802800F20DB4D6DA34",
INIT_0B => X"6824911331CA84D346A964F0125CD7AB1938A00AEFDD567DE480116848C9426A",
INIT_0C => X"01AD7016D701ED7012D701ED7016D701AAB8096B80F5A21828041846620F5AB8",
INIT_0D => X"847B053F48A8308A644A412BCA8470FF0209019081C706EABDAAC0DC0AF012D7",
INIT_0E => X"2194FFC044FF84B08FC862A2CD8F0A89014080A2425422151870500544991292",
INIT_0F => X"038ABBCBC7C7802F86FF87C002F87F002F86FF87C002F87F2000804821021004",
INIT_10 => X"0380230F2FFC002F94FF87C002F87F002F94FF87C002F87F2201BFFEBC2BA0C2",
INIT_11 => X"BFFE7C69E01804E1E7EABE3F000FF97D7C4BC0E008C7C3FE58FC029FEF5CD9A7",
INIT_12 => X"EC9C8120C4DFC802808B2EB22E777ADDE6F8A47CC0600C2683E0FFAAE3F1F001",
INIT_13 => X"FC14DFC5186104C6FE5037FFF00FC0000FC0FEE487A7066FA38C3082637F83BD",
INIT_14 => X"072FFF41C1C0C2038A7CED87A7D109FBBA5070380131CBFB2477BF919024189B",
INIT_15 => X"9F46DFBEB1B7F0380C4A80092E0FC1FDE607A7C077FFE828F0080AE1DFAA1E9F",
INIT_16 => X"5594254A10A03446128898494C09402081F83200A9442217159880640942320E",
INIT_17 => X"1940509465014251140519445094251142511445094451942511425014451940",
INIT_18 => X"9405094450944511425114650146501425194450944509405194250146501405",
INIT_19 => X"0A983124B2DA6924965B4D509445094051940501465014251142501465094451",
INIT_1A => X"BE5FDFF3F7F773CF3CF7D79FA8F5BB4E7F7B9DB7FF3A7E0FF4807F1B6DB7ED43",
INIT_1B => X"F77BBDDEEF77BBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEF",
INIT_1C => X"EF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEE",
INIT_1D => X"FFBFFE00000000000000000000000000000000000000000000001007FE1BFB5E",
INIT_1E => X"FFAE821FF552E820105500155555D2AA8A00AA843FFFFF78002155AAAE974AAF",
INIT_1F => X"0FFAE80000AAAE974BAFFAEAAB45AAAEBDEAAA2FFEAA00AAFFC21FFF7D542000",
INIT_20 => X"000055574BA557FFFF55087BEABFF552ABDF45A2D16AAAAF7D56AA00AA840000",
INIT_21 => X"0BA550015400087FD74BAFFD540000F780155555D7BE8B45085168BFFA2D17FE",
INIT_22 => X"AA10005140145FFFBC01EFAAFFD75FF002E97555A2AABDEAAAAAAAAA00AAAE82",
INIT_23 => X"174BA5D043FF45AAAA974AAF7AEBFF55082AAAA10F7FFEAB455500175FF5D2AA",
INIT_24 => X"000000A2FFC21555551554005D2EA8AAAF78015545FFD555410552EA8BEFAA84",
INIT_25 => X"8E0217DBEA4954AAE3FBFDE00000000000000000000000000000000000000000",
INIT_26 => X"2F1C01D7F7D142028EBAA801EF492087A10490A171455D2EADA28B6803FFFFFF",
INIT_27 => X"FFD56FA10AA8417428E3AE87010A2A4974AAE3AEAFB6DAAA4BDEAAA2F1EDA28A",
INIT_28 => X"D14516DBD7BEDB7DE381451554AA497FFFF451C75EABEF4124BAF55B6DF6FABA",
INIT_29 => X"AAAAA0AFA28A2A4850925D0010400087FD24AAE3DF47010E38E0516D5D7BE8B6",
INIT_2A => X"B7D5500155FF552AAFA10007155545F7F1C21D7AAF1D55FF082A9057DA2AABDE",
INIT_2B => X"70384124ADBFFBE84174AA55043FF6DBEAE950AAEB8ABDF7D1C2AAFA28EBF5E8",
INIT_2C => X"00000000000000000000010A2FBC01555D51524004920ADA82EB8A12410EBFB4",
INIT_2D => X"EBFEBAF7843DFEFF7AE801EFF780174AAAAFBFEE000000000000000000000000",
INIT_2E => X"803FEBAAAD17CEAAAAD140155FFD5420BAA2AA821FF080415410002A96555552",
INIT_2F => X"80028B55FFFFFDEBAFFD57FE00A280144AAA2AA97400A280174AAA2AEBDFEFA2",
INIT_30 => X"A2AE965FF557FE8BFF55557FF55FFFBFFEAA5D51554AA087BFEF555D556ABEF0",
INIT_31 => X"F0004821FFAAAEBDEAAAA843CEAAAA80174105D0402000087FC00BAA2FBD7410",
INIT_32 => X"FF5D2EBDEAAA2D16ABEF5500175EF552ABDE00005554545F7D140145A2D5555F",
INIT_33 => X"E00AAAA81114AAFFD64BA00043FFFFFF80174AA55043DFFFFFAE974BAA2AEBEF",
INIT_34 => X"0000000000000000000000000000000000000000AAFBC015555554001008003F",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000180",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(5),        -- Port A data input
DOA(0)   => data_read_a_lo(5),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(5),        -- Port B data input
DOB(0)   => data_read_b_lo(5),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_6_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10804B0061A010A2840012C030028180004003220200403302301C0381A0086",
INIT_01 => X"870041CA3839684D18A160000C52424841000000090800090210010008110204",
INIT_02 => X"080108200C1000004464480400C0080100000000010432400800800009882050",
INIT_03 => X"040001008C2340D0840208624210002182800584488000103080010E08C10000",
INIT_04 => X"00101611A029B08410044800000000040088102A440814040400900500001800",
INIT_05 => X"02800000400C820934E4A0002900404400820004000A00824004085011200A00",
INIT_06 => X"2210001A12100830434040870BFE004044420322C00812900308010000829400",
INIT_07 => X"00000860400108C22000A103090074120044800040001103005180911FE0C134",
INIT_08 => X"FD01C0120484C0580020C10000000000087C0800209100004228000110000C10",
INIT_09 => X"88FC08362240404100228080D200DFC1610200E40AA050000040D0C463008083",
INIT_0A => X"29561B22D77C720D2522400000400882091210008440005F8BF4C00002900004",
INIT_0B => X"7E25D11A200024541100342A5A2886285502A880C00107FD355E022005026BCA",
INIT_0C => X"D8282D8A82D8A82D8682D8682D8E82D8A016C1416C15A01D68209A127208A6B1",
INIT_0D => X"807888180A80910A1460150900013400410CB5C9D96236883460B60B602D8282",
INIT_0E => X"0062003C10002442006429124290034E85A742D1A368D0DA2004696884851806",
INIT_0F => X"000000157000604050000000028000D04050000000028000CE80004C00000000",
INIT_10 => X"000000000483D04042000000028000D04042000000028000C508000100000000",
INIT_11 => X"000100000000000000078000A40006000000000000000019A003080010200000",
INIT_12 => X"1001000000093490308001408000000200020000000000000000900518000508",
INIT_13 => X"23490002400000004993C000080000000000001FC000C8804020000000246800",
INIT_14 => X"C05000802000000000001740002256004100000000000000FD00000220000001",
INIT_15 => X"00A000404A000200020000000000002099C000330000040000000000001F0000",
INIT_16 => X"68DA308D09D0804880089A49461032040C07C1440C8190800020530865400540",
INIT_17 => X"9DA7695A1685A369DA7685A168DA369DA5685A168DA7695A5685A368DA7695A5",
INIT_18 => X"5A168DA7695A168DA1695A769DA1685A3695A569DA3685A169DA769DA1685A16",
INIT_19 => X"00046638C31C71C718638E68DA7695A568DA3685A769DA5685A368DA569DA368",
INIT_1A => X"8E76DDB3B7B377DF7DF7D7CEE7F78BCE7F8FF0F4FA957FC7F37F3F5F7CF7F108",
INIT_1B => X"7F3F9FCFE7F3F8E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E3",
INIT_1C => X"E7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE",
INIT_1D => X"AAABFE00000000000000000000000000000000000000000000181007FFDE534F",
INIT_1E => X"F78002155AAAE974AAFFFBFFE10F7FBE8BEF552E95555552EAABEF082E975EFA",
INIT_1F => X"0A2AAAAA10087FC01EF552EAAB45F7AE821550851555555D2AA8A00AA843FFFF",
INIT_20 => X"EFA2AEBDFFF552AAAA00AAFFC21FFF7D542000FFAE821FF552E8001055001541",
INIT_21 => X"000AAAE974BAFFAEAAB45AAAEBDEAAA2FFEAB45552E800AA555568A105D002AB",
INIT_22 => X"AA00AA8400000007BC21FFAA803FFEF5551420105D5568B45FF8400000FFAE80",
INIT_23 => X"C2155007FC20BAA2D5575FF087FFFF55087BEABFF552ABDF45A2D16AAAAF7D56",
INIT_24 => X"0001555D7BE8B45085168BFFA2D17FE000055574BA557FFFE10F7AAA8A00F7FB",
INIT_25 => X"24ADBD70820975FFA2A4BFE00000000000000000000000000000000000000000",
INIT_26 => X"D2EADA28B6803FFFFFF8E0217DBEA4954AAE3FBFDE38F7FFEABFF412A9056D49",
INIT_27 => X"492087010490A07038B6A0AFA38007BC51EF4920AFB55EBA4851450855555455",
INIT_28 => X"2555F68A3855002FBC7BEA4BFFFF492EADA28A2F1C01D7F7D142028EBAA801EF",
INIT_29 => X"45E38A07028E3AE87010A2A4974AAE3AEAFB6DAAA4BDEAAA2F1EDB55492A8508",
INIT_2A => X"F55B6DF6FABAFFD56FA10AA84174381C7FC01C7B68E3DFC75555400105D516DB",
INIT_2B => X"FE38F7A0AFA38E3FFC21450071C2092A2D5571FF0851FDF451C75EABEF4124BA",
INIT_2C => X"0000000000000000000016D5D7BE8B6D14516DBD7BEDB7DE381451554AA497FF",
INIT_2D => X"BEABEF002E801EF00003FF550800155FFA2803CE000000000000000000000000",
INIT_2E => X"8417555085154555552EBFEBAF7843DFEFF7AE801EFF780174AAAAFBFEEAAF7F",
INIT_2F => X"FD5420BAA2AA821FF080415410002A964AAFF803DEAA087FD55FF00043DF45A2",
INIT_30 => X"AAD17CF55002E95410557BEAABA55043DF55F7803FFEF002ABEEAAAAD140155F",
INIT_31 => X"55D51420105D517DF55AAAA964AAA2AA97400A280174AAA2AEBDFEFA2803FEBA",
INIT_32 => X"555D556ABEF080028B55FFFFFDEBAFFD57FE00A280144BA5D7FC2155FFAABDF4",
INIT_33 => X"EAA5D51554AA087BFEEAAF7803DEAAAAFBC0155085540000A2D5575FF08517CF",
INIT_34 => X"00000000000000000000000000000000000001FF557FE8BFF55557FF55FFFBFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000120",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(6),        -- Port A data input
DOA(0)   => data_read_a_lo(6),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(6),        -- Port B data input
DOB(0)   => data_read_b_lo(6),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_7_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10804B00482010A2842012C024500188000003000000003302300C018180002",
INIT_01 => X"0200084020084048040080000201024040000000080000080200010008110204",
INIT_02 => X"4801082248100000444008000080000041000000002222400800000009008010",
INIT_03 => X"0401008108A1444000020A400000002902006400088000003080040408C10000",
INIT_04 => X"0000100022418000000C80C00400000400201839040000050001140400201820",
INIT_05 => X"02000000400041092C80C0214144004400000000000800045004000020220800",
INIT_06 => X"0000300000000830435150020003004060000000080800801100000030829001",
INIT_07 => X"00000840000008C02000A503010002928040800062481919047140D40008C000",
INIT_08 => X"0A0002120484C0580850810000000000487C000000910000402A800110024810",
INIT_09 => X"8802083624504000022680A1DA20800164000400112284000004D404022A8800",
INIT_0A => X"30014050280040180020400011640CC72E029000084800503004C40100D21024",
INIT_0B => X"3801078228010454210028240082200081140800900220000000002011440009",
INIT_0C => X"40022400224002240822408224082240C1120211202008900800100242428280",
INIT_0D => X"807802988294900A00451109006230006E000800001280110050902901240022",
INIT_0E => X"0042C000C0002000000020020490000400020001020080401010813094801146",
INIT_0F => X"807144102420700052000003C00780B00052000003C007808450484C00000000",
INIT_10 => X"2C0E00E0D003300052000003C00780B00052000003C00780890800010000130C",
INIT_11 => X"000100000661801E18042100E000060100000B03803838012403800010240000",
INIT_12 => X"10111848322020512000414400000002000A1001058300C0741C005412080908",
INIT_13 => X"029F008240864231013BF00008000C3C003F00184040EF8041204321188053E0",
INIT_14 => X"F770008060130C8071821040403F5600411004C2600E3400C27C020223090644",
INIT_15 => X"00B8CA406A0002C812240B0201F038021140403F740004010472041E20110100",
INIT_16 => X"0080228011010042802890484040000008004945000100008844430060198941",
INIT_17 => X"0000000000000600802008020000400000000000080200802008000000000000",
INIT_18 => X"8020100000000008020080000000000020080200000000040080200802008060",
INIT_19 => X"0A14584104000208208000018020080200000010020080200800010000080200",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000442",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"82AAAA00000000000000000000000000000000000000000000001007FEBC3240",
INIT_1E => X"552EAABEF082E975EFAAAABFFEF002ABDF555D5157555F7FBC00AAAAD5400BA0",
INIT_1F => X"AAAAABDF55FFFBFDF55555568ABAAAD5401FF5D2AAAA10F7FBE8BEF552E95555",
INIT_20 => X"005D55554105D51401555D2AA8A00AA843FFFFF78002155AAAE974AAFFFBFFEA",
INIT_21 => X"A10087FC01EF552EAAB45F7AE821550851554AAF7FBFFEAA007BFFFEFF7D5400",
INIT_22 => X"00105500155EF5D2EBFF450000020AA5D7BC0000F7D555545A28000010A2AAAA",
INIT_23 => X"A8A10FFD568ABAA2D56AAAAF7AABFE00AAFFC21FFF7D542000FFAE821FF552E8",
INIT_24 => X"000145552E800AA555568A105D002ABEFA2AEBDFFF552AAAABAA2AE95555FFAA",
INIT_25 => X"F5C20BAAAD5420821C2EAAA00000000000000000000000000000000000000000",
INIT_26 => X"7FFEABFF412A9056D4924ADBD70820975FFA2A4BFFFF1C2EB8F45555550545E3",
INIT_27 => X"BEA4954AAE3FBFDE82B6AEBAF55E3FFFAF55555F6FA92BED5421C75D20AAA38F",
INIT_28 => X"20075FDFD7F7D5400385D51504385D55401455D2EADA28B6803FFFFFF8E0217D",
INIT_29 => X"7DB68E02038B6A0AFA38007BC51EF4920AFB55EBA485145085555492F7F5FFE9",
INIT_2A => X"028EBAA801EF492087010490A071EF4920B8F45140E07082417BC2000EBD5505",
INIT_2B => X"DA92A2A09257DE3A4AAA10F7D16FAAABED56AE82F780BAE28A2F1C01D7F7D142",
INIT_2C => X"00000000000000000000155492A85082555F68A3855002FBC7BEA4BFFFF492EA",
INIT_2D => X"EAAB455D5142155AAD1400AAA2D1420005D2EA9A000000000000000000000000",
INIT_2E => X"D1421555D042BAAAF7FBEABEF002E801EF00003FF550800155FFA2803CFFF552",
INIT_2F => X"7843DFEFF7AE801EFF780174AAAAFBFEE00F7AAAAB55AAFBEAB555D7BFDE00F7",
INIT_30 => X"085154400FFD17FE1000517FF55FFD5420BA5D55400BA555543155552EBFEBAF",
INIT_31 => X"0087BC0000A2D5421EFF7AE810AAFF803DEAA087FD55FF00043DF45A28417555",
INIT_32 => X"AAAAD140155FFD5420BAA2AA821FF080415410002A965FF080428B45552A9540",
INIT_33 => X"F55F7803FFEF002ABEE00A280001FFA28028A00FFD17DEAAF7D56AA10FF842BA",
INIT_34 => X"0000000000000000000000000000000000000155002E95410557BEAABA55043D",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"FFFFFFFE00000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000000000000000000001F",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(7),        -- Port A data input
DOA(0)   => data_read_a_lo(7),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(7),        -- Port B data input
DOB(0)   => data_read_b_lo(7),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_8_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10004B00000400E2840012C0000001800000070000000033022000000000082",
INIT_01 => X"000009C0183808481C0160000E02424040000000180800080200010048110204",
INIT_02 => X"080108000090000004400C000080000051000000000002400800000009000010",
INIT_03 => X"0000000004300840000200000000000002800504488000103080880008800000",
INIT_04 => X"00009410A028A084000440C00400000400001032040800150400008500221800",
INIT_05 => X"4280008040048A09302420202804400400800010200A00000204080011014A00",
INIT_06 => X"2B02000A32114192434010001FFC004240428122000800000008012000821400",
INIT_07 => X"00000840000008402001A50200000630404080006248381B000080837FF88114",
INIT_08 => X"0A000210040440480000090000000000087C0000009100000002000110000090",
INIT_09 => X"08020A322000400102260021DA2080114502002409A04400004282C4E1228800",
INIT_0A => X"904A4522920052012120400011641C4601005000041100002004800100C21024",
INIT_0B => X"78051792A8000454104020001280008845022000900000010444000000020009",
INIT_0C => X"000000000000000000000000000000000800040000452A9008001002424A8002",
INIT_0D => X"807880508202100A1000810B2020340041248548490004800400000008000800",
INIT_0E => X"20020000C000044214240932000001428CA14650A128508A2004284024840022",
INIT_0F => X"80000000001020404000783FC0000010404000783FC000000880084C01041008",
INIT_10 => X"FC7E0000000010404000783FC0000010404000783FC000000500000103D45F3D",
INIT_11 => X"000103961FE78000000000402400020003B43F1F800000002201080000202658",
INIT_12 => X"01617CD8000000803000804080000020090659833F9F03C00000000000040500",
INIT_13 => X"00400018639EC000000000000FE03FFC00000000400840000C31CF6000000800",
INIT_14 => X"4000001E2A3F3D80000000400802000401AA8FC7E00000000100002C2F5B0000",
INIT_15 => X"4020000104480DC372B47F060000000000400802000017570FF6000000010020",
INIT_16 => X"28CA30051851A0C0002890484600320408004444048090800022130864000540",
INIT_17 => X"84A1284A1284A328CA328CA328CA328CA328CA3284A1284A1284A1284A1284A1",
INIT_18 => X"CA328CA328CA3284A1284A1284A1284A328CA328CA328CA3284A1284A1284A12",
INIT_19 => X"080440000000000000000028CA328CA328CA328CA1284A1284A1284A128CA328",
INIT_1A => X"9EDFC8F33637D6CB6CB2900DA6128A0A543EBC57A10A244257C5051E75D64108",
INIT_1B => X"1F0F87C3E1F0F9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7",
INIT_1C => X"E1F4F87D3E1F4F87D3E1F4F87D3E1F4F87D3E1F4F87D3E1F4F87D3E1F0F87C3E",
INIT_1D => X"02ABFE00000000000000000000000000000000000000000000001007FE8A8913",
INIT_1E => X"F7FBC00AAAAD5400BA082AAAA10000000010F7D5421EF007BC01FF5D7FFFE100",
INIT_1F => X"A5551554AAFF80021EF002A820BAFF8428A00A2AAAABEF002ABDF555D5157555",
INIT_20 => X"EFFFFFEAB55002ABFE10F7FBE8BEF552E95555552EAABEF082E975EFAAAABFEA",
INIT_21 => X"F55FFFBFDF55555568ABAAAD5401FF5D2AAAB55FFD1400AA5D7FC01EFA2FFE8B",
INIT_22 => X"74AAFFFBFFEAA08001555555516ABEFA280020AA5D043DF55557BEAAAAAAAABD",
INIT_23 => X"2AB55005140145AAFFE8AAAF7D1401555D2AA8A00AA843FFFFF78002155AAAE9",
INIT_24 => X"0000AAF7FBFFEAA007BFFFEFF7D5400005D55554105D51400005551421EF0804",
INIT_25 => X"7FC21EF5D75FFE10142EBAE00000000000000000000000000000000000000000",
INIT_26 => X"C2EB8F45555550545E3F5C20BAAAD5420821C2EAAA101C0005000E3D1401D71C",
INIT_27 => X"0820975FFA2A4BFE925D51554AAE384001FF142E800AAFF802AA28AAAEAFBFF1",
INIT_28 => X"2557BC21D7BEF5EDBC7FFF1EFB6D1420BAE38F7FFEABFF412A9056D4924ADBD7",
INIT_29 => X"55417BEDA82B6AEBAF55E3FFFAF55555F6FA92BED5421C75D20AAB45F7D14709",
INIT_2A => X"FFFFF8E0217DBEA4954AAE3FBFDEAA1C001056D415F6ABEFA2840208249043AF",
INIT_2B => X"00385D51401EF00002FB45085F4016DAAF1EDAAAFFFB401455D2EADA28B6803F",
INIT_2C => X"00000000000000000000092F7F5FFE920075FDFD7F7D5400385D51504385D554",
INIT_2D => X"417410AAD540155557FC01EF5D557DE105D2AA8A000000000000000000000000",
INIT_2E => X"842AABAA2AEBDFFF552EAAB455D5142155AAD1400AAA2D1420005D2EA9A105D0",
INIT_2F => X"02E801EF00003FF550800155FFA2803CE105D55574BAA280021EF5D2E820BAF7",
INIT_30 => X"5D042BB45FFD157410557FC0155F7D57FF55F7D57FFEF550028AAAF7FBEABEF0",
INIT_31 => X"FAA8000000080428B55087FFFE00F7AAAAB55AAFBEAB555D7BFDE00F7D142155",
INIT_32 => X"55552EBFEBAF7843DFEFF7AE801EFF780174AAAAFBFEEBA5D04021EF087BE8BF",
INIT_33 => X"0BA5D55400BA5555430BA5555421EF00043FF45007BC21FFA2D57FEBAF7FBC21",
INIT_34 => X"0000000000000000000000000000000000000000FFD17FE1000517FF55FFD542",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000080",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(8),        -- Port A data input
DOA(0)   => data_read_a_lo(8),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(8),        -- Port B data input
DOB(0)   => data_read_b_lo(8),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_9_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10004B00018000A2840012C0000281800000030000000033022000000000006",
INIT_01 => X"000008000000004C0020000000100268413C0A61590001D90213C10008110204",
INIT_02 => X"680108200010000054400C000080000041000000010002400800800009082011",
INIT_03 => X"0004000000002040000200100000000042800584488000103081880008800000",
INIT_04 => X"00001610A00AB084000400C00600000400001030040010050020020400001880",
INIT_05 => X"02000200400C8A09206420000C00410400000000000800000804000000000800",
INIT_06 => X"2A10201A12104010435051000801004040000322980800000080000100821000",
INIT_07 => X"000018400000086020002502000002000040800062C8081B0000008000088034",
INIT_08 => X"0A000610040440480000010000000000187C0000009100002046000110000010",
INIT_09 => X"4802082220084001002400214A2080014400006400A000000000015421800800",
INIT_0A => X"4B505008020032032320400011640447000010040000000020048409004A9020",
INIT_0B => X"280005922000045400002001100000000D0000008000000041C48000002003EA",
INIT_0C => X"2080020000208002000020800200002080010000104100800000100202420142",
INIT_0D => X"C06800100240180A0010010921003400432C8CC8D80044000000080080020800",
INIT_0E => X"2002C000C000240004641932041403428DA146D0A36850DA3200684004800403",
INIT_0F => X"0000000144002000420000000280001000420000000280000000084C01041008",
INIT_10 => X"0000000004801000500000000280001000500000000280001100000100000000",
INIT_11 => X"00010000000000000002A0002000020100000000000000182001000000240000",
INIT_12 => X"00110000000900003000004000000000000A0000000000000000900002000100",
INIT_13 => X"205D0080400000004803F0000800000000000004E0004E800120000000240BA0",
INIT_14 => X"4770000060000000000005600013560001100000000000002574020020000001",
INIT_15 => X"0020CA406A0000080200000000000020806000137400040000000000000B8000",
INIT_16 => X"68DA320D19D1A0CA8028984D46543600080040440C8090800000130061400140",
INIT_17 => X"8DA368DA368DA1685A1685A1685A1685A1685A1685A1685A1685A1685A1685A1",
INIT_18 => X"5A1685A1685A1685A1685A1685A1685A368DA368DA368DA368DA368DA368DA36",
INIT_19 => X"801010000000000000000068DA368DA368DA368DA368DA368DA368DA3685A168",
INIT_1A => X"344A2D840100E492082405548817344CCCF48DE68A89004F98614C5C38E2540A",
INIT_1B => X"1A0D068341A0D14514514514514514514514514514514514514534D34D34D34D",
INIT_1C => X"41A4D268341A0D069349A0D069349A0D068341A4D268341A4D268341A0D06834",
INIT_1D => X"FD557400000000000000000000000000000000000000000000001FFFFE2CAD83",
INIT_1E => X"007BC01FF5D7FFFE10002ABFF55F7D168A00552E95555007BFFF55087BE8BFFF",
INIT_1F => X"0F7FBC0145F7AE801EFF7FBFFF455D7BC0155F7D557410000000010F7D5421EF",
INIT_20 => X"00AA803FFEF5D55421EF002ABDF555D5157555F7FBC00AAAAD5400BA082AAAA1",
INIT_21 => X"4AAFF80021EF002A820BAFF8428A00A2AAAAAAAF7D17DE00FFFBD5555A2AABDE",
INIT_22 => X"75EFAAAABFFEF002A954BA5551421EF552E954105D00021455555420AA555155",
INIT_23 => X"575EFA2FFD75455D7BE8A005D5557410F7FBE8BEF552E95555552EAABEF082E9",
INIT_24 => X"000155FFD1400AA5D7FC01EFA2FFE8BEFFFFFEAB55002ABFE10080028BFFF7D5",
INIT_25 => X"71F8F7D147BEFBEFEBD152400000000000000000000000000000000000000000",
INIT_26 => X"C0005000E3D1401D71C7FC21EF5D75FFE10142EBAF7DE3D16DA0041209056D1C",
INIT_27 => X"AAD5420821C2EAAA10E3FFC0145F7A0801FFEBFBF8F6D417BC716DEBD1524101",
INIT_28 => X"8F7F5D0545B6AAB8E38B68A3AFFF5551471FF1C2EB8F45555550545E3F5C20BA",
INIT_29 => X"455D5B470925D51554AAE384001FF142E800AAFF802AA28AAAEAFABAE3D17DE2",
INIT_2A => X"56D4924ADBD70820975FFA2A4BFFFF082E974BA4155401C7552097428550E021",
INIT_2B => X"AE0008002ABFFF7DB505FFAAFBD7555417FEFA00495B52438F7FFEABFF412A90",
INIT_2C => X"00000000000000000000145F7D147092557BC21D7BEF5EDBC7FFF1EFB6D1420B",
INIT_2D => X"17DE100804001EF55516ABFF557BFDFEFA2D5400000000000000000000000000",
INIT_2E => X"7FD55FFA2D5400105D0417410AAD540155557FC01EF5D557DE105D2AA8BEFAAD",
INIT_2F => X"D5142155AAD1400AAA2D1420005D2EA9A00A2FBC0145FF84001EFA2FFEABFF00",
INIT_30 => X"A2AEBDEAAAAD17DEBAFFD142155FFAAAAABAFFAAAABFF5551555FF552EAAB455",
INIT_31 => X"55D00154AA552E801455D7BD54105D55574BAA280021EF5D2E820BAF7842AABA",
INIT_32 => X"AAF7FBEABEF002E801EF00003FF550800155FFA2803CFFF002E954BA00514015",
INIT_33 => X"F55F7D57FFEF550028A10000428BEFF7FFC01FFA2FFD5545007BFDE10087FC00",
INIT_34 => X"0000000000000000000000000000000000000145FFD157410557FC0155F7D57F",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000100",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(9),        -- Port A data input
DOA(0)   => data_read_a_lo(9),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(9),        -- Port B data input
DOB(0)   => data_read_b_lo(9),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_10_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10040B0001824802840102C00002C18000202300500030B3132000400992006",
INIT_01 => X"A140098018300848180060000C00424040000000080000080200010008110200",
INIT_02 => X"0801080200100000046558040080000041000000002402400800000009008010",
INIT_03 => X"00010100840000D0842242024210810802006400088000003080054288C10000",
INIT_04 => X"0000100022008000000C08C00C00000400A83A3044200C840000800400101820",
INIT_05 => X"0200000040000000248080210044000402000025000800020004207010100800",
INIT_06 => X"0800200000004010435040A14001004844000800CC0812541020008230829000",
INIT_07 => X"00000860408108502000250208000600004080006248081B0040808000088000",
INIT_08 => X"0A000210040440480060010000000000087C0810209900000002000110020010",
INIT_09 => X"08020A2222004040000484214A2080110108C280022210020240000401080880",
INIT_0A => X"000000000200000C042040001164044609101000840000802004800100421020",
INIT_0B => X"782415809888A45010082408028010080110280800001001051A124810410800",
INIT_0C => X"0089000890000900009000890008900008800048004420910800120242488000",
INIT_0D => X"4110000006008820020010010001300040000100014000808C48004008800090",
INIT_0E => X"2002000040002000040020020490080400020001000482000010012080008005",
INIT_0F => X"0000010140002040100000000280401040100000000280400000204801041008",
INIT_10 => X"0000000006801040020000000280401040020000000280400500000000000000",
INIT_11 => X"0000000000000000010280002400040000000000000001182001080010000000",
INIT_12 => X"10000000000D0000808000408000000200000000000000000000902000000500",
INIT_13 => X"A000000200000000681000000000000000008004A00040004000000000340000",
INIT_14 => X"4000008000000000000085200002000040000000000001002400000200000001",
INIT_15 => X"00200000000002000000000000000021802000020000000000000000020A8000",
INIT_16 => X"040006E00100044200289048085D402008000040000100000000020065400000",
INIT_17 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_18 => X"0000000000000000000000000000000020080200802008020080200802008020",
INIT_19 => X"8290100000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"8A355950666151451453D5006F86890A940FE0D39712614261D20E4355520542",
INIT_1B => X"6532994CA65328A28A28A28A28A28A28A28A28A28A28A28A28A28A28A28A28A2",
INIT_1C => X"AE532994CA6532995CAE572B94CA6532994CA6572B95CAE532994CA6532994CA",
INIT_1D => X"FFBC2000000000000000000000000000000000000000000000001007FECF31DC",
INIT_1E => X"007BFFF55087BE8BFFFFD557400FF842ABEFA2AAA8B5500003DF55F7D568AAAF",
INIT_1F => X"008556ABFFA2D16AB550000021FFF7D17FFEF08042AB55F7D168A00552E95555",
INIT_20 => X"55A2D557400557BC2010000000010F7D5421EF007BC01FF5D7FFFE10002ABFE0",
INIT_21 => X"145F7AE801EFF7FBFFF455D7BC0155F7D557545FFAE820AA007BFDFEF55003FF",
INIT_22 => X"00BA082AAAA00FFAE820AAAAAABDFEFF78028BEF005140145A2842AA10F7FBC0",
INIT_23 => X"6AB55A2D157400552EBFFEF5D7BD75EF002ABDF555D5157555F7FBC00AAAAD54",
INIT_24 => X"0000AAF7D17DE00FFFBD5555A2AABDE00AA803FFEF5D55420BA08557FEBAAAD5",
INIT_25 => X"0E3AF55F7DF68ABAE3F1C0000000000000000000000000000000000000000000",
INIT_26 => X"3D16DA0041209056D1C71F8F7D147BEFBEFEBD152400F7842FBD7B6AAAAB551C",
INIT_27 => X"5D75FFE10142EBAE0008556FBD7B6DB6AB7D1C0A001D7FFD178FC71C0E28B7DE",
INIT_28 => X"2147BFAFEF49043AF45A2DF504285D71C00101C0005000E3D1401D71C7FC21EF",
INIT_29 => X"7DA28428A10E3FFC0145F7A0801FFEBFBF8F6D417BC716DEBD15256DF7AA8209",
INIT_2A => X"545E3F5C20BAAAD5420821C2EAAA00E3AA82092A2AABAFD7EB8A2ABC70855401",
INIT_2B => X"70821C557AE92A2DF6AB7DA2DF50410412ABDFC75D7BD55FF1C2EB8F45555550",
INIT_2C => X"000000000000000000000BAE3D17DE28F7F5D0545B6AAB8E38B68A3AFFF55514",
INIT_2D => X"03DF45FFAEA8B555D2EAAB45F7FBE8ABAAAD5400000000000000000000000000",
INIT_2E => X"D168B55552AA8BEFAAD17DE100804001EF55516ABFF557BFDFEFA2D540010FF8",
INIT_2F => X"AD540155557FC01EF5D557DE105D2AA8A0008557FF45FFFFE8BEF5D2E80155FF",
INIT_30 => X"A2D5401FFF7AA800105D7FE8BEF08002AB45AAFFC00AA5D51400105D0417410A",
INIT_31 => X"5AAAEAAB450055421FFAA8428A00A2FBC0145FF84001EFA2FFEABFF007FD55FF",
INIT_32 => X"FF552EAAB455D5142155AAD1400AAA2D1420005D2EA9A10A2AA82010AAAEAAB5",
INIT_33 => X"ABAFFAAAABFF555155400555568A10AAFBEABEFA2FFC0010082ABFF55557BD55",
INIT_34 => X"00000000000000000000000000000000000000AAAAD17DEBAFFD142155FFAAAA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"FFFFFFFE00000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000000000000000000011F",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(10),        -- Port A data input
DOA(0)   => data_read_a_lo(10),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(10),        -- Port B data input
DOB(0)   => data_read_b_lo(10),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_11_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10180B05A0010402840602C2D001019000000300000000330A20080EC180002",
INIT_01 => X"AB400986B830284D1820E0000C36424840000000080000088200080802512220",
INIT_02 => X"8801081438106400A4F55800008000004100000040CCE24208005000C9060032",
INIT_03 => X"000406A492E6E440842254D002108153432004800880000030C0315688C00006",
INIT_04 => X"00001201200090001205400000000094108C322644240C840008030440111800",
INIT_05 => X"222000444008010028404002A002009402400025080880000C04223000170900",
INIT_06 => X"01080C1020002810436532AB4003004864200A00540816544522008200821100",
INIT_07 => X"6400E96C488108502001295BA100022E4340800062D82819435143F20008C0A0",
INIT_08 => X"0A0012160585C1D809A3810000000000C8FD0B1420992419034A0221116C3810",
INIT_09 => X"4902083E2CB0400002020480C2008009000ACEC06B25500202988C84C0220028",
INIT_0A => X"004040000203600E06204000116C14474A36500499C49C802004C00800088000",
INIT_0B => X"6804110230CBA4576708201C0212100B492A2008000A1001C49A9348498B0808",
INIT_0C => X"410E5418E5410E5418E5418E5410E5418B2A0872A08428010000120202085000",
INIT_0D => X"41110244066C0820221480010AA7300042080980919580808C9A5002880A18E5",
INIT_0E => X"2022C000C0002020094030220C960A0409020481024482501A00401410088521",
INIT_0F => X"836090540355D86C046619A54052A5B86A046619694063168280004801041008",
INIT_10 => X"A2C60289802AB86A046619A54052A5B86C04661969406316AC018B0E2936DA02",
INIT_11 => X"CB0E1076D4A200B2AC611A3D0405886C6EB211550815A8A2686EC81E2A48B68A",
INIT_12 => X"8CE0C5E8F650E48000892B37885620C1E1A06D7016A90A4626D82B10F1B1FC09",
INIT_13 => X"4E02144D335546F28724001B030A56140A184483000C410A2699A2E32AC9C041",
INIT_14 => X"E8018A0A01B2990242E278056AAA203920E0BAE2012C08281808319C186F1E16",
INIT_15 => X"44F9051C049B18A12CB481042AD140C227002A0A02066954E7540CCDB58415AA",
INIT_16 => X"409024681181044080809A490C0964200800200108010003A02272400C19B80D",
INIT_17 => X"0902409024090240902409024090240902409024090240902409024090240902",
INIT_18 => X"1004010040100401004010040100401024090240902409024090240902409024",
INIT_19 => X"0284000000000000000000401004010040100401004010040100401004010040",
INIT_1A => X"20A069105251C0000001541148062608804180C0B10A04CA0900474210420140",
INIT_1B => X"0000000000000000000000000000000000000000000000000000208208208208",
INIT_1C => X"0000000000004020000000000000000000100800000000000000000000000000",
INIT_1D => X"00015400000000000000000000000000000000000000000000001007FE0FC1C0",
INIT_1E => X"00003DF55F7D568AAAFFFBC2010557BEAA10AAFBE8A00557BFFFEF007BC21550",
INIT_1F => X"55D7FE8BFF5D7FD540055003FFEFFFD142145000000000FF842ABEFA2AAA8B55",
INIT_20 => X"45557FC2010557FFDF55F7D168A00552E95555007BFFF55087BE8BFFFFD55754",
INIT_21 => X"BFFA2D16AB550000021FFF7D17FFEF08042AB55A2AAAAB4508517FE00557BC01",
INIT_22 => X"FE10002ABFE00AAFFE8AAAFF8402000550002145085555400F7FFE8A0008556A",
INIT_23 => X"3FEBA002A975EFF7D17DFFFAA8000010000000010F7D5421EF007BC01FF5D7FF",
INIT_24 => X"000145FFAE820AA007BFDFEF55003FF55A2D557400557BC2145A2D1421450804",
INIT_25 => X"7BF8FEF1C7FC516D080E15400000000000000000000000000000000000000000",
INIT_26 => X"7842FBD7B6AAAAB551C0E3AF55F7DF68ABAE3F1C00005D7BEDA00B6F1EFA2855",
INIT_27 => X"147BEFBEFEBD15257D5D7FEFBD7417BD5438550038FC7FFDF4216D080E07000F",
INIT_28 => X"514517FE105575C216D5571C50104171FDF7DE3D16DA0041209056D1C71F8F7D",
INIT_29 => X"00FFF1EFA0008556FBD7B6DB6AB7D1C0A001D7FFD178FC71C0E28B6DA2AEADB4",
INIT_2A => X"1D71C7FC21EF5D75FFE10142EBAE10A2FBEFA92F78A05028550E001451455524",
INIT_2B => X"016DB6D54514500003FEBA1420905FFFFDF78FC7BE84050101C0005000E3D140",
INIT_2C => X"0000000000000000000016DF7AA82092147BFAFEF49043AF45A2DF504285D71C",
INIT_2D => X"FFDE00F7D17FEBA557BEABEF557BD55EF082A974000000000000000000000000",
INIT_2E => X"FBC01FF082A97410FF803DF45FFAEA8B555D2EAAB45F7FBE8ABAAAD5400105D7",
INIT_2F => X"804001EF55516ABFF557BFDFEFA2D5401FF5D7FFDF55007BD74BA5D042AB45F7",
INIT_30 => X"552AA8BEFAAAABFF5555517FE005555401FF55515541000517FFEFAAD17DE100",
INIT_31 => X"A5D2A801455D5140000FFD57FE0008557FF45FFFFE8BEF5D2E80155FFD168B55",
INIT_32 => X"105D0417410AAD540155557FC01EF5D557DE105D2AA8A10AAFBFFE00F7AA974B",
INIT_33 => X"B45AAFFC00AA5D51401FFFFD15555500003FEBA5D04001EFFFFFE8B55FF84174",
INIT_34 => X"00000000000000000000000000000000000001FFF7AA800105D7FE8BEF08002A",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000100",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(11),        -- Port A data input
DOA(0)   => data_read_a_lo(11),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(11),        -- Port B data input
DOB(0)   => data_read_b_lo(11),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_12_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50080B01BC002006940202C0DE041196A83183000000023322287E0FC000006",
INIT_01 => X"0E000C048000C048400380000007026040000000080000088200002802153231",
INIT_02 => X"2809AD0E7D180040945008040090000061800000C0E2F66009DA3D11CB148015",
INIT_03 => X"210D050012F6F8D2108216E24842005B8A20640008800000B8E0141C28851006",
INIT_04 => X"0080100022408000060DE0000066630C70241827041000040800820480001AA4",
INIT_05 => X"0240000C400000003C808003E0C8001401000000040900020904004000070800",
INIT_06 => X"00006C00000008784B4D210E0001006050800000100804005784000130821200",
INIT_07 => X"A64019490A044860300FA3968B20028FC06080106249F819A19143FE00088200",
INIT_08 => X"0A002610240D494A0753D1810240000038FC234480B1709A81C67325B31EFD18",
INIT_09 => X"090209222EB84000010000104200802180210C007827C000009DBE040800008C",
INIT_0A => X"0000000002000030003040081164FC469227D20019F413503004900020000200",
INIT_0B => X"28200100004304D267C06CC500566003C13E0000000460000000000010CE0000",
INIT_0C => X"E1865E1065E1065E1865E1065E1065E1832F0C32F08000000004100202015940",
INIT_0D => X"0403CFE7E03E8080382FD0018FE670004000000000D5C023009278B7835E1065",
INIT_0E => X"01EA0000440000800A0040028108000000000000000000000A74812DF00E0BF4",
INIT_0F => X"8362F658A7E5F82CD23B6B0E403DBBE82C563B6A4E403DBB88C0E04820020004",
INIT_10 => X"BE5403AB992F282C563B6B0E403DBBE82CD23B6A4E403DBBB1084E4B25AC48DF",
INIT_11 => X"0E4B1D32BAB504BB74AD3F3FE04A8E0D0C319A7988B6F0C75CFD801A962454CF",
INIT_12 => X"18D994B866E2E8C3808B6B63040328E7A33AF99B0AC20DE634D06C437BF85100",
INIT_13 => X"5F6214CA5991C6A7177402C49CA354D808D358A927EAD10A652CC8E3538BEC41",
INIT_14 => X"E80083C3EAEB2003695430A7CDAA289553922990C11A4E494988231B32570CDC",
INIT_15 => X"D5B304AD05A946D81616970A225658940BA7CDAA0A312666BD600E5550B49F36",
INIT_16 => X"00000100000010420000904C0040000008003B81000000021CFEE02E2803BC0F",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"8020080200802008020080200802008000000000000000000000000000000000",
INIT_19 => X"0210100000000000000000008020080200802008020080200802008020080200",
INIT_1A => X"24481C040000B5145144015085C1B946088881360A95118D90215C090CB05442",
INIT_1B => X"32190C8643219041041041041041041041041041041041041041249249249249",
INIT_1C => X"4B2592C964B2592C964B2592C964B2592C964B2592C964B2592C964B2190C864",
INIT_1D => X"AFBC2000000000000000000000000000000000000000000000001007FEF001D6",
INIT_1E => X"557BFFFEF007BC2155000015555087FC0010AAFBFFE100004020BAAAFFD5400A",
INIT_1F => X"5AA8400000A2AABFF45550400000AAFBFFFEF550000010557BEAA10AAFBE8A00",
INIT_20 => X"10555155555FF8017400FF842ABEFA2AAA8B5500003DF55F7D568AAAFFFBC215",
INIT_21 => X"BFF5D7FD540055003FFEFFFD142145000000145A2AA821EFFFFFD7410007FC00",
INIT_22 => X"8BFFFFD5574000051420BA557FC2145557FC20AAA2D57DEBAA2FBD55455D7FE8",
INIT_23 => X"AAA00550415410AAFBFFFEF55042AB55F7D168A00552E95555007BFFF55087BE",
INIT_24 => X"000155A2AAAAB4508517FE00557BC0145557FC2010557FFDE10AA8400000082E",
INIT_25 => X"0A02092B6F5D2438A2FBC2000000000000000000000000000000000000000000",
INIT_26 => X"D7BEDA00B6F1EFA28557BF8FEF1C7FC516D080E1557D0075C7028B6F1FAE0000",
INIT_27 => X"F7DF68ABAE3F1C017DAA8E07028B6A0BFF6D490E00000BEF5FAFEF4904070005",
INIT_28 => X"FE3FBD0438007FC00385D555556DEB8410400F7842FBD7B6AAAAB551C0E3AF55",
INIT_29 => X"BAA2FBD557D5D7FEFBD7417BD5438550038FC7FFDF4216D080E0716DAAA0851F",
INIT_2A => X"56D1C71F8F7D147BEFBEFEBD152400005F450BA417BC51454971C20AAB6D17DE",
INIT_2B => X"DE10BE8E070280020AAA28410410400BEFBFAFEF49042AB7DE3D16DA00412090",
INIT_2C => X"0000000000000000000016DA2AEADB4514517FE105575C216D5571C50104171F",
INIT_2D => X"5574BAFFD568A10002A82000FFD5400AAA2FBC00000000000000000000000000",
INIT_2E => X"D568BEF0004174105D7FFDE00F7D17FEBA557BEABEF557BD55EF082A975EF005",
INIT_2F => X"FAEA8B555D2EAAB45F7FBE8ABAAAD5401EFA2AA974BAF7803FFFF002A82000FF",
INIT_30 => X"082A975EFA280175FFAAFFC00BA087FC20AA5D55555FFA28000010FF803DF45F",
INIT_31 => X"50851420BAFFD57DEAAAAFBD75FF5D7FFDF55007BD74BA5D042AB45F7FBC01FF",
INIT_32 => X"EFAAD17DE100804001EF55516ABFF557BFDFEFA2D540010007FD74AA007BD754",
INIT_33 => X"1FF55515541000517FE10F7AA954AA080428AAA000002010FFFFE8BEF080428B",
INIT_34 => X"00000000000000000000000000000000000001EFAAAABFF5555517FE00555540",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"FFFFFFFE00000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000000000000000000001F",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(12),        -- Port A data input
DOA(0)   => data_read_a_lo(12),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(12),        -- Port B data input
DOB(0)   => data_read_b_lo(12),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_13_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10110A0441812402840402822007818000E00700000000330A3000000008042",
INIT_01 => X"A1400984B830C848180260000C0042404001000008220008A200100802110200",
INIT_02 => X"88010C02801040002475580400800000410000000064024608134C0CC9018034",
INIT_03 => X"00010100926220D084234212421085084300648A0880000630C0654288C10000",
INIT_04 => X"0004122122029100100C00001200009C40A83A2044360C84190BAC04E0101820",
INIT_05 => X"027000004009050064C8C00104C10184034010250089C00EB004327064B60900",
INIT_06 => X"910000152500A050436A10A14003004864B00A50440812541027008230821380",
INIT_07 => X"640029605091495020002B8AAA000AF003408000E258081963F100C00008C2E8",
INIT_08 => X"0A001210040441C802E0010084000000AAFC09142899000B20020001105A0010",
INIT_09 => X"4A02096A62004000020004104200802D9838C2C80322100202020194408000A0",
INIT_0A => X"000000000203240E46204000516C04468C101005800E95802004B20020080200",
INIT_0B => X"28200101118BA4510008241D005211000910000A000A1000809A93485D610000",
INIT_0C => X"0000000800000000000000800000000000000400000000000000100202055040",
INIT_0D => X"0100000006C0802042501001C8017000C2190890904000508908000000000800",
INIT_0E => X"0010C000C00081A08BC832A209AB0A85094284A14254A2551010513080109404",
INIT_0F => X"01293C0F5012906A96DCD13042CE0C206E92DCD07042CE0C40D0204800000000",
INIT_10 => X"71CA2168ACB0E06E92DCD13042CE0C206A96DCD07042CE0C4408632C39530BA9",
INIT_11 => X"632C30D522CE80239CC2806AC44E954939AB299E000738F88296CA13B444CA42",
INIT_12 => X"D5306028F01990C080808494A64708B265CC4052B0F30302E060965EA0058408",
INIT_13 => X"28A2CA9722094650CCAC0629112BA89C04A228568547B1654B9104A32865145C",
INIT_14 => X"B80D4D8D48CB54012290470562EC29E44050B1DC60132282B68B9AA60C051E03",
INIT_15 => X"0A5C11B9008FE2FA38F87804251CB0FAD40562EC0B426149D17E0044B10A158B",
INIT_16 => X"5094246A10A10441010090480C0964201800044109012001A000726E45428000",
INIT_17 => X"0942509425094250942509425094250942509425094250942509425094250942",
INIT_18 => X"9425094250942509425094250942509425094250942509425094250942509425",
INIT_19 => X"02A8000000000000000000509425094250942509425094250942509425094250",
INIT_1A => X"BAFFD7F7F7F775555557DF9FE0FFBBEEFF3F7DF7FF3E7E2FF0087B9F7DF7E245",
INIT_1B => X"FD7EBF5FAFD7EBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAE",
INIT_1C => X"AFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FA",
INIT_1D => X"0557DE00000000000000000000000000000000000000000000001007FE0001DF",
INIT_1E => X"0004020BAAAFFD5400AAFBC2155AAAA97410FFFFEAAAAF7AA955EFF7803FF450",
INIT_1F => X"0F7AEBDE10FFFFFDEAAF7D568AAA5D002AB55005568B55087FC0010AAFBFFE10",
INIT_20 => X"FF5D04154BAAAAEAAA10557BEAA10AAFBE8A00557BFFFEF007BC215500001541",
INIT_21 => X"000A2AABFF45550400000AAFBFFFEF550000155A28415410F7AEAABFFA2D1555",
INIT_22 => X"8AAAFFFBC21555D517FF45F7AEA8BFFA2AEAAA10A280021EF5D557FF55AA8400",
INIT_23 => X"974AAF7D142145082A975FF555568A00FF842ABEFA2AAA8B5500003DF55F7D56",
INIT_24 => X"000145A2AA821EFFFFFD7410007FC0010555155555FF80174000055555EFAAAE",
INIT_25 => X"A0925C7E38E38F7D14557AE00000000000000000000000000000000000000000",
INIT_26 => X"075C7028B6F1FAE00000A02092B6F5D2438A2FBC2145B6A090428FFF5EAA92E3",
INIT_27 => X"1C7FC516D080E15438E3A4BAE00FFF5FAE92F7D16AAAA41042FB7D145568B7D0",
INIT_28 => X"8FFA4AFBFFAAD1505FF490E174AABEA0ADA005D7BEDA00B6F1EFA28557BF8FEF",
INIT_29 => X"FF555F7FF7DAA8E07028B6A0BFF6D490E00000BEF5FAFEF490407155BE8E1242",
INIT_2A => X"B551C0E3AF55F7DF68ABAE3F1C0145415B78F45FFA4AFBC7BEA4AAA10A284001",
INIT_2B => X"04380055525FFBEAE90482E3D54216D0024975FF555F68A00F7842FBD7B6AAAA",
INIT_2C => X"0000000000000000000016DAAA0851FFE3FBD0438007FC00385D555556DEB841",
INIT_2D => X"0020BAF7D16AA10A28402155A2AEA8BEF5D516AA000000000000000000000000",
INIT_2E => X"003DFEF55516ABEF0055574BAFFD568A10002A82000FFD5400AAA2FBC0145FF8",
INIT_2F => X"7D17FEBA557BEABEF557BD55EF082A974BAA28028A00F7D16AA10F7D56AABA08",
INIT_30 => X"000417545FFAA820BAFF843DFFFA2D5421FF002E954AAFF843DE105D7FFDE00F",
INIT_31 => X"5F7802AA10AA80001FF5D7FFDFEFA2AA974BAF7803FFFF002A82000FFD568BEF",
INIT_32 => X"10FF803DF45FFAEA8B555D2EAAB45F7FBE8ABAAAD540145007FE8B55FF843DF5",
INIT_33 => X"0AA5D55555FFA280000BA0855401EFF7AA82010AAD1421FF0004155FF557FEAA",
INIT_34 => X"00000000000000000000000000000000000001EFA280175FFAAFFC00BA087FC2",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"FFFFFFFE00000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000000000000000000019F",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(13),        -- Port A data input
DOA(0)   => data_read_a_lo(13),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(13),        -- Port B data input
DOB(0)   => data_read_b_lo(13),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_14_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10020A000180000284008280000281800000030000000033022000000580002",
INIT_01 => X"A140098018300848184860000C20C24040000000084000084200000000110200",
INIT_02 => X"88010C5A8010A600A4F558040080000041000000022C024008003CCCC9028030",
INIT_03 => X"000103A7A00904D0842242024210810803006480088000003081054288C10000",
INIT_04 => X"0000120122009000100C00000000000400A83A2044200C840000800400101820",
INIT_05 => X"020000004008010024C0C0010040000402000025000800020004207000100800",
INIT_06 => X"010000102000005043403AA14003004864000A00440812541020008230821000",
INIT_07 => X"2400A96850A16854200021DA2A0002000340800062C80819EBC402800008C020",
INIT_08 => X"0A0012140404414814E001000000000029FD0A10289924810182000110028010",
INIT_09 => X"080208222200400002000400420080010008C2C0032210020200008440000080",
INIT_0A => X"000000000203200E0620400011640446DA101004800005802004800000000000",
INIT_0B => X"282001001088A45000082408000010000910000800001000009A924810410000",
INIT_0C => X"0080000000000000080000000000000080000000000000000000100202000000",
INIT_0D => X"0100000004408020021010010001700042080880904000008808000000000800",
INIT_0E => X"00000000C00000000040302200800A0409020481024482501010413080008404",
INIT_0F => X"8090008142014840100002C38280000840100003838280000640204800000000",
INIT_10 => X"072C000444C00840020002C38280000840020003838280002C09D01086839746",
INIT_11 => X"D0104B01C57100440202900184414430534605E3804802180022480419183514",
INIT_12 => X"594C194000090450808802008830024F0E248C902AEF0024170CF18001003C09",
INIT_13 => X"20020E5A08E6000048200196264BCF1C030C0604800001076C04730000240049",
INIT_14 => X"2003DEDE82C78900902A0D0000080019FAAA32D9602490302409292B83280001",
INIT_15 => X"049100021171F6C34080240108AB292CA000000800AD1A19F6F000AA0C0A0000",
INIT_16 => X"4090246810810440000090480C0964200800000108010016000012004542800D",
INIT_17 => X"0902409024090240902409024090240902409024090240902409024090240902",
INIT_18 => X"9024090240902409024090240902409024090240902409024090240902409024",
INIT_19 => X"0280000000000000000000409024090240902409024090240902409024090240",
INIT_1A => X"9E7FDDF77777F3CF3CF7D54CEFD79B4E5C8FF0F7BE9D75C7F7B71F5F7DF65040",
INIT_1B => X"7F3F9FCFE7F3F9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7",
INIT_1C => X"E7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE",
INIT_1D => X"28417400000000000000000000000000000000000000000000001007FEFFFE0F",
INIT_1E => X"F7AA955EFF7803FF4500557DF45F7D16AB455D00001EFAAAAAAABA555557555A",
INIT_1F => X"555003FF450804001555D2AA8AAA002ABDE10082ABDF55AAAA97410FFFFEAAAA",
INIT_20 => X"EF5D5168A10082E80155087FC0010AAFBFFE100004020BAAAFFD5400AAFBC214",
INIT_21 => X"E10FFFFFDEAAF7D568AAA5D002AB55005568A00A2D5401455D00175FFFF84175",
INIT_22 => X"2155000015400AAD157545080402145087FD75FFF7AE82145A2D17FE10F7AEBD",
INIT_23 => X"000BAFFFBE8AAAA2FBFDE00087FD5410557BEAA10AAFBE8A00557BFFFEF007BC",
INIT_24 => X"000155A28415410F7AEAABFFA2D1555FF5D04154BAAAAEAAA005D002AB450000",
INIT_25 => X"A0AAA82555157555B68012400000000000000000000000000000000000000000",
INIT_26 => X"6A090428FFF5EAA92E3A0925C7E38E38F7D14557AF45FFDB6AB6D4100071C7B6",
INIT_27 => X"B6F5D2438A2FBC21455D0A3FF6D080407155552AAAA920020BFE10002EBAF45B",
INIT_28 => X"54100175C7E380125D7555B6DA1014248217D0075C7028B6F1FAE00000A02092",
INIT_29 => X"45AAD178E38E3A4BAE00FFF5FAE92F7D16AAAA41042FB7D145568A38AADF4014",
INIT_2A => X"A28557BF8FEF1C7FC516D080E15400A2DB5754508040716D007BD05EFEBAA821",
INIT_2B => X"DA0055002AB6D0000020BAFFF1E8ABABEF1FAE001C7FD54005D7BEDA00B6F1EF",
INIT_2C => X"00000000000000000000155BE8E12428FFA4AFBFFAAD1505FF490E174AABEA0A",
INIT_2D => X"FEABFF080015555F78028A00555155555FF84000000000000000000000000000",
INIT_2E => X"003DE10082EAAB45FF80020BAF7D16AA10A28402155A2AEA8BEF5D516AB45F7F",
INIT_2F => X"FD568A10002A82000FFD5400AAA2FBC0145552ABFFFF000417555552EA8A1000",
INIT_30 => X"55516AABAAAFFC0145000417555A280001455D7FFDE105504021EF0055574BAF",
INIT_31 => X"F007BC01FFAAAE80155AAD568ABAA28028A00F7D16AA10F7D56AABA08003DFEF",
INIT_32 => X"105D7FFDE00F7D17FEBA557BEABEF557BD55EF082A97410AAFFD55450800155F",
INIT_33 => X"1FF002E954AAFF843DE10550028BEF0004020BAF7D568AAAF7D168A105D7FD74",
INIT_34 => X"0000000000000000000000000000000000000145FFAA820BAFF843DFFFA2D542",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"FFFFFFFE00000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000000000000000000001F",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(14),        -- Port A data input
DOA(0)   => data_read_a_lo(14),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(14),        -- Port B data input
DOB(0)   => data_read_b_lo(14),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_15_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000A000000000284000280000001800020030000000033022000000180002",
INIT_01 => X"A140098018300848180060000C00424040000000080000080200000000110200",
INIT_02 => X"080108000010E60004E55800008000004100000000040240080000C009170016",
INIT_03 => X"0000000080000040842240000210810002000400888000003080014288C00000",
INIT_04 => X"0001100024A0800000440000000000040088322044200C840000011400151800",
INIT_05 => X"A200014C4000000020000000000B8094020000254C8800000514203000108800",
INIT_06 => X"000821000000A050434010A14001004844000801540812540020008600831000",
INIT_07 => X"C2000864489128502000210222000200034080006248081958C0008000088000",
INIT_08 => X"0A001214050540C800200101860000000B7C0910209900000002000110000010",
INIT_09 => X"0B0208222004400000000400420080010008C28002201002020001140800002C",
INIT_0A => X"000000000203000C04204000116404460810100080000F802004800000000000",
INIT_0B => X"280001001088A45000082008000010000100000800001000001A124800010000",
INIT_0C => X"0080000800008000000000000000000080000400004000000000100202000008",
INIT_0D => X"0100000004C00020025000018801600040000000000000008808000000000800",
INIT_0E => X"00108000C0000000000020020080080000000000000402000000000000009400",
INIT_0F => X"00000000000000404200000000000000404200000000000008C0004800000000",
INIT_10 => X"0000000000000040500000000000000040500000000000000400000100000000",
INIT_11 => X"0001000000000000000000000400020100000000000000000000080000240000",
INIT_12 => X"00110000000000C00080010180000000001A1024050000000000000000000400",
INIT_13 => X"0002008040000000002000000804002000000000000001000120000000000040",
INIT_14 => X"2000000061100280000000000008000001104422000000000008020020000000",
INIT_15 => X"00100000000009080E2E0A000000000000000008000004000000000000000000",
INIT_16 => X"0000046000000440000090480809402008000001000000000000000004188000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0280000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000040000000000040",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"8517DE00000000000000000000000000000000000000000000001007FE000000",
INIT_1E => X"AAAAAAABA555557555A284175FF000002010552A97400007BFDE10A2AA801EF0",
INIT_1F => X"F5D2AAAB45F7D17DF45087BC0155002A801FF08003DF45F7D16AB455D00001EF",
INIT_20 => X"45F7D568BEFAAD557555AAAA97410FFFFEAAAAF7AA955EFF7803FF4500557DFE",
INIT_21 => X"F450804001555D2AA8AAA002ABDE10082ABDFFFF7D17FE10002E954AAF7FBC21",
INIT_22 => X"5400AAFBC21EFA2AE95545A2D56ABFFAAD17DE10FFD1420AA007FC014555003F",
INIT_23 => X"801550055401555D00174BA002AA8B55087FC0010AAFBFFE100004020BAAAFFD",
INIT_24 => X"000000A2D5401455D00175FFFF84175EF5D5168A10082E801FFFF8428A10002A",
INIT_25 => X"71FAE00A2A0871EF145B7FE00000000000000000000000000000000000000000",
INIT_26 => X"FDB6AB6D4100071C7B6A0AAA82555157555B680125C71C0E0500049209543808",
INIT_27 => X"E38E38F7D14557AFC75524AFB45FFD178F7D1C71C2145002E801C7140A3FF45F",
INIT_28 => X"00024954AAFFFBC2145F7DB6DBEFA2D557545B6A090428FFF5EAA92E3A0925C7",
INIT_29 => X"820071C71455D0A3FF6D080407155552AAAA920020BFE10002EBAFC7FFDF7AE0",
INIT_2A => X"E00000A02092B6F5D2438A2FBC21FFBEA090545B6D568BFFAADB7AE10F7D5470",
INIT_2B => X"21FFE3802FA2808208017D1C5142155410A104AA1420AFB7D0075C7028B6F1FA",
INIT_2C => X"00000000000000000000038AADF401454100175C7E380125D7555B6DA1014248",
INIT_2D => X"E954100004174AA00516AA10AA80155EF5D7BFDE000000000000000000000000",
INIT_2E => X"2E801555D2EBDF45F7FFEABFF080015555F78028A00555155555FF8400155552",
INIT_2F => X"7D16AA10A28402155A2AEA8BEF5D516AB555D043DF55F7D56ABEF55514015508",
INIT_30 => X"082EAAB55FFFBE8A100804154AAF7FFC2145FFFFFDFEFAAD157545FF80020BAF",
INIT_31 => X"FA2FBE8A00FFD155410005555545552ABFFFF000417555552EA8A1000003DE10",
INIT_32 => X"EF0055574BAFFD568A10002A82000FFD5400AAA2FBC01FFF78400155F7D16ABE",
INIT_33 => X"1455D7FFDE105504021FFAA843DEBA0000021EF555142155002E800AA55003DF",
INIT_34 => X"00000000000000000000000000000000000000BAAAFFC0145000417555A28000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000180",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(15),        -- Port A data input
DOA(0)   => data_read_a_lo(15),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(15),        -- Port B data input
DOB(0)   => data_read_b_lo(15),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_16_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"DA22C618B1000482B688B186588884862A400438255FC38381441205BA803003",
INIT_01 => X"8645A80028404C211203A952A90341080B173340412000E1005D628000820484",
INIT_02 => X"A101A9006DC1084833011850AAC55001349B10881802821808B4110007005E11",
INIT_03 => X"010108A802BB00080080006020020001A61036202800000D2410104200404550",
INIT_04 => X"8BFA58800005C40A46240252145148B38248030356415A4E62B6FC660F287240",
INIT_05 => X"0F05EA11E570000D610000000710296E542B6E3A825C15FB30A643695BFC2D56",
INIT_06 => X"408003200040202B8584112645554B029006000140BCC0460050690A95C8383D",
INIT_07 => X"00480A2140040BE1480FA004342AA6F12000054004867415401DCDCF2AA10800",
INIT_08 => X"B32A8819064E48288012D45000005050247AA85220700009C06206C48080EDEA",
INIT_09 => X"445B2081340B6596594800400413CAC020894480000008C54C00311002000002",
INIT_0A => X"000000004B240028000342A00002FE00A3A1F06E491800AA29588181040A0020",
INIT_0B => X"2400848002912300200092BA80325A20000000000A8A5AA80018120E00066000",
INIT_0C => X"00220002200022000220002200022000210001100010000A40450100210072A0",
INIT_0D => X"002815014B90000205DA00880100095A648000000010006AC23000C7B69EC220",
INIT_0E => X"80922554515512174000000490009000000000000004010042A204A0C5817680",
INIT_0F => X"63EAA9C238B2D4C800632B266E828EE4C800632AAAB6830D0FC6B06C04102800",
INIT_10 => X"A149339E8FB964C800632B266E82B2E4C800632AAAB683310872800EDA52DA00",
INIT_11 => X"800EB090D4AAC91268FFCBE81397826C4A20D2B6C510E8624792A4A30A40839A",
INIT_12 => X"8849D5C532408DD6E004C90C06AC019D88B9795012CA96902C799912BC3C087A",
INIT_13 => X"531C74485BD42A30906057FADAA456218FD8E3ED83B60E3A242DC0F18983638E",
INIT_14 => X"A06FB555793057C444CF45C5C9E89543B8BC6E80193DC36F6C71D1093A478706",
INIT_15 => X"45DC02B331650CA8ACB4007E00D1C6A6A58395C917F7E74D936F650D69B51727",
INIT_16 => X"0000012000081500008A422150884081ACAAC0542054004FC588464050810DCD",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"147A7797E1E1A79E79E1560EEFBD11544C690DA64C1C69A9916D7E4F68A36040",
INIT_1B => X"7A7D1E9F47A7D345345345345345345345345345345345345345145145145145",
INIT_1C => X"4FA7D3E9F4FA3D1E8F47A3D1E8F47A3D1E9F4FA7D3E9F4FA7D3E9F4FA7D1E9F4",
INIT_1D => X"F8015400000000000000000000000000000000000000000000001007FE00001F",
INIT_1E => X"007BFDE10A2AA801EF08517DE10FFFFFDFEFA2D16AB55A2FFFFEAA5D7FC0000F",
INIT_1F => X"A5D2EBDFEFAAD17FFFF002EBDE000800174AA55043FFFF000002010552A97400",
INIT_20 => X"AAAA80000105D557FF45F7D16AB455D00001EFAAAAAAABA555557555A284174B",
INIT_21 => X"B45F7D17DF45087BC0155002A801FF08003DE000004154BA002A800BA087FE8A",
INIT_22 => X"FF4500557DEAAF7D57DEBA082A82010FFAE975555D7FFDEAAFF80155EF5D2AAA",
INIT_23 => X"7FFFF557FD55FF08003FE0055043FF55AAAA97410FFFFEAAAAF7AA955EFF7803",
INIT_24 => X"0001FFF7D17FE10002E954AAF7FBC2145F7D568BEFAAD557410552EA8BEFA2D5",
INIT_25 => X"FFFDEAA5571C7010FF8412400000000000000000000000000000000000000000",
INIT_26 => X"C0E050004920954380871FAE00A2A0871EF145B7FE10E3F1F8FC7AAD56DB7DB6",
INIT_27 => X"555157555B680124924124BDFEFA2D57FFC71C2EBDE280000174825D0E3FFC71",
INIT_28 => X"21424800AA007FEDAAAA284020385D5F7AF45FFDB6AB6D4100071C7B6A0AAA82",
INIT_29 => X"AAFF80175C75524AFB45FFD178F7D1C71C2145002E801C7140A3FE10080A1748",
INIT_2A => X"A92E3A0925C7E38E38F7D14557AE92EBDB78EAA1C2482010FFAE9556D557FF8E",
INIT_2B => X"7410492EADBEFA2D178FEF5575D55EF000A38E10490A3AF45B6A090428FFF5EA",
INIT_2C => X"000000000000000000001C7FFDF7AE000024954AAFFFBC2145F7DB6DBEFA2D55",
INIT_2D => X"56AB45A2D57DFFFF7FBFFEAA555555400F780000000000000000000000000000",
INIT_2E => X"0415400552ABDF55552E954100004174AA00516AA10AA80155EF5D7BFDE10A2D",
INIT_2F => X"80015555F78028A00555155555FF840000000043DFEFAAD17FF45552ABFEBA08",
INIT_30 => X"5D2EBDE10002E974005D04020BA007BFDEBAA284000BA557FE8B45F7FFEABFF0",
INIT_31 => X"0F7AE955EF5D7BE8ABAF784175555D043DF55F7D56ABEF555140155082E80155",
INIT_32 => X"45FF80020BAF7D16AA10A28402155A2AEA8BEF5D516AA00AAFBE8AAA55040000",
INIT_33 => X"145FFFFFDFEFAAD157410082ABFFEFAAD16ABFF5555575FF082AA8A00002AAAB",
INIT_34 => X"0000000000000000000000000000000000000155FFFBE8A100804154AAF7FFC2",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000080",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(16),        -- Port A data input
DOA(0)   => data_read_a_lo(16),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(16),        -- Port B data input
DOB(0)   => data_read_b_lo(16),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_17_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"5284CE4FB7BD2C8994A13392DBD02E14006B82AC7E800D44D3DD2FD5F9B961C0",
INIT_01 => X"F8ACD01F7E03FC6793F2199B39FC233C11D93AE6F3BB92B32091DBC339B24542",
INIT_02 => X"8F333007FD6808092A2AFA6667033DB50853379C10BFF70F1BD011110F205F18",
INIT_03 => X"294ADB4AFFCBF0DAD63ABF836B58EAFE060478202022234B2E0303FDC9E18339",
INIT_04 => X"DB7A40806FE4040840EBC563A0150A0926146FECB04196482236FC2005282AE1",
INIT_05 => X"0403DA0383200831C68206D7E6D0250834336D1E81500FDB306045255BFC2076",
INIT_06 => X"4470716040413D29AAC69F5FE33C072F06062C003670497AFF00291B3C0E2015",
INIT_07 => X"0849147160448EBB9537A0022DC67987042EE976ABEA77684653547819FF2000",
INIT_08 => X"E019C0C82A4E4820C15B089C380110002446045A31345000A84432409207F02D",
INIT_09 => X"983838A3BFF1030C397C060B4254064302042F803A69DB931FF4391C00002CC0",
INIT_0A => X"FB1F1F7BC81C003C001674BB55B5FBB4BB4F26A1BEE004F9D0DE08F7DE336DB2",
INIT_0B => X"28302F800633F1D0A7CC9AE74117FE01D34E82AC0CE8FCCC200A59BDD2FFE3E3",
INIT_0C => X"E9F79E9F79E9F79E9F79E9F79E9F79E9F7CF4FBCF4F000C2E225C8DE0BA05BB0",
INIT_0D => X"A5A99FD6D3FEF4BEB5FF994F0FEFFCCF8430000000D9D147E0D57AE7B79E9F79",
INIT_0E => X"0593F33FA0CF170F40006001B1A05C0000000000000008004BA78428C7AD7FE4",
INIT_0F => X"E46444357B3950A9BFBAC94CFA8581E0A9BFBAC8CCFA8580C7CAF51EF68B2976",
INIT_10 => X"B5DB54A09003E0A9BFBAC94CFA8581E0A9BFBAC8CCFA8580E46FBFCB0CBEDA57",
INIT_11 => X"BFCB1D5CFEB56A1A100D5345C1BFFE8FBDB892DB463034198E2881F3F787DF76",
INIT_12 => X"D39387F92B2935DFEAADDF38EBCFB9E3D636DCDF9B90F966BF92966D5D9E7467",
INIT_13 => X"27055EB6D555CB294981B7FB5B2954CD3013013FDF5E82AF5B6AAAE594A4E0AD",
INIT_14 => X"835C67E655BAA868610117575EA1C34BD6975D48B44A0405FC15BA7270FF2565",
INIT_15 => X"6CD2A47D0CBA96252756D7217E5E1C61DBDF5FA167F7AE5D3D21A414007F7D7E",
INIT_16 => X"000005F08000179C16DECF67F08BC02F9067ED55805600545DFE45A80E7BD07F",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"00C0000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"9A919261A1A6075D75D10DDF2F82003009EDCC4052E92E0826462117114F9818",
INIT_1B => X"8D068351A8D069A6BAE9A69A6BAE9A6BAE9A69A6BAE9A6BAE9A69A69A69A69A6",
INIT_1C => X"A8D46A351A8D46A351A8D46A351A8D46A341A0D068341A0D068341A0D068351A",
INIT_1D => X"AFFD5400000000000000000000000000000000000000000000001FFFFE000011",
INIT_1E => X"A2FFFFEAA5D7FC0000FF8015410FFFFFFFFFFFFFFDFEFF7D568A1008003DF55A",
INIT_1F => X"5A2D1400000804154BAF7D168A00A2803DE10FFAE95410FFFFFDFEFA2D16AB55",
INIT_20 => X"BAFFD56ABFF002EBDFFF000002010552A97400007BFDE10A2AA801EF08517DF5",
INIT_21 => X"FEFAAD17FFFF002EBDE000800174AA55043FEBA0004174AA5504000AA55042AA",
INIT_22 => X"7555A284175FFFFFBE8B55A2FFFFF55F7803DEBA002AAAAAAF7FBD74BA5D2EBD",
INIT_23 => X"17400FFD57DE00AAAAAAB45A2AA97545F7D16AB455D00001EFAAAAAAABA55555",
INIT_24 => X"0000000004154BA002A800BA087FE8AAAAA80000105D557FE00A2D5420AA5D04",
INIT_25 => X"D16AA00000E3DF6DBEF5D2400000000000000000000000000000000000000000",
INIT_26 => X"3F1F8FC7AAD56DB7DB6FFFDEAA5571C7010FF8412428FFFFFFFFFF7FBF8FD7EB",
INIT_27 => X"A2A0871EF145B7FF7DA2D547038140E10492FFDF6DA28A28E3DE00F7A092410E",
INIT_28 => X"2550A020BA55002AA82F7DF6DBD71C2EBFFC71C0E050004920954380871FAE00",
INIT_29 => X"BAF7F5D74924124BDFEFA2D57FFC71C2EBDE280000174825D0E3FEAA14001249",
INIT_2A => X"1C7B6A0AAA82555157555B680125FFEBFFEDB55BEFFFAF6DE38E3DEAA002EADA",
INIT_2B => X"AE28B6D545092490E10400FFDB7AE00A2AAADB45BEA092545FFDB6AB6D410007",
INIT_2C => X"00000000000000000000010080A174821424800AA007FEDAAAA284020385D5F7",
INIT_2D => X"BFDFEFF7FFEAB45A2D56AA00002EBDFFFF7D5400000000000000000000000000",
INIT_2E => X"AABDE10FF8400010A2D56AB45A2D57DFFFF7FBFFEAA555555400F780000AAFFF",
INIT_2F => X"004174AA00516AA10AA80155EF5D7BFDFEFAAD1554BA552E82000F7FFFFEAAA2",
INIT_30 => X"552ABDEBA5D0002000552A800BA55042AA10FFFFFDF55552EBDF55552E954100",
INIT_31 => X"FA2AEBFEAA082EBDEBAFFD55540000043DFEFAAD17FF45552ABFEBA080415400",
INIT_32 => X"45F7FFEABFF080015555F78028A00555155555FF84001FFAAFBFFF55FFFBEABF",
INIT_33 => X"EBAA284000BA557FE8AAAFFD155400082A82000F7FFE8A00A2AABDF45F780001",
INIT_34 => X"0000000000000000000000000000000000000010002E974005D04020BA007BFD",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"FFFFFFFE00000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000000000000000000019F",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(17),        -- Port A data input
DOA(0)   => data_read_a_lo(17),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(17),        -- Port B data input
DOB(0)   => data_read_b_lo(17),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_18_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"69844019080000A21A611406840014122A641074155FC28A2024001001801003",
INIT_01 => X"A643D920034004180005E9E3C90360C0041C0181002001602025800008440084",
INIT_02 => X"B7333980808408103F2000F81FC0FEDEAC2161B0B84D0002188011110C018041",
INIT_03 => X"0405D434003F2C020081587008020561E55116B0290000042B71240C800440F8",
INIT_04 => X"50805AC31007D6125724029216554A9847669903D640EC8E2001002604503004",
INIT_05 => X"07008000E0EA11803850C800010022660C1C0065003C0404002646DC20A02D40",
INIT_06 => X"0100001028040C093D0491A640FFC10028000280002C44D620F0228454C83810",
INIT_07 => X"08501620028007500CE801241021FE78E40486014006009044359DC707F55C20",
INIT_08 => X"9307CC082A0A4A6A01ECDCC40850001630080002A5CA500344040108120080AB",
INIT_09 => X"A0172083200B6186128040600C10C1C02009505081100088080BC6A052802001",
INIT_0A => X"002020000F0CA8428642430080438408A510185A40000008B83181C000141040",
INIT_0B => X"2E00C04C44C92A88DC42215C882E82240880000060D7030C30B885200D274404",
INIT_0C => X"10006100061000610006100061000610003080030800800C0540310130006E21",
INIT_0D => X"10202021000780004200408C1002003F66CA18A1B62622381B2B841840614006",
INIT_0E => X"806400FC503F08180050942E4200020C1B060D8306C182701404C19730108010",
INIT_0F => X"ABAF377DF1CA160820520EB3057E70E60820520F33057E72E915415900002900",
INIT_10 => X"5D48F37FAFEFE60820520EB3057E7CE60820520F33057E7EC658BF2DA7822AAB",
INIT_11 => X"BF2D4B2A80BF8FE39FD78EB0D882014A62C568FFAFC73FFDD9C2B30E0468A2AD",
INIT_12 => X"800DFC06F59F710107533C0C4E37619440FBFBAB2400AFC1600361D798F32658",
INIT_13 => X"EB9454005BAA36DEFF894823A3D1A88A2FE29D5FC6DCAA2A002DD51B6E7C728C",
INIT_14 => X"92A78606A28A5427AAB9FF4EDD251C7123E291660733EBF6FE519001BF40DEBB",
INIT_15 => X"AB58AFBFD5DE200A8EBE3A3EC110339E1DCEDC2590495BB2112E2BE4BF5F3B70",
INIT_16 => X"C1B06808348340000020301805002D008C1F92000A5F421B8000DB4910382202",
INIT_17 => X"1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06",
INIT_18 => X"B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C",
INIT_19 => X"000000000000000000000041B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1",
INIT_1A => X"8A244C16454170410412CA064A9BBECEB80EE173C2300FE3F1A3550F7DF16000",
INIT_1B => X"A552A944A2512AAA8A28A28A2AAAAAA8A28A28A2AAAAAA8A28A28A28A28A28A2",
INIT_1C => X"A25128944A25128944A25128944A25128944A25128944A25128944A25128954A",
INIT_1D => X"D2A80000000000000000000000000000000000000000000000001007FE000004",
INIT_1E => X"F7D568A1008003DF55AAFFD5410FFFFFFFFFFFFFFFFFFFFFBFDEBA552E974105",
INIT_1F => X"0FFFFFFFFFF7FBE8B55AAD16AA1000516AA005D0400010FFFFFFFFFFFFFFDFEF",
INIT_20 => X"00087BC2155087BC0010FFFFFDFEFA2D16AB55A2FFFFEAA5D7FC0000FF801541",
INIT_21 => X"0000804154BAF7D168A00A2803DE10FFAE95555FFFBE8B45A2D56ABEFFFFFFFE",
INIT_22 => X"01EF08517DF55000000010082A974AA08557DEBAFFAEBFF55AA8028B55A2D140",
INIT_23 => X"800105D2AAAA10A2D1420AAFFAEA8BFF000002010552A97400007BFDE10A2AA8",
INIT_24 => X"0000BA0004174AA5504000AA55042AABAFFD56ABFF002EBDEBA0004020BA552E",
INIT_25 => X"FBFFEBA552A95410552485000000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFF7FBF8FD7EBD16AA00000E3DF6DBEF5D2438FFFFFFFFFFFFFFFFEFF7",
INIT_27 => X"5571C7010FF8412410FFFBF8FC7E3F5EAB45BEDB6FA3800556FA00550405028F",
INIT_28 => X"5BEDB6FBC7EBF5F8E10007BC516D1C71C5010E3F1F8FC7AAD56DB7DB6FFFDEAA",
INIT_29 => X"55BE8A2DB7DA2D547038140E10492FFDF6DA28A28E3DE00F7A09256DE3F1EAB5",
INIT_2A => X"4380871FAE00A2A0871EF145B7FF45080E070280820924AA145578E92F7A4BFF",
INIT_2B => X"FEBA1C0A00092412E850005D2AAFA38A2DF45082F7AAA8BC71C0E05000492095",
INIT_2C => X"000000000000000000000AA140012492550A020BA55002AA82F7DF6DBD71C2EB",
INIT_2D => X"FFFFFFFFFBFDFEFF7FFFDEAA5D2E954105504154000000000000000000000000",
INIT_2E => X"557DE005500154AAFFFBFDFEFF7FFEAB45A2D56AA00002EBDFFFF7D5400AAFFF",
INIT_2F => X"2D57DFFFF7FBFFEAA555555400F78000010F7FBE8B55AAD16AB55F7FBFDEAA08",
INIT_30 => X"FF84001FFAAD568B45FFFBFFF55A2D568A00087BD55FF5D5555410A2D56AB45A",
INIT_31 => X"A555168A10FF803DF45FFAABDFEFAAD1554BA552E82000F7FFFFEAAA2AABDE10",
INIT_32 => X"55552E954100004174AA00516AA10AA80155EF5D7BFDF45002A974AA0800000A",
INIT_33 => X"A10FFFFFDF55552EBDEBA5D2E80010082A97410552EBDEBAA2FBD5400F7AAA8B",
INIT_34 => X"00000000000000000000000000000000000000BA5D0002000552A800BA55042A",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000080",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(18),        -- Port A data input
DOA(0)   => data_read_a_lo(18),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(18),        -- Port B data input
DOB(0)   => data_read_b_lo(18),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_19_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"042200000000000041088001001AA00000000000000000000000500802000003",
INIT_01 => X"200048000024000000000404000000000A22000800000800004A200000000001",
INIT_02 => X"032210008DEF00400060000001C008002489E0F0004037B00010101010000000",
INIT_03 => X"0000008128000000000000000000000024001620280000000000354200004008",
INIT_04 => X"000058800004C4024024001210001054B1C822009640000E2000002604003000",
INIT_05 => X"07008000E0200000000000000000200604000000001C04000026400000002C40",
INIT_06 => X"000000000000002600859AA1000D410000000000002C42010010200004C83810",
INIT_07 => X"0040380142810010564C41001140120024020280448088050008108100640000",
INIT_08 => X"83004C390242006200000868000040001020A850040AD0080426006933800DC4",
INIT_09 => X"0013200000016186100000000010C04002C00000000000707000000000000000",
INIT_0A => X"000000000B0C0000000101400040C0408100000000000008A810000000000000",
INIT_0B => X"00000000000400020000440000000000000000002F0001F00002024B20002000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"000210001D800000000000000002000964000000000000000000000000000000",
INIT_0E => X"0000000C50030008000000000000000000000000000000000000000000000000",
INIT_0F => X"101088A37034E156600D740022800EC156600D740022800D01E0412D06904000",
INIT_10 => X"0224081044914156600D7400228002C156600D7400228001098F00D0FB750500",
INIT_11 => X"00D0F2DD014010046037814EA63DBB31CE7605001008C41A061F0E7D693E6170",
INIT_12 => X"6D600000004089E12350C0E01FF23315422BABB46FEF5019146C0800380CC98F",
INIT_13 => X"130AA3592000000000629C03F3E60330C00C628908214551AC90000001036152",
INIT_14 => X"65C006070845039014460088235ACC3123E2A29148841008482A4DAC00000000",
INIT_15 => X"53A66BE7A5040018D8A8AD9090A1EC20A188235AC509FB50C2D0500B4094208D",
INIT_16 => X"000000000000000000000000000000008C01800270000061100084046086CD49",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"861A2882313054D34D301C862AA08BBA3F0C7010C6600A00200251C744192000",
INIT_1B => X"130984C261309861861861A69861861861861A69861861861861861861861861",
INIT_1C => X"6130984C26130984C26130984C26130984C26130984C26130984C261349A4C26",
INIT_1D => X"82E97400000000000000000000000000000000000000000000001007FE000002",
INIT_1E => X"FFFBFDEBA552E974105D2A801EFFFFFFFFFFFFFFFFFFFFFFFFFEAA552E954000",
INIT_1F => X"FFFFFFFFFFFFFFFFFEFF7FBFFEAA5D2E97545FFFFC2010FFFFFFFFFFFFFFFFFF",
INIT_20 => X"0008003DF555D5157410FFFFFFFFFFFFFFDFEFF7D568A1008003DF55AAFFD55E",
INIT_21 => X"FFFF7FBE8B55AAD16AA1000516AA005D04001EFFFFFFFFFFFFFBFDF45AAD16AA",
INIT_22 => X"0000FF80155EFFFFFFFFEFF7D16AB55A2D57DEBA557FEAA10080402010FFFFFF",
INIT_23 => X"6AB45FFFBFDEBA5D7FC0155FFFFD7410FFFFFDFEFA2D16AB55A2FFFFEAA5D7FC",
INIT_24 => X"000155FFFBE8B45A2D56ABEFFFFFFFE00087BC2155087BC00AAFFFBFDF45A2D5",
INIT_25 => X"FFFDEAA552E95400002095400000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFEFF7FBFFEBA552A954105524851C7FFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"000E3DF6DBEF5D25D7FFFFFFFFFFFFBFDFEFEBF5F8E92552E9556DEBF1C2038F",
INIT_28 => X"FE3F1FAF55A2D568A0000003FF7D495155428FFFFFFFFFF7FBF8FD7EBD16AA00",
INIT_29 => X"00000002010FFFBF8FC7E3F5EAB45BEDB6FA3800556FA005504051FFFFFFFDFE",
INIT_2A => X"B7DB6FFFDEAA5571C7010FF84125EFF7F1F8FC7EBD568B6DBEDF7DEBA5571EFA",
INIT_2B => X"5092E3F1F8F55AADB6DB7DEBF1FAE82557FC516DEBF1D0410E3F1F8FC7AAD56D",
INIT_2C => X"0000000000000000000016DE3F1EAB55BEDB6FBC7EBF5F8E10007BC516D1C71C",
INIT_2D => X"FFFFFFFFFFFFFFFFFFBFDEAA5D2A954000800154000000000000000000000000",
INIT_2E => X"2A955EFAAD1400AAFFFFFFFFFFFFBFDFEFF7FFFDEAA5D2E95410550415545FFF",
INIT_2F => X"7FFEAB45A2D56AA00002EBDFFFF7D540145FFFFFFFEFF7FBFFFFFAAD16AA0055",
INIT_30 => X"5500155EFF7FBFDFEFAAD568B55AAD568A0008003DFFF0855554AAFFFBFDFEFF",
INIT_31 => X"FFFFFFFEAA55517DE10080400010F7FBE8B55AAD16AB55F7FBFDEAA08557DE00",
INIT_32 => X"10A2D56AB45A2D57DFFFF7FBFFEAA555555400F780001FFF7D16AB55A2D16ABE",
INIT_33 => X"A00087BD55FF5D5555410AAD56AB45AAFFFFFEFAAD168A00557BD55FFA2D5400",
INIT_34 => X"00000000000000000000000000000000000001FFAAD568B45FFFBFFF55A2D568",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000100",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(19),        -- Port A data input
DOA(0)   => data_read_a_lo(19),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(19),        -- Port B data input
DOB(0)   => data_read_b_lo(19),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_20_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000003",
INIT_01 => X"A75FF80000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"14088080800008400F655001FFCFF80018FA8044000000000000011000000007",
INIT_03 => X"0000000000000000000000000000000024001660380000000000000000004FF8",
INIT_04 => X"000079800014CC02C034001600000000000000101EC0012EE0C0026E1E80F000",
INIT_05 => X"1F0FF433EFF0440C3902100002203F2EFC040388137C3E20C8EEC00284033CC0",
INIT_06 => X"4400080040440C000000000017FD5F239108000155FDC0000010E40087D8787A",
INIT_07 => X"08000EE00000000000000002101FF2002C00000004018001000030817FF50C00",
INIT_08 => X"FF7FCA302C0C00082148000008405550087C0000000000000002412489808000",
INIT_09 => X"44FF60000001EFBEF0040008023FDFC00000000040062A040001071004000013",
INIT_0A => X"000000002B7C0000008000000200000200A0C0040118400FABF9000000480002",
INIT_0B => X"0000000000000000000000000000004200310000000000000000200000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000400040",
INIT_0D => X"000000200000020000004000100203FF6C000000000000000000000000000000",
INIT_0E => X"00600FFC53FF001800000002004080000000000000040900005C848538000010",
INIT_0F => X"00009A9C300020080000800000003CC0080000800000003CC020007800000000",
INIT_10 => X"000000012963C0080000800000003CC0080000800000003CC100800000080000",
INIT_11 => X"800004000000000066C5000020020000000800000000C2E18001000200000800",
INIT_12 => X"000000000052B0200000014200040C2829000400000000000860F98798000100",
INIT_13 => X"4B00400000000002958000240400000000007E1B000040200000000001496004",
INIT_14 => X"4004181800000000005C5A00000200C40808000000000AF0D80080000000000A",
INIT_15 => X"0020141812737DC3020100400001C19C1D80000200400000000000015D140000",
INIT_16 => X"04010080800801810100000000000093EDFF8020000000000001001001000080",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0020000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0C8192608486879E79E681D903000030038200010089054D460400120104D204",
INIT_1B => X"86432190C86432CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB0C30C30C30C3",
INIT_1C => X"C86432190C86432190C86432190C86432190C86432190C86432190C86432190C",
INIT_1D => X"80402000000000000000000000000000000000000000000000001007FE000010",
INIT_1E => X"FFFFFFEAA552E95400082E975FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2A954100",
INIT_1F => X"0FFFFFFFFFFFFFFFFFFFFFFFDEAA5D2A954000800001EFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"BA5D2A97400FF8017410FFFFFFFFFFFFFFFFFFFFFBFDEBA552E974105D2A8000",
INIT_21 => X"FFFFFFFFFFEFF7FBFFEAA5D2E97545FFFFC21FFFFFFFFFFFFFFFFFFFFF7FBFFE",
INIT_22 => X"DF55AAFFD5400FFFFFFFFFFFFFFDFEFF7FFEAA10000417555AAD5555EFFFFFFF",
INIT_23 => X"FDFEFAAD568A0000043DF45AAFBC2010FFFFFFFFFFFFFFDFEFF7D568A1008003",
INIT_24 => X"0001EFFFFFFFFFFFFFBFDF45AAD16AA0008003DF555D51574BAFFFFFFFFFFFFB",
INIT_25 => X"FFFFEBA5D2A95410000A00000000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFDEAA552E954000020955FFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"552A95410552485010FFFFFFFFFFFFFFFFFFF7FBFDEBA5D2E95400140E001C7F",
INIT_28 => X"FFFFFFDFEFF7FFFFEAA5D2E95400E38A17438FFFFFFFFFFFFFFFFEFF7FBFFEBA",
INIT_29 => X"7DBEDF575D7FFFFFFFFFFFFBFDFEFEBF5F8E92552E9556DEBF1C21C7FFFFFFFF",
INIT_2A => X"FD7EBD16AA00000E3DF6DBEF5D2438FFFFFFFFFF7FBFDFC7EBF1E8A00080A155",
INIT_2B => X"5492FFFFFFFEFF7F1F8FD7A2D168A1008043FF6DAAFBC5028FFFFFFFFFF7FBF8",
INIT_2C => X"000000000000000000001FFFFFFFDFEFE3F1FAF55A2D568A0000003FF7D49515",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFEBA552A95410002E820000000000000000000000000",
INIT_2E => X"2E954005D2A82145FFFFFFFFFFFFFFFFFFFFFBFDEAA5D2A954000800155FFFFF",
INIT_2F => X"FFBFDFEFF7FFFDEAA5D2E95410550415410FFFFFFFFFFFFFFDFEFF7FBFFEBA55",
INIT_30 => X"AAD140155FFFFFFFFFF7FBFDFFFFFFBFDEBA5D2A95400A2AA974AAFFFFFFFFFF",
INIT_31 => X"5A2D568A10082E955FFFFFFD7545FFFFFFFEFF7FBFFFFFAAD16AA00552A955EF",
INIT_32 => X"AAFFFBFDFEFF7FFEAB45A2D56AA00002EBDFFFF7D5400BAFFFFFDFEFF7FBFFF5",
INIT_33 => X"A0008003DFFF085555410F7FBFDFEFFFD568B45AAD16AA1008003DFEFAAFBD74",
INIT_34 => X"00000000000000000000000000000000000001EFF7FBFDFEFAAD568B55AAD568",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"FFFFFFFE00000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000000000000000000001F",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(20),        -- Port A data input
DOA(0)   => data_read_a_lo(20),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(20),        -- Port B data input
DOB(0)   => data_read_b_lo(20),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_21_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"4A302428B824900A128C090A5C1800261500213C005FE812D10420054085A202",
INIT_01 => X"081FFE3440B609703B0427F801A40B8115BC4F655300340288A40D30040E4DD8",
INIT_02 => X"0109095C30C98809800000F9FFFFFFFF149FF1FCA4C0421B182E3490DF145FE4",
INIT_03 => X"084A76341244919000099486400026523C041660BA000100CC12701015007FF8",
INIT_04 => X"000079800014CC03C075161E001118653D2408041FC004AEF000816E1C11F541",
INIT_05 => X"3F0F807BFFE000240100004683103E7FFE02482553FC3C0204EFC25010143CC0",
INIT_06 => X"C42040304101118B84E4880817FD7F028000000101FFE4036450E08247F87870",
INIT_07 => X"0A09000D00204A855B000A08A61FF20C3D004D331D3400805984B7A1FFF00860",
INIT_08 => X"F7FFC08D234B4002030314D0001104500000034089902D0901A021E4015410EA",
INIT_09 => X"B4FFE10158E1FFBEF0440021083DFFCE22DC2880E24D1BFA7C98480802000023",
INIT_0A => X"A31514636FFC00080013029811240444A82422A85180778FAFF82A04B6356DD0",
INIT_0B => X"0600E20806520398C682157A49389667126880806FF917FC30010107688862A2",
INIT_0C => X"1B2451B2451B2451B2451B2451B2451B3228D9228D90800C6120881034003631",
INIT_0D => X"0403000A01282088624001201A8C43FF7C00100102A53208B2A246406081B245",
INIT_0E => X"C4053FFD5BFF00A04A00200602CA520011000880044402104803400400189000",
INIT_0F => X"63009140094D81A5040605800B506901A3040605401360562027218196506102",
INIT_10 => X"02811209062801A3040605800B506901A50406054013605604350B812822A002",
INIT_11 => X"0B811068C00049A0A5820A3C1725A8006C0A40404D058320496C2C9C600890A2",
INIT_12 => X"AC808127C454402483153A3A895BB3C1E2E820704020381702C1AAA2C4B3F435",
INIT_13 => X"CC1B154510413CC2A200501B400A40018A00C80400040D8AA288209AA2198361",
INIT_14 => X"0141AA00418080460678A4012288463B2050302019200B00206C35901024D910",
INIT_15 => X"2440470C8A9310280C0180302A01427D060022011606E800E00169C19A00048A",
INIT_16 => X"40100448008004000000E07008010003EFFFE0373056024B0111801198823314",
INIT_17 => X"0100401004010040100401004010040100401004010040100401004010040100",
INIT_18 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_19 => X"0000000000000000000000401004010040100401004010040100401004010040",
INIT_1A => X"BEFFFFF7F7FFF3CF3CFFFF9FE0FF9FEEFF7FFDF7FF3EFC2FF8107F3DFDF7E000",
INIT_1B => X"FF7FBFDFEFF7FBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEF",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FBFDFE",
INIT_1D => X"80002000000000000000000000000000000000000000000000001007FE00003F",
INIT_1E => X"FFFFFFEBA5D2A954100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974000",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFEBA552A97400082A975FFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"AA5D2E974100800155EFFFFFFFFFFFFFFFFFFFFFFFFFEAA552E95400082E975F",
INIT_21 => X"FFFFFFFFFFFFFFFFFDEAA5D2A95400080000000FFFFFFFFFFFFFFFFFFFFFFFDE",
INIT_22 => X"74105D2A80000FFFFFFFFFFFFFFFFFFFFFBFDEBA5D2E974005D2E80000FFFFFF",
INIT_23 => X"FFFFFF7FBFDEBA552A954005D2E97410FFFFFFFFFFFFFFFFFFFFFBFDEBA552E9",
INIT_24 => X"0001FFFFFFFFFFFFFFFFFFFFF7FBFFEBA5D2A97400FF80174BAFFFFFFFFFFFFF",
INIT_25 => X"FFFFEBA5D2E97400000400000000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFEBA5D2A95410000A001FFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"552E954000020955EFFFFFFFFFFFFFFFFFFFFFFFFFEAA552E97400002E955FFF",
INIT_28 => X"FFFFFFFFFFFFFBFDEAA5D2A974101400155C7FFFFFFFFFFFFFFFFFFFFFFFDEAA",
INIT_29 => X"00552A80010FFFFFFFFFFFFFFFFFFF7FBFDEBA5D2E95400140E00000FFFFFFFF",
INIT_2A => X"FEFF7FBFFEBA552A95410552485038FFFFFFFFFFFFFFFFFFF7FBFDEBA552E974",
INIT_2B => X"74AAFFFFFFFFFFFFFFFFEFF7FBFFEAA5D2E97400412497438FFFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000001C7FFFFFFFFFFFFFFDFEFF7FFFFEAA5D2E95400E38A1",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974000004000000000000000000000000000",
INIT_2E => X"2E97400002E975FFFFFFFFFFFFFFFFFFFFFFFFFFEBA552A95410002E821FFFFF",
INIT_2F => X"FFFFFFFFFFFBFDEAA5D2A954000800155EFFFFFFFFFFFFFFFFFFFFFFFFDEAA55",
INIT_30 => X"5D2A82010FFFFFFFFFFFFFFFFEFF7FBFDEBA552A974105D0015545FFFFFFFFFF",
INIT_31 => X"FF7FFFFEAA5D2A974005D2E82010FFFFFFFFFFFFFFDFEFF7FBFFEBA552E95400",
INIT_32 => X"AAFFFFFFFFFFFFBFDFEFF7FFFDEAA5D2E954105504154AAFFFFFFFFFFFFFFDFE",
INIT_33 => X"EBA5D2A95400A2AA974BAFFFFFFFFFF7FBFDFEFFFFFFDEBA552E974000004154",
INIT_34 => X"0000000000000000000000000000000000000155FFFFFFFFFF7FBFDFFFFFFBFD",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(21),        -- Port A data input
DOA(0)   => data_read_a_lo(21),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(21),        -- Port B data input
DOB(0)   => data_read_b_lo(21),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_22_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"5290F4CDE914905A14A43D33F488243E17122300F55FEB189B343A1140548380",
INIT_01 => X"A94007B259F6A975386262000C344BA9573C6FF57B18A5FB0ABFCD3C2C5F4F0C",
INIT_02 => X"877FE30EB378008D202551040030071869D0040180AC4B685F6E26FAA0810006",
INIT_03 => X"431965109E4481D6B5AAD6875AD6AB5A1815600802888808DEA83552954D3000",
INIT_04 => X"492C0020220001010E4916C884DCD607E5EC2A344103E48003D0800023D0072C",
INIT_05 => X"00107C441001100D620A06D683018001023D37E5088043620101179092540112",
INIT_06 => X"9108E1550544A451E0CE1AA94000206B541C08414402365774611E047020008E",
INIT_07 => X"809DA02F56A92FD7247E10305C40040D136E6A023F7FCF780C4C0528800C8028",
INIT_08 => X"00803A884B5B5206B7C3391F288551002401E993AF59012740A2E4F65586923D",
INIT_09 => X"040081C91AA010000560141801002028A83D2A08E06D0002FED9680A0E002A94",
INIT_0A => X"A71514E700838460402635019FBFE7FCA13520F8D580A08044081201206334A0",
INIT_0B => X"00A0220103D2A512C6A8C4F0011550070368000A0004D0000002126F30C902A2",
INIT_0C => X"0385503855038550385503855038550392A81C2A81C00280000C200006405A08",
INIT_0D => X"0D0E153941A8B1A262CA542A9A8D6C0010A1001002C500268ACA419412503855",
INIT_0E => X"089180008800143D83888281A2034A85014280A14050A01509E050854498B294",
INIT_0F => X"6706B3C189CD84ACD20B03001E387D04AC560B02401E387E1028AC0450080410",
INIT_10 => X"0201570B036C04AC560B03001E387D04ACD20B02401E387E24708E7E242000C2",
INIT_11 => X"8E7E1C20A0106EA167C84EBF052A8E010C0180606E86C3F459DC08DA90245887",
INIT_12 => X"189980254CDEC22A98032A22C50EAC462030A01800407C2700C2ACA2C0F04470",
INIT_13 => X"CC1154C258012D86F601A2E49003400138C0DA2443A208AA612C0096C3798225",
INIT_14 => X"025483C1E0C0006B085CEC03858958D15310201015504B512044A3133004A99B",
INIT_15 => X"9512C6FC01A1421006028038720640310643858162712020B001AA415F290E16",
INIT_16 => X"110445E22022365034A8EA754008004C0200323001182122548881649D16B046",
INIT_17 => X"1044110441104411044110441104411044110441104411044110441104411044",
INIT_18 => X"0401004010040100401004010040100401004010040100441104411044110441",
INIT_19 => X"22890000000003FFFFFFFF900401004010040100401004010040100401004010",
INIT_1A => X"9EFFDFF7F5F777DF7DF7DF5FEFBFBFDEFE8FF1F7DEBD6FEFF7EF6FDF7DF7D051",
INIT_1B => X"7F3F9FCFE7F3F9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7",
INIT_1C => X"E7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE",
INIT_1D => X"00000000000000000000000000000000000000000000000000001007FE00000F",
INIT_1E => X"FFFFFFEBA5D2E974000800021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E954000004001FFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"BA552A97400002A801FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2A954100804021F",
INIT_21 => X"FFFFFFFFFFFFFFFFFFEBA552A97400082A975FFFFFFFFFFFFFFFFFFFFFFFFFFE",
INIT_22 => X"5400082E975FFFFFFFFFFFFFFFFFFFFFFFFFFEAA552E95410002A955FFFFFFFF",
INIT_23 => X"FFFFFFFFFFFEAA552E95400002E975EFFFFFFFFFFFFFFFFFFFFFFFFFEAA552E9",
INIT_24 => X"000000FFFFFFFFFFFFFFFFFFFFFFFDEAA5D2E97410080015545FFFFFFFFFFFFF",
INIT_25 => X"FFFFEBA5D2E97410080002000000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974000004001FFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"5D2A95410000A001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2A954000804021FFF",
INIT_28 => X"FFFFFFFFFFFFFFFFEBA552A97400082E821FFFFFFFFFFFFFFFFFFFFFFFFFFEBA",
INIT_29 => X"10082A975EFFFFFFFFFFFFFFFFFFFFFFFFFEAA552E97400002E955FFFFFFFFFF",
INIT_2A => X"FFFFFFFFDEAA552E954000020955C7FFFFFFFFFFFFFFFFFFFFFFFFEAA552E954",
INIT_2B => X"5545FFFFFFFFFFFFFFFFFFFFFFFDEAA5D2A974001C24975C7FFFFFFFFFFFFFFF",
INIT_2C => X"00000000000000000000000FFFFFFFFFFFFFFFFFFFFFBFDEAA5D2A9741014001",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800020000000000000000000000000",
INIT_2E => X"2A954000800021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974000004001FFFFF",
INIT_2F => X"FFFFFFFFFFFFFFEBA552A95410002E821FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_30 => X"002E975EFFFFFFFFFFFFFFFFFFFFFFFFFEAA552A97400082A801FFFFFFFFFFFF",
INIT_31 => X"FFFFBFDEAA5D2E95410082E955EFFFFFFFFFFFFFFFFFFFFFFFFDEAA552E97400",
INIT_32 => X"45FFFFFFFFFFFFFFFFFFFFFBFDEAA5D2A95400080015545FFFFFFFFFFFFFFFFF",
INIT_33 => X"EBA552A974105D0015555FFFFFFFFFFFFFFFFFFF7FBFDEBA5D2A974005504175",
INIT_34 => X"0000000000000000000000000000000000000010FFFFFFFFFFFFFFFFEFF7FBFD",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"FFFFFFFE00000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000000000000000000001F",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(22),        -- Port A data input
DOA(0)   => data_read_a_lo(22),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(22),        -- Port B data input
DOB(0)   => data_read_b_lo(22),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_23_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"EF20906D902424807BC8241BC81801B97D38AD3C0800103362A6741C80A12A02",
INIT_01 => X"001FFF8409F089003B4422000D80C80106804A7951C5B9D1C828043EA28838F9",
INIT_02 => X"073B8858218C2C50801000F9FFEFF8E72CA7F5FC2E048026496834D84721DFE0",
INIT_03 => X"2C4360101A4001001005080400401420350016E0BB222341C312000014006FF8",
INIT_04 => X"00017B810015DC03D034201E14000036486008101FC0002EE006297E1C05F561",
INIT_05 => X"BF0F817FFFE80100004044800080BEFFFC0248005FFC3C18A5FFC2444484BCC0",
INIT_06 => X"00000070604191C93F02800017FF7F002000020001FFC0832050E00047F97870",
INIT_07 => X"AE4080091A0071070FA07A1CB23FFA403F0C4D23BF7C0EF85788B681FFFC6C20",
INIT_08 => X"F7FFD8880A034AC096620C46AC5055508401A24684227DB880000008B05001A3",
INIT_09 => X"21FFE0004047FFBEF2000000001DFFC612C0C04001000BF8000000804000003F",
INIT_0A => X"000000006FFEA002020626995FBE077430001E734020DF0FAFF5080496044B51",
INIT_0B => X"0600C48907120AC81083315A49388660180082A06FF907FC3081812048006000",
INIT_0C => X"182021820218202182021820218202182010C1010C10800C6120885430003631",
INIT_0D => X"80600020040030090000012A500003FF7E081881902233483828864860A18202",
INIT_0E => X"C7043FFD5FFF00A04BC010A7724B100008000400020000415003001000400002",
INIT_0F => X"290C2909080A872BC4FC8500054840072FC0FC8440054840200705F986106542",
INIT_10 => X"0180F1082E00072FC0FC8500054840072BC4FC84400548402214A380380B2080",
INIT_11 => X"A380344920080B21810240AB182EB37C380B40800707011001B43253EE50C822",
INIT_12 => X"E4000026C00C00042BD4149067465910640A0050C060A0028063672A00019214",
INIT_13 => X"800CCB050001344060211629580B80022480A444111706658280009A2030019C",
INIT_14 => X"232D6D0100C040250200845132C10BE200403018061101A220339C800004D801",
INIT_15 => X"2A5493B8E287E03808480060E40C83C1405132C90742E408D0082140820944CB",
INIT_16 => X"00802000100100000000000004002403EFFF8002385F03490101946500140210",
INIT_17 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_18 => X"8020080200802008020080200802008020080200802008020080200802008020",
INIT_19 => X"0000000000000000000000008020080200802008020080200802008020080200",
INIT_1A => X"0000000000000000000000000000000000000000000000000040000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"80400000000000000000000000000000000000000000000000001007FE000000",
INIT_1E => X"FFFFFFEBA5D2E974100000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100004021FFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"BA5D2E954000800001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974000800021F",
INIT_21 => X"FFFFFFFFFFFFFFFFFFEBA5D2E954000004001FFFFFFFFFFFFFFFFFFFFFFFFFFE",
INIT_22 => X"54100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2A954100000021FFFFFFFF",
INIT_23 => X"FFFFFFFFFFFEBA5D2A954100800021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2A9",
INIT_24 => X"0001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA552A97400002A801FFFFFFFFFFFFFFF",
INIT_25 => X"FFFFEBA5D2E97410080400000000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800021FFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"5D2E974000004001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100004021FFF",
INIT_28 => X"FFFFFFFFFFFFFFFFEBA5D2E954000800001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA",
INIT_29 => X"100004021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2A954000804021FFFFFFFFFF",
INIT_2A => X"FFFFFFFFFEBA5D2A95410000A001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2A954",
INIT_2B => X"21FFFFFFFFFFFFFFFFFFFFFFFFFFEBA552A97410080E001FFFFFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA552A97400082E8",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804000000000000000000000000000",
INIT_2E => X"2E974100000021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800021FFFFF",
INIT_2F => X"FFFFFFFFFFFFFFEBA5D2E974000004001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_30 => X"0800021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E954000804021FFFFFFFFFFFF",
INIT_31 => X"FFFFFFFEBA552A954100004001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2A95400",
INIT_32 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA552A95410002E821FFFFFFFFFFFFFFFFFFF",
INIT_33 => X"EAA552A97400082A801EFFFFFFFFFFFFFFFFFFFFFFFFFEAA552A97410002A821",
INIT_34 => X"00000000000000000000000000000000000001EFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"FFFFFFFE00000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000000000000000000001F",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(23),        -- Port A data input
DOA(0)   => data_read_a_lo(23),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(23),        -- Port B data input
DOB(0)   => data_read_b_lo(23),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_24_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100600007FFF000080108004000800020000840041000080808",
INIT_02 => X"172A00D000EF8210000000F9FFEFF8E7240FF1FC224087B1000639401D005FC0",
INIT_03 => X"00003A2E200811000000000400000000340016603A0000004860400014006FFF",
INIT_04 => X"000079800014CC03C034001E04010850300000101FC0002EE000006E1C00F500",
INIT_05 => X"1F0F8033FFE000000000000000003E2FFC024800137C3C0000EFC00000003CC0",
INIT_06 => X"00000040004111CE08AA800017FD7F000000000001FFC0000010E00007F87870",
INIT_07 => X"001080040814210254000A00B21FF2003F2A80D5000006E461803081FFF40000",
INIT_08 => X"F7FFD88D2B4A02C0940018EB0A1000058400810205E2D8030900004D925821CC",
INIT_09 => X"20FFE0000001FFBEF0000000001DFFC002C0000000000BF80000000000000003",
INIT_0A => X"000000006FFE80000015406A80000338800002500000470FAFF0080496044950",
INIT_0B => X"0600C008140800080000100248288660100080806FD107FC3000000000006000",
INIT_0C => X"182001820018200182001820018200182000C1000C10800C6020881030002431",
INIT_0D => X"000900160000000000000000000003FF7C001001002032083020060060018200",
INIT_0E => X"C4043FFD5BFF0000410000000041100000000000000000004003000000000000",
INIT_0F => X"1080012302010049400086C02200420049400087802200412027059996516100",
INIT_10 => X"0300081406100049400086C0220042004940008780220041248190818403A042",
INIT_11 => X"90814C09C01010400132100106836001504240E01040051200200D06410C1924",
INIT_12 => X"680C0100010408240BD80008983596CD86EA84104060503C0B00002025023481",
INIT_13 => X"90164F40086000082062C1B6600BC000C300818044000B27A0043000041202CD",
INIT_14 => X"2577FE4080C08010842180C40018545BBA00301808A0810C0059AD0180200020",
INIT_15 => X"04100852B931F00800010081980B042D2044001850ED8808F00050A002C11000",
INIT_16 => X"00000000000000000000000000000003EFFF80037046031E0110001100A4820C",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"BEC99E61848655D75D7FCB598CC0AEEAF6E7CC1132CD73C8261273B444199000",
INIT_1B => X"0F0783C1E0F07BEFBEFBEF9E79E79E79E79E7BEFBEFBEFBEFBEFBE7BE7BE7BE7",
INIT_1C => X"E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E",
INIT_1D => X"80402000000000000000000000000000000000000000000000001007FE000001",
INIT_1E => X"FFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800021FFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"BA5D2E974100000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100000001F",
INIT_21 => X"FFFFFFFFFFFFFFFFFFEBA5D2E974100004021FFFFFFFFFFFFFFFFFFFFFFFFFFE",
INIT_22 => X"74000800021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974000004001FFFFFFFF",
INIT_23 => X"FFFFFFFFFFFEBA5D2E974000800001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9",
INIT_24 => X"0001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E954000800001FFFFFFFFFFFFFFF",
INIT_25 => X"FFFFEBA5D2E97410080402000000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"5D2E974100800021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800021FFF",
INIT_28 => X"FFFFFFFFFFFFFFFFEBA5D2E974100000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA",
INIT_29 => X"000004001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100004021FFFFFFFFFF",
INIT_2A => X"FFFFFFFFFEBA5D2E974000004001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_2B => X"01FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E954000800021FFFFFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9540008000",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804020000000000000000000000000",
INIT_2E => X"2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFF",
INIT_2F => X"FFFFFFFFFFFFFFEBA5D2E974100800021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_30 => X"0000021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100000001FFFFFFFFFFFF",
INIT_31 => X"FFFFFFFEBA5D2E974000004021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E97410",
INIT_32 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974000004001FFFFFFFFFFFFFFFFFFF",
INIT_33 => X"EBA5D2E954000804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E954000004021",
INIT_34 => X"00000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(24),        -- Port A data input
DOA(0)   => data_read_a_lo(24),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(24),        -- Port B data input
DOB(0)   => data_read_b_lo(24),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_25_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100200002000000080100004000000020000800041000080808",
INIT_02 => X"1000218000000800000000F9FFEFF8E738FFF1FC20400400000004455A375FE0",
INIT_03 => X"00002000000001000000000400000000340016623A0000004000000014006FFF",
INIT_04 => X"924279824C94CC1BE0B4001F20000000020380401FE0082EF000106E1C00F500",
INIT_05 => X"1F0F8033FFF048202582800100523E2FFE024820137C3C0040EFE02000003CE4",
INIT_06 => X"D4A00671414191800000800017FD7F038100201101FFC0000010E08A07FC7870",
INIT_07 => X"080000000000000000000A00B21FF2003E0000000000066041803081FFFC2C60",
INIT_08 => X"F7FFFA0008000200A0400002280000050400800204000000000201202B800000",
INIT_09 => X"B4FFF0008001FFBEF80C40630C7DFFEEBAF0008002021BF80000400A02000003",
INIT_0A => X"000000006FFF800C0400000000000330080000500006470FAFFD29F7DE565971",
INIT_0B => X"0600C008040000080000100248688760101080806FD107FC3018000000006000",
INIT_0C => X"182001820018200182001820018200182000C1000C10800EE6618911398524B1",
INIT_0D => X"000000000000000000000002500003FF7C001001002032083120060060018200",
INIT_0E => X"C6043FFD5BFF00A04B80608003CB120C11060883044582114013412080000000",
INIT_0F => X"000000200200000900000400200000000900000400200000200701E186106140",
INIT_10 => X"0000001000000009000004002000000009000004002000000000808000002000",
INIT_11 => X"8080000800000000001010000002200000004000000004000000000240000020",
INIT_12 => X"2000000001000004031802000004100000100024400000000800800001000000",
INIT_13 => X"0000410000000008000000204004000000000100040000208000000004000004",
INIT_14 => X"0004200001000200000100040000004200004020000000040000840000000020",
INIT_15 => X"00000010800000000C0A00000000040000040000004080000000000000401000",
INIT_16 => X"451044C82082068C0200000008014023EFFFC006304602080100000100000308",
INIT_17 => X"1104411044110441104411044110441104411044110441104411044110441104",
INIT_18 => X"1044110441104411044110441104411044110441104411044110441104411044",
INIT_19 => X"00002FFFFFFFFFFFFFFFFFC11044110441104411044110441104411044110441",
INIT_1A => X"042824014C48569A69AFEE9E50B2894A196A8C5A2932F7C8086034EC15DA0808",
INIT_1B => X"6231188C46231249249249249249249249249041041041041041041249041249",
INIT_1C => X"562B158AC562B158AC562B158AC562B158AC562B158AC562B158AC56231188C4",
INIT_1D => X"80400000000000000000000000000000000000000000000000001FFFFE00002C",
INIT_1E => X"FFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"BA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001F",
INIT_21 => X"FFFFFFFFFFFFFFFFFFEBA5D2E974100800021FFFFFFFFFFFFFFFFFFFFFFFFFFE",
INIT_22 => X"74100000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800001FFFFFFFF",
INIT_23 => X"FFFFFFFFFFFEBA5D2E974100000021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9",
INIT_24 => X"0001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100000001FFFFFFFFFFFFFFF",
INIT_25 => X"FFFFEBA5D2E97410080400000000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFF",
INIT_28 => X"FFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA",
INIT_29 => X"100800001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800021FFFFFFFFFF",
INIT_2A => X"FFFFFFFFFEBA5D2E974100800021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_2B => X"01FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100000021FFFFFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741000000",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804000000000000000000000000000",
INIT_2E => X"2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFF",
INIT_2F => X"FFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_30 => X"0804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFF",
INIT_31 => X"FFFFFFFEBA5D2E974100800001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E97410",
INIT_32 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800021FFFFFFFFFFFFFFFFFFF",
INIT_33 => X"EBA5D2E974100000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800021",
INIT_34 => X"00000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"FFFFFFFE00000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000000000000000000001F",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(25),        -- Port A data input
DOA(0)   => data_read_a_lo(25),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(25),        -- Port B data input
DOB(0)   => data_read_b_lo(25),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_26_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"E9264EAB20190CA3BA4997AA9002AE9C001006B0778015CFA17E0811039879C7",
INIT_01 => X"F1FFF9BB1F773C7F9BB07DFFFDD863FC5FFF3FEFFBBF9FFB22FFFBC7B9F30686",
INIT_02 => X"1B33188302E708180F6FFBFFFFCFFFFF9C7FF7FC24350B99082400001D00DFD8",
INIT_03 => X"4A53D958C50000DCE7366303739CD98C27C57EF57980014F271807E3C9E9CFF8",
INIT_04 => X"DBFAFBD7FB1CDEBEF1BE17F7AC88042787FBFFF8FEE9FF7EE6F4C0EE1FFAF869",
INIT_05 => X"5F0FFEB3EFFEFFBDA7F7FED508707E2EFEBF6FFEB37C3FF302EEEDFF9B487CF6",
INIT_06 => X"67F2B27AFAD11587B7C094F1FFFFDF0FAF4E8FAA67FDDB7FB870FF30FFDEF87F",
INIT_07 => X"08180EF060C18E5BEFB051225CDFF7002C4EEDE77F6E0EFD044ABC817FFFDD35",
INIT_08 => X"FF7FC8790E46426CE06C2C7E381041460C7E8C1A35DF80000C0084C9188302E7",
INIT_09 => X"2CFF7A27B303EFBEFAFCC2E35E7FDFD147CCF3F583FA3FFF7D6000EC75088ED3",
INIT_0A => X"5A3A3B5AFF7CFACFAFE776F39FF7077E29D83CFAE601602FEBFFCDF7DEE77DF7",
INIT_0B => X"3EB1EDDCDEBCFF589807B70AD9A99EE41FD18884FFF19FFC71FEFED7B251E747",
INIT_0C => X"1AF181AF181AF181AF181AF181AF181AF4C0D78C0D718ADEEE61D99B7BE2A433",
INIT_0D => X"B9EC20181CC1F73F87501DED3409BFFFEFFEBCEBFE68370CFA6D07407481EF18",
INIT_0E => X"CE04FFFFF3FF1F5F5475BD7F72E4D75EBFAF5FD7AFEFDFFAF59B6FF28FE1D406",
INIT_0F => X"7C040101480807D17B0004001F804007D17B0004001F8040212F35FFC6D86D70",
INIT_10 => X"0001DC00068007D17B0004001F804007D17B0004001F804006F6008140002000",
INIT_11 => X"0081800800007B000102C0801FB02683800040007700011801003DE050A70020",
INIT_12 => X"32130207080D012CEFF41008D188D502100B02004000F01900039020040206F6",
INIT_13 => X"A01F21A2C40039006823F80048100003F0008004D8100F90D162001C803403E2",
INIT_14 => X"27F020A07400007C040085581019D602451500001EC00100247C46426080E101",
INIT_15 => X"2010EA40EA00020C830100F0D000022180581019F40084800001F100020B6040",
INIT_16 => X"EFFBFEFDFDDFE7DD87FEFF7FF796FFFFFDFFC017FEFFD7E841001D8197DCC3F0",
INIT_17 => X"BFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAF",
INIT_18 => X"FAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFE",
INIT_19 => X"88646FFFFFFFFFFFFFFFFFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEB",
INIT_1A => X"86EBCAF55357E1C71C751D53C44B15BCF491E166CC853E8117696853F86EDB5C",
INIT_1B => X"130984C261309861861861861861861861861861861861861861861A69A69861",
INIT_1C => X"6130984C26130984C26130984C26130984C26130984C26130984C26130984C26",
INIT_1D => X"80400000000000000000000000000000000000000000000000001007FE000002",
INIT_1E => X"FFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"BA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021F",
INIT_21 => X"FFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFE",
INIT_22 => X"74100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFF",
INIT_23 => X"FFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9",
INIT_24 => X"0001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFF",
INIT_25 => X"FFFFEBA5D2E97410080400000000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFF",
INIT_28 => X"FFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA",
INIT_29 => X"100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFF",
INIT_2A => X"FFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_2B => X"21FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008040",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804000000000000000000000000000",
INIT_2E => X"2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFF",
INIT_2F => X"FFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_30 => X"0804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFF",
INIT_31 => X"FFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E97410",
INIT_32 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFF",
INIT_33 => X"EBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001",
INIT_34 => X"00000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(26),        -- Port A data input
DOA(0)   => data_read_a_lo(26),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(26),        -- Port B data input
DOB(0)   => data_read_b_lo(26),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_27_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"00080A40000A41248002029000050A088000008242A0004404480002000A1155",
INIT_01 => X"F1FFF1C11F781C129C107DFFFE0860941E81258CA2B71C2220EC1B86E1A00002",
INIT_02 => X"4000002100000014400FF6FFFF0FFFFF8007F1FC211100014200800000887FC0",
INIT_03 => X"0842D85841000098C63061026318C18404C459757000015F00088BE3C0618FF8",
INIT_04 => X"DBEAE5D6D91C2EBCE1B21EA72C00000007FBE7C8F8E9EF79E6D440E91FDAE061",
INIT_05 => X"5C8FFCB38FF6B68984B5BCE408347E28FEBF6FEEB3723F7102E8EDBF8A4872F6",
INIT_06 => X"6E62106ADAD14180035044F1FFFC9F0C0E4C8DAAEFF1DB7FA868FE30EF1CE47E",
INIT_07 => X"0014401060C180190310540118DFF1000C0849673F6C06FE000A38007FF13115",
INIT_08 => X"F47FC80208808210880C00020814000044008C1A340C00000A08000000210000",
INIT_09 => X"04FC721491038F7DF8BEC2E39C5F1FD047CEF1B582D83FF779200062B12A8EC3",
INIT_0A => X"02606042787C5AC5ADC424B39FB6073D00D8048A6201002F83F04DFFDE83FDD6",
INIT_0B => X"56B5F0DEFABC705488069302DBA98EAC16C1A884FFE18FFD757E7ED7A211EC0C",
INIT_0C => X"186881868818688186881868818688187840C3440C35A8DFEE61CB9979AAA433",
INIT_0D => X"D1F820101441DA3A8310198C34089BFF8DD6B56B6F28378C7E2D07007801C688",
INIT_0E => X"E4047FFD23FF315D54358D593474955AB6AD5B56ADAB5FAAE58B2F628EA0C407",
INIT_0F => X"7C0400004C080791290004001D80001791290004001D8000210F15879715710A",
INIT_10 => X"0001DC0000801791290004001D80001791290004001D800012F6008040002000",
INIT_11 => X"0080800800007B000000E0801BB020828000400077000008210035E040830020",
INIT_12 => X"220202070801010C6F1410085188D500100102004000F01900031000060202F6",
INIT_13 => X"205D2120840039000813F80040100003F0000000F8100E909042001C80040BA2",
INIT_14 => X"07F020201400007C040001781011D602040500001EC00000057444404080E100",
INIT_15 => X"2000EA40EA000004810100F0D000020080781011F40080800001F1000003E040",
INIT_16 => X"AB6BDE75ED5EC71385FC2512E3565BBBF1FFC00636EED7E841000D81924C43F0",
INIT_17 => X"B6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6AD",
INIT_18 => X"6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADA",
INIT_19 => X"88747FFFFFFFFFFFFFFFFFAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB",
INIT_1A => X"00780401CBC8400000052412F84E2168100481CA8604368008402F02104A4716",
INIT_1B => X"4020100804020000000000000000000000000000000000000000208000000000",
INIT_1C => X"140A05028140A05028140A05028140A05028140A05028140A050281402010080",
INIT_1D => X"80400000000000000000000000000000000000000000000000001007FE000028",
INIT_1E => X"FFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"BA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001F",
INIT_21 => X"FFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFE",
INIT_22 => X"74100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFF",
INIT_23 => X"FFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9",
INIT_24 => X"0001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFF",
INIT_25 => X"FFFFEBA5D2E97410080400000000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFF",
INIT_28 => X"FFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA",
INIT_29 => X"100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFF",
INIT_2A => X"FFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_2B => X"21FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008040",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804000000000000000000000000000",
INIT_2E => X"2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFF",
INIT_2F => X"FFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_30 => X"0804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFF",
INIT_31 => X"FFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E97410",
INIT_32 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFF",
INIT_33 => X"EBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021",
INIT_34 => X"00000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"FFFFFFFE00000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000000000000000000001F",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(27),        -- Port A data input
DOA(0)   => data_read_a_lo(27),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(27),        -- Port B data input
DOB(0)   => data_read_b_lo(27),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_28_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"02200AA400180030808802A900002A08001280A08A801044104A1000001818C3",
INIT_01 => X"50A00011460214428114180000882214413D0A71592A01D92213D28005210202",
INIT_02 => X"1444428102100884000AA30200000000C1000401041108404400022220800000",
INIT_03 => X"461080404900000C6314A900318C52A40051081000888806108802A141288001",
INIT_04 => X"00800040110102000902002000888400081045A8A00003C00000500000080008",
INIT_05 => X"0000000000024CA0A0101800032000400000000B800000014000000B08180000",
INIT_06 => X"0040B0000804001040000450A00080444A002480220009A88800009A88000000",
INIT_07 => X"088400122448908A204020004080010000408200000001000002080000099000",
INIT_08 => X"0000028040101004200C21002084555500004489120509244022801244810210",
INIT_09 => X"9000008101400000049016080102000220001110001020058320402A16002650",
INIT_0A => X"A53534A50000080080E041000000008000C81000220020A00004000000300003",
INIT_0B => X"0090024440245400082D0220800008000081022C0000080000206CB0821086A6",
INIT_0C => X"02C0A02C0A02C0A02C0A02C0A02C0A02C050160501600240010860CC04200280",
INIT_0D => X"1884200810C1631181500CA60400B40080720020240A00004005800800206C0A",
INIT_0E => X"0A00C000200005000010040A0020CC000200010000800920040804020A605400",
INIT_0F => X"0000000140000010290000000280000010290000000280000100180210410442",
INIT_10 => X"0000000004800010290000000280000010290000000280000002000040000000",
INIT_11 => X"0000800000000000000280000010008280000000000000180000002000830000",
INIT_12 => X"0202020000090100548000000080000010010200000000000000900000000002",
INIT_13 => X"2000202084000000480008000010000000000004880000101042000000240002",
INIT_14 => X"0080002014000000000005080000800004050000000000002400404040800001",
INIT_15 => X"00002000000000048100000000000020800800008000008000000000000A2000",
INIT_16 => X"80210810840861CD33548542A10209D4100000010200400000000880035840A0",
INIT_17 => X"0200802008020080200802008020080200802008020080200802008020080200",
INIT_18 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_19 => X"22E1000000000000000000002008020080200802008020080200802008020080",
INIT_1A => X"200360D4141D630C30C7788C0211102C110A00246972C0C19D0154BD89A40A0C",
INIT_1B => X"6030180C06030208208208208208208208208208208208208208208208208208",
INIT_1C => X"160B0582C160B0582C160B0582C160B0582C160B0582C160B0582C16030180C0",
INIT_1D => X"80400000000000000000000000000000000000000000000000001007FE00002C",
INIT_1E => X"FFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"BA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001F",
INIT_21 => X"FFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFE",
INIT_22 => X"74100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFF",
INIT_23 => X"FFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9",
INIT_24 => X"0001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFF",
INIT_25 => X"FFFFEBA5D2E97410080400000000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFF",
INIT_28 => X"FFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA",
INIT_29 => X"100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFF",
INIT_2A => X"FFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_2B => X"01FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008040",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804000000000000000000000000000",
INIT_2E => X"2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFF",
INIT_2F => X"FFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_30 => X"0804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFF",
INIT_31 => X"FFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E97410",
INIT_32 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFF",
INIT_33 => X"EBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001",
INIT_34 => X"00000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"FFFFFFFE00000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000000000000000000001F",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(28),        -- Port A data input
DOA(0)   => data_read_a_lo(28),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(28),        -- Port B data input
DOB(0)   => data_read_b_lo(28),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_29_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"79964E4BA01DACAB9E659792D00AAE160002829C7FDFEFCEE97C2815039D70C3",
INIT_01 => X"50BFF9AB0775343F9AB01DF80D5821FC0FFF3FEFD1AF9FF1207FFBC7B9720586",
INIT_02 => X"0B33180300E700080F6AAA7BFFC007189C7FF2FC003503980A0000001D00DFD8",
INIT_03 => X"0401D940CD0000C8421A2B03210868AC23403E903900010E271006A148A0C000",
INIT_04 => X"49B87A417315D20A313E17F1800000058013DDF8BE21F36E02F0D06E03E8F800",
INIT_05 => X"1F007E33E01A4D9C87525E5101603E6E023D27DA937C03E340EE25CB9B483C12",
INIT_06 => X"4570301028001487B7809450B7FFC007AB0E068023FC3BFC98101F109FC6780F",
INIT_07 => X"00080EF020408EC8CFA01122149FF700200665A35D260B250442BC8100177C20",
INIT_08 => X"FF00007906464068406C0C7E100000020C7E840A15D6800044200049180300E7",
INIT_09 => X"A8FF18222341E0820AD40201423FC00122C4935001722BFD056040A452000443",
INIT_0A => X"5A2A2B5AAF00A80A82C332D18ED301D229C82C7AA600402FE80B8813485534A2",
INIT_0B => X"28102D445624DB481806A628810018400B9100042FF0180000ABFEF892508545",
INIT_0C => X"00D1A00D1A00D1A00D1A00D1A00D1A00D4D0068D006000428200508A0A600280",
INIT_0D => X"B0E8201018C1561E855008C50401B7FFE27A08A0B64A0100CA45814814A04D1A",
INIT_0E => X"4400DFFFF0001F1F0050342D42A086040B02058102C48970541944B20FA15402",
INIT_0F => X"00000101480000507B00000002804000507B000000028040212034FAD2892832",
INIT_10 => X"00000000068000507B00000002804000507B0000000280400402000140000000",
INIT_11 => X"00018000000000000102C0000410068380000000000001180000082010A70000",
INIT_12 => X"12130200000D0120ED64000080800002100B0200000000000000902004000402",
INIT_13 => X"A00220A2C4000000682008000810000000008004D80001105162000000340042",
INIT_14 => X"208000A074000000000085580008800045150000000001002408424260800001",
INIT_15 => X"001020000000020C8300000000000021805800088000048000000000020B6000",
INIT_16 => X"C4B12C989489418D13FE7F3FFD8BADB7FC004012CA5141600000198087D8C0F0",
INIT_17 => X"0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02",
INIT_18 => X"B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C",
INIT_19 => X"00602FFFFFFFFFFFFFFFFFC0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0",
INIT_1A => X"AEFFFFF7E7EFBFFFFFFAEF1DE1EF9F96EE7FFDF7FE78FC2FE8847F3FFDFFEA0C",
INIT_1B => X"F7FBFDFEFF7FBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBAEBAEBAEBAEB",
INIT_1C => X"FF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEF",
INIT_1D => X"80400000000000000000000000000000000000000000000000001007FE00003E",
INIT_1E => X"FFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"BA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001F",
INIT_21 => X"FFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFE",
INIT_22 => X"74100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFF",
INIT_23 => X"FFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9",
INIT_24 => X"0001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFF",
INIT_25 => X"FFFFEBA5D2E97410080400000000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFF",
INIT_28 => X"FFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA",
INIT_29 => X"100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFF",
INIT_2A => X"FFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_2B => X"01FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008040",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804000000000000000000000000000",
INIT_2E => X"2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFF",
INIT_2F => X"FFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_30 => X"0804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFF",
INIT_31 => X"FFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E97410",
INIT_32 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFF",
INIT_33 => X"EBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001",
INIT_34 => X"00000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(29),        -- Port A data input
DOA(0)   => data_read_a_lo(29),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(29),        -- Port B data input
DOB(0)   => data_read_b_lo(29),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_30_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"9EEBFEF5D7D7F7DF7DFFDFDFCEFFBFFEFF9FE1F7FFBFEFC9B77B7FFFFDFFD000",
INIT_1B => X"7F3F9FCFE7F3F9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7",
INIT_1C => X"E7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE",
INIT_1D => X"80400000000000000000000000000000000000000000000000001007FE00000F",
INIT_1E => X"FFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"BA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001F",
INIT_21 => X"FFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFE",
INIT_22 => X"74100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFF",
INIT_23 => X"FFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9",
INIT_24 => X"0001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFF",
INIT_25 => X"FFFFEBA5D2E97410080400000000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFF",
INIT_28 => X"FFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA",
INIT_29 => X"100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFF",
INIT_2A => X"FFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_2B => X"01FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008040",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804000000000000000000000000000",
INIT_2E => X"2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFF",
INIT_2F => X"FFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_30 => X"0804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFF",
INIT_31 => X"FFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E97410",
INIT_32 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFF",
INIT_33 => X"EBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001",
INIT_34 => X"00000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(30),        -- Port A data input
DOA(0)   => data_read_a_lo(30),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(30),        -- Port B data input
DOB(0)   => data_read_b_lo(30),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_31_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"129000008004A00804A40000400800020000000C005FEA005800200400050100",
INIT_01 => X"A15FF18019700810180065FFFC0040801E80258CA2951C2200EC0906A0804140",
INIT_02 => X"0000000000000011000550FDFF0FFFFF0007F1FC200000011000000000205FC0",
INIT_03 => X"08425818000000908428C0024210A30004045060302223490002014280410FF8",
INIT_04 => X"DB6A618248140C18E0B016872400000007EBA24058E1ECA8E2D400681FD0E061",
INIT_05 => X"1C0FFC338FF01009048084C400103E28FE3F6FE513703F7000E8E5B4825030F6",
INIT_06 => X"4420006040410180034000A157FC1F08040C080045F1F2572060FE82671C607E",
INIT_07 => X"001100004081001103107000185FF0000C0849673F6C06FC000830007FF00000",
INIT_08 => X"F47FC80008000200800000020811000004008812240800000800000000000000",
INIT_09 => X"04FC700090038F3CF82C44630C5D1FC002CCE08082481BF27A00000000000883",
INIT_0A => X"00000000687C0044040424B39FB6073C0010048A4000008F83F009F7DE037DD0",
INIT_0B => X"0620E08812982050800A910249298624124080886FE187FC301B124F20016000",
INIT_0C => X"182001820018200182001820018200183000C1000C10808EE661891139802431",
INIT_0D => X"816800100400902A0200110810080BFF0C8010010220330C3A28070070018200",
INIT_0E => X"C4043FFD03FF101D400080013040180810040802040102004183012084808006",
INIT_0F => X"7C04000008080781000004001D00000781000004001D0000200F018586106100",
INIT_10 => X"0001DC0000000781000004001D00000781000004001D000002F4008000002000",
INIT_11 => X"0080000800007B00000040801BA020000000400077000000010035C040000020",
INIT_12 => X"200000070800000C231410085108D500000000004000F01900030000040202F4",
INIT_13 => X"001D0100000039000003F00040000003F000000050100E808000001C800003A0",
INIT_14 => X"077020000000007C0400005010115602000000001EC00000007404000000E100",
INIT_15 => X"2000CA40EA000000000100F0D000020000501011740080000001F10000014040",
INIT_16 => X"010044602002061004A820104809402BE1FFC006304E03684100050190040350",
INIT_17 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_18 => X"0040100401004010040100401004010040100401004010040100401004010040",
INIT_19 => X"00802FFFFFFFFFFFFFFFFF810040100401004010040100401004010040100401",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000010",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"80400000000000000000000000000000000000000000000000001007FE000000",
INIT_1E => X"FFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"BA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001F",
INIT_21 => X"FFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFE",
INIT_22 => X"74100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFF",
INIT_23 => X"FFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9",
INIT_24 => X"0001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFF",
INIT_25 => X"FFFFEBA5D2E97410080400000000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFF",
INIT_28 => X"FFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA",
INIT_29 => X"100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFF",
INIT_2A => X"FFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_2B => X"01FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008040",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804000000000000000000000000000",
INIT_2E => X"2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFF",
INIT_2F => X"FFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_30 => X"0804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFF",
INIT_31 => X"FFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E97410",
INIT_32 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFF",
INIT_33 => X"EBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001",
INIT_34 => X"00000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(31),        -- Port A data input
DOA(0)   => data_read_a_lo(31),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(31),        -- Port B data input
DOB(0)   => data_read_b_lo(31),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_0_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"ED39BA795990D275FB4A6E96ACC4731DEA4598B0AFB54867F6EE4618C3749807",
INIT_01 => X"58A0047D8607944AC7DA180001ECA2544042106208408208C20022E9173734B3",
INIT_02 => X"9F775E7CB273E6CCA7DAAF00001000000478020113C9C38E09FB7CCCDD9F203E",
INIT_03 => X"441406267B4CB04443163C91110C58F24A31000B8028A810A3D0F8B169A01006",
INIT_04 => X"0005802424830120024121209088809DF81454ACA01E03501D0A3B91E00F0A00",
INIT_05 => X"E0F001CC00012034C20B0232838F80D001C0100AEC83C008EF101A034C8CC300",
INIT_06 => X"908A0D058584A45164BE6E58A000000583F08459A2000DA8C40F003C80030780",
INIT_07 => X"E6CCAFDC3870EEEEC44E2BDFE220094D03022210C011C103FB860B28000007C9",
INIT_08 => X"080032BF07C7C1FC3F87253D96C45557ABFF070C19D62C9065EAF36919FCB273",
INIT_09 => X"DB0009EF68EC0000045082984202002DB93119096025040581B9691E8A88262C",
INIT_0A => X"8014546E000344A0488111084048E082D0ED020133A6BF200005F60820B88206",
INIT_0B => X"28000947E16656074EA560F08054490B01280A26900C4800814069B0C8888008",
INIT_0C => X"03DCF03CCF03DCF03CCF03DCF03CCF038E780C6781C008500804708A42255A88",
INIT_0D => X"7095352BD2A90515A1CA44E7EA84B00001010012008700624187C09C0E707CCF",
INIT_0E => X"0B92800224008AE09F8942C48D1BC49120489024481225058860128543287291",
INIT_0F => X"038ABACB83C7E03EA5FF83C002783F103EA5FF83C002783F0120847A70470C7E",
INIT_10 => X"0380230F2D7C103EACFF83C002783F103EACFF83C002783F310BBF7EFC2B80C2",
INIT_11 => X"BF7EFC61E01804E1E6EA1E3FA01FD97EFC4B80E008C7C2F678FF023FAF5BD987",
INIT_12 => X"CC8E8320C4DAC9220C6B2FF22EF72ADDE6F1A67C80600C2683E0EF8AE1F1F10B",
INIT_13 => X"5C00FE651C6104C6D6400FFFB01FC0000FC07EE42FA7C07F22CE3082636B801F",
INIT_14 => X"C08FDF4195C0C2038A7C6CAFA7E289F9BA4570380131CAFB2003F9D190A4189B",
INIT_15 => X"9FE635BE11B7F0308D4A80092E0FC1FC662FA7E283FF68A8F0080AE1DDA8BE9F",
INIT_16 => X"12058312C1241140A056954AB0D680D000003350013024179498C2EC6B9270AE",
INIT_17 => X"2048120481204812048120481204812048120481204812048120481204812048",
INIT_18 => X"0481204812048120481204812048120481204812048120481204812048120481",
INIT_19 => X"2859400000000000000000120481204812048120481204812048120481204812",
INIT_1A => X"082218821390771C71C557C449F3898E09B56C74DAB16787E0760E5D1CF13043",
INIT_1B => X"7C3E1F0F87C3E082082082082082082082082082082082082082082082082082",
INIT_1C => X"87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F8",
INIT_1D => X"D7BD7400000000000000000000000000000000000000000000061007FE00000F",
INIT_1E => X"A2D1574005D0428A10A2AAA8BEF552EBDFFF557BC01FF5D7BFFEBA5D55555EF5",
INIT_1F => X"AFFFFC2000AA8428AAAFFAAA8BFF00002AA10FF802ABEFA2D16AA00F7FBE8A10",
INIT_20 => X"EFFF8002010002EAAAAAAAD1555FFFFAEA8B550051401450055575FF00517DEB",
INIT_21 => X"5FF0855575455D2AA8BFFA2D1575EF5D5555545FFFBE8A00087FC20BA5D2A975",
INIT_22 => X"8A00FFAE800AA082A820005D2E974BAA2D140145A2842AA00A284021FF5D0415",
INIT_23 => X"7FFEF000017400FFD1555FF007FFFEBA55042AA00000017400FFAABFEBAFF802",
INIT_24 => X"000155F7D540000F7FBFFE105D7BE8ABAA284000105D0428BFFA2FBFDFFFA2D1",
INIT_25 => X"7BFAEBA5551501D51C5FC7E00000000000000000000000000000000000000000",
INIT_26 => X"6D16AA28EBF5EDA38AADE1543849557D492BF8E2DE00552EBFFC7552BC01D75D",
INIT_27 => X"A85400E00E38A175FDE3F5C002DAAD42DAAAF784AFA82BC042DF47E3D1F8028B",
INIT_28 => X"50021C0092490E904BAFFD550A90FFA495FC7A05B555C257AAA8B45007540000",
INIT_29 => X"02402ABD4AD1D0E175D7140B455D516A1EAB45E2A000B4748717A095F571EAA1",
INIT_2A => X"4A8BC0ABFF7D03A17D1D5147540B454AA080038E9748542AE3D0051C7B6F02DA",
INIT_2B => X"D4B8FC7BFFFD2168B68F57492F505FF5FA550490BFA482B420B8428A3DA85400",
INIT_2C => X"0000000000000000000016ABD554201543A1EDE9016D4AAB454AF400547ABFB6",
INIT_2D => X"EBDF55556BC35E7557FE8AB25D11415FD0151614000000000000000000000000",
INIT_2E => X"6CBEA41D7D3DECFAF7D43FABAAAD57DEBAAAFFD74AA04547EE18D680BE9A55D2",
INIT_2F => X"78228E5000EA422E10439C1FBCD282351BDAAF9C20AAAABCBEB1DFF803FC5959",
INIT_30 => X"284683ABBDD7DEAA100069C14B25495A00F38EBAC0E198B9760501805357547D",
INIT_31 => X"8FE6A755ED8EFEFE41B2D17EAF02552BC0545556BD61E501001DF5DD3EBA31E6",
INIT_32 => X"F922ACA8AB8283C8310FAB1588916D3861C0422C44082B52A81550A828141440",
INIT_33 => X"DBCD7D262E5AFAC4B6AADDD562AF57D7C369AF25495A23068A8301BA7FB95556",
INIT_34 => X"FE0000003FE0000003FE0000003FE0000003FE03D5789700282E9FEFB501EA5F",
INIT_35 => X"3FE0000003FE0000003FE0000003FE0000003FE0000003FE0000003FE0000003",
INIT_36 => X"00000000000000000000000000000000000000000000000000000003FE000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000020",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(0),        -- Port A data input
DOA(0)   => data_read_a_hi(0),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(0),        -- Port B data input
DOB(0)   => data_read_b_hi(0),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_1_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"212C001411984004084D000508C53810A03D1450E839B003342114428A000807",
INIT_01 => X"08000010400A0008010600000084004000400002000000000000000000140000",
INIT_02 => X"484DEBA0111800C004400D000000000028800001CC404E6008B4933336880010",
INIT_03 => X"650C00000848A0423183089008C604224200000100A200002C280810098C0001",
INIT_04 => X"00000004208B00200E010800006667BE7000102C00080000040012010000080C",
INIT_05 => X"0080000000002020600100208D04414000800000000200004800080000800200",
INIT_06 => X"0000CB008084001C481040080000006050402008080000800488000000020400",
INIT_07 => X"00C00843060C19E2300221036000004400208000400041034001042000000101",
INIT_08 => X"08000290248CC84E0801318000C45555087C60C182B1592FE26AD7B7F7A01118",
INIT_09 => X"D8000AA220480040050080085200001161020001202100008008611687A28000",
INIT_0A => X"2640440000000080081040000040208300041000008004104006840000B80004",
INIT_0B => X"78051112A80000840200202112800001010828008000000105400020082800A8",
INIT_0C => X"2358323483234832358323583234832340190AC191A52801000C1002020883C2",
INIT_0D => X"4417882F82C00181707044212080300001002102010244800400C80C80323183",
INIT_0E => X"0B92C000000000400001004200004010200810040802040080200284401C1C11",
INIT_0F => X"00000043C2016000000F03C00280030000000F03C00280030000004860C60C0C",
INIT_10 => X"03800000049C0000000F03C00280030000000F03C002800321080000BC2380C2",
INIT_11 => X"00007861E0180000002A9001A00000007C4380E00000001E002300000008D187",
INIT_12 => X"4C0C81200009480010280340000008082430A07C80600C000000900861001108",
INIT_13 => X"34400241186100004A500007B00FC000000000E4A402C001208C308000268800",
INIT_14 => X"C0001E0181C0C200000025A400A200812A4070380000000B2500098190240001",
INIT_15 => X"04A0002410A170300C4A800800000020E22400A200096828F008000000AA9002",
INIT_16 => X"0200820040041002000010080014000000002340002004118010C22861400008",
INIT_17 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_18 => X"0080200802008020080200802008020080200802008020080200802008020080",
INIT_19 => X"0A04000000000000000000020080200802008020080200802008020080200802",
INIT_1A => X"8AB2048634B03249249604C061028A46BABEFC54A08170062002340C7452B500",
INIT_1B => X"DD6EB75BADD6EAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA8A28A28A28A2",
INIT_1C => X"A5D2E974BA5D2E974BA5D2E974BA5D2E974BA5D2E974BA5D2E974BA5D6EB75BA",
INIT_1D => X"AAAAAA00000000000000000000000000000000000000000000181FFFFF00000B",
INIT_1E => X"5D7BE8ABA5D557DFEFFFD17FEBA00042AAAAFFFFFFE00FF843DF45FFAE95555A",
INIT_1F => X"F552A800AA5555575FFA2AE820BAFFAEBFF555500155EF552E975FFF7D168BEF",
INIT_20 => X"00A2FBEAABA5D55420AA00002AA00AAFBE8B55A280175455D002AA00A2AABDFE",
INIT_21 => X"5FFAA802AAAAFFAA801EF00517FFFFF7D56ABEF0004155550004154105D556AA",
INIT_22 => X"75FF08557DEBAA2FBEAAAA552E955EF5D0415410A2AE97545A2AE954BAF7FBD7",
INIT_23 => X"7DF55A2AEBDEAAFFFFC20AAFFFFFFFFFAAD5555FFFFAEAAB55A2D168B555D555",
INIT_24 => X"0000BAFFFBE8A00087FC20BA5D2A975EF5D0002010552E820AAFFD57FF55F7D1",
INIT_25 => X"8A38F45F7AA9217FA380AD400000000000000000000000000000000000000000",
INIT_26 => X"52E975EFFFDF68BFF557BEAA925551785D7BFD5EFE3F08002FA92EBA5FDE28FF",
INIT_27 => X"41017DE92BF8E3AA824924870BF5551555C7A28A821EFE3AABAE38005B575D75",
INIT_28 => X"8005A1041055716DB7DB6FBEFEA81C55D0A0516802AA28BEF5EDB7DAA8A15438",
INIT_29 => X"EF1C043FE28E3FBD55FFAADE2DAAAE3A5C51C71C042DF45A3D1D00281E8A1056",
INIT_2A => X"B45B47F6FB55A95555E90F78E17F52FEF5EDA82FD249057F080417492AAAFC7F",
INIT_2B => X"8AAAA95B7AF45FF8F7DFEDFFAFF8E005FAE92A3AE3DBFF57FA2DF555D257AAA8",
INIT_2C => X"000000000000000000000A8F571EAA150021C0092490E905FFFD0550BD75C5FF",
INIT_2D => X"43DE00A2C57DE08FFAAA8B55F7EE801F7F2849EE000000000000000000000000",
INIT_2E => X"AE29F067155543A15D2E955EFFFFBEABEF557FEAA10595169BED83D1EBCA8000",
INIT_2F => X"FD57DEEAAA15976EB0444BFEB086808A8E3082C954BA5D7DD6145AAAA821A6AA",
INIT_30 => X"FFD55D6107782001FF0812000A255D57FFBEF3B97EEAB2C40217B9778428ABAF",
INIT_31 => X"F003F17418AEE817B540D11CA80BAAFA825EFAABEBCA18FE803755D08079EB47",
INIT_32 => X"EBA2D757547D7862AF57ABFFCABE5553FD5FBEFE86353EFFFD03FE027500035F",
INIT_33 => X"1F70C6AA04537957D6FB4807FFFB45F7EFFDA58FF2AA88A0F3C5014018AC28BD",
INIT_34 => X"00000000000000000000000000000000000000B2DD7DEAA100069C14B25495A0",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000020",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(1),        -- Port A data input
DOA(0)   => data_read_a_hi(1),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(1),        -- Port B data input
DOB(0)   => data_read_b_hi(1),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_2_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10E44660018259B2843913100062C98004802322D3E030235201006009B2812",
INIT_01 => X"8005A188084900481C8024A542400340404000720885800802000906E4910204",
INIT_02 => X"5C010802020408040C640850AA055254090541A111240A104A0000000908B510",
INIT_03 => X"0C1101108800004481060A001204102802156020218808002440850008C80550",
INIT_04 => X"8840C08022050400482812C21C0804040968987810688899444090C10A124A69",
INIT_05 => X"4885109105400029210000010340086856B141212252142242A068A080106372",
INIT_06 => X"0082006020044004C240108005540A400440880000908281302852A6710AA420",
INIT_07 => X"08040860400008C022402502100AA00004404B5075460111044014002AAA2100",
INIT_08 => X"382A885244145048C860214020040505487C0800049000004220000110820204",
INIT_09 => X"88582833A24105145404D4694E710A832488C000002205C23600408C872A2A12",
INIT_0A => X"A211100D0828800A022025A81AE3048228002A7080012082C15C859D5073D520",
INIT_0B => X"3E00659A308809540009202A5820068019108A88B1D007285082002B10416820",
INIT_0C => X"1A0021A5021A1021A5021A1021A4021A0010C2010D010887470912171342A683",
INIT_0D => X"89180010084038220410042B2000715A0400200080623400380886086021A002",
INIT_0E => X"40000554015500481000300000C4480810000002040000000913000004C18402",
INIT_0F => X"00000001440002C052000400028000154052000400028000200501CCD28D206A",
INIT_10 => X"00000000048015405200040002800012C05200040002800014E0000100002000",
INIT_11 => X"00010008000000000002A0000D80060100004000000000180000294010240020",
INIT_12 => X"1011000000090000A310000881080102000A0000400000000000900002000684",
INIT_13 => X"204E008240000000483250000800000000000004E00007004120000000240A60",
INIT_14 => X"254000806000000000000560000942004110000000000000254C020220000001",
INIT_15 => X"00108840600002080200000000000020806000093000040000000000000B8000",
INIT_16 => X"008022200100000020A89068084D402120AAC005C00000000000000005408140",
INIT_17 => X"0802008020080601806018060180200802008020080601806018060180200802",
INIT_18 => X"8040080000800008000180401804018040080000800008060180601806018020",
INIT_19 => X"A2852F81F81F83F03F03F0018040180401804008000080000800018040180401",
INIT_1A => X"04609D21808205965965D64CC5B60040138D70C030B54284722B291C50C7D100",
INIT_1B => X"4A25128944A25041041041041041041041041041041041041041041041041041",
INIT_1C => X"44A25128944A25128944A25128944A25128944A25128944A25128944A2512894",
INIT_1D => X"055400000000000000000000000000000000000000000000001E1007FFE3F009",
INIT_1E => X"FF843DF45FFAEBDF55082A82155082AAAA10F7FFEAB455500175FF5D2A800100",
INIT_1F => X"F082ABDF455D7BD5545F7D5574BAFFD16AAAAA28428ABA000428AAA5D7FD7400",
INIT_20 => X"455D7BEAABA5D2A97545552E975FFFFD168AAA5D7BE8BFF5D557FFEFFFD16ABE",
INIT_21 => X"5555555555FFA2AE820BAFFFFEAABA5555554BA5D0417545F7D56AAAAAAFBEAB",
INIT_22 => X"AA00AAAEBDFFF08042AABA087BD54BA08043DEAAFF843FF5508517FF55552A95",
INIT_23 => X"82010AAD1401FF002EBFF45A2FBFDFEF00042AA00AAFBEAB5500003FF5500002",
INIT_24 => X"0000BA0004155550004154105D556AA00A2FBEAABA085542145082A800BA002A",
INIT_25 => X"00155FF552A87410007145400000000000000000000000000000000000000000",
INIT_26 => X"8002FABA4171D5400FF8A38F45F7AABA57D0000855FD1C2AAFA00EBA5E8B7D55",
INIT_27 => X"555178FD7BFD5FDFFA0020BFF78417BD5545F7F1554AAF7D16DABABFF57DE920",
INIT_28 => X"DFFDF6DAAAAAF1EFB6D417BEFA901C2E97F40552E975EFEBDF68ABA557BEAA92",
INIT_29 => X"7DA3FBD21C7492E9256D555B555C7A2ABC20AAE3AABAE38005B574AA49041756",
INIT_2A => X"B7D1E803AF6D400028E02AB8A3A012540E2AABABC75D043A00003FE10E3802DB",
INIT_2B => X"8B7D0AAA800AA147085000FFDA001C7B47BFABC7BFFF7AB4714042AA38BEF5ED",
INIT_2C => X"000000000000000000000821E8A10568005A1041055716DA38B6FBEFFEF1C0EB",
INIT_2D => X"EBDE00AAC16ABEF5500155EF552A954000855544000000000000000000000000",
INIT_2E => X"D57DE0AFAD1EBEB400043DEAA085555400FFAAAAB55F7AEA8BF77004147EF5D2",
INIT_2F => X"AFBEABAF557FEA8515951E8B4D83D1EBDFF082CBDFEF005756145FFD5574AAF7",
INIT_30 => X"5951550100004155EFF7FFFDE08AA557FFFF083FFCEB95104210405D2E955EFA",
INIT_31 => X"A002A3FE18AE803CBE7A3C014351082E951FF5D7FD6145AAAA820A2AAAD29E00",
INIT_32 => X"45550028ABAFFD17FFED01001FFEF5542ABEB2AA848AAA2552EA8ABA7551400A",
INIT_33 => X"EBAF3F95EEE95C00B7CF12AAA800BA551417105FFFFC21555556EAB4CD6D5EAD",
INIT_34 => X"00000000000000000000000000000000000000187782001FF0812000A255D57F",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000040",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(2),        -- Port A data input
DOA(0)   => data_read_a_hi(2),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(2),        -- Port B data input
DOB(0)   => data_read_b_hi(2),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_3_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"210C00A20020000108430020001600B815602110494074133520400E02B92206",
INIT_01 => X"A00C9BC048800168240442C99E004B61404040028804A0080A000D16A0990A08",
INIT_02 => X"4809A902031800444445089866E331352180D468B8200E600C0081110B80ACD0",
INIT_03 => X"6D0A60100C000142B1A30A040AC68428320006010A80881068A80D401C846330",
INIT_04 => X"482218076809C03B24841CD92CDD5A440209127847294C042640102107102D04",
INIT_05 => X"0583180353202129000104E40B04644B32A86D24014A0D204063297092000E34",
INIT_06 => X"0120D000808040181B5000A014CC662814442808805A52C03068280004629414",
INIT_07 => X"00444841428409C038B02523041994001C644C82732001190000B400E6640901",
INIT_08 => X"E8E64010248C4A5AA040308000440005487C285284B1D00BC22AC005B2820318",
INIT_09 => X"A8D588362040534C3B0E80A9DB742641620AC281826816925040408483008A10",
INIT_0A => X"040450A1439800840C32264119D004860110104004010001E732C0DF80F3B174",
INIT_0B => X"7C8575909088A4D010202422520090840B4028209AC1111954DA902230010002",
INIT_0C => X"032920329203692036920329203392036C900BC9019528100A0D30024BC8A283",
INIT_0D => X"446A101C05C0088A42D001032000333931001902010234888C68804808A03692",
INIT_0E => X"8601CCCC8B33004C0001004240140018380818040A0706009000028000903401",
INIT_0F => X"00000120000006000000000020004011000000000020004010072CC92416414C",
INIT_10 => X"0000001002001400000000002000401380000000002000401070000000000000",
INIT_11 => X"00000000000000000110000001A0000000000000000005002000244000000000",
INIT_12 => X"00000000010402049910000011000500000000000000000008000020000002C0",
INIT_13 => X"805500000000000820133000000000000000810000000C000000000004100B20",
INIT_14 => X"0530000000000000000180000011060000000000000001040154000000000020",
INIT_15 => X"0000820062000000000000000000040100000010700000000000000002400000",
INIT_16 => X"0680C2A05104100280A8D06C004044230B998021002004000001011000380000",
INIT_17 => X"280C0280C0280803808038080380803808038080380C0280C0280C0280C0280C",
INIT_18 => X"00C0280E0200C0280E030080380A030080380A030080380C0280C0280C0280C0",
INIT_19 => X"8A145D54AAB556AA9556AA830080380A030080380A030080380A0200C0280E02",
INIT_1A => X"04A20E858000049249240540430303C0C78C706428A141046016224C58629502",
INIT_1B => X"EA753A9D4EA75249249249249249249249249249249249249249041041041041",
INIT_1C => X"46A351A8D46A351A8D46A351A8D46A351A8D46A351A8D46A351A8D46A753A9D4",
INIT_1D => X"A8400000000000000000000000000000000000000000000000001007FEB6FECD",
INIT_1E => X"5500175FF5D2AA8A10005540155087BEABFF552ABDF45A2D16AAAAF7D540000A",
INIT_1F => X"000556AB55552ABDE00AAD140010F7D17FF45A2AA82155082AAAA10F7FFEAB45",
INIT_20 => X"55557FEAA10007FEAABA000428AAA557FD7400FF843DE00FFAEBFF55082A8201",
INIT_21 => X"A105D7BD5545F7D5574BAFF802AA00A2D168ABA085568BEFFFAE820000855421",
INIT_22 => X"FFEFF7D56ABEF557BD74BAFF8402145A2AEBFFEF552EAAABA5D0028BEF082AA8",
INIT_23 => X"3DEAAAAAA95410F7803FFFF55556AAAA552A975FFFFD16AAAA5D7BC01EF5D557",
INIT_24 => X"0000105D0417545F7D56AAAAAAFBEAB455D7BEAABA5D2A974005D55574005504",
INIT_25 => X"DF6FABAFFD547010AA8407400000000000000000000000000000000000000000",
INIT_26 => X"C2AAFA28EBF5E8B7D5500155FF552AAF0100071455451C75EABC74174BAF55B6",
INIT_27 => X"F7AABAF7D00009543D1C556AB6D4124BAE10BED542010FFD57AF55AAF5D756D1",
INIT_28 => X"FEBA0870281C5F4716D5D7FEDA3A0955FF48208002FABA4171D5400FF8A38F45",
INIT_29 => X"BA15203FFFF002AAFA384171D5545F7D0154AAF7D16DABABFF57DE92005F6ABF",
INIT_2A => X"ABA417BC01D7555178FD7BFD5FDF571575D24BA438E021D5B6A4BAFFF5D2EB8E",
INIT_2B => X"FE005D5B52428410E3AE92E3A490410EB843ABD71551FFE02552A975FFEBDF68",
INIT_2C => X"0000000000000000000003849041756DFFDF6DAAAAAF1EFB6D417BEFBD71C24B",
INIT_2D => X"56AB45081028B55FFFFFFEBAFFD557400A280144000000000000000000000000",
INIT_2E => X"D56ABF5AAD15455F5D2EBDEAAA2D16ABEF5500175EF552ABDE000855545455D5",
INIT_2F => X"85555400FFAAAAB14F7AE28BF77004146BA557DEABEF00002BE10FFD540000FF",
INIT_30 => X"F2D1EAEBA007FEABEFAA84174BA557FD55EF5D3BFEEB35055DEE1000043DEAA0",
INIT_31 => X"5FFAA28BF7592EABE0A0804ABFFB082EBDEAA005556145FFD5574AAF7D47DE0A",
INIT_32 => X"105D2E955EFAAFBE8AAA547FE21550853E8B4FABD5EBFF75D55420AA82AA8015",
INIT_33 => X"FFF087FFCEF90104B780A557FC20AA082AAAE10AA8000000A2AC2ABFD2151EB8",
INIT_34 => X"00000000000000000000000000000000000000AA0004155EFF7FFFDE08AA557F",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000020",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(3),        -- Port A data input
DOA(0)   => data_read_a_hi(3),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(3),        -- Port B data input
DOB(0)   => data_read_b_hi(3),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_4_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10804002061080A284201081034809800A00230350007833422C82904204006",
INIT_01 => X"204398001038084C0420050E12100368403008418984014902030906A0910204",
INIT_02 => X"480108A000000000446118E01E80F00A41043118680402000800000009882390",
INIT_03 => X"065140108C0000400026480000009120270072E03000000030808840888100F0",
INIT_04 => X"9100EB826A155C1AF0B81C160033B9440222BA281AE0D8B8E02010E81C22E821",
INIT_05 => X"5C0F20B36F08010924C084C501441C4CF21C48B133483C8042EAE1E0101074C4",
INIT_06 => X"010290102005118043508020543C1E480002820085D9C0C70000F2AA375A6071",
INIT_07 => X"00000860008008D200102502000786000C00C8025C00091B0400B00061F84020",
INIT_08 => X"991E02100C84C0480020010000004404087C8010009800004022800110000000",
INIT_09 => X"B83D6A2620418F7CF8084082425D01D123C2C040816A00708840408483000011",
INIT_0A => X"BB1B585C1304E002000064010E4007F7210010500400400800F0CC249C1401C1",
INIT_0B => X"7A04331814080458100134201A2086441B50A088078106C14540906D004068A0",
INIT_0C => X"186921829218692182921829218692182090D3490C352296CC60B11357088682",
INIT_0D => X"411050002500A9200A8014010001370F03080980912204883C28864860A18A92",
INIT_0E => X"C40903C1430F20025040102200441A040906008300418050501341208002A005",
INIT_0F => X"0000012004000BC01200000020004008C012000000200040000721CD86146108",
INIT_10 => X"0000001002000A40120000002000400DC01200000020004004D4400000000000",
INIT_11 => X"40000000000000000110200007600401000000000000050020005D4010040000",
INIT_12 => X"1010000001040004A3B000018008850200080000000000000800002002000650",
INIT_13 => X"80360082000000082034300000000000000081004000170041000000041005E0",
INIT_14 => X"2B200080400000000001804000192000401000000000010400F8020200000020",
INIT_15 => X"00114A00200002080000000000000401004000085C0000000000000002410000",
INIT_16 => X"459040281181004A8088986D045C24436C7840A6180300082001211304208140",
INIT_17 => X"1106409004110240904411024090040106419004010640900411064090440102",
INIT_18 => X"9024010041104409024190240104411004190240906411024190440102419004",
INIT_19 => X"021074B261934D964C3269C09064110040104409064190240104401004190640",
INIT_1A => X"8A74C1323433345145130282E6228A063807E05000143842130115063450454A",
INIT_1B => X"8D46A351A8D46AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA8A28A28A28A2",
INIT_1C => X"A0D068341A0D068341A0D068341A0D068341A0D068341A0D068341A0D46A351A",
INIT_1D => X"50015400000000000000000000000000000000000000000000001007FEA73FC1",
INIT_1E => X"A2D16AAAAF7D568A00AA8400000AAFFC21FFF7D542000FFAE821FF552EAAA105",
INIT_1F => X"0AAAE820BA550015400087FD74BAFFD540000F7D155555087BEABFF552ABDF45",
INIT_20 => X"AAF78015545FFD555555082AAAA10F7FFEAB455500175FF5D2AAAA1000554000",
INIT_21 => X"B45552ABDE00AAD140010F7D17FF45A2FBC2000A2FFC21555551554005D2EA8A",
INIT_22 => X"FF55082E82145A280001EFF78402145A2AE801555D2E95555552E9741000556A",
INIT_23 => X"7DF45557BD5410F7D555545F7AA97410000428AAA557FD5400FF843DE00FFAEB",
INIT_24 => X"0000AA085568BEFFFAE82000085542155557FEAA10007FEABEFAAD1400AA5D51",
INIT_25 => X"AA801EF4920AFA10490A17000000000000000000000000000000000000000000",
INIT_26 => X"C75EABEF4124BAF55B6DF6FABAFFD56F010AA8407428A2F1C01FFF7D142028EB",
INIT_27 => X"552AAFA10007155428A2AE850925D0010400087FD24AAE3DF47010E38E051451",
INIT_28 => X"55D51524004920ADA82EB8A12555EBFB4717D1C2AAFA28EBF5E8B7D5500155FF",
INIT_29 => X"55492A850381C5F6AB6D4124BAE10BED542010FFD57AF55AAF5D7410A2FBC015",
INIT_2A => X"400FF8A38E00F7AABAF7D0000955FDB684051D7F7840517DA2A4871554124925",
INIT_2B => X"75EFBED5400825D557FF55007BD7410EBDB5017DE38E8708008002FAAA4171D5",
INIT_2C => X"00000000000000000000082005F6ABFFEBA0870281C5F4716D5D7FEDB7D0955D",
INIT_2D => X"1401FFFFD5420BAA2AA821FF08043DE10002A964000000000000000000000000",
INIT_2E => X"FBD7410A2AE965555D556ABEF080028B55FFFFFDEBAFFD57FE00A280144BAAAD",
INIT_2F => X"2D16ABEF5500175EF552ABDE000855544AAAA82174105D0402000087FC00BAA2",
INIT_30 => X"AAD154400AAFBC015555554001008003FE00AAEA81154AAFFD65FF5D2EBDEAAA",
INIT_31 => X"FA2AA155550004021E5582A964BE557FEABEF00002BE10FFD540000FFD56ABF5",
INIT_32 => X"1000043DEAA085555400FFAAAAA10F7AC28BF558001454DF78017555F780175E",
INIT_33 => X"5EF5D7BFEEF35055487EFF7D1400105D517FF55087FD7410A2FBC01E7F2AE966",
INIT_34 => X"0000000000000000000000000000000000000010007FEABEFAA84174BA557FD5",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000040",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(4),        -- Port A data input
DOA(0)   => data_read_a_hi(4),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(4),        -- Port B data input
DOB(0)   => data_read_b_hi(4),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_5_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50DB4A0791B1B4B694369283C81F9996A091832102004AB37B20E07C0C1E006",
INIT_01 => X"285FBC448000804C446A00000034824841280A00084000C8C212892EE2953235",
INIT_02 => X"C809AD5CB118E640A4D118FC011FF0002080000082C8C66609DB7DDDCB1F2036",
INIT_03 => X"250907263A4C90D210A35C82484285720B20648A88800000B8E0F850A8C4500E",
INIT_04 => X"4005122126899100064D20001044429C78243A2C0436C887198AB916E0551A24",
INIT_05 => X"A370C14CA0E900004048002389CFE2F20F7D7A314CB5C20AE51437E044948912",
INIT_06 => X"90184D150505A1D84B7E2A285401412870B20A51842404C44437118630839B88",
INIT_07 => X"E640A94D1AB469D6300E2FFFAA7F8A4D23248130E259C903FBC403A9601A62E8",
INIT_08 => X"0A7E3016250D49CA3F83108186400000EBFD235488B9749BC1AAF325B35CB118",
INIT_09 => X"9B020B7E6AE46082032004904200C03DBC3BCA4860270BFA829968040B0800AC",
INIT_0A => X"22181A2B9203642840124098516CE0C3D825124111A79F802800F20DB4D6DA34",
INIT_0B => X"6824911331CA84D346A964F0125CD7AB1938A00AEFDD567DE480116848C9426A",
INIT_0C => X"01AD7016D701ED7012D701ED7016D701AAB8096B80F5A21828041846620F5AB8",
INIT_0D => X"847B053F48A8308A644A412BCA8470FF0209019081C706EABDAAC0DC0AF012D7",
INIT_0E => X"2194FFC044FF84B08FC862A2CD8F0A89014080A2425422151870500544991292",
INIT_0F => X"038ABBCBC7C7802F86FF87C002F87F002F86FF87C002F87F2000804821021004",
INIT_10 => X"0380230F2FFC002F94FF87C002F87F002F94FF87C002F87F2201BFFEBC2BA0C2",
INIT_11 => X"BFFE7C69E01804E1E7EABE3F000FF97D7C4BC0E008C7C3FE58FC029FEF5CD9A7",
INIT_12 => X"EC9C8120C4DFC802808B2EB22E777ADDE6F8A47CC0600C2683E0FFAAE3F1F001",
INIT_13 => X"FC14DFC5186104C6FE5037FFF00FC0000FC0FEE487A7066FA38C3082637F83BD",
INIT_14 => X"072FFF41C1C0C2038A7CED87A7D109FBBA5070380131CBFB2477BF919024189B",
INIT_15 => X"9F46DFBEB1B7F0380C4A80092E0FC1FDE607A7C077FFE828F0080AE1DFAA1E9F",
INIT_16 => X"5594254A10A03446128898494C09402081F83200A9442217159880640942320E",
INIT_17 => X"1940509465014251140519445094251142511445094451942511425014451940",
INIT_18 => X"9405094450944511425114650146501425194450944509405194250146501405",
INIT_19 => X"0A983124B2DA6924965B4D509445094051940501465014251142501465094451",
INIT_1A => X"BE5FDFF3F7F773CF3CF7D79FA8F5BB4E7F7B9DB7FF3A7E0FF4807F1B6DB7ED43",
INIT_1B => X"F77BBDDEEF77BBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEF",
INIT_1C => X"EF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEE",
INIT_1D => X"FFBFFE00000000000000000000000000000000000000000000001007FE1BFB5E",
INIT_1E => X"FFAE821FF552E820105500155555D2AA8A00AA843FFFFF78002155AAAE974AAF",
INIT_1F => X"0FFAE80000AAAE974BAFFAEAAB45AAAEBDEAAA2FFEAA00AAFFC21FFF7D542000",
INIT_20 => X"000055574BA557FFFF55087BEABFF552ABDF45A2D16AAAAF7D56AA00AA840000",
INIT_21 => X"0BA550015400087FD74BAFFD540000F780155555D7BE8B45085168BFFA2D17FE",
INIT_22 => X"AA10005140145FFFBC01EFAAFFD75FF002E97555A2AABDEAAAAAAAAA00AAAE82",
INIT_23 => X"174BA5D043FF45AAAA974AAF7AEBFF55082AAAA10F7FFEAB455500175FF5D2AA",
INIT_24 => X"000000A2FFC21555551554005D2EA8AAAF78015545FFD555410552EA8BEFAA84",
INIT_25 => X"8E0217DBEA4954AAE3FBFDE00000000000000000000000000000000000000000",
INIT_26 => X"2F1C01D7F7D142028EBAA801EF492087A10490A171455D2EADA28B6803FFFFFF",
INIT_27 => X"FFD56FA10AA8417428E3AE87010A2A4974AAE3AEAFB6DAAA4BDEAAA2F1EDA28A",
INIT_28 => X"D14516DBD7BEDB7DE381451554AA497FFFF451C75EABEF4124BAF55B6DF6FABA",
INIT_29 => X"AAAAA0AFA28A2A4850925D0010400087FD24AAE3DF47010E38E0516D5D7BE8B6",
INIT_2A => X"B7D5500155FF552AAFA10007155545F7F1C21D7AAF1D55FF082A9057DA2AABDE",
INIT_2B => X"70384124ADBFFBE84174AA55043FF6DBEAE950AAEB8ABDF7D1C2AAFA28EBF5E8",
INIT_2C => X"00000000000000000000010A2FBC01555D51524004920ADA82EB8A12410EBFB4",
INIT_2D => X"EBFEBAF7843DFEFF7AE801EFF780174AAAAFBFEE000000000000000000000000",
INIT_2E => X"803FEBAAAD17CEAAAAD140155FFD5420BAA2AA821FF080415410002A96555552",
INIT_2F => X"80028B55FFFFFDEBAFFD57FE00A280144AAA2AA97400A280174AAA2AEBDFEFA2",
INIT_30 => X"A2AE965FF557FE8BFF55557FF55FFFBFFEAA5D51554AA087BFEF555D556ABEF0",
INIT_31 => X"F0004821FFAAAEBDEAAAA843CEAAAA80174105D0402000087FC00BAA2FBD7410",
INIT_32 => X"FF5D2EBDEAAA2D16ABEF5500175EF552ABDE00005554545F7D140145A2D5555F",
INIT_33 => X"E00AAAA81114AAFFD64BA00043FFFFFF80174AA55043DFFFFFAE974BAA2AEBEF",
INIT_34 => X"0000000000000000000000000000000000000000AAFBC015555554001008003F",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000180",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(5),        -- Port A data input
DOA(0)   => data_read_a_hi(5),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(5),        -- Port B data input
DOB(0)   => data_read_b_hi(5),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_6_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10804B0061A010A2840012C030028180004003220200403302301C0381A0086",
INIT_01 => X"870041CA3839684D18A160000C52424841000000090800090210010008110204",
INIT_02 => X"080108200C1000004464480400C0080100000000010432400800800009882050",
INIT_03 => X"040001008C2340D0840208624210002182800584488000103080010E08C10000",
INIT_04 => X"00101611A029B08410044800000000040088102A440814040400900500001800",
INIT_05 => X"02800000400C820934E4A0002900404400820004000A00824004085011200A00",
INIT_06 => X"2210001A12100830434040870BFE004044420322C00812900308010000829400",
INIT_07 => X"00000860400108C22000A103090074120044800040001103005180911FE0C134",
INIT_08 => X"FD01C0120484C0580020C10000000000087C0800209100004228000110000C10",
INIT_09 => X"88FC08362240404100228080D200DFC1610200E40AA050000040D0C463008083",
INIT_0A => X"29561B22D77C720D2522400000400882091210008440005F8BF4C00002900004",
INIT_0B => X"7E25D11A200024541100342A5A2886285502A880C00107FD355E022005026BCA",
INIT_0C => X"D8282D8A82D8A82D8682D8682D8E82D8A016C1416C15A01D68209A127208A6B1",
INIT_0D => X"807888180A80910A1460150900013400410CB5C9D96236883460B60B602D8282",
INIT_0E => X"0062003C10002442006429124290034E85A742D1A368D0DA2004696884851806",
INIT_0F => X"000000157000604050000000028000D04050000000028000CE80004C00000000",
INIT_10 => X"000000000483D04042000000028000D04042000000028000C508000100000000",
INIT_11 => X"000100000000000000078000A40006000000000000000019A003080010200000",
INIT_12 => X"1001000000093490308001408000000200020000000000000000900518000508",
INIT_13 => X"23490002400000004993C000080000000000001FC000C8804020000000246800",
INIT_14 => X"C05000802000000000001740002256004100000000000000FD00000220000001",
INIT_15 => X"00A000404A000200020000000000002099C000330000040000000000001F0000",
INIT_16 => X"68DA308D09D0804880089A49461032040C07C1440C8190800020530865400540",
INIT_17 => X"9DA7695A1685A369DA7685A168DA369DA5685A168DA7695A5685A368DA7695A5",
INIT_18 => X"5A168DA7695A168DA1695A769DA1685A3695A569DA3685A169DA769DA1685A16",
INIT_19 => X"00046638C31C71C718638E68DA7695A568DA3685A769DA5685A368DA569DA368",
INIT_1A => X"8E76DDB3B7B377DF7DF7D7CEE7F78BCE7F8FF0F4FA957FC7F37F3F5F7CF7F108",
INIT_1B => X"7F3F9FCFE7F3F8E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E3",
INIT_1C => X"E7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE",
INIT_1D => X"AAABFE00000000000000000000000000000000000000000000181007FFDE534F",
INIT_1E => X"F78002155AAAE974AAFFFBFFE10F7FBE8BEF552E95555552EAABEF082E975EFA",
INIT_1F => X"0A2AAAAA10087FC01EF552EAAB45F7AE821550851555555D2AA8A00AA843FFFF",
INIT_20 => X"EFA2AEBDFFF552AAAA00AAFFC21FFF7D542000FFAE821FF552E8001055001541",
INIT_21 => X"000AAAE974BAFFAEAAB45AAAEBDEAAA2FFEAB45552E800AA555568A105D002AB",
INIT_22 => X"AA00AA8400000007BC21FFAA803FFEF5551420105D5568B45FF8400000FFAE80",
INIT_23 => X"C2155007FC20BAA2D5575FF087FFFF55087BEABFF552ABDF45A2D16AAAAF7D56",
INIT_24 => X"0001555D7BE8B45085168BFFA2D17FE000055574BA557FFFE10F7AAA8A00F7FB",
INIT_25 => X"24ADBD70820975FFA2A4BFE00000000000000000000000000000000000000000",
INIT_26 => X"D2EADA28B6803FFFFFF8E0217DBEA4954AAE3FBFDE38F7FFEABFF412A9056D49",
INIT_27 => X"492087010490A07038B6A0AFA38007BC51EF4920AFB55EBA4851450855555455",
INIT_28 => X"2555F68A3855002FBC7BEA4BFFFF492EADA28A2F1C01D7F7D142028EBAA801EF",
INIT_29 => X"45E38A07028E3AE87010A2A4974AAE3AEAFB6DAAA4BDEAAA2F1EDB55492A8508",
INIT_2A => X"F55B6DF6FABAFFD56FA10AA84174381C7FC01C7B68E3DFC75555400105D516DB",
INIT_2B => X"FE38F7A0AFA38E3FFC21450071C2092A2D5571FF0851FDF451C75EABEF4124BA",
INIT_2C => X"0000000000000000000016D5D7BE8B6D14516DBD7BEDB7DE381451554AA497FF",
INIT_2D => X"BEABEF002E801EF00003FF550800155FFA2803CE000000000000000000000000",
INIT_2E => X"8417555085154555552EBFEBAF7843DFEFF7AE801EFF780174AAAAFBFEEAAF7F",
INIT_2F => X"FD5420BAA2AA821FF080415410002A964AAFF803DEAA087FD55FF00043DF45A2",
INIT_30 => X"AAD17CF55002E95410557BEAABA55043DF55F7803FFEF002ABEEAAAAD140155F",
INIT_31 => X"55D51420105D517DF55AAAA964AAA2AA97400A280174AAA2AEBDFEFA2803FEBA",
INIT_32 => X"555D556ABEF080028B55FFFFFDEBAFFD57FE00A280144BA5D7FC2155FFAABDF4",
INIT_33 => X"EAA5D51554AA087BFEEAAF7803DEAAAAFBC0155085540000A2D5575FF08517CF",
INIT_34 => X"00000000000000000000000000000000000001FF557FE8BFF55557FF55FFFBFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000120",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(6),        -- Port A data input
DOA(0)   => data_read_a_hi(6),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(6),        -- Port B data input
DOB(0)   => data_read_b_hi(6),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_7_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10804B00482010A2842012C024500188000003000000003302300C018180002",
INIT_01 => X"0200084020084048040080000201024040000000080000080200010008110204",
INIT_02 => X"4801082248100000444008000080000041000000002222400800000009008010",
INIT_03 => X"0401008108A1444000020A400000002902006400088000003080040408C10000",
INIT_04 => X"0000100022418000000C80C00400000400201839040000050001140400201820",
INIT_05 => X"02000000400041092C80C0214144004400000000000800045004000020220800",
INIT_06 => X"0000300000000830435150020003004060000000080800801100000030829001",
INIT_07 => X"00000840000008C02000A503010002928040800062481919047140D40008C000",
INIT_08 => X"0A0002120484C0580850810000000000487C000000910000402A800110024810",
INIT_09 => X"8802083624504000022680A1DA20800164000400112284000004D404022A8800",
INIT_0A => X"30014050280040180020400011640CC72E029000084800503004C40100D21024",
INIT_0B => X"3801078228010454210028240082200081140800900220000000002011440009",
INIT_0C => X"40022400224002240822408224082240C1120211202008900800100242428280",
INIT_0D => X"807802988294900A00451109006230006E000800001280110050902901240022",
INIT_0E => X"0042C000C0002000000020020490000400020001020080401010813094801146",
INIT_0F => X"807144102420700052000003C00780B00052000003C007808450484C00000000",
INIT_10 => X"2C0E00E0D003300052000003C00780B00052000003C00780890800010000130C",
INIT_11 => X"000100000661801E18042100E000060100000B03803838012403800010240000",
INIT_12 => X"10111848322020512000414400000002000A1001058300C0741C005412080908",
INIT_13 => X"029F008240864231013BF00008000C3C003F00184040EF8041204321188053E0",
INIT_14 => X"F770008060130C8071821040403F5600411004C2600E3400C27C020223090644",
INIT_15 => X"00B8CA406A0002C812240B0201F038021140403F740004010472041E20110100",
INIT_16 => X"0080228011010042802890484040000008004945000100008844430060198941",
INIT_17 => X"0000000000000600802008020000400000000000080200802008000000000000",
INIT_18 => X"8020100000000008020080000000000020080200000000040080200802008060",
INIT_19 => X"0A14584104000208208000018020080200000010020080200800010000080200",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000442",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"82AAAA00000000000000000000000000000000000000000000001007FEBC3240",
INIT_1E => X"552EAABEF082E975EFAAAABFFEF002ABDF555D5157555F7FBC00AAAAD5400BA0",
INIT_1F => X"AAAAABDF55FFFBFDF55555568ABAAAD5401FF5D2AAAA10F7FBE8BEF552E95555",
INIT_20 => X"005D55554105D51401555D2AA8A00AA843FFFFF78002155AAAE974AAFFFBFFEA",
INIT_21 => X"A10087FC01EF552EAAB45F7AE821550851554AAF7FBFFEAA007BFFFEFF7D5400",
INIT_22 => X"00105500155EF5D2EBFF450000020AA5D7BC0000F7D555545A28000010A2AAAA",
INIT_23 => X"A8A10FFD568ABAA2D56AAAAF7AABFE00AAFFC21FFF7D542000FFAE821FF552E8",
INIT_24 => X"000145552E800AA555568A105D002ABEFA2AEBDFFF552AAAABAA2AE95555FFAA",
INIT_25 => X"F5C20BAAAD5420821C2EAAA00000000000000000000000000000000000000000",
INIT_26 => X"7FFEABFF412A9056D4924ADBD70820975FFA2A4BFFFF1C2EB8F45555550545E3",
INIT_27 => X"BEA4954AAE3FBFDE82B6AEBAF55E3FFFAF55555F6FA92BED5421C75D20AAA38F",
INIT_28 => X"20075FDFD7F7D5400385D51504385D55401455D2EADA28B6803FFFFFF8E0217D",
INIT_29 => X"7DB68E02038B6A0AFA38007BC51EF4920AFB55EBA485145085555492F7F5FFE9",
INIT_2A => X"028EBAA801EF492087010490A071EF4920B8F45140E07082417BC2000EBD5505",
INIT_2B => X"DA92A2A09257DE3A4AAA10F7D16FAAABED56AE82F780BAE28A2F1C01D7F7D142",
INIT_2C => X"00000000000000000000155492A85082555F68A3855002FBC7BEA4BFFFF492EA",
INIT_2D => X"EAAB455D5142155AAD1400AAA2D1420005D2EA9A000000000000000000000000",
INIT_2E => X"D1421555D042BAAAF7FBEABEF002E801EF00003FF550800155FFA2803CFFF552",
INIT_2F => X"7843DFEFF7AE801EFF780174AAAAFBFEE00F7AAAAB55AAFBEAB555D7BFDE00F7",
INIT_30 => X"085154400FFD17FE1000517FF55FFD5420BA5D55400BA555543155552EBFEBAF",
INIT_31 => X"0087BC0000A2D5421EFF7AE810AAFF803DEAA087FD55FF00043DF45A28417555",
INIT_32 => X"AAAAD140155FFD5420BAA2AA821FF080415410002A965FF080428B45552A9540",
INIT_33 => X"F55F7803FFEF002ABEE00A280001FFA28028A00FFD17DEAAF7D56AA10FF842BA",
INIT_34 => X"0000000000000000000000000000000000000155002E95410557BEAABA55043D",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"FFFFFFFE00000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000000000000000000001F",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(7),        -- Port A data input
DOA(0)   => data_read_a_hi(7),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(7),        -- Port B data input
DOB(0)   => data_read_b_hi(7),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_8_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10004B00000400E2840012C0000001800000070000000033022000000000082",
INIT_01 => X"000009C0183808481C0160000E02424040000000180800080200010048110204",
INIT_02 => X"080108000090000004400C000080000051000000000002400800000009000010",
INIT_03 => X"0000000004300840000200000000000002800504488000103080880008800000",
INIT_04 => X"00009410A028A084000440C00400000400001032040800150400008500221800",
INIT_05 => X"4280008040048A09302420202804400400800010200A00000204080011014A00",
INIT_06 => X"2B02000A32114192434010001FFC004240428122000800000008012000821400",
INIT_07 => X"00000840000008402001A50200000630404080006248381B000080837FF88114",
INIT_08 => X"0A000210040440480000090000000000087C0000009100000002000110000090",
INIT_09 => X"08020A322000400102260021DA2080114502002409A04400004282C4E1228800",
INIT_0A => X"904A4522920052012120400011641C4601005000041100002004800100C21024",
INIT_0B => X"78051792A8000454104020001280008845022000900000010444000000020009",
INIT_0C => X"000000000000000000000000000000000800040000452A9008001002424A8002",
INIT_0D => X"807880508202100A1000810B2020340041248548490004800400000008000800",
INIT_0E => X"20020000C000044214240932000001428CA14650A128508A2004284024840022",
INIT_0F => X"80000000001020404000783FC0000010404000783FC000000880084C01041008",
INIT_10 => X"FC7E0000000010404000783FC0000010404000783FC000000500000103D45F3D",
INIT_11 => X"000103961FE78000000000402400020003B43F1F800000002201080000202658",
INIT_12 => X"01617CD8000000803000804080000020090659833F9F03C00000000000040500",
INIT_13 => X"00400018639EC000000000000FE03FFC00000000400840000C31CF6000000800",
INIT_14 => X"4000001E2A3F3D80000000400802000401AA8FC7E00000000100002C2F5B0000",
INIT_15 => X"4020000104480DC372B47F060000000000400802000017570FF6000000010020",
INIT_16 => X"28CA30051851A0C0002890484600320408004444048090800022130864000540",
INIT_17 => X"84A1284A1284A328CA328CA328CA328CA328CA3284A1284A1284A1284A1284A1",
INIT_18 => X"CA328CA328CA3284A1284A1284A1284A328CA328CA328CA3284A1284A1284A12",
INIT_19 => X"080440000000000000000028CA328CA328CA328CA1284A1284A1284A128CA328",
INIT_1A => X"9EDFC8F33637D6CB6CB2900DA6128A0A543EBC57A10A244257C5051E75D64108",
INIT_1B => X"1F0F87C3E1F0F9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7",
INIT_1C => X"E1F4F87D3E1F4F87D3E1F4F87D3E1F4F87D3E1F4F87D3E1F4F87D3E1F0F87C3E",
INIT_1D => X"02ABFE00000000000000000000000000000000000000000000001007FE8A8913",
INIT_1E => X"F7FBC00AAAAD5400BA082AAAA10000000010F7D5421EF007BC01FF5D7FFFE100",
INIT_1F => X"A5551554AAFF80021EF002A820BAFF8428A00A2AAAABEF002ABDF555D5157555",
INIT_20 => X"EFFFFFEAB55002ABFE10F7FBE8BEF552E95555552EAABEF082E975EFAAAABFEA",
INIT_21 => X"F55FFFBFDF55555568ABAAAD5401FF5D2AAAB55FFD1400AA5D7FC01EFA2FFE8B",
INIT_22 => X"74AAFFFBFFEAA08001555555516ABEFA280020AA5D043DF55557BEAAAAAAAABD",
INIT_23 => X"2AB55005140145AAFFE8AAAF7D1401555D2AA8A00AA843FFFFF78002155AAAE9",
INIT_24 => X"0000AAF7FBFFEAA007BFFFEFF7D5400005D55554105D51400005551421EF0804",
INIT_25 => X"7FC21EF5D75FFE10142EBAE00000000000000000000000000000000000000000",
INIT_26 => X"C2EB8F45555550545E3F5C20BAAAD5420821C2EAAA101C0005000E3D1401D71C",
INIT_27 => X"0820975FFA2A4BFE925D51554AAE384001FF142E800AAFF802AA28AAAEAFBFF1",
INIT_28 => X"2557BC21D7BEF5EDBC7FFF1EFB6D1420BAE38F7FFEABFF412A9056D4924ADBD7",
INIT_29 => X"55417BEDA82B6AEBAF55E3FFFAF55555F6FA92BED5421C75D20AAB45F7D14709",
INIT_2A => X"FFFFF8E0217DBEA4954AAE3FBFDEAA1C001056D415F6ABEFA2840208249043AF",
INIT_2B => X"00385D51401EF00002FB45085F4016DAAF1EDAAAFFFB401455D2EADA28B6803F",
INIT_2C => X"00000000000000000000092F7F5FFE920075FDFD7F7D5400385D51504385D554",
INIT_2D => X"417410AAD540155557FC01EF5D557DE105D2AA8A000000000000000000000000",
INIT_2E => X"842AABAA2AEBDFFF552EAAB455D5142155AAD1400AAA2D1420005D2EA9A105D0",
INIT_2F => X"02E801EF00003FF550800155FFA2803CE105D55574BAA280021EF5D2E820BAF7",
INIT_30 => X"5D042BB45FFD157410557FC0155F7D57FF55F7D57FFEF550028AAAF7FBEABEF0",
INIT_31 => X"FAA8000000080428B55087FFFE00F7AAAAB55AAFBEAB555D7BFDE00F7D142155",
INIT_32 => X"55552EBFEBAF7843DFEFF7AE801EFF780174AAAAFBFEEBA5D04021EF087BE8BF",
INIT_33 => X"0BA5D55400BA5555430BA5555421EF00043FF45007BC21FFA2D57FEBAF7FBC21",
INIT_34 => X"0000000000000000000000000000000000000000FFD17FE1000517FF55FFD542",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000080",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(8),        -- Port A data input
DOA(0)   => data_read_a_hi(8),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(8),        -- Port B data input
DOB(0)   => data_read_b_hi(8),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_9_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10004B00018000A2840012C0000281800000030000000033022000000000006",
INIT_01 => X"000008000000004C0020000000100268413C0A61590001D90213C10008110204",
INIT_02 => X"680108200010000054400C000080000041000000010002400800800009082011",
INIT_03 => X"0004000000002040000200100000000042800584488000103081880008800000",
INIT_04 => X"00001610A00AB084000400C00600000400001030040010050020020400001880",
INIT_05 => X"02000200400C8A09206420000C00410400000000000800000804000000000800",
INIT_06 => X"2A10201A12104010435051000801004040000322980800000080000100821000",
INIT_07 => X"000018400000086020002502000002000040800062C8081B0000008000088034",
INIT_08 => X"0A000610040440480000010000000000187C0000009100002046000110000010",
INIT_09 => X"4802082220084001002400214A2080014400006400A000000000015421800800",
INIT_0A => X"4B505008020032032320400011640447000010040000000020048409004A9020",
INIT_0B => X"280005922000045400002001100000000D0000008000000041C48000002003EA",
INIT_0C => X"2080020000208002000020800200002080010000104100800000100202420142",
INIT_0D => X"C06800100240180A0010010921003400432C8CC8D80044000000080080020800",
INIT_0E => X"2002C000C000240004641932041403428DA146D0A36850DA3200684004800403",
INIT_0F => X"0000000144002000420000000280001000420000000280000000084C01041008",
INIT_10 => X"0000000004801000500000000280001000500000000280001100000100000000",
INIT_11 => X"00010000000000000002A0002000020100000000000000182001000000240000",
INIT_12 => X"00110000000900003000004000000000000A0000000000000000900002000100",
INIT_13 => X"205D0080400000004803F0000800000000000004E0004E800120000000240BA0",
INIT_14 => X"4770000060000000000005600013560001100000000000002574020020000001",
INIT_15 => X"0020CA406A0000080200000000000020806000137400040000000000000B8000",
INIT_16 => X"68DA320D19D1A0CA8028984D46543600080040440C8090800000130061400140",
INIT_17 => X"8DA368DA368DA1685A1685A1685A1685A1685A1685A1685A1685A1685A1685A1",
INIT_18 => X"5A1685A1685A1685A1685A1685A1685A368DA368DA368DA368DA368DA368DA36",
INIT_19 => X"801010000000000000000068DA368DA368DA368DA368DA368DA368DA3685A168",
INIT_1A => X"344A2D840100E492082405548817344CCCF48DE68A89004F98614C5C38E2540A",
INIT_1B => X"1A0D068341A0D14514514514514514514514514514514514514534D34D34D34D",
INIT_1C => X"41A4D268341A0D069349A0D069349A0D068341A4D268341A4D268341A0D06834",
INIT_1D => X"FD557400000000000000000000000000000000000000000000001FFFFE2CAD83",
INIT_1E => X"007BC01FF5D7FFFE10002ABFF55F7D168A00552E95555007BFFF55087BE8BFFF",
INIT_1F => X"0F7FBC0145F7AE801EFF7FBFFF455D7BC0155F7D557410000000010F7D5421EF",
INIT_20 => X"00AA803FFEF5D55421EF002ABDF555D5157555F7FBC00AAAAD5400BA082AAAA1",
INIT_21 => X"4AAFF80021EF002A820BAFF8428A00A2AAAAAAAF7D17DE00FFFBD5555A2AABDE",
INIT_22 => X"75EFAAAABFFEF002A954BA5551421EF552E954105D00021455555420AA555155",
INIT_23 => X"575EFA2FFD75455D7BE8A005D5557410F7FBE8BEF552E95555552EAABEF082E9",
INIT_24 => X"000155FFD1400AA5D7FC01EFA2FFE8BEFFFFFEAB55002ABFE10080028BFFF7D5",
INIT_25 => X"71F8F7D147BEFBEFEBD152400000000000000000000000000000000000000000",
INIT_26 => X"C0005000E3D1401D71C7FC21EF5D75FFE10142EBAF7DE3D16DA0041209056D1C",
INIT_27 => X"AAD5420821C2EAAA10E3FFC0145F7A0801FFEBFBF8F6D417BC716DEBD1524101",
INIT_28 => X"8F7F5D0545B6AAB8E38B68A3AFFF5551471FF1C2EB8F45555550545E3F5C20BA",
INIT_29 => X"455D5B470925D51554AAE384001FF142E800AAFF802AA28AAAEAFABAE3D17DE2",
INIT_2A => X"56D4924ADBD70820975FFA2A4BFFFF082E974BA4155401C7552097428550E021",
INIT_2B => X"AE0008002ABFFF7DB505FFAAFBD7555417FEFA00495B52438F7FFEABFF412A90",
INIT_2C => X"00000000000000000000145F7D147092557BC21D7BEF5EDBC7FFF1EFB6D1420B",
INIT_2D => X"17DE100804001EF55516ABFF557BFDFEFA2D5400000000000000000000000000",
INIT_2E => X"7FD55FFA2D5400105D0417410AAD540155557FC01EF5D557DE105D2AA8BEFAAD",
INIT_2F => X"D5142155AAD1400AAA2D1420005D2EA9A00A2FBC0145FF84001EFA2FFEABFF00",
INIT_30 => X"A2AEBDEAAAAD17DEBAFFD142155FFAAAAABAFFAAAABFF5551555FF552EAAB455",
INIT_31 => X"55D00154AA552E801455D7BD54105D55574BAA280021EF5D2E820BAF7842AABA",
INIT_32 => X"AAF7FBEABEF002E801EF00003FF550800155FFA2803CFFF002E954BA00514015",
INIT_33 => X"F55F7D57FFEF550028A10000428BEFF7FFC01FFA2FFD5545007BFDE10087FC00",
INIT_34 => X"0000000000000000000000000000000000000145FFD157410557FC0155F7D57F",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000100",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(9),        -- Port A data input
DOA(0)   => data_read_a_hi(9),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(9),        -- Port B data input
DOB(0)   => data_read_b_hi(9),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_10_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10040B0001824802840102C00002C18000202300500030B3132000400992006",
INIT_01 => X"A140098018300848180060000C00424040000000080000080200010008110200",
INIT_02 => X"0801080200100000046558040080000041000000002402400800000009008010",
INIT_03 => X"00010100840000D0842242024210810802006400088000003080054288C10000",
INIT_04 => X"0000100022008000000C08C00C00000400A83A3044200C840000800400101820",
INIT_05 => X"0200000040000000248080210044000402000025000800020004207010100800",
INIT_06 => X"0800200000004010435040A14001004844000800CC0812541020008230829000",
INIT_07 => X"00000860408108502000250208000600004080006248081B0040808000088000",
INIT_08 => X"0A000210040440480060010000000000087C0810209900000002000110020010",
INIT_09 => X"08020A2222004040000484214A2080110108C280022210020240000401080880",
INIT_0A => X"000000000200000C042040001164044609101000840000802004800100421020",
INIT_0B => X"782415809888A45010082408028010080110280800001001051A124810410800",
INIT_0C => X"0089000890000900009000890008900008800048004420910800120242488000",
INIT_0D => X"4110000006008820020010010001300040000100014000808C48004008800090",
INIT_0E => X"2002000040002000040020020490080400020001000482000010012080008005",
INIT_0F => X"0000010140002040100000000280401040100000000280400000204801041008",
INIT_10 => X"0000000006801040020000000280401040020000000280400500000000000000",
INIT_11 => X"0000000000000000010280002400040000000000000001182001080010000000",
INIT_12 => X"10000000000D0000808000408000000200000000000000000000902000000500",
INIT_13 => X"A000000200000000681000000000000000008004A00040004000000000340000",
INIT_14 => X"4000008000000000000085200002000040000000000001002400000200000001",
INIT_15 => X"00200000000002000000000000000021802000020000000000000000020A8000",
INIT_16 => X"040006E00100044200289048085D402008000040000100000000020065400000",
INIT_17 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_18 => X"0000000000000000000000000000000020080200802008020080200802008020",
INIT_19 => X"8290100000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"8A355950666151451453D5006F86890A940FE0D39712614261D20E4355520542",
INIT_1B => X"6532994CA65328A28A28A28A28A28A28A28A28A28A28A28A28A28A28A28A28A2",
INIT_1C => X"AE532994CA6532995CAE572B94CA6532994CA6572B95CAE532994CA6532994CA",
INIT_1D => X"FFBC2000000000000000000000000000000000000000000000001007FECF31DC",
INIT_1E => X"007BFFF55087BE8BFFFFD557400FF842ABEFA2AAA8B5500003DF55F7D568AAAF",
INIT_1F => X"008556ABFFA2D16AB550000021FFF7D17FFEF08042AB55F7D168A00552E95555",
INIT_20 => X"55A2D557400557BC2010000000010F7D5421EF007BC01FF5D7FFFE10002ABFE0",
INIT_21 => X"145F7AE801EFF7FBFFF455D7BC0155F7D557545FFAE820AA007BFDFEF55003FF",
INIT_22 => X"00BA082AAAA00FFAE820AAAAAABDFEFF78028BEF005140145A2842AA10F7FBC0",
INIT_23 => X"6AB55A2D157400552EBFFEF5D7BD75EF002ABDF555D5157555F7FBC00AAAAD54",
INIT_24 => X"0000AAF7D17DE00FFFBD5555A2AABDE00AA803FFEF5D55420BA08557FEBAAAD5",
INIT_25 => X"0E3AF55F7DF68ABAE3F1C0000000000000000000000000000000000000000000",
INIT_26 => X"3D16DA0041209056D1C71F8F7D147BEFBEFEBD152400F7842FBD7B6AAAAB551C",
INIT_27 => X"5D75FFE10142EBAE0008556FBD7B6DB6AB7D1C0A001D7FFD178FC71C0E28B7DE",
INIT_28 => X"2147BFAFEF49043AF45A2DF504285D71C00101C0005000E3D1401D71C7FC21EF",
INIT_29 => X"7DA28428A10E3FFC0145F7A0801FFEBFBF8F6D417BC716DEBD15256DF7AA8209",
INIT_2A => X"545E3F5C20BAAAD5420821C2EAAA00E3AA82092A2AABAFD7EB8A2ABC70855401",
INIT_2B => X"70821C557AE92A2DF6AB7DA2DF50410412ABDFC75D7BD55FF1C2EB8F45555550",
INIT_2C => X"000000000000000000000BAE3D17DE28F7F5D0545B6AAB8E38B68A3AFFF55514",
INIT_2D => X"03DF45FFAEA8B555D2EAAB45F7FBE8ABAAAD5400000000000000000000000000",
INIT_2E => X"D168B55552AA8BEFAAD17DE100804001EF55516ABFF557BFDFEFA2D540010FF8",
INIT_2F => X"AD540155557FC01EF5D557DE105D2AA8A0008557FF45FFFFE8BEF5D2E80155FF",
INIT_30 => X"A2D5401FFF7AA800105D7FE8BEF08002AB45AAFFC00AA5D51400105D0417410A",
INIT_31 => X"5AAAEAAB450055421FFAA8428A00A2FBC0145FF84001EFA2FFEABFF007FD55FF",
INIT_32 => X"FF552EAAB455D5142155AAD1400AAA2D1420005D2EA9A10A2AA82010AAAEAAB5",
INIT_33 => X"ABAFFAAAABFF555155400555568A10AAFBEABEFA2FFC0010082ABFF55557BD55",
INIT_34 => X"00000000000000000000000000000000000000AAAAD17DEBAFFD142155FFAAAA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"FFFFFFFE00000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000000000000000000011F",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(10),        -- Port A data input
DOA(0)   => data_read_a_hi(10),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(10),        -- Port B data input
DOB(0)   => data_read_b_hi(10),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_11_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10180B05A0010402840602C2D001019000000300000000330A20080EC180002",
INIT_01 => X"AB400986B830284D1820E0000C36424840000000080000088200080802512220",
INIT_02 => X"8801081438106400A4F55800008000004100000040CCE24208005000C9060032",
INIT_03 => X"000406A492E6E440842254D002108153432004800880000030C0315688C00006",
INIT_04 => X"00001201200090001205400000000094108C322644240C840008030440111800",
INIT_05 => X"222000444008010028404002A002009402400025080880000C04223000170900",
INIT_06 => X"01080C1020002810436532AB4003004864200A00540816544522008200821100",
INIT_07 => X"6400E96C488108502001295BA100022E4340800062D82819435143F20008C0A0",
INIT_08 => X"0A0012160585C1D809A3810000000000C8FD0B1420992419034A0221116C3810",
INIT_09 => X"4902083E2CB0400002020480C2008009000ACEC06B25500202988C84C0220028",
INIT_0A => X"004040000203600E06204000116C14474A36500499C49C802004C00800088000",
INIT_0B => X"6804110230CBA4576708201C0212100B492A2008000A1001C49A9348498B0808",
INIT_0C => X"410E5418E5410E5418E5418E5410E5418B2A0872A08428010000120202085000",
INIT_0D => X"41110244066C0820221480010AA7300042080980919580808C9A5002880A18E5",
INIT_0E => X"2022C000C0002020094030220C960A0409020481024482501A00401410088521",
INIT_0F => X"836090540355D86C046619A54052A5B86A046619694063168280004801041008",
INIT_10 => X"A2C60289802AB86A046619A54052A5B86C04661969406316AC018B0E2936DA02",
INIT_11 => X"CB0E1076D4A200B2AC611A3D0405886C6EB211550815A8A2686EC81E2A48B68A",
INIT_12 => X"8CE0C5E8F650E48000892B37885620C1E1A06D7016A90A4626D82B10F1B1FC09",
INIT_13 => X"4E02144D335546F28724001B030A56140A184483000C410A2699A2E32AC9C041",
INIT_14 => X"E8018A0A01B2990242E278056AAA203920E0BAE2012C08281808319C186F1E16",
INIT_15 => X"44F9051C049B18A12CB481042AD140C227002A0A02066954E7540CCDB58415AA",
INIT_16 => X"409024681181044080809A490C0964200800200108010003A02272400C19B80D",
INIT_17 => X"0902409024090240902409024090240902409024090240902409024090240902",
INIT_18 => X"1004010040100401004010040100401024090240902409024090240902409024",
INIT_19 => X"0284000000000000000000401004010040100401004010040100401004010040",
INIT_1A => X"20A069105251C0000001541148062608804180C0B10A04CA0900474210420140",
INIT_1B => X"0000000000000000000000000000000000000000000000000000208208208208",
INIT_1C => X"0000000000004020000000000000000000100800000000000000000000000000",
INIT_1D => X"00015400000000000000000000000000000000000000000000001007FE0FC1C0",
INIT_1E => X"00003DF55F7D568AAAFFFBC2010557BEAA10AAFBE8A00557BFFFEF007BC21550",
INIT_1F => X"55D7FE8BFF5D7FD540055003FFEFFFD142145000000000FF842ABEFA2AAA8B55",
INIT_20 => X"45557FC2010557FFDF55F7D168A00552E95555007BFFF55087BE8BFFFFD55754",
INIT_21 => X"BFFA2D16AB550000021FFF7D17FFEF08042AB55A2AAAAB4508517FE00557BC01",
INIT_22 => X"FE10002ABFE00AAFFE8AAAFF8402000550002145085555400F7FFE8A0008556A",
INIT_23 => X"3FEBA002A975EFF7D17DFFFAA8000010000000010F7D5421EF007BC01FF5D7FF",
INIT_24 => X"000145FFAE820AA007BFDFEF55003FF55A2D557400557BC2145A2D1421450804",
INIT_25 => X"7BF8FEF1C7FC516D080E15400000000000000000000000000000000000000000",
INIT_26 => X"7842FBD7B6AAAAB551C0E3AF55F7DF68ABAE3F1C00005D7BEDA00B6F1EFA2855",
INIT_27 => X"147BEFBEFEBD15257D5D7FEFBD7417BD5438550038FC7FFDF4216D080E07000F",
INIT_28 => X"514517FE105575C216D5571C50104171FDF7DE3D16DA0041209056D1C71F8F7D",
INIT_29 => X"00FFF1EFA0008556FBD7B6DB6AB7D1C0A001D7FFD178FC71C0E28B6DA2AEADB4",
INIT_2A => X"1D71C7FC21EF5D75FFE10142EBAE10A2FBEFA92F78A05028550E001451455524",
INIT_2B => X"016DB6D54514500003FEBA1420905FFFFDF78FC7BE84050101C0005000E3D140",
INIT_2C => X"0000000000000000000016DF7AA82092147BFAFEF49043AF45A2DF504285D71C",
INIT_2D => X"FFDE00F7D17FEBA557BEABEF557BD55EF082A974000000000000000000000000",
INIT_2E => X"FBC01FF082A97410FF803DF45FFAEA8B555D2EAAB45F7FBE8ABAAAD5400105D7",
INIT_2F => X"804001EF55516ABFF557BFDFEFA2D5401FF5D7FFDF55007BD74BA5D042AB45F7",
INIT_30 => X"552AA8BEFAAAABFF5555517FE005555401FF55515541000517FFEFAAD17DE100",
INIT_31 => X"A5D2A801455D5140000FFD57FE0008557FF45FFFFE8BEF5D2E80155FFD168B55",
INIT_32 => X"105D0417410AAD540155557FC01EF5D557DE105D2AA8A10AAFBFFE00F7AA974B",
INIT_33 => X"B45AAFFC00AA5D51401FFFFD15555500003FEBA5D04001EFFFFFE8B55FF84174",
INIT_34 => X"00000000000000000000000000000000000001FFF7AA800105D7FE8BEF08002A",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000100",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(11),        -- Port A data input
DOA(0)   => data_read_a_hi(11),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(11),        -- Port B data input
DOB(0)   => data_read_b_hi(11),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_12_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50080B01BC002006940202C0DE041196A83183000000023322287E0FC000006",
INIT_01 => X"0E000C048000C048400380000007026040000000080000088200002802153231",
INIT_02 => X"2809AD0E7D180040945008040090000061800000C0E2F66009DA3D11CB148015",
INIT_03 => X"210D050012F6F8D2108216E24842005B8A20640008800000B8E0141C28851006",
INIT_04 => X"0080100022408000060DE0000066630C70241827041000040800820480001AA4",
INIT_05 => X"0240000C400000003C808003E0C8001401000000040900020904004000070800",
INIT_06 => X"00006C00000008784B4D210E0001006050800000100804005784000130821200",
INIT_07 => X"A64019490A044860300FA3968B20028FC06080106249F819A19143FE00088200",
INIT_08 => X"0A002610240D494A0753D1810240000038FC234480B1709A81C67325B31EFD18",
INIT_09 => X"090209222EB84000010000104200802180210C007827C000009DBE040800008C",
INIT_0A => X"0000000002000030003040081164FC469227D20019F413503004900020000200",
INIT_0B => X"28200100004304D267C06CC500566003C13E0000000460000000000010CE0000",
INIT_0C => X"E1865E1065E1065E1865E1065E1065E1832F0C32F08000000004100202015940",
INIT_0D => X"0403CFE7E03E8080382FD0018FE670004000000000D5C023009278B7835E1065",
INIT_0E => X"01EA0000440000800A0040028108000000000000000000000A74812DF00E0BF4",
INIT_0F => X"8362F658A7E5F82CD23B6B0E403DBBE82C563B6A4E403DBB88C0E04820020004",
INIT_10 => X"BE5403AB992F282C563B6B0E403DBBE82CD23B6A4E403DBBB1084E4B25AC48DF",
INIT_11 => X"0E4B1D32BAB504BB74AD3F3FE04A8E0D0C319A7988B6F0C75CFD801A962454CF",
INIT_12 => X"18D994B866E2E8C3808B6B63040328E7A33AF99B0AC20DE634D06C437BF85100",
INIT_13 => X"5F6214CA5991C6A7177402C49CA354D808D358A927EAD10A652CC8E3538BEC41",
INIT_14 => X"E80083C3EAEB2003695430A7CDAA289553922990C11A4E494988231B32570CDC",
INIT_15 => X"D5B304AD05A946D81616970A225658940BA7CDAA0A312666BD600E5550B49F36",
INIT_16 => X"00000100000010420000904C0040000008003B81000000021CFEE02E2803BC0F",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"8020080200802008020080200802008000000000000000000000000000000000",
INIT_19 => X"0210100000000000000000008020080200802008020080200802008020080200",
INIT_1A => X"24481C040000B5145144015085C1B946088881360A95118D90215C090CB05442",
INIT_1B => X"32190C8643219041041041041041041041041041041041041041249249249249",
INIT_1C => X"4B2592C964B2592C964B2592C964B2592C964B2592C964B2592C964B2190C864",
INIT_1D => X"AFBC2000000000000000000000000000000000000000000000001007FEF001D6",
INIT_1E => X"557BFFFEF007BC2155000015555087FC0010AAFBFFE100004020BAAAFFD5400A",
INIT_1F => X"5AA8400000A2AABFF45550400000AAFBFFFEF550000010557BEAA10AAFBE8A00",
INIT_20 => X"10555155555FF8017400FF842ABEFA2AAA8B5500003DF55F7D568AAAFFFBC215",
INIT_21 => X"BFF5D7FD540055003FFEFFFD142145000000145A2AA821EFFFFFD7410007FC00",
INIT_22 => X"8BFFFFD5574000051420BA557FC2145557FC20AAA2D57DEBAA2FBD55455D7FE8",
INIT_23 => X"AAA00550415410AAFBFFFEF55042AB55F7D168A00552E95555007BFFF55087BE",
INIT_24 => X"000155A2AAAAB4508517FE00557BC0145557FC2010557FFDE10AA8400000082E",
INIT_25 => X"0A02092B6F5D2438A2FBC2000000000000000000000000000000000000000000",
INIT_26 => X"D7BEDA00B6F1EFA28557BF8FEF1C7FC516D080E1557D0075C7028B6F1FAE0000",
INIT_27 => X"F7DF68ABAE3F1C017DAA8E07028B6A0BFF6D490E00000BEF5FAFEF4904070005",
INIT_28 => X"FE3FBD0438007FC00385D555556DEB8410400F7842FBD7B6AAAAB551C0E3AF55",
INIT_29 => X"BAA2FBD557D5D7FEFBD7417BD5438550038FC7FFDF4216D080E0716DAAA0851F",
INIT_2A => X"56D1C71F8F7D147BEFBEFEBD152400005F450BA417BC51454971C20AAB6D17DE",
INIT_2B => X"DE10BE8E070280020AAA28410410400BEFBFAFEF49042AB7DE3D16DA00412090",
INIT_2C => X"0000000000000000000016DA2AEADB4514517FE105575C216D5571C50104171F",
INIT_2D => X"5574BAFFD568A10002A82000FFD5400AAA2FBC00000000000000000000000000",
INIT_2E => X"D568BEF0004174105D7FFDE00F7D17FEBA557BEABEF557BD55EF082A975EF005",
INIT_2F => X"FAEA8B555D2EAAB45F7FBE8ABAAAD5401EFA2AA974BAF7803FFFF002A82000FF",
INIT_30 => X"082A975EFA280175FFAAFFC00BA087FC20AA5D55555FFA28000010FF803DF45F",
INIT_31 => X"50851420BAFFD57DEAAAAFBD75FF5D7FFDF55007BD74BA5D042AB45F7FBC01FF",
INIT_32 => X"EFAAD17DE100804001EF55516ABFF557BFDFEFA2D540010007FD74AA007BD754",
INIT_33 => X"1FF55515541000517FE10F7AA954AA080428AAA000002010FFFFE8BEF080428B",
INIT_34 => X"00000000000000000000000000000000000001EFAAAABFF5555517FE00555540",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"FFFFFFFE00000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000000000000000000001F",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(12),        -- Port A data input
DOA(0)   => data_read_a_hi(12),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(12),        -- Port B data input
DOB(0)   => data_read_b_hi(12),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_13_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10110A0441812402840402822007818000E00700000000330A3000000008042",
INIT_01 => X"A1400984B830C848180260000C0042404001000008220008A200100802110200",
INIT_02 => X"88010C02801040002475580400800000410000000064024608134C0CC9018034",
INIT_03 => X"00010100926220D084234212421085084300648A0880000630C0654288C10000",
INIT_04 => X"0004122122029100100C00001200009C40A83A2044360C84190BAC04E0101820",
INIT_05 => X"027000004009050064C8C00104C10184034010250089C00EB004327064B60900",
INIT_06 => X"910000152500A050436A10A14003004864B00A50440812541027008230821380",
INIT_07 => X"640029605091495020002B8AAA000AF003408000E258081963F100C00008C2E8",
INIT_08 => X"0A001210040441C802E0010084000000AAFC09142899000B20020001105A0010",
INIT_09 => X"4A02096A62004000020004104200802D9838C2C80322100202020194408000A0",
INIT_0A => X"000000000203240E46204000516C04468C101005800E95802004B20020080200",
INIT_0B => X"28200101118BA4510008241D005211000910000A000A1000809A93485D610000",
INIT_0C => X"0000000800000000000000800000000000000400000000000000100202055040",
INIT_0D => X"0100000006C0802042501001C8017000C2190890904000508908000000000800",
INIT_0E => X"0010C000C00081A08BC832A209AB0A85094284A14254A2551010513080109404",
INIT_0F => X"01293C0F5012906A96DCD13042CE0C206E92DCD07042CE0C40D0204800000000",
INIT_10 => X"71CA2168ACB0E06E92DCD13042CE0C206A96DCD07042CE0C4408632C39530BA9",
INIT_11 => X"632C30D522CE80239CC2806AC44E954939AB299E000738F88296CA13B444CA42",
INIT_12 => X"D5306028F01990C080808494A64708B265CC4052B0F30302E060965EA0058408",
INIT_13 => X"28A2CA9722094650CCAC0629112BA89C04A228568547B1654B9104A32865145C",
INIT_14 => X"B80D4D8D48CB54012290470562EC29E44050B1DC60132282B68B9AA60C051E03",
INIT_15 => X"0A5C11B9008FE2FA38F87804251CB0FAD40562EC0B426149D17E0044B10A158B",
INIT_16 => X"5094246A10A10441010090480C0964201800044109012001A000726E45428000",
INIT_17 => X"0942509425094250942509425094250942509425094250942509425094250942",
INIT_18 => X"9425094250942509425094250942509425094250942509425094250942509425",
INIT_19 => X"02A8000000000000000000509425094250942509425094250942509425094250",
INIT_1A => X"BAFFD7F7F7F775555557DF9FE0FFBBEEFF3F7DF7FF3E7E2FF0087B9F7DF7E245",
INIT_1B => X"FD7EBF5FAFD7EBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAE",
INIT_1C => X"AFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FA",
INIT_1D => X"0557DE00000000000000000000000000000000000000000000001007FE0001DF",
INIT_1E => X"0004020BAAAFFD5400AAFBC2155AAAA97410FFFFEAAAAF7AA955EFF7803FF450",
INIT_1F => X"0F7AEBDE10FFFFFDEAAF7D568AAA5D002AB55005568B55087FC0010AAFBFFE10",
INIT_20 => X"FF5D04154BAAAAEAAA10557BEAA10AAFBE8A00557BFFFEF007BC215500001541",
INIT_21 => X"000A2AABFF45550400000AAFBFFFEF550000155A28415410F7AEAABFFA2D1555",
INIT_22 => X"8AAAFFFBC21555D517FF45F7AEA8BFFA2AEAAA10A280021EF5D557FF55AA8400",
INIT_23 => X"974AAF7D142145082A975FF555568A00FF842ABEFA2AAA8B5500003DF55F7D56",
INIT_24 => X"000145A2AA821EFFFFFD7410007FC0010555155555FF80174000055555EFAAAE",
INIT_25 => X"A0925C7E38E38F7D14557AE00000000000000000000000000000000000000000",
INIT_26 => X"075C7028B6F1FAE00000A02092B6F5D2438A2FBC2145B6A090428FFF5EAA92E3",
INIT_27 => X"1C7FC516D080E15438E3A4BAE00FFF5FAE92F7D16AAAA41042FB7D145568B7D0",
INIT_28 => X"8FFA4AFBFFAAD1505FF490E174AABEA0ADA005D7BEDA00B6F1EFA28557BF8FEF",
INIT_29 => X"FF555F7FF7DAA8E07028B6A0BFF6D490E00000BEF5FAFEF490407155BE8E1242",
INIT_2A => X"B551C0E3AF55F7DF68ABAE3F1C0145415B78F45FFA4AFBC7BEA4AAA10A284001",
INIT_2B => X"04380055525FFBEAE90482E3D54216D0024975FF555F68A00F7842FBD7B6AAAA",
INIT_2C => X"0000000000000000000016DAAA0851FFE3FBD0438007FC00385D555556DEB841",
INIT_2D => X"0020BAF7D16AA10A28402155A2AEA8BEF5D516AA000000000000000000000000",
INIT_2E => X"003DFEF55516ABEF0055574BAFFD568A10002A82000FFD5400AAA2FBC0145FF8",
INIT_2F => X"7D17FEBA557BEABEF557BD55EF082A974BAA28028A00F7D16AA10F7D56AABA08",
INIT_30 => X"000417545FFAA820BAFF843DFFFA2D5421FF002E954AAFF843DE105D7FFDE00F",
INIT_31 => X"5F7802AA10AA80001FF5D7FFDFEFA2AA974BAF7803FFFF002A82000FFD568BEF",
INIT_32 => X"10FF803DF45FFAEA8B555D2EAAB45F7FBE8ABAAAD540145007FE8B55FF843DF5",
INIT_33 => X"0AA5D55555FFA280000BA0855401EFF7AA82010AAD1421FF0004155FF557FEAA",
INIT_34 => X"00000000000000000000000000000000000001EFA280175FFAAFFC00BA087FC2",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"FFFFFFFE00000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000000000000000000019F",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(13),        -- Port A data input
DOA(0)   => data_read_a_hi(13),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(13),        -- Port B data input
DOB(0)   => data_read_b_hi(13),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_14_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10020A000180000284008280000281800000030000000033022000000580002",
INIT_01 => X"A140098018300848184860000C20C24040000000084000084200000000110200",
INIT_02 => X"88010C5A8010A600A4F558040080000041000000022C024008003CCCC9028030",
INIT_03 => X"000103A7A00904D0842242024210810803006480088000003081054288C10000",
INIT_04 => X"0000120122009000100C00000000000400A83A2044200C840000800400101820",
INIT_05 => X"020000004008010024C0C0010040000402000025000800020004207000100800",
INIT_06 => X"010000102000005043403AA14003004864000A00440812541020008230821000",
INIT_07 => X"2400A96850A16854200021DA2A0002000340800062C80819EBC402800008C020",
INIT_08 => X"0A0012140404414814E001000000000029FD0A10289924810182000110028010",
INIT_09 => X"080208222200400002000400420080010008C2C0032210020200008440000080",
INIT_0A => X"000000000203200E0620400011640446DA101004800005802004800000000000",
INIT_0B => X"282001001088A45000082408000010000910000800001000009A924810410000",
INIT_0C => X"0080000000000000080000000000000080000000000000000000100202000000",
INIT_0D => X"0100000004408020021010010001700042080880904000008808000000000800",
INIT_0E => X"00000000C00000000040302200800A0409020481024482501010413080008404",
INIT_0F => X"8090008142014840100002C38280000840100003838280000640204800000000",
INIT_10 => X"072C000444C00840020002C38280000840020003838280002C09D01086839746",
INIT_11 => X"D0104B01C57100440202900184414430534605E3804802180022480419183514",
INIT_12 => X"594C194000090450808802008830024F0E248C902AEF0024170CF18001003C09",
INIT_13 => X"20020E5A08E6000048200196264BCF1C030C0604800001076C04730000240049",
INIT_14 => X"2003DEDE82C78900902A0D0000080019FAAA32D9602490302409292B83280001",
INIT_15 => X"049100021171F6C34080240108AB292CA000000800AD1A19F6F000AA0C0A0000",
INIT_16 => X"4090246810810440000090480C0964200800000108010016000012004542800D",
INIT_17 => X"0902409024090240902409024090240902409024090240902409024090240902",
INIT_18 => X"9024090240902409024090240902409024090240902409024090240902409024",
INIT_19 => X"0280000000000000000000409024090240902409024090240902409024090240",
INIT_1A => X"9E7FDDF77777F3CF3CF7D54CEFD79B4E5C8FF0F7BE9D75C7F7B71F5F7DF65040",
INIT_1B => X"7F3F9FCFE7F3F9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7",
INIT_1C => X"E7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE",
INIT_1D => X"28417400000000000000000000000000000000000000000000001007FEFFFE0F",
INIT_1E => X"F7AA955EFF7803FF4500557DF45F7D16AB455D00001EFAAAAAAABA555557555A",
INIT_1F => X"555003FF450804001555D2AA8AAA002ABDE10082ABDF55AAAA97410FFFFEAAAA",
INIT_20 => X"EF5D5168A10082E80155087FC0010AAFBFFE100004020BAAAFFD5400AAFBC214",
INIT_21 => X"E10FFFFFDEAAF7D568AAA5D002AB55005568A00A2D5401455D00175FFFF84175",
INIT_22 => X"2155000015400AAD157545080402145087FD75FFF7AE82145A2D17FE10F7AEBD",
INIT_23 => X"000BAFFFBE8AAAA2FBFDE00087FD5410557BEAA10AAFBE8A00557BFFFEF007BC",
INIT_24 => X"000155A28415410F7AEAABFFA2D1555FF5D04154BAAAAEAAA005D002AB450000",
INIT_25 => X"A0AAA82555157555B68012400000000000000000000000000000000000000000",
INIT_26 => X"6A090428FFF5EAA92E3A0925C7E38E38F7D14557AF45FFDB6AB6D4100071C7B6",
INIT_27 => X"B6F5D2438A2FBC21455D0A3FF6D080407155552AAAA920020BFE10002EBAF45B",
INIT_28 => X"54100175C7E380125D7555B6DA1014248217D0075C7028B6F1FAE00000A02092",
INIT_29 => X"45AAD178E38E3A4BAE00FFF5FAE92F7D16AAAA41042FB7D145568A38AADF4014",
INIT_2A => X"A28557BF8FEF1C7FC516D080E15400A2DB5754508040716D007BD05EFEBAA821",
INIT_2B => X"DA0055002AB6D0000020BAFFF1E8ABABEF1FAE001C7FD54005D7BEDA00B6F1EF",
INIT_2C => X"00000000000000000000155BE8E12428FFA4AFBFFAAD1505FF490E174AABEA0A",
INIT_2D => X"FEABFF080015555F78028A00555155555FF84000000000000000000000000000",
INIT_2E => X"003DE10082EAAB45FF80020BAF7D16AA10A28402155A2AEA8BEF5D516AB45F7F",
INIT_2F => X"FD568A10002A82000FFD5400AAA2FBC0145552ABFFFF000417555552EA8A1000",
INIT_30 => X"55516AABAAAFFC0145000417555A280001455D7FFDE105504021EF0055574BAF",
INIT_31 => X"F007BC01FFAAAE80155AAD568ABAA28028A00F7D16AA10F7D56AABA08003DFEF",
INIT_32 => X"105D7FFDE00F7D17FEBA557BEABEF557BD55EF082A97410AAFFD55450800155F",
INIT_33 => X"1FF002E954AAFF843DE10550028BEF0004020BAF7D568AAAF7D168A105D7FD74",
INIT_34 => X"0000000000000000000000000000000000000145FFAA820BAFF843DFFFA2D542",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"FFFFFFFE00000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000000000000000000001F",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(14),        -- Port A data input
DOA(0)   => data_read_a_hi(14),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(14),        -- Port B data input
DOB(0)   => data_read_b_hi(14),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_15_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000A000000000284000280000001800020030000000033022000000180002",
INIT_01 => X"A140098018300848180060000C00424040000000080000080200000000110200",
INIT_02 => X"080108000010E60004E55800008000004100000000040240080000C009170016",
INIT_03 => X"0000000080000040842240000210810002000400888000003080014288C00000",
INIT_04 => X"0001100024A0800000440000000000040088322044200C840000011400151800",
INIT_05 => X"A200014C4000000020000000000B8094020000254C8800000514203000108800",
INIT_06 => X"000821000000A050434010A14001004844000801540812540020008600831000",
INIT_07 => X"C2000864489128502000210222000200034080006248081958C0008000088000",
INIT_08 => X"0A001214050540C800200101860000000B7C0910209900000002000110000010",
INIT_09 => X"0B0208222004400000000400420080010008C28002201002020001140800002C",
INIT_0A => X"000000000203000C04204000116404460810100080000F802004800000000000",
INIT_0B => X"280001001088A45000082008000010000100000800001000001A124800010000",
INIT_0C => X"0080000800008000000000000000000080000400004000000000100202000008",
INIT_0D => X"0100000004C00020025000018801600040000000000000008808000000000800",
INIT_0E => X"00108000C0000000000020020080080000000000000402000000000000009400",
INIT_0F => X"00000000000000404200000000000000404200000000000008C0004800000000",
INIT_10 => X"0000000000000040500000000000000040500000000000000400000100000000",
INIT_11 => X"0001000000000000000000000400020100000000000000000000080000240000",
INIT_12 => X"00110000000000C00080010180000000001A1024050000000000000000000400",
INIT_13 => X"0002008040000000002000000804002000000000000001000120000000000040",
INIT_14 => X"2000000061100280000000000008000001104422000000000008020020000000",
INIT_15 => X"00100000000009080E2E0A000000000000000008000004000000000000000000",
INIT_16 => X"0000046000000440000090480809402008000001000000000000000004188000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0280000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000040000000000040",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"8517DE00000000000000000000000000000000000000000000001007FE000000",
INIT_1E => X"AAAAAAABA555557555A284175FF000002010552A97400007BFDE10A2AA801EF0",
INIT_1F => X"F5D2AAAB45F7D17DF45087BC0155002A801FF08003DF45F7D16AB455D00001EF",
INIT_20 => X"45F7D568BEFAAD557555AAAA97410FFFFEAAAAF7AA955EFF7803FF4500557DFE",
INIT_21 => X"F450804001555D2AA8AAA002ABDE10082ABDFFFF7D17FE10002E954AAF7FBC21",
INIT_22 => X"5400AAFBC21EFA2AE95545A2D56ABFFAAD17DE10FFD1420AA007FC014555003F",
INIT_23 => X"801550055401555D00174BA002AA8B55087FC0010AAFBFFE100004020BAAAFFD",
INIT_24 => X"000000A2D5401455D00175FFFF84175EF5D5168A10082E801FFFF8428A10002A",
INIT_25 => X"71FAE00A2A0871EF145B7FE00000000000000000000000000000000000000000",
INIT_26 => X"FDB6AB6D4100071C7B6A0AAA82555157555B680125C71C0E0500049209543808",
INIT_27 => X"E38E38F7D14557AFC75524AFB45FFD178F7D1C71C2145002E801C7140A3FF45F",
INIT_28 => X"00024954AAFFFBC2145F7DB6DBEFA2D557545B6A090428FFF5EAA92E3A0925C7",
INIT_29 => X"820071C71455D0A3FF6D080407155552AAAA920020BFE10002EBAFC7FFDF7AE0",
INIT_2A => X"E00000A02092B6F5D2438A2FBC21FFBEA090545B6D568BFFAADB7AE10F7D5470",
INIT_2B => X"21FFE3802FA2808208017D1C5142155410A104AA1420AFB7D0075C7028B6F1FA",
INIT_2C => X"00000000000000000000038AADF401454100175C7E380125D7555B6DA1014248",
INIT_2D => X"E954100004174AA00516AA10AA80155EF5D7BFDE000000000000000000000000",
INIT_2E => X"2E801555D2EBDF45F7FFEABFF080015555F78028A00555155555FF8400155552",
INIT_2F => X"7D16AA10A28402155A2AEA8BEF5D516AB555D043DF55F7D56ABEF55514015508",
INIT_30 => X"082EAAB55FFFBE8A100804154AAF7FFC2145FFFFFDFEFAAD157545FF80020BAF",
INIT_31 => X"FA2FBE8A00FFD155410005555545552ABFFFF000417555552EA8A1000003DE10",
INIT_32 => X"EF0055574BAFFD568A10002A82000FFD5400AAA2FBC01FFF78400155F7D16ABE",
INIT_33 => X"1455D7FFDE105504021FFAA843DEBA0000021EF555142155002E800AA55003DF",
INIT_34 => X"00000000000000000000000000000000000000BAAAFFC0145000417555A28000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000180",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(15),        -- Port A data input
DOA(0)   => data_read_a_hi(15),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(15),        -- Port B data input
DOB(0)   => data_read_b_hi(15),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_16_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"DA22C618B1000482B688B186588884862A400438255FC38381441205BA803003",
INIT_01 => X"8645A80028404C211203A952A90341080B173340412000E1005D628000820484",
INIT_02 => X"A101A9006DC1084833011850AAC55001349B10881802821808B4110007005E11",
INIT_03 => X"010108A802BB00080080006020020001A61036202800000D2410104200404550",
INIT_04 => X"8BFA58800005C40A46240252145148B38248030356415A4E62B6FC660F287240",
INIT_05 => X"0F05EA11E570000D610000000710296E542B6E3A825C15FB30A643695BFC2D56",
INIT_06 => X"408003200040202B8584112645554B029006000140BCC0460050690A95C8383D",
INIT_07 => X"00480A2140040BE1480FA004342AA6F12000054004867415401DCDCF2AA10800",
INIT_08 => X"B32A8819064E48288012D45000005050247AA85220700009C06206C48080EDEA",
INIT_09 => X"445B2081340B6596594800400413CAC020894480000008C54C00311002000002",
INIT_0A => X"000000004B240028000342A00002FE00A3A1F06E491800AA29588181040A0020",
INIT_0B => X"2400848002912300200092BA80325A20000000000A8A5AA80018120E00066000",
INIT_0C => X"00220002200022000220002200022000210001100010000A40450100210072A0",
INIT_0D => X"002815014B90000205DA00880100095A648000000010006AC23000C7B69EC220",
INIT_0E => X"80922554515512174000000490009000000000000004010042A204A0C5817680",
INIT_0F => X"63EAA9C238B2D4C800632B266E828EE4C800632AAAB6830D0FC6B06C04102800",
INIT_10 => X"A149339E8FB964C800632B266E82B2E4C800632AAAB683310872800EDA52DA00",
INIT_11 => X"800EB090D4AAC91268FFCBE81397826C4A20D2B6C510E8624792A4A30A40839A",
INIT_12 => X"8849D5C532408DD6E004C90C06AC019D88B9795012CA96902C799912BC3C087A",
INIT_13 => X"531C74485BD42A30906057FADAA456218FD8E3ED83B60E3A242DC0F18983638E",
INIT_14 => X"A06FB555793057C444CF45C5C9E89543B8BC6E80193DC36F6C71D1093A478706",
INIT_15 => X"45DC02B331650CA8ACB4007E00D1C6A6A58395C917F7E74D936F650D69B51727",
INIT_16 => X"0000012000081500008A422150884081ACAAC0542054004FC588464050810DCD",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"147A7797E1E1A79E79E1560EEFBD11544C690DA64C1C69A9916D7E4F68A36040",
INIT_1B => X"7A7D1E9F47A7D345345345345345345345345345345345345345145145145145",
INIT_1C => X"4FA7D3E9F4FA3D1E8F47A3D1E8F47A3D1E9F4FA7D3E9F4FA7D3E9F4FA7D1E9F4",
INIT_1D => X"F8015400000000000000000000000000000000000000000000001007FE00001F",
INIT_1E => X"007BFDE10A2AA801EF08517DE10FFFFFDFEFA2D16AB55A2FFFFEAA5D7FC0000F",
INIT_1F => X"A5D2EBDFEFAAD17FFFF002EBDE000800174AA55043FFFF000002010552A97400",
INIT_20 => X"AAAA80000105D557FF45F7D16AB455D00001EFAAAAAAABA555557555A284174B",
INIT_21 => X"B45F7D17DF45087BC0155002A801FF08003DE000004154BA002A800BA087FE8A",
INIT_22 => X"FF4500557DEAAF7D57DEBA082A82010FFAE975555D7FFDEAAFF80155EF5D2AAA",
INIT_23 => X"7FFFF557FD55FF08003FE0055043FF55AAAA97410FFFFEAAAAF7AA955EFF7803",
INIT_24 => X"0001FFF7D17FE10002E954AAF7FBC2145F7D568BEFAAD557410552EA8BEFA2D5",
INIT_25 => X"FFFDEAA5571C7010FF8412400000000000000000000000000000000000000000",
INIT_26 => X"C0E050004920954380871FAE00A2A0871EF145B7FE10E3F1F8FC7AAD56DB7DB6",
INIT_27 => X"555157555B680124924124BDFEFA2D57FFC71C2EBDE280000174825D0E3FFC71",
INIT_28 => X"21424800AA007FEDAAAA284020385D5F7AF45FFDB6AB6D4100071C7B6A0AAA82",
INIT_29 => X"AAFF80175C75524AFB45FFD178F7D1C71C2145002E801C7140A3FE10080A1748",
INIT_2A => X"A92E3A0925C7E38E38F7D14557AE92EBDB78EAA1C2482010FFAE9556D557FF8E",
INIT_2B => X"7410492EADBEFA2D178FEF5575D55EF000A38E10490A3AF45B6A090428FFF5EA",
INIT_2C => X"000000000000000000001C7FFDF7AE000024954AAFFFBC2145F7DB6DBEFA2D55",
INIT_2D => X"56AB45A2D57DFFFF7FBFFEAA555555400F780000000000000000000000000000",
INIT_2E => X"0415400552ABDF55552E954100004174AA00516AA10AA80155EF5D7BFDE10A2D",
INIT_2F => X"80015555F78028A00555155555FF840000000043DFEFAAD17FF45552ABFEBA08",
INIT_30 => X"5D2EBDE10002E974005D04020BA007BFDEBAA284000BA557FE8B45F7FFEABFF0",
INIT_31 => X"0F7AE955EF5D7BE8ABAF784175555D043DF55F7D56ABEF555140155082E80155",
INIT_32 => X"45FF80020BAF7D16AA10A28402155A2AEA8BEF5D516AA00AAFBE8AAA55040000",
INIT_33 => X"145FFFFFDFEFAAD157410082ABFFEFAAD16ABFF5555575FF082AA8A00002AAAB",
INIT_34 => X"0000000000000000000000000000000000000155FFFBE8A100804154AAF7FFC2",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000080",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(16),        -- Port A data input
DOA(0)   => data_read_a_hi(16),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(16),        -- Port B data input
DOB(0)   => data_read_b_hi(16),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_17_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"5284CE4FB7BD2C8994A13392DBD02E14006B82AC7E800D44D3DD2FD5F9B961C0",
INIT_01 => X"F8ACD01F7E03FC6793F2199B39FC233C11D93AE6F3BB92B32091DBC339B24542",
INIT_02 => X"8F333007FD6808092A2AFA6667033DB50853379C10BFF70F1BD011110F205F18",
INIT_03 => X"294ADB4AFFCBF0DAD63ABF836B58EAFE060478202022234B2E0303FDC9E18339",
INIT_04 => X"DB7A40806FE4040840EBC563A0150A0926146FECB04196482236FC2005282AE1",
INIT_05 => X"0403DA0383200831C68206D7E6D0250834336D1E81500FDB306045255BFC2076",
INIT_06 => X"4470716040413D29AAC69F5FE33C072F06062C003670497AFF00291B3C0E2015",
INIT_07 => X"0849147160448EBB9537A0022DC67987042EE976ABEA77684653547819FF2000",
INIT_08 => X"E019C0C82A4E4820C15B089C380110002446045A31345000A84432409207F02D",
INIT_09 => X"983838A3BFF1030C397C060B4254064302042F803A69DB931FF4391C00002CC0",
INIT_0A => X"FB1F1F7BC81C003C001674BB55B5FBB4BB4F26A1BEE004F9D0DE08F7DE336DB2",
INIT_0B => X"28302F800633F1D0A7CC9AE74117FE01D34E82AC0CE8FCCC200A59BDD2FFE3E3",
INIT_0C => X"E9F79E9F79E9F79E9F79E9F79E9F79E9F7CF4FBCF4F000C2E225C8DE0BA05BB0",
INIT_0D => X"A5A99FD6D3FEF4BEB5FF994F0FEFFCCF8430000000D9D147E0D57AE7B79E9F79",
INIT_0E => X"0593F33FA0CF170F40006001B1A05C0000000000000008004BA78428C7AD7FE4",
INIT_0F => X"E46444357B3950A9BFBAC94CFA8581E0A9BFBAC8CCFA8580C7CAF51EF68B2976",
INIT_10 => X"B5DB54A09003E0A9BFBAC94CFA8581E0A9BFBAC8CCFA8580E46FBFCB0CBEDA57",
INIT_11 => X"BFCB1D5CFEB56A1A100D5345C1BFFE8FBDB892DB463034198E2881F3F787DF76",
INIT_12 => X"D39387F92B2935DFEAADDF38EBCFB9E3D636DCDF9B90F966BF92966D5D9E7467",
INIT_13 => X"27055EB6D555CB294981B7FB5B2954CD3013013FDF5E82AF5B6AAAE594A4E0AD",
INIT_14 => X"835C67E655BAA868610117575EA1C34BD6975D48B44A0405FC15BA7270FF2565",
INIT_15 => X"6CD2A47D0CBA96252756D7217E5E1C61DBDF5FA167F7AE5D3D21A414007F7D7E",
INIT_16 => X"000005F08000179C16DECF67F08BC02F9067ED55805600545DFE45A80E7BD07F",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"00C0000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"9A919261A1A6075D75D10DDF2F82003009EDCC4052E92E0826462117114F9818",
INIT_1B => X"8D068351A8D069A6BAE9A69A6BAE9A6BAE9A69A6BAE9A6BAE9A69A69A69A69A6",
INIT_1C => X"A8D46A351A8D46A351A8D46A351A8D46A341A0D068341A0D068341A0D068351A",
INIT_1D => X"AFFD5400000000000000000000000000000000000000000000001FFFFE000011",
INIT_1E => X"A2FFFFEAA5D7FC0000FF8015410FFFFFFFFFFFFFFDFEFF7D568A1008003DF55A",
INIT_1F => X"5A2D1400000804154BAF7D168A00A2803DE10FFAE95410FFFFFDFEFA2D16AB55",
INIT_20 => X"BAFFD56ABFF002EBDFFF000002010552A97400007BFDE10A2AA801EF08517DF5",
INIT_21 => X"FEFAAD17FFFF002EBDE000800174AA55043FEBA0004174AA5504000AA55042AA",
INIT_22 => X"7555A284175FFFFFBE8B55A2FFFFF55F7803DEBA002AAAAAAF7FBD74BA5D2EBD",
INIT_23 => X"17400FFD57DE00AAAAAAB45A2AA97545F7D16AB455D00001EFAAAAAAABA55555",
INIT_24 => X"0000000004154BA002A800BA087FE8AAAAA80000105D557FE00A2D5420AA5D04",
INIT_25 => X"D16AA00000E3DF6DBEF5D2400000000000000000000000000000000000000000",
INIT_26 => X"3F1F8FC7AAD56DB7DB6FFFDEAA5571C7010FF8412428FFFFFFFFFF7FBF8FD7EB",
INIT_27 => X"A2A0871EF145B7FF7DA2D547038140E10492FFDF6DA28A28E3DE00F7A092410E",
INIT_28 => X"2550A020BA55002AA82F7DF6DBD71C2EBFFC71C0E050004920954380871FAE00",
INIT_29 => X"BAF7F5D74924124BDFEFA2D57FFC71C2EBDE280000174825D0E3FEAA14001249",
INIT_2A => X"1C7B6A0AAA82555157555B680125FFEBFFEDB55BEFFFAF6DE38E3DEAA002EADA",
INIT_2B => X"AE28B6D545092490E10400FFDB7AE00A2AAADB45BEA092545FFDB6AB6D410007",
INIT_2C => X"00000000000000000000010080A174821424800AA007FEDAAAA284020385D5F7",
INIT_2D => X"BFDFEFF7FFEAB45A2D56AA00002EBDFFFF7D5400000000000000000000000000",
INIT_2E => X"AABDE10FF8400010A2D56AB45A2D57DFFFF7FBFFEAA555555400F780000AAFFF",
INIT_2F => X"004174AA00516AA10AA80155EF5D7BFDFEFAAD1554BA552E82000F7FFFFEAAA2",
INIT_30 => X"552ABDEBA5D0002000552A800BA55042AA10FFFFFDF55552EBDF55552E954100",
INIT_31 => X"FA2AEBFEAA082EBDEBAFFD55540000043DFEFAAD17FF45552ABFEBA080415400",
INIT_32 => X"45F7FFEABFF080015555F78028A00555155555FF84001FFAAFBFFF55FFFBEABF",
INIT_33 => X"EBAA284000BA557FE8AAAFFD155400082A82000F7FFE8A00A2AABDF45F780001",
INIT_34 => X"0000000000000000000000000000000000000010002E974005D04020BA007BFD",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"FFFFFFFE00000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000000000000000000019F",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(17),        -- Port A data input
DOA(0)   => data_read_a_hi(17),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(17),        -- Port B data input
DOB(0)   => data_read_b_hi(17),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_18_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"69844019080000A21A611406840014122A641074155FC28A2024001001801003",
INIT_01 => X"A643D920034004180005E9E3C90360C0041C0181002001602025800008440084",
INIT_02 => X"B7333980808408103F2000F81FC0FEDEAC2161B0B84D0002188011110C018041",
INIT_03 => X"0405D434003F2C020081587008020561E55116B0290000042B71240C800440F8",
INIT_04 => X"50805AC31007D6125724029216554A9847669903D640EC8E2001002604503004",
INIT_05 => X"07008000E0EA11803850C800010022660C1C0065003C0404002646DC20A02D40",
INIT_06 => X"0100001028040C093D0491A640FFC10028000280002C44D620F0228454C83810",
INIT_07 => X"08501620028007500CE801241021FE78E40486014006009044359DC707F55C20",
INIT_08 => X"9307CC082A0A4A6A01ECDCC40850001630080002A5CA500344040108120080AB",
INIT_09 => X"A0172083200B6186128040600C10C1C02009505081100088080BC6A052802001",
INIT_0A => X"002020000F0CA8428642430080438408A510185A40000008B83181C000141040",
INIT_0B => X"2E00C04C44C92A88DC42215C882E82240880000060D7030C30B885200D274404",
INIT_0C => X"10006100061000610006100061000610003080030800800C0540310130006E21",
INIT_0D => X"10202021000780004200408C1002003F66CA18A1B62622381B2B841840614006",
INIT_0E => X"806400FC503F08180050942E4200020C1B060D8306C182701404C19730108010",
INIT_0F => X"ABAF377DF1CA160820520EB3057E70E60820520F33057E72E915415900002900",
INIT_10 => X"5D48F37FAFEFE60820520EB3057E7CE60820520F33057E7EC658BF2DA7822AAB",
INIT_11 => X"BF2D4B2A80BF8FE39FD78EB0D882014A62C568FFAFC73FFDD9C2B30E0468A2AD",
INIT_12 => X"800DFC06F59F710107533C0C4E37619440FBFBAB2400AFC1600361D798F32658",
INIT_13 => X"EB9454005BAA36DEFF894823A3D1A88A2FE29D5FC6DCAA2A002DD51B6E7C728C",
INIT_14 => X"92A78606A28A5427AAB9FF4EDD251C7123E291660733EBF6FE519001BF40DEBB",
INIT_15 => X"AB58AFBFD5DE200A8EBE3A3EC110339E1DCEDC2590495BB2112E2BE4BF5F3B70",
INIT_16 => X"C1B06808348340000020301805002D008C1F92000A5F421B8000DB4910382202",
INIT_17 => X"1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06",
INIT_18 => X"B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C",
INIT_19 => X"000000000000000000000041B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1",
INIT_1A => X"8A244C16454170410412CA064A9BBECEB80EE173C2300FE3F1A3550F7DF16000",
INIT_1B => X"A552A944A2512AAA8A28A28A2AAAAAA8A28A28A2AAAAAA8A28A28A28A28A28A2",
INIT_1C => X"A25128944A25128944A25128944A25128944A25128944A25128944A25128954A",
INIT_1D => X"D2A80000000000000000000000000000000000000000000000001007FE000004",
INIT_1E => X"F7D568A1008003DF55AAFFD5410FFFFFFFFFFFFFFFFFFFFFBFDEBA552E974105",
INIT_1F => X"0FFFFFFFFFF7FBE8B55AAD16AA1000516AA005D0400010FFFFFFFFFFFFFFDFEF",
INIT_20 => X"00087BC2155087BC0010FFFFFDFEFA2D16AB55A2FFFFEAA5D7FC0000FF801541",
INIT_21 => X"0000804154BAF7D168A00A2803DE10FFAE95555FFFBE8B45A2D56ABEFFFFFFFE",
INIT_22 => X"01EF08517DF55000000010082A974AA08557DEBAFFAEBFF55AA8028B55A2D140",
INIT_23 => X"800105D2AAAA10A2D1420AAFFAEA8BFF000002010552A97400007BFDE10A2AA8",
INIT_24 => X"0000BA0004174AA5504000AA55042AABAFFD56ABFF002EBDEBA0004020BA552E",
INIT_25 => X"FBFFEBA552A95410552485000000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFF7FBF8FD7EBD16AA00000E3DF6DBEF5D2438FFFFFFFFFFFFFFFFEFF7",
INIT_27 => X"5571C7010FF8412410FFFBF8FC7E3F5EAB45BEDB6FA3800556FA00550405028F",
INIT_28 => X"5BEDB6FBC7EBF5F8E10007BC516D1C71C5010E3F1F8FC7AAD56DB7DB6FFFDEAA",
INIT_29 => X"55BE8A2DB7DA2D547038140E10492FFDF6DA28A28E3DE00F7A09256DE3F1EAB5",
INIT_2A => X"4380871FAE00A2A0871EF145B7FF45080E070280820924AA145578E92F7A4BFF",
INIT_2B => X"FEBA1C0A00092412E850005D2AAFA38A2DF45082F7AAA8BC71C0E05000492095",
INIT_2C => X"000000000000000000000AA140012492550A020BA55002AA82F7DF6DBD71C2EB",
INIT_2D => X"FFFFFFFFFBFDFEFF7FFFDEAA5D2E954105504154000000000000000000000000",
INIT_2E => X"557DE005500154AAFFFBFDFEFF7FFEAB45A2D56AA00002EBDFFFF7D5400AAFFF",
INIT_2F => X"2D57DFFFF7FBFFEAA555555400F78000010F7FBE8B55AAD16AB55F7FBFDEAA08",
INIT_30 => X"FF84001FFAAD568B45FFFBFFF55A2D568A00087BD55FF5D5555410A2D56AB45A",
INIT_31 => X"A555168A10FF803DF45FFAABDFEFAAD1554BA552E82000F7FFFFEAAA2AABDE10",
INIT_32 => X"55552E954100004174AA00516AA10AA80155EF5D7BFDF45002A974AA0800000A",
INIT_33 => X"A10FFFFFDF55552EBDEBA5D2E80010082A97410552EBDEBAA2FBD5400F7AAA8B",
INIT_34 => X"00000000000000000000000000000000000000BA5D0002000552A800BA55042A",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000080",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(18),        -- Port A data input
DOA(0)   => data_read_a_hi(18),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(18),        -- Port B data input
DOB(0)   => data_read_b_hi(18),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_19_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"042200000000000041088001001AA00000000000000000000000500802000003",
INIT_01 => X"200048000024000000000404000000000A22000800000800004A200000000001",
INIT_02 => X"032210008DEF00400060000001C008002489E0F0004037B00010101010000000",
INIT_03 => X"0000008128000000000000000000000024001620280000000000354200004008",
INIT_04 => X"000058800004C4024024001210001054B1C822009640000E2000002604003000",
INIT_05 => X"07008000E0200000000000000000200604000000001C04000026400000002C40",
INIT_06 => X"000000000000002600859AA1000D410000000000002C42010010200004C83810",
INIT_07 => X"0040380142810010564C41001140120024020280448088050008108100640000",
INIT_08 => X"83004C390242006200000868000040001020A850040AD0080426006933800DC4",
INIT_09 => X"0013200000016186100000000010C04002C00000000000707000000000000000",
INIT_0A => X"000000000B0C0000000101400040C0408100000000000008A810000000000000",
INIT_0B => X"00000000000400020000440000000000000000002F0001F00002024B20002000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"000210001D800000000000000002000964000000000000000000000000000000",
INIT_0E => X"0000000C50030008000000000000000000000000000000000000000000000000",
INIT_0F => X"101088A37034E156600D740022800EC156600D740022800D01E0412D06904000",
INIT_10 => X"0224081044914156600D7400228002C156600D7400228001098F00D0FB750500",
INIT_11 => X"00D0F2DD014010046037814EA63DBB31CE7605001008C41A061F0E7D693E6170",
INIT_12 => X"6D600000004089E12350C0E01FF23315422BABB46FEF5019146C0800380CC98F",
INIT_13 => X"130AA3592000000000629C03F3E60330C00C628908214551AC90000001036152",
INIT_14 => X"65C006070845039014460088235ACC3123E2A29148841008482A4DAC00000000",
INIT_15 => X"53A66BE7A5040018D8A8AD9090A1EC20A188235AC509FB50C2D0500B4094208D",
INIT_16 => X"000000000000000000000000000000008C01800270000061100084046086CD49",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"861A2882313054D34D301C862AA08BBA3F0C7010C6600A00200251C744192000",
INIT_1B => X"130984C261309861861861A69861861861861A69861861861861861861861861",
INIT_1C => X"6130984C26130984C26130984C26130984C26130984C26130984C261349A4C26",
INIT_1D => X"82E97400000000000000000000000000000000000000000000001007FE000002",
INIT_1E => X"FFFBFDEBA552E974105D2A801EFFFFFFFFFFFFFFFFFFFFFFFFFEAA552E954000",
INIT_1F => X"FFFFFFFFFFFFFFFFFEFF7FBFFEAA5D2E97545FFFFC2010FFFFFFFFFFFFFFFFFF",
INIT_20 => X"0008003DF555D5157410FFFFFFFFFFFFFFDFEFF7D568A1008003DF55AAFFD55E",
INIT_21 => X"FFFF7FBE8B55AAD16AA1000516AA005D04001EFFFFFFFFFFFFFBFDF45AAD16AA",
INIT_22 => X"0000FF80155EFFFFFFFFEFF7D16AB55A2D57DEBA557FEAA10080402010FFFFFF",
INIT_23 => X"6AB45FFFBFDEBA5D7FC0155FFFFD7410FFFFFDFEFA2D16AB55A2FFFFEAA5D7FC",
INIT_24 => X"000155FFFBE8B45A2D56ABEFFFFFFFE00087BC2155087BC00AAFFFBFDF45A2D5",
INIT_25 => X"FFFDEAA552E95400002095400000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFEFF7FBFFEBA552A954105524851C7FFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"000E3DF6DBEF5D25D7FFFFFFFFFFFFBFDFEFEBF5F8E92552E9556DEBF1C2038F",
INIT_28 => X"FE3F1FAF55A2D568A0000003FF7D495155428FFFFFFFFFF7FBF8FD7EBD16AA00",
INIT_29 => X"00000002010FFFBF8FC7E3F5EAB45BEDB6FA3800556FA005504051FFFFFFFDFE",
INIT_2A => X"B7DB6FFFDEAA5571C7010FF84125EFF7F1F8FC7EBD568B6DBEDF7DEBA5571EFA",
INIT_2B => X"5092E3F1F8F55AADB6DB7DEBF1FAE82557FC516DEBF1D0410E3F1F8FC7AAD56D",
INIT_2C => X"0000000000000000000016DE3F1EAB55BEDB6FBC7EBF5F8E10007BC516D1C71C",
INIT_2D => X"FFFFFFFFFFFFFFFFFFBFDEAA5D2A954000800154000000000000000000000000",
INIT_2E => X"2A955EFAAD1400AAFFFFFFFFFFFFBFDFEFF7FFFDEAA5D2E95410550415545FFF",
INIT_2F => X"7FFEAB45A2D56AA00002EBDFFFF7D540145FFFFFFFEFF7FBFFFFFAAD16AA0055",
INIT_30 => X"5500155EFF7FBFDFEFAAD568B55AAD568A0008003DFFF0855554AAFFFBFDFEFF",
INIT_31 => X"FFFFFFFEAA55517DE10080400010F7FBE8B55AAD16AB55F7FBFDEAA08557DE00",
INIT_32 => X"10A2D56AB45A2D57DFFFF7FBFFEAA555555400F780001FFF7D16AB55A2D16ABE",
INIT_33 => X"A00087BD55FF5D5555410AAD56AB45AAFFFFFEFAAD168A00557BD55FFA2D5400",
INIT_34 => X"00000000000000000000000000000000000001FFAAD568B45FFFBFFF55A2D568",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000100",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(19),        -- Port A data input
DOA(0)   => data_read_a_hi(19),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(19),        -- Port B data input
DOB(0)   => data_read_b_hi(19),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_20_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000003",
INIT_01 => X"A75FF80000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"14088080800008400F655001FFCFF80018FA8044000000000000011000000007",
INIT_03 => X"0000000000000000000000000000000024001660380000000000000000004FF8",
INIT_04 => X"000079800014CC02C034001600000000000000101EC0012EE0C0026E1E80F000",
INIT_05 => X"1F0FF433EFF0440C3902100002203F2EFC040388137C3E20C8EEC00284033CC0",
INIT_06 => X"4400080040440C000000000017FD5F239108000155FDC0000010E40087D8787A",
INIT_07 => X"08000EE00000000000000002101FF2002C00000004018001000030817FF50C00",
INIT_08 => X"FF7FCA302C0C00082148000008405550087C0000000000000002412489808000",
INIT_09 => X"44FF60000001EFBEF0040008023FDFC00000000040062A040001071004000013",
INIT_0A => X"000000002B7C0000008000000200000200A0C0040118400FABF9000000480002",
INIT_0B => X"0000000000000000000000000000004200310000000000000000200000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000400040",
INIT_0D => X"000000200000020000004000100203FF6C000000000000000000000000000000",
INIT_0E => X"00600FFC53FF001800000002004080000000000000040900005C848538000010",
INIT_0F => X"00009A9C300020080000800000003CC0080000800000003CC020007800000000",
INIT_10 => X"000000012963C0080000800000003CC0080000800000003CC100800000080000",
INIT_11 => X"800004000000000066C5000020020000000800000000C2E18001000200000800",
INIT_12 => X"000000000052B0200000014200040C2829000400000000000860F98798000100",
INIT_13 => X"4B00400000000002958000240400000000007E1B000040200000000001496004",
INIT_14 => X"4004181800000000005C5A00000200C40808000000000AF0D80080000000000A",
INIT_15 => X"0020141812737DC3020100400001C19C1D80000200400000000000015D140000",
INIT_16 => X"04010080800801810100000000000093EDFF8020000000000001001001000080",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0020000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0C8192608486879E79E681D903000030038200010089054D460400120104D204",
INIT_1B => X"86432190C86432CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB0C30C30C30C3",
INIT_1C => X"C86432190C86432190C86432190C86432190C86432190C86432190C86432190C",
INIT_1D => X"80402000000000000000000000000000000000000000000000001007FE000010",
INIT_1E => X"FFFFFFEAA552E95400082E975FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2A954100",
INIT_1F => X"0FFFFFFFFFFFFFFFFFFFFFFFDEAA5D2A954000800001EFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"BA5D2A97400FF8017410FFFFFFFFFFFFFFFFFFFFFBFDEBA552E974105D2A8000",
INIT_21 => X"FFFFFFFFFFEFF7FBFFEAA5D2E97545FFFFC21FFFFFFFFFFFFFFFFFFFFF7FBFFE",
INIT_22 => X"DF55AAFFD5400FFFFFFFFFFFFFFDFEFF7FFEAA10000417555AAD5555EFFFFFFF",
INIT_23 => X"FDFEFAAD568A0000043DF45AAFBC2010FFFFFFFFFFFFFFDFEFF7D568A1008003",
INIT_24 => X"0001EFFFFFFFFFFFFFBFDF45AAD16AA0008003DF555D51574BAFFFFFFFFFFFFB",
INIT_25 => X"FFFFEBA5D2A95410000A00000000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFDEAA552E954000020955FFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"552A95410552485010FFFFFFFFFFFFFFFFFFF7FBFDEBA5D2E95400140E001C7F",
INIT_28 => X"FFFFFFDFEFF7FFFFEAA5D2E95400E38A17438FFFFFFFFFFFFFFFFEFF7FBFFEBA",
INIT_29 => X"7DBEDF575D7FFFFFFFFFFFFBFDFEFEBF5F8E92552E9556DEBF1C21C7FFFFFFFF",
INIT_2A => X"FD7EBD16AA00000E3DF6DBEF5D2438FFFFFFFFFF7FBFDFC7EBF1E8A00080A155",
INIT_2B => X"5492FFFFFFFEFF7F1F8FD7A2D168A1008043FF6DAAFBC5028FFFFFFFFFF7FBF8",
INIT_2C => X"000000000000000000001FFFFFFFDFEFE3F1FAF55A2D568A0000003FF7D49515",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFEBA552A95410002E820000000000000000000000000",
INIT_2E => X"2E954005D2A82145FFFFFFFFFFFFFFFFFFFFFBFDEAA5D2A954000800155FFFFF",
INIT_2F => X"FFBFDFEFF7FFFDEAA5D2E95410550415410FFFFFFFFFFFFFFDFEFF7FBFFEBA55",
INIT_30 => X"AAD140155FFFFFFFFFF7FBFDFFFFFFBFDEBA5D2A95400A2AA974AAFFFFFFFFFF",
INIT_31 => X"5A2D568A10082E955FFFFFFD7545FFFFFFFEFF7FBFFFFFAAD16AA00552A955EF",
INIT_32 => X"AAFFFBFDFEFF7FFEAB45A2D56AA00002EBDFFFF7D5400BAFFFFFDFEFF7FBFFF5",
INIT_33 => X"A0008003DFFF085555410F7FBFDFEFFFD568B45AAD16AA1008003DFEFAAFBD74",
INIT_34 => X"00000000000000000000000000000000000001EFF7FBFDFEFAAD568B55AAD568",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"FFFFFFFE00000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000000000000000000001F",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(20),        -- Port A data input
DOA(0)   => data_read_a_hi(20),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(20),        -- Port B data input
DOB(0)   => data_read_b_hi(20),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_21_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"4A302428B824900A128C090A5C1800261500213C005FE812D10420054085A202",
INIT_01 => X"081FFE3440B609703B0427F801A40B8115BC4F655300340288A40D30040E4DD8",
INIT_02 => X"0109095C30C98809800000F9FFFFFFFF149FF1FCA4C0421B182E3490DF145FE4",
INIT_03 => X"084A76341244919000099486400026523C041660BA000100CC12701015007FF8",
INIT_04 => X"000079800014CC03C075161E001118653D2408041FC004AEF000816E1C11F541",
INIT_05 => X"3F0F807BFFE000240100004683103E7FFE02482553FC3C0204EFC25010143CC0",
INIT_06 => X"C42040304101118B84E4880817FD7F028000000101FFE4036450E08247F87870",
INIT_07 => X"0A09000D00204A855B000A08A61FF20C3D004D331D3400805984B7A1FFF00860",
INIT_08 => X"F7FFC08D234B4002030314D0001104500000034089902D0901A021E4015410EA",
INIT_09 => X"B4FFE10158E1FFBEF0440021083DFFCE22DC2880E24D1BFA7C98480802000023",
INIT_0A => X"A31514636FFC00080013029811240444A82422A85180778FAFF82A04B6356DD0",
INIT_0B => X"0600E20806520398C682157A49389667126880806FF917FC30010107688862A2",
INIT_0C => X"1B2451B2451B2451B2451B2451B2451B3228D9228D90800C6120881034003631",
INIT_0D => X"0403000A01282088624001201A8C43FF7C00100102A53208B2A246406081B245",
INIT_0E => X"C4053FFD5BFF00A04A00200602CA520011000880044402104803400400189000",
INIT_0F => X"63009140094D81A5040605800B506901A3040605401360562027218196506102",
INIT_10 => X"02811209062801A3040605800B506901A50406054013605604350B812822A002",
INIT_11 => X"0B811068C00049A0A5820A3C1725A8006C0A40404D058320496C2C9C600890A2",
INIT_12 => X"AC808127C454402483153A3A895BB3C1E2E820704020381702C1AAA2C4B3F435",
INIT_13 => X"CC1B154510413CC2A200501B400A40018A00C80400040D8AA288209AA2198361",
INIT_14 => X"0141AA00418080460678A4012288463B2050302019200B00206C35901024D910",
INIT_15 => X"2440470C8A9310280C0180302A01427D060022011606E800E00169C19A00048A",
INIT_16 => X"40100448008004000000E07008010003EFFFE0373056024B0111801198823314",
INIT_17 => X"0100401004010040100401004010040100401004010040100401004010040100",
INIT_18 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_19 => X"0000000000000000000000401004010040100401004010040100401004010040",
INIT_1A => X"BEFFFFF7F7FFF3CF3CFFFF9FE0FF9FEEFF7FFDF7FF3EFC2FF8107F3DFDF7E000",
INIT_1B => X"FF7FBFDFEFF7FBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEF",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FBFDFE",
INIT_1D => X"80002000000000000000000000000000000000000000000000001007FE00003F",
INIT_1E => X"FFFFFFEBA5D2A954100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974000",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFEBA552A97400082A975FFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"AA5D2E974100800155EFFFFFFFFFFFFFFFFFFFFFFFFFEAA552E95400082E975F",
INIT_21 => X"FFFFFFFFFFFFFFFFFDEAA5D2A95400080000000FFFFFFFFFFFFFFFFFFFFFFFDE",
INIT_22 => X"74105D2A80000FFFFFFFFFFFFFFFFFFFFFBFDEBA5D2E974005D2E80000FFFFFF",
INIT_23 => X"FFFFFF7FBFDEBA552A954005D2E97410FFFFFFFFFFFFFFFFFFFFFBFDEBA552E9",
INIT_24 => X"0001FFFFFFFFFFFFFFFFFFFFF7FBFFEBA5D2A97400FF80174BAFFFFFFFFFFFFF",
INIT_25 => X"FFFFEBA5D2E97400000400000000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFEBA5D2A95410000A001FFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"552E954000020955EFFFFFFFFFFFFFFFFFFFFFFFFFEAA552E97400002E955FFF",
INIT_28 => X"FFFFFFFFFFFFFBFDEAA5D2A974101400155C7FFFFFFFFFFFFFFFFFFFFFFFDEAA",
INIT_29 => X"00552A80010FFFFFFFFFFFFFFFFFFF7FBFDEBA5D2E95400140E00000FFFFFFFF",
INIT_2A => X"FEFF7FBFFEBA552A95410552485038FFFFFFFFFFFFFFFFFFF7FBFDEBA552E974",
INIT_2B => X"74AAFFFFFFFFFFFFFFFFEFF7FBFFEAA5D2E97400412497438FFFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000001C7FFFFFFFFFFFFFFDFEFF7FFFFEAA5D2E95400E38A1",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974000004000000000000000000000000000",
INIT_2E => X"2E97400002E975FFFFFFFFFFFFFFFFFFFFFFFFFFEBA552A95410002E821FFFFF",
INIT_2F => X"FFFFFFFFFFFBFDEAA5D2A954000800155EFFFFFFFFFFFFFFFFFFFFFFFFDEAA55",
INIT_30 => X"5D2A82010FFFFFFFFFFFFFFFFEFF7FBFDEBA552A974105D0015545FFFFFFFFFF",
INIT_31 => X"FF7FFFFEAA5D2A974005D2E82010FFFFFFFFFFFFFFDFEFF7FBFFEBA552E95400",
INIT_32 => X"AAFFFFFFFFFFFFBFDFEFF7FFFDEAA5D2E954105504154AAFFFFFFFFFFFFFFDFE",
INIT_33 => X"EBA5D2A95400A2AA974BAFFFFFFFFFF7FBFDFEFFFFFFDEBA552E974000004154",
INIT_34 => X"0000000000000000000000000000000000000155FFFFFFFFFF7FBFDFFFFFFBFD",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(21),        -- Port A data input
DOA(0)   => data_read_a_hi(21),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(21),        -- Port B data input
DOB(0)   => data_read_b_hi(21),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_22_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"5290F4CDE914905A14A43D33F488243E17122300F55FEB189B343A1140548380",
INIT_01 => X"A94007B259F6A975386262000C344BA9573C6FF57B18A5FB0ABFCD3C2C5F4F0C",
INIT_02 => X"877FE30EB378008D202551040030071869D0040180AC4B685F6E26FAA0810006",
INIT_03 => X"431965109E4481D6B5AAD6875AD6AB5A1815600802888808DEA83552954D3000",
INIT_04 => X"492C0020220001010E4916C884DCD607E5EC2A344103E48003D0800023D0072C",
INIT_05 => X"00107C441001100D620A06D683018001023D37E5088043620101179092540112",
INIT_06 => X"9108E1550544A451E0CE1AA94000206B541C08414402365774611E047020008E",
INIT_07 => X"809DA02F56A92FD7247E10305C40040D136E6A023F7FCF780C4C0528800C8028",
INIT_08 => X"00803A884B5B5206B7C3391F288551002401E993AF59012740A2E4F65586923D",
INIT_09 => X"040081C91AA010000560141801002028A83D2A08E06D0002FED9680A0E002A94",
INIT_0A => X"A71514E700838460402635019FBFE7FCA13520F8D580A08044081201206334A0",
INIT_0B => X"00A0220103D2A512C6A8C4F0011550070368000A0004D0000002126F30C902A2",
INIT_0C => X"0385503855038550385503855038550392A81C2A81C00280000C200006405A08",
INIT_0D => X"0D0E153941A8B1A262CA542A9A8D6C0010A1001002C500268ACA419412503855",
INIT_0E => X"089180008800143D83888281A2034A85014280A14050A01509E050854498B294",
INIT_0F => X"6706B3C189CD84ACD20B03001E387D04AC560B02401E387E1028AC0450080410",
INIT_10 => X"0201570B036C04AC560B03001E387D04ACD20B02401E387E24708E7E242000C2",
INIT_11 => X"8E7E1C20A0106EA167C84EBF052A8E010C0180606E86C3F459DC08DA90245887",
INIT_12 => X"189980254CDEC22A98032A22C50EAC462030A01800407C2700C2ACA2C0F04470",
INIT_13 => X"CC1154C258012D86F601A2E49003400138C0DA2443A208AA612C0096C3798225",
INIT_14 => X"025483C1E0C0006B085CEC03858958D15310201015504B512044A3133004A99B",
INIT_15 => X"9512C6FC01A1421006028038720640310643858162712020B001AA415F290E16",
INIT_16 => X"110445E22022365034A8EA754008004C0200323001182122548881649D16B046",
INIT_17 => X"1044110441104411044110441104411044110441104411044110441104411044",
INIT_18 => X"0401004010040100401004010040100401004010040100441104411044110441",
INIT_19 => X"22890000000003FFFFFFFF900401004010040100401004010040100401004010",
INIT_1A => X"9EFFDFF7F5F777DF7DF7DF5FEFBFBFDEFE8FF1F7DEBD6FEFF7EF6FDF7DF7D051",
INIT_1B => X"7F3F9FCFE7F3F9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7",
INIT_1C => X"E7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE",
INIT_1D => X"00000000000000000000000000000000000000000000000000001007FE00000F",
INIT_1E => X"FFFFFFEBA5D2E974000800021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E954000004001FFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"BA552A97400002A801FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2A954100804021F",
INIT_21 => X"FFFFFFFFFFFFFFFFFFEBA552A97400082A975FFFFFFFFFFFFFFFFFFFFFFFFFFE",
INIT_22 => X"5400082E975FFFFFFFFFFFFFFFFFFFFFFFFFFEAA552E95410002A955FFFFFFFF",
INIT_23 => X"FFFFFFFFFFFEAA552E95400002E975EFFFFFFFFFFFFFFFFFFFFFFFFFEAA552E9",
INIT_24 => X"000000FFFFFFFFFFFFFFFFFFFFFFFDEAA5D2E97410080015545FFFFFFFFFFFFF",
INIT_25 => X"FFFFEBA5D2E97410080002000000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974000004001FFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"5D2A95410000A001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2A954000804021FFF",
INIT_28 => X"FFFFFFFFFFFFFFFFEBA552A97400082E821FFFFFFFFFFFFFFFFFFFFFFFFFFEBA",
INIT_29 => X"10082A975EFFFFFFFFFFFFFFFFFFFFFFFFFEAA552E97400002E955FFFFFFFFFF",
INIT_2A => X"FFFFFFFFDEAA552E954000020955C7FFFFFFFFFFFFFFFFFFFFFFFFEAA552E954",
INIT_2B => X"5545FFFFFFFFFFFFFFFFFFFFFFFDEAA5D2A974001C24975C7FFFFFFFFFFFFFFF",
INIT_2C => X"00000000000000000000000FFFFFFFFFFFFFFFFFFFFFBFDEAA5D2A9741014001",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800020000000000000000000000000",
INIT_2E => X"2A954000800021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974000004001FFFFF",
INIT_2F => X"FFFFFFFFFFFFFFEBA552A95410002E821FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_30 => X"002E975EFFFFFFFFFFFFFFFFFFFFFFFFFEAA552A97400082A801FFFFFFFFFFFF",
INIT_31 => X"FFFFBFDEAA5D2E95410082E955EFFFFFFFFFFFFFFFFFFFFFFFFDEAA552E97400",
INIT_32 => X"45FFFFFFFFFFFFFFFFFFFFFBFDEAA5D2A95400080015545FFFFFFFFFFFFFFFFF",
INIT_33 => X"EBA552A974105D0015555FFFFFFFFFFFFFFFFFFF7FBFDEBA5D2A974005504175",
INIT_34 => X"0000000000000000000000000000000000000010FFFFFFFFFFFFFFFFEFF7FBFD",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"FFFFFFFE00000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000000000000000000001F",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(22),        -- Port A data input
DOA(0)   => data_read_a_hi(22),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(22),        -- Port B data input
DOB(0)   => data_read_b_hi(22),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_23_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"EF20906D902424807BC8241BC81801B97D38AD3C0800103362A6741C80A12A02",
INIT_01 => X"001FFF8409F089003B4422000D80C80106804A7951C5B9D1C828043EA28838F9",
INIT_02 => X"073B8858218C2C50801000F9FFEFF8E72CA7F5FC2E048026496834D84721DFE0",
INIT_03 => X"2C4360101A4001001005080400401420350016E0BB222341C312000014006FF8",
INIT_04 => X"00017B810015DC03D034201E14000036486008101FC0002EE006297E1C05F561",
INIT_05 => X"BF0F817FFFE80100004044800080BEFFFC0248005FFC3C18A5FFC2444484BCC0",
INIT_06 => X"00000070604191C93F02800017FF7F002000020001FFC0832050E00047F97870",
INIT_07 => X"AE4080091A0071070FA07A1CB23FFA403F0C4D23BF7C0EF85788B681FFFC6C20",
INIT_08 => X"F7FFD8880A034AC096620C46AC5055508401A24684227DB880000008B05001A3",
INIT_09 => X"21FFE0004047FFBEF2000000001DFFC612C0C04001000BF8000000804000003F",
INIT_0A => X"000000006FFEA002020626995FBE077430001E734020DF0FAFF5080496044B51",
INIT_0B => X"0600C48907120AC81083315A49388660180082A06FF907FC3081812048006000",
INIT_0C => X"182021820218202182021820218202182010C1010C10800C6120885430003631",
INIT_0D => X"80600020040030090000012A500003FF7E081881902233483828864860A18202",
INIT_0E => X"C7043FFD5FFF00A04BC010A7724B100008000400020000415003001000400002",
INIT_0F => X"290C2909080A872BC4FC8500054840072FC0FC8440054840200705F986106542",
INIT_10 => X"0180F1082E00072FC0FC8500054840072BC4FC84400548402214A380380B2080",
INIT_11 => X"A380344920080B21810240AB182EB37C380B40800707011001B43253EE50C822",
INIT_12 => X"E4000026C00C00042BD4149067465910640A0050C060A0028063672A00019214",
INIT_13 => X"800CCB050001344060211629580B80022480A444111706658280009A2030019C",
INIT_14 => X"232D6D0100C040250200845132C10BE200403018061101A220339C800004D801",
INIT_15 => X"2A5493B8E287E03808480060E40C83C1405132C90742E408D0082140820944CB",
INIT_16 => X"00802000100100000000000004002403EFFF8002385F03490101946500140210",
INIT_17 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_18 => X"8020080200802008020080200802008020080200802008020080200802008020",
INIT_19 => X"0000000000000000000000008020080200802008020080200802008020080200",
INIT_1A => X"0000000000000000000000000000000000000000000000000040000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"80400000000000000000000000000000000000000000000000001007FE000000",
INIT_1E => X"FFFFFFEBA5D2E974100000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100004021FFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"BA5D2E954000800001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974000800021F",
INIT_21 => X"FFFFFFFFFFFFFFFFFFEBA5D2E954000004001FFFFFFFFFFFFFFFFFFFFFFFFFFE",
INIT_22 => X"54100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2A954100000021FFFFFFFF",
INIT_23 => X"FFFFFFFFFFFEBA5D2A954100800021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2A9",
INIT_24 => X"0001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA552A97400002A801FFFFFFFFFFFFFFF",
INIT_25 => X"FFFFEBA5D2E97410080400000000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800021FFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"5D2E974000004001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100004021FFF",
INIT_28 => X"FFFFFFFFFFFFFFFFEBA5D2E954000800001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA",
INIT_29 => X"100004021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2A954000804021FFFFFFFFFF",
INIT_2A => X"FFFFFFFFFEBA5D2A95410000A001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2A954",
INIT_2B => X"21FFFFFFFFFFFFFFFFFFFFFFFFFFEBA552A97410080E001FFFFFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA552A97400082E8",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804000000000000000000000000000",
INIT_2E => X"2E974100000021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800021FFFFF",
INIT_2F => X"FFFFFFFFFFFFFFEBA5D2E974000004001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_30 => X"0800021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E954000804021FFFFFFFFFFFF",
INIT_31 => X"FFFFFFFEBA552A954100004001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2A95400",
INIT_32 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA552A95410002E821FFFFFFFFFFFFFFFFFFF",
INIT_33 => X"EAA552A97400082A801EFFFFFFFFFFFFFFFFFFFFFFFFFEAA552A97410002A821",
INIT_34 => X"00000000000000000000000000000000000001EFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"FFFFFFFE00000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000000000000000000001F",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(23),        -- Port A data input
DOA(0)   => data_read_a_hi(23),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(23),        -- Port B data input
DOB(0)   => data_read_b_hi(23),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_24_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100600007FFF000080108004000800020000840041000080808",
INIT_02 => X"172A00D000EF8210000000F9FFEFF8E7240FF1FC224087B1000639401D005FC0",
INIT_03 => X"00003A2E200811000000000400000000340016603A0000004860400014006FFF",
INIT_04 => X"000079800014CC03C034001E04010850300000101FC0002EE000006E1C00F500",
INIT_05 => X"1F0F8033FFE000000000000000003E2FFC024800137C3C0000EFC00000003CC0",
INIT_06 => X"00000040004111CE08AA800017FD7F000000000001FFC0000010E00007F87870",
INIT_07 => X"001080040814210254000A00B21FF2003F2A80D5000006E461803081FFF40000",
INIT_08 => X"F7FFD88D2B4A02C0940018EB0A1000058400810205E2D8030900004D925821CC",
INIT_09 => X"20FFE0000001FFBEF0000000001DFFC002C0000000000BF80000000000000003",
INIT_0A => X"000000006FFE80000015406A80000338800002500000470FAFF0080496044950",
INIT_0B => X"0600C008140800080000100248288660100080806FD107FC3000000000006000",
INIT_0C => X"182001820018200182001820018200182000C1000C10800C6020881030002431",
INIT_0D => X"000900160000000000000000000003FF7C001001002032083020060060018200",
INIT_0E => X"C4043FFD5BFF0000410000000041100000000000000000004003000000000000",
INIT_0F => X"1080012302010049400086C02200420049400087802200412027059996516100",
INIT_10 => X"0300081406100049400086C0220042004940008780220041248190818403A042",
INIT_11 => X"90814C09C01010400132100106836001504240E01040051200200D06410C1924",
INIT_12 => X"680C0100010408240BD80008983596CD86EA84104060503C0B00002025023481",
INIT_13 => X"90164F40086000082062C1B6600BC000C300818044000B27A0043000041202CD",
INIT_14 => X"2577FE4080C08010842180C40018545BBA00301808A0810C0059AD0180200020",
INIT_15 => X"04100852B931F00800010081980B042D2044001850ED8808F00050A002C11000",
INIT_16 => X"00000000000000000000000000000003EFFF80037046031E0110001100A4820C",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"BEC99E61848655D75D7FCB598CC0AEEAF6E7CC1132CD73C8261273B444199000",
INIT_1B => X"0F0783C1E0F07BEFBEFBEF9E79E79E79E79E7BEFBEFBEFBEFBEFBE7BE7BE7BE7",
INIT_1C => X"E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E",
INIT_1D => X"80402000000000000000000000000000000000000000000000001007FE000001",
INIT_1E => X"FFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800021FFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"BA5D2E974100000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100000001F",
INIT_21 => X"FFFFFFFFFFFFFFFFFFEBA5D2E974100004021FFFFFFFFFFFFFFFFFFFFFFFFFFE",
INIT_22 => X"74000800021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974000004001FFFFFFFF",
INIT_23 => X"FFFFFFFFFFFEBA5D2E974000800001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9",
INIT_24 => X"0001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E954000800001FFFFFFFFFFFFFFF",
INIT_25 => X"FFFFEBA5D2E97410080402000000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"5D2E974100800021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800021FFF",
INIT_28 => X"FFFFFFFFFFFFFFFFEBA5D2E974100000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA",
INIT_29 => X"000004001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100004021FFFFFFFFFF",
INIT_2A => X"FFFFFFFFFEBA5D2E974000004001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_2B => X"01FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E954000800021FFFFFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9540008000",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804020000000000000000000000000",
INIT_2E => X"2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFF",
INIT_2F => X"FFFFFFFFFFFFFFEBA5D2E974100800021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_30 => X"0000021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100000001FFFFFFFFFFFF",
INIT_31 => X"FFFFFFFEBA5D2E974000004021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E97410",
INIT_32 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974000004001FFFFFFFFFFFFFFFFFFF",
INIT_33 => X"EBA5D2E954000804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E954000004021",
INIT_34 => X"00000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(24),        -- Port A data input
DOA(0)   => data_read_a_hi(24),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(24),        -- Port B data input
DOB(0)   => data_read_b_hi(24),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_25_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100200002000000080100004000000020000800041000080808",
INIT_02 => X"1000218000000800000000F9FFEFF8E738FFF1FC20400400000004455A375FE0",
INIT_03 => X"00002000000001000000000400000000340016623A0000004000000014006FFF",
INIT_04 => X"924279824C94CC1BE0B4001F20000000020380401FE0082EF000106E1C00F500",
INIT_05 => X"1F0F8033FFF048202582800100523E2FFE024820137C3C0040EFE02000003CE4",
INIT_06 => X"D4A00671414191800000800017FD7F038100201101FFC0000010E08A07FC7870",
INIT_07 => X"080000000000000000000A00B21FF2003E0000000000066041803081FFFC2C60",
INIT_08 => X"F7FFFA0008000200A0400002280000050400800204000000000201202B800000",
INIT_09 => X"B4FFF0008001FFBEF80C40630C7DFFEEBAF0008002021BF80000400A02000003",
INIT_0A => X"000000006FFF800C0400000000000330080000500006470FAFFD29F7DE565971",
INIT_0B => X"0600C008040000080000100248688760101080806FD107FC3018000000006000",
INIT_0C => X"182001820018200182001820018200182000C1000C10800EE6618911398524B1",
INIT_0D => X"000000000000000000000002500003FF7C001001002032083120060060018200",
INIT_0E => X"C6043FFD5BFF00A04B80608003CB120C11060883044582114013412080000000",
INIT_0F => X"000000200200000900000400200000000900000400200000200701E186106140",
INIT_10 => X"0000001000000009000004002000000009000004002000000000808000002000",
INIT_11 => X"8080000800000000001010000002200000004000000004000000000240000020",
INIT_12 => X"2000000001000004031802000004100000100024400000000800800001000000",
INIT_13 => X"0000410000000008000000204004000000000100040000208000000004000004",
INIT_14 => X"0004200001000200000100040000004200004020000000040000840000000020",
INIT_15 => X"00000010800000000C0A00000000040000040000004080000000000000401000",
INIT_16 => X"451044C82082068C0200000008014023EFFFC006304602080100000100000308",
INIT_17 => X"1104411044110441104411044110441104411044110441104411044110441104",
INIT_18 => X"1044110441104411044110441104411044110441104411044110441104411044",
INIT_19 => X"00002FFFFFFFFFFFFFFFFFC11044110441104411044110441104411044110441",
INIT_1A => X"042824014C48569A69AFEE9E50B2894A196A8C5A2932F7C8086034EC15DA0808",
INIT_1B => X"6231188C46231249249249249249249249249041041041041041041249041249",
INIT_1C => X"562B158AC562B158AC562B158AC562B158AC562B158AC562B158AC56231188C4",
INIT_1D => X"80400000000000000000000000000000000000000000000000001FFFFE00002C",
INIT_1E => X"FFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"BA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001F",
INIT_21 => X"FFFFFFFFFFFFFFFFFFEBA5D2E974100800021FFFFFFFFFFFFFFFFFFFFFFFFFFE",
INIT_22 => X"74100000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800001FFFFFFFF",
INIT_23 => X"FFFFFFFFFFFEBA5D2E974100000021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9",
INIT_24 => X"0001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100000001FFFFFFFFFFFFFFF",
INIT_25 => X"FFFFEBA5D2E97410080400000000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFF",
INIT_28 => X"FFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA",
INIT_29 => X"100800001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800021FFFFFFFFFF",
INIT_2A => X"FFFFFFFFFEBA5D2E974100800021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_2B => X"01FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100000021FFFFFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741000000",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804000000000000000000000000000",
INIT_2E => X"2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFF",
INIT_2F => X"FFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_30 => X"0804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFF",
INIT_31 => X"FFFFFFFEBA5D2E974100800001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E97410",
INIT_32 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800021FFFFFFFFFFFFFFFFFFF",
INIT_33 => X"EBA5D2E974100000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800021",
INIT_34 => X"00000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"FFFFFFFE00000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000000000000000000001F",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(25),        -- Port A data input
DOA(0)   => data_read_a_hi(25),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(25),        -- Port B data input
DOB(0)   => data_read_b_hi(25),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_26_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"E9264EAB20190CA3BA4997AA9002AE9C001006B0778015CFA17E0811039879C7",
INIT_01 => X"F1FFF9BB1F773C7F9BB07DFFFDD863FC5FFF3FEFFBBF9FFB22FFFBC7B9F30686",
INIT_02 => X"1B33188302E708180F6FFBFFFFCFFFFF9C7FF7FC24350B99082400001D00DFD8",
INIT_03 => X"4A53D958C50000DCE7366303739CD98C27C57EF57980014F271807E3C9E9CFF8",
INIT_04 => X"DBFAFBD7FB1CDEBEF1BE17F7AC88042787FBFFF8FEE9FF7EE6F4C0EE1FFAF869",
INIT_05 => X"5F0FFEB3EFFEFFBDA7F7FED508707E2EFEBF6FFEB37C3FF302EEEDFF9B487CF6",
INIT_06 => X"67F2B27AFAD11587B7C094F1FFFFDF0FAF4E8FAA67FDDB7FB870FF30FFDEF87F",
INIT_07 => X"08180EF060C18E5BEFB051225CDFF7002C4EEDE77F6E0EFD044ABC817FFFDD35",
INIT_08 => X"FF7FC8790E46426CE06C2C7E381041460C7E8C1A35DF80000C0084C9188302E7",
INIT_09 => X"2CFF7A27B303EFBEFAFCC2E35E7FDFD147CCF3F583FA3FFF7D6000EC75088ED3",
INIT_0A => X"5A3A3B5AFF7CFACFAFE776F39FF7077E29D83CFAE601602FEBFFCDF7DEE77DF7",
INIT_0B => X"3EB1EDDCDEBCFF589807B70AD9A99EE41FD18884FFF19FFC71FEFED7B251E747",
INIT_0C => X"1AF181AF181AF181AF181AF181AF181AF4C0D78C0D718ADEEE61D99B7BE2A433",
INIT_0D => X"B9EC20181CC1F73F87501DED3409BFFFEFFEBCEBFE68370CFA6D07407481EF18",
INIT_0E => X"CE04FFFFF3FF1F5F5475BD7F72E4D75EBFAF5FD7AFEFDFFAF59B6FF28FE1D406",
INIT_0F => X"7C040101480807D17B0004001F804007D17B0004001F8040212F35FFC6D86D70",
INIT_10 => X"0001DC00068007D17B0004001F804007D17B0004001F804006F6008140002000",
INIT_11 => X"0081800800007B000102C0801FB02683800040007700011801003DE050A70020",
INIT_12 => X"32130207080D012CEFF41008D188D502100B02004000F01900039020040206F6",
INIT_13 => X"A01F21A2C40039006823F80048100003F0008004D8100F90D162001C803403E2",
INIT_14 => X"27F020A07400007C040085581019D602451500001EC00100247C46426080E101",
INIT_15 => X"2010EA40EA00020C830100F0D000022180581019F40084800001F100020B6040",
INIT_16 => X"EFFBFEFDFDDFE7DD87FEFF7FF796FFFFFDFFC017FEFFD7E841001D8197DCC3F0",
INIT_17 => X"BFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAF",
INIT_18 => X"FAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFE",
INIT_19 => X"88646FFFFFFFFFFFFFFFFFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEB",
INIT_1A => X"86EBCAF55357E1C71C751D53C44B15BCF491E166CC853E8117696853F86EDB5C",
INIT_1B => X"130984C261309861861861861861861861861861861861861861861A69A69861",
INIT_1C => X"6130984C26130984C26130984C26130984C26130984C26130984C26130984C26",
INIT_1D => X"80400000000000000000000000000000000000000000000000001007FE000002",
INIT_1E => X"FFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"BA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021F",
INIT_21 => X"FFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFE",
INIT_22 => X"74100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFF",
INIT_23 => X"FFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9",
INIT_24 => X"0001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFF",
INIT_25 => X"FFFFEBA5D2E97410080400000000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFF",
INIT_28 => X"FFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA",
INIT_29 => X"100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFF",
INIT_2A => X"FFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_2B => X"21FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008040",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804000000000000000000000000000",
INIT_2E => X"2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFF",
INIT_2F => X"FFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_30 => X"0804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFF",
INIT_31 => X"FFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E97410",
INIT_32 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFF",
INIT_33 => X"EBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001",
INIT_34 => X"00000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(26),        -- Port A data input
DOA(0)   => data_read_a_hi(26),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(26),        -- Port B data input
DOB(0)   => data_read_b_hi(26),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_27_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"00080A40000A41248002029000050A088000008242A0004404480002000A1155",
INIT_01 => X"F1FFF1C11F781C129C107DFFFE0860941E81258CA2B71C2220EC1B86E1A00002",
INIT_02 => X"4000002100000014400FF6FFFF0FFFFF8007F1FC211100014200800000887FC0",
INIT_03 => X"0842D85841000098C63061026318C18404C459757000015F00088BE3C0618FF8",
INIT_04 => X"DBEAE5D6D91C2EBCE1B21EA72C00000007FBE7C8F8E9EF79E6D440E91FDAE061",
INIT_05 => X"5C8FFCB38FF6B68984B5BCE408347E28FEBF6FEEB3723F7102E8EDBF8A4872F6",
INIT_06 => X"6E62106ADAD14180035044F1FFFC9F0C0E4C8DAAEFF1DB7FA868FE30EF1CE47E",
INIT_07 => X"0014401060C180190310540118DFF1000C0849673F6C06FE000A38007FF13115",
INIT_08 => X"F47FC80208808210880C00020814000044008C1A340C00000A08000000210000",
INIT_09 => X"04FC721491038F7DF8BEC2E39C5F1FD047CEF1B582D83FF779200062B12A8EC3",
INIT_0A => X"02606042787C5AC5ADC424B39FB6073D00D8048A6201002F83F04DFFDE83FDD6",
INIT_0B => X"56B5F0DEFABC705488069302DBA98EAC16C1A884FFE18FFD757E7ED7A211EC0C",
INIT_0C => X"186881868818688186881868818688187840C3440C35A8DFEE61CB9979AAA433",
INIT_0D => X"D1F820101441DA3A8310198C34089BFF8DD6B56B6F28378C7E2D07007801C688",
INIT_0E => X"E4047FFD23FF315D54358D593474955AB6AD5B56ADAB5FAAE58B2F628EA0C407",
INIT_0F => X"7C0400004C080791290004001D80001791290004001D8000210F15879715710A",
INIT_10 => X"0001DC0000801791290004001D80001791290004001D800012F6008040002000",
INIT_11 => X"0080800800007B000000E0801BB020828000400077000008210035E040830020",
INIT_12 => X"220202070801010C6F1410085188D500100102004000F01900031000060202F6",
INIT_13 => X"205D2120840039000813F80040100003F0000000F8100E909042001C80040BA2",
INIT_14 => X"07F020201400007C040001781011D602040500001EC00000057444404080E100",
INIT_15 => X"2000EA40EA000004810100F0D000020080781011F40080800001F1000003E040",
INIT_16 => X"AB6BDE75ED5EC71385FC2512E3565BBBF1FFC00636EED7E841000D81924C43F0",
INIT_17 => X"B6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6AD",
INIT_18 => X"6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADA",
INIT_19 => X"88747FFFFFFFFFFFFFFFFFAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB",
INIT_1A => X"00780401CBC8400000052412F84E2168100481CA8604368008402F02104A4716",
INIT_1B => X"4020100804020000000000000000000000000000000000000000208000000000",
INIT_1C => X"140A05028140A05028140A05028140A05028140A05028140A050281402010080",
INIT_1D => X"80400000000000000000000000000000000000000000000000001007FE000028",
INIT_1E => X"FFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"BA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001F",
INIT_21 => X"FFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFE",
INIT_22 => X"74100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFF",
INIT_23 => X"FFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9",
INIT_24 => X"0001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFF",
INIT_25 => X"FFFFEBA5D2E97410080400000000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFF",
INIT_28 => X"FFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA",
INIT_29 => X"100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFF",
INIT_2A => X"FFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_2B => X"21FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008040",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804000000000000000000000000000",
INIT_2E => X"2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFF",
INIT_2F => X"FFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_30 => X"0804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFF",
INIT_31 => X"FFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E97410",
INIT_32 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFF",
INIT_33 => X"EBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021",
INIT_34 => X"00000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"FFFFFFFE00000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000000000000000000001F",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(27),        -- Port A data input
DOA(0)   => data_read_a_hi(27),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(27),        -- Port B data input
DOB(0)   => data_read_b_hi(27),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_28_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"02200AA400180030808802A900002A08001280A08A801044104A1000001818C3",
INIT_01 => X"50A00011460214428114180000882214413D0A71592A01D92213D28005210202",
INIT_02 => X"1444428102100884000AA30200000000C1000401041108404400022220800000",
INIT_03 => X"461080404900000C6314A900318C52A40051081000888806108802A141288001",
INIT_04 => X"00800040110102000902002000888400081045A8A00003C00000500000080008",
INIT_05 => X"0000000000024CA0A0101800032000400000000B800000014000000B08180000",
INIT_06 => X"0040B0000804001040000450A00080444A002480220009A88800009A88000000",
INIT_07 => X"088400122448908A204020004080010000408200000001000002080000099000",
INIT_08 => X"0000028040101004200C21002084555500004489120509244022801244810210",
INIT_09 => X"9000008101400000049016080102000220001110001020058320402A16002650",
INIT_0A => X"A53534A50000080080E041000000008000C81000220020A00004000000300003",
INIT_0B => X"0090024440245400082D0220800008000081022C0000080000206CB0821086A6",
INIT_0C => X"02C0A02C0A02C0A02C0A02C0A02C0A02C050160501600240010860CC04200280",
INIT_0D => X"1884200810C1631181500CA60400B40080720020240A00004005800800206C0A",
INIT_0E => X"0A00C000200005000010040A0020CC000200010000800920040804020A605400",
INIT_0F => X"0000000140000010290000000280000010290000000280000100180210410442",
INIT_10 => X"0000000004800010290000000280000010290000000280000002000040000000",
INIT_11 => X"0000800000000000000280000010008280000000000000180000002000830000",
INIT_12 => X"0202020000090100548000000080000010010200000000000000900000000002",
INIT_13 => X"2000202084000000480008000010000000000004880000101042000000240002",
INIT_14 => X"0080002014000000000005080000800004050000000000002400404040800001",
INIT_15 => X"00002000000000048100000000000020800800008000008000000000000A2000",
INIT_16 => X"80210810840861CD33548542A10209D4100000010200400000000880035840A0",
INIT_17 => X"0200802008020080200802008020080200802008020080200802008020080200",
INIT_18 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_19 => X"22E1000000000000000000002008020080200802008020080200802008020080",
INIT_1A => X"200360D4141D630C30C7788C0211102C110A00246972C0C19D0154BD89A40A0C",
INIT_1B => X"6030180C06030208208208208208208208208208208208208208208208208208",
INIT_1C => X"160B0582C160B0582C160B0582C160B0582C160B0582C160B0582C16030180C0",
INIT_1D => X"80400000000000000000000000000000000000000000000000001007FE00002C",
INIT_1E => X"FFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"BA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001F",
INIT_21 => X"FFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFE",
INIT_22 => X"74100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFF",
INIT_23 => X"FFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9",
INIT_24 => X"0001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFF",
INIT_25 => X"FFFFEBA5D2E97410080400000000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFF",
INIT_28 => X"FFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA",
INIT_29 => X"100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFF",
INIT_2A => X"FFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_2B => X"01FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008040",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804000000000000000000000000000",
INIT_2E => X"2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFF",
INIT_2F => X"FFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_30 => X"0804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFF",
INIT_31 => X"FFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E97410",
INIT_32 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFF",
INIT_33 => X"EBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001",
INIT_34 => X"00000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"FFFFFFFE00000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000000000000000000001F",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(28),        -- Port A data input
DOA(0)   => data_read_a_hi(28),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(28),        -- Port B data input
DOB(0)   => data_read_b_hi(28),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_29_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"79964E4BA01DACAB9E659792D00AAE160002829C7FDFEFCEE97C2815039D70C3",
INIT_01 => X"50BFF9AB0775343F9AB01DF80D5821FC0FFF3FEFD1AF9FF1207FFBC7B9720586",
INIT_02 => X"0B33180300E700080F6AAA7BFFC007189C7FF2FC003503980A0000001D00DFD8",
INIT_03 => X"0401D940CD0000C8421A2B03210868AC23403E903900010E271006A148A0C000",
INIT_04 => X"49B87A417315D20A313E17F1800000058013DDF8BE21F36E02F0D06E03E8F800",
INIT_05 => X"1F007E33E01A4D9C87525E5101603E6E023D27DA937C03E340EE25CB9B483C12",
INIT_06 => X"4570301028001487B7809450B7FFC007AB0E068023FC3BFC98101F109FC6780F",
INIT_07 => X"00080EF020408EC8CFA01122149FF700200665A35D260B250442BC8100177C20",
INIT_08 => X"FF00007906464068406C0C7E100000020C7E840A15D6800044200049180300E7",
INIT_09 => X"A8FF18222341E0820AD40201423FC00122C4935001722BFD056040A452000443",
INIT_0A => X"5A2A2B5AAF00A80A82C332D18ED301D229C82C7AA600402FE80B8813485534A2",
INIT_0B => X"28102D445624DB481806A628810018400B9100042FF0180000ABFEF892508545",
INIT_0C => X"00D1A00D1A00D1A00D1A00D1A00D1A00D4D0068D006000428200508A0A600280",
INIT_0D => X"B0E8201018C1561E855008C50401B7FFE27A08A0B64A0100CA45814814A04D1A",
INIT_0E => X"4400DFFFF0001F1F0050342D42A086040B02058102C48970541944B20FA15402",
INIT_0F => X"00000101480000507B00000002804000507B000000028040212034FAD2892832",
INIT_10 => X"00000000068000507B00000002804000507B0000000280400402000140000000",
INIT_11 => X"00018000000000000102C0000410068380000000000001180000082010A70000",
INIT_12 => X"12130200000D0120ED64000080800002100B0200000000000000902004000402",
INIT_13 => X"A00220A2C4000000682008000810000000008004D80001105162000000340042",
INIT_14 => X"208000A074000000000085580008800045150000000001002408424260800001",
INIT_15 => X"001020000000020C8300000000000021805800088000048000000000020B6000",
INIT_16 => X"C4B12C989489418D13FE7F3FFD8BADB7FC004012CA5141600000198087D8C0F0",
INIT_17 => X"0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02",
INIT_18 => X"B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C",
INIT_19 => X"00602FFFFFFFFFFFFFFFFFC0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0",
INIT_1A => X"AEFFFFF7E7EFBFFFFFFAEF1DE1EF9F96EE7FFDF7FE78FC2FE8847F3FFDFFEA0C",
INIT_1B => X"F7FBFDFEFF7FBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBAEBAEBAEBAEB",
INIT_1C => X"FF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEF",
INIT_1D => X"80400000000000000000000000000000000000000000000000001007FE00003E",
INIT_1E => X"FFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"BA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001F",
INIT_21 => X"FFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFE",
INIT_22 => X"74100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFF",
INIT_23 => X"FFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9",
INIT_24 => X"0001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFF",
INIT_25 => X"FFFFEBA5D2E97410080400000000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFF",
INIT_28 => X"FFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA",
INIT_29 => X"100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFF",
INIT_2A => X"FFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_2B => X"01FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008040",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804000000000000000000000000000",
INIT_2E => X"2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFF",
INIT_2F => X"FFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_30 => X"0804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFF",
INIT_31 => X"FFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E97410",
INIT_32 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFF",
INIT_33 => X"EBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001",
INIT_34 => X"00000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(29),        -- Port A data input
DOA(0)   => data_read_a_hi(29),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(29),        -- Port B data input
DOB(0)   => data_read_b_hi(29),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_30_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"9EEBFEF5D7D7F7DF7DFFDFDFCEFFBFFEFF9FE1F7FFBFEFC9B77B7FFFFDFFD000",
INIT_1B => X"7F3F9FCFE7F3F9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7",
INIT_1C => X"E7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE",
INIT_1D => X"80400000000000000000000000000000000000000000000000001007FE00000F",
INIT_1E => X"FFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"BA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001F",
INIT_21 => X"FFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFE",
INIT_22 => X"74100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFF",
INIT_23 => X"FFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9",
INIT_24 => X"0001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFF",
INIT_25 => X"FFFFEBA5D2E97410080400000000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFF",
INIT_28 => X"FFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA",
INIT_29 => X"100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFF",
INIT_2A => X"FFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_2B => X"01FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008040",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804000000000000000000000000000",
INIT_2E => X"2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFF",
INIT_2F => X"FFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_30 => X"0804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFF",
INIT_31 => X"FFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E97410",
INIT_32 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFF",
INIT_33 => X"EBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001",
INIT_34 => X"00000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(30),        -- Port A data input
DOA(0)   => data_read_a_hi(30),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(30),        -- Port B data input
DOB(0)   => data_read_b_hi(30),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_31_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"129000008004A00804A40000400800020000000C005FEA005800200400050100",
INIT_01 => X"A15FF18019700810180065FFFC0040801E80258CA2951C2200EC0906A0804140",
INIT_02 => X"0000000000000011000550FDFF0FFFFF0007F1FC200000011000000000205FC0",
INIT_03 => X"08425818000000908428C0024210A30004045060302223490002014280410FF8",
INIT_04 => X"DB6A618248140C18E0B016872400000007EBA24058E1ECA8E2D400681FD0E061",
INIT_05 => X"1C0FFC338FF01009048084C400103E28FE3F6FE513703F7000E8E5B4825030F6",
INIT_06 => X"4420006040410180034000A157FC1F08040C080045F1F2572060FE82671C607E",
INIT_07 => X"001100004081001103107000185FF0000C0849673F6C06FC000830007FF00000",
INIT_08 => X"F47FC80008000200800000020811000004008812240800000800000000000000",
INIT_09 => X"04FC700090038F3CF82C44630C5D1FC002CCE08082481BF27A00000000000883",
INIT_0A => X"00000000687C0044040424B39FB6073C0010048A4000008F83F009F7DE037DD0",
INIT_0B => X"0620E08812982050800A910249298624124080886FE187FC301B124F20016000",
INIT_0C => X"182001820018200182001820018200183000C1000C10808EE661891139802431",
INIT_0D => X"816800100400902A0200110810080BFF0C8010010220330C3A28070070018200",
INIT_0E => X"C4043FFD03FF101D400080013040180810040802040102004183012084808006",
INIT_0F => X"7C04000008080781000004001D00000781000004001D0000200F018586106100",
INIT_10 => X"0001DC0000000781000004001D00000781000004001D000002F4008000002000",
INIT_11 => X"0080000800007B00000040801BA020000000400077000000010035C040000020",
INIT_12 => X"200000070800000C231410085108D500000000004000F01900030000040202F4",
INIT_13 => X"001D0100000039000003F00040000003F000000050100E808000001C800003A0",
INIT_14 => X"077020000000007C0400005010115602000000001EC00000007404000000E100",
INIT_15 => X"2000CA40EA000000000100F0D000020000501011740080000001F10000014040",
INIT_16 => X"010044602002061004A820104809402BE1FFC006304E03684100050190040350",
INIT_17 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_18 => X"0040100401004010040100401004010040100401004010040100401004010040",
INIT_19 => X"00802FFFFFFFFFFFFFFFFF810040100401004010040100401004010040100401",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000010",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"80400000000000000000000000000000000000000000000000001007FE000000",
INIT_1E => X"FFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"BA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001F",
INIT_21 => X"FFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFE",
INIT_22 => X"74100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFF",
INIT_23 => X"FFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9",
INIT_24 => X"0001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFF",
INIT_25 => X"FFFFEBA5D2E97410080400000000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFF",
INIT_28 => X"FFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA",
INIT_29 => X"100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFF",
INIT_2A => X"FFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_2B => X"01FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008040",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804000000000000000000000000000",
INIT_2E => X"2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFF",
INIT_2F => X"FFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_30 => X"0804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFF",
INIT_31 => X"FFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E97410",
INIT_32 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFF",
INIT_33 => X"EBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001",
INIT_34 => X"00000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(31),        -- Port A data input
DOA(0)   => data_read_a_hi(31),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(31),        -- Port B data input
DOB(0)   => data_read_b_hi(31),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_0_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"ED39BA795990D275FB4A6E96ACC4731DEA4598B0AFB54867F6EE4618C3749807",
INIT_01 => X"58A0047D8607944AC7DA180001ECA2544042106208408208C20022E9173734B3",
INIT_02 => X"9F775E7CB273E6CCA7DAAF00001000000478020113C9C38E09FB7CCCDD9F203E",
INIT_03 => X"441406267B4CB04443163C91110C58F24A31000B8028A810A3D0F8B169A01006",
INIT_04 => X"0005802424830120024121209088809DF81454ACA01E03501D0A3B91E00F0A00",
INIT_05 => X"E0F001CC00012034C20B0232838F80D001C0100AEC83C008EF101A034C8CC300",
INIT_06 => X"908A0D058584A45164BE6E58A000000583F08459A2000DA8C40F003C80030780",
INIT_07 => X"E6CCAFDC3870EEEEC44E2BDFE220094D03022210C011C103FB860B28000007C9",
INIT_08 => X"080032BF07C7C1FC3F87253D96C45557ABFF070C19D62C9065EAF36919FCB273",
INIT_09 => X"DB0009EF68EC0000045082984202002DB93119096025040581B9691E8A88262C",
INIT_0A => X"8014546E000344A0488111084048E082D0ED020133A6BF200005F60820B88206",
INIT_0B => X"28000947E16656074EA560F08054490B01280A26900C4800814069B0C8888008",
INIT_0C => X"03DCF03CCF03DCF03CCF03DCF03CCF038E780C6781C008500804708A42255A88",
INIT_0D => X"7095352BD2A90515A1CA44E7EA84B00001010012008700624187C09C0E707CCF",
INIT_0E => X"0B92800224008AE09F8942C48D1BC49120489024481225058860128543287291",
INIT_0F => X"038ABACB83C7E03EA5FF83C002783F103EA5FF83C002783F0120847A70470C7E",
INIT_10 => X"0380230F2D7C103EACFF83C002783F103EACFF83C002783F310BBF7EFC2B80C2",
INIT_11 => X"BF7EFC61E01804E1E6EA1E3FA01FD97EFC4B80E008C7C2F678FF023FAF5BD987",
INIT_12 => X"CC8E8320C4DAC9220C6B2FF22EF72ADDE6F1A67C80600C2683E0EF8AE1F1F10B",
INIT_13 => X"5C00FE651C6104C6D6400FFFB01FC0000FC07EE42FA7C07F22CE3082636B801F",
INIT_14 => X"C08FDF4195C0C2038A7C6CAFA7E289F9BA4570380131CAFB2003F9D190A4189B",
INIT_15 => X"9FE635BE11B7F0308D4A80092E0FC1FC662FA7E283FF68A8F0080AE1DDA8BE9F",
INIT_16 => X"12058312C1241140A056954AB0D680D000003350013024179498C2EC6B9270AE",
INIT_17 => X"2048120481204812048120481204812048120481204812048120481204812048",
INIT_18 => X"0481204812048120481204812048120481204812048120481204812048120481",
INIT_19 => X"2859400000000000000000120481204812048120481204812048120481204812",
INIT_1A => X"082218821390771C71C557C449F3898E09B56C74DAB16787E0760E5D1CF13043",
INIT_1B => X"7C3E1F0F87C3E082082082082082082082082082082082082082082082082082",
INIT_1C => X"87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F8",
INIT_1D => X"D7BD7400000000000000000000000000000000000000000000061007FE00000F",
INIT_1E => X"A2D1574005D0428A10A2AAA8BEF552EBDFFF557BC01FF5D7BFFEBA5D55555EF5",
INIT_1F => X"AFFFFC2000AA8428AAAFFAAA8BFF00002AA10FF802ABEFA2D16AA00F7FBE8A10",
INIT_20 => X"EFFF8002010002EAAAAAAAD1555FFFFAEA8B550051401450055575FF00517DEB",
INIT_21 => X"5FF0855575455D2AA8BFFA2D1575EF5D5555545FFFBE8A00087FC20BA5D2A975",
INIT_22 => X"8A00FFAE800AA082A820005D2E974BAA2D140145A2842AA00A284021FF5D0415",
INIT_23 => X"7FFEF000017400FFD1555FF007FFFEBA55042AA00000017400FFAABFEBAFF802",
INIT_24 => X"000155F7D540000F7FBFFE105D7BE8ABAA284000105D0428BFFA2FBFDFFFA2D1",
INIT_25 => X"7BFAEBA5551501D51C5FC7E00000000000000000000000000000000000000000",
INIT_26 => X"6D16AA28EBF5EDA38AADE1543849557D492BF8E2DE00552EBFFC7552BC01D75D",
INIT_27 => X"A85400E00E38A175FDE3F5C002DAAD42DAAAF784AFA82BC042DF47E3D1F8028B",
INIT_28 => X"50021C0092490E904BAFFD550A90FFA495FC7A05B555C257AAA8B45007540000",
INIT_29 => X"02402ABD4AD1D0E175D7140B455D516A1EAB45E2A000B4748717A095F571EAA1",
INIT_2A => X"4A8BC0ABFF7D03A17D1D5147540B454AA080038E9748542AE3D0051C7B6F02DA",
INIT_2B => X"D4B8FC7BFFFD2168B68F57492F505FF5FA550490BFA482B420B8428A3DA85400",
INIT_2C => X"0000000000000000000016ABD554201543A1EDE9016D4AAB454AF400547ABFB6",
INIT_2D => X"EBDF55556BC35E7557FE8AB25D11415FD0151614000000000000000000000000",
INIT_2E => X"6CBEA41D7D3DECFAF7D43FABAAAD57DEBAAAFFD74AA04547EE18D680BE9A55D2",
INIT_2F => X"78228E5000EA422E10439C1FBCD282351BDAAF9C20AAAABCBEB1DFF803FC5959",
INIT_30 => X"284683ABBDD7DEAA100069C14B25495A00F38EBAC0E198B9760501805357547D",
INIT_31 => X"8FE6A755ED8EFEFE41B2D17EAF02552BC0545556BD61E501001DF5DD3EBA31E6",
INIT_32 => X"F922ACA8AB8283C8310FAB1588916D3861C0422C44082B52A81550A828141440",
INIT_33 => X"DBCD7D262E5AFAC4B6AADDD562AF57D7C369AF25495A23068A8301BA7FB95556",
INIT_34 => X"FE0000003FE0000003FE0000003FE0000003FE03D5789700282E9FEFB501EA5F",
INIT_35 => X"3FE0000003FE0000003FE0000003FE0000003FE0000003FE0000003FE0000003",
INIT_36 => X"00000000000000000000000000000000000000000000000000000003FE000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000020",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(0),        -- Port A data input
DOA(0)   => data_read_a_lo_256(0),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(0),        -- Port B data input
DOB(0)   => data_read_b_lo_256(0),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_1_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"212C001411984004084D000508C53810A03D1450E839B003342114428A000807",
INIT_01 => X"08000010400A0008010600000084004000400002000000000000000000140000",
INIT_02 => X"484DEBA0111800C004400D000000000028800001CC404E6008B4933336880010",
INIT_03 => X"650C00000848A0423183089008C604224200000100A200002C280810098C0001",
INIT_04 => X"00000004208B00200E010800006667BE7000102C00080000040012010000080C",
INIT_05 => X"0080000000002020600100208D04414000800000000200004800080000800200",
INIT_06 => X"0000CB008084001C481040080000006050402008080000800488000000020400",
INIT_07 => X"00C00843060C19E2300221036000004400208000400041034001042000000101",
INIT_08 => X"08000290248CC84E0801318000C45555087C60C182B1592FE26AD7B7F7A01118",
INIT_09 => X"D8000AA220480040050080085200001161020001202100008008611687A28000",
INIT_0A => X"2640440000000080081040000040208300041000008004104006840000B80004",
INIT_0B => X"78051112A80000840200202112800001010828008000000105400020082800A8",
INIT_0C => X"2358323483234832358323583234832340190AC191A52801000C1002020883C2",
INIT_0D => X"4417882F82C00181707044212080300001002102010244800400C80C80323183",
INIT_0E => X"0B92C000000000400001004200004010200810040802040080200284401C1C11",
INIT_0F => X"00000043C2016000000F03C00280030000000F03C00280030000004860C60C0C",
INIT_10 => X"03800000049C0000000F03C00280030000000F03C002800321080000BC2380C2",
INIT_11 => X"00007861E0180000002A9001A00000007C4380E00000001E002300000008D187",
INIT_12 => X"4C0C81200009480010280340000008082430A07C80600C000000900861001108",
INIT_13 => X"34400241186100004A500007B00FC000000000E4A402C001208C308000268800",
INIT_14 => X"C0001E0181C0C200000025A400A200812A4070380000000B2500098190240001",
INIT_15 => X"04A0002410A170300C4A800800000020E22400A200096828F008000000AA9002",
INIT_16 => X"0200820040041002000010080014000000002340002004118010C22861400008",
INIT_17 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_18 => X"0080200802008020080200802008020080200802008020080200802008020080",
INIT_19 => X"0A04000000000000000000020080200802008020080200802008020080200802",
INIT_1A => X"8AB2048634B03249249604C061028A46BABEFC54A08170062002340C7452B500",
INIT_1B => X"DD6EB75BADD6EAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA8A28A28A28A2",
INIT_1C => X"A5D2E974BA5D2E974BA5D2E974BA5D2E974BA5D2E974BA5D2E974BA5D6EB75BA",
INIT_1D => X"AAAAAA00000000000000000000000000000000000000000000181FFFFF00000B",
INIT_1E => X"5D7BE8ABA5D557DFEFFFD17FEBA00042AAAAFFFFFFE00FF843DF45FFAE95555A",
INIT_1F => X"F552A800AA5555575FFA2AE820BAFFAEBFF555500155EF552E975FFF7D168BEF",
INIT_20 => X"00A2FBEAABA5D55420AA00002AA00AAFBE8B55A280175455D002AA00A2AABDFE",
INIT_21 => X"5FFAA802AAAAFFAA801EF00517FFFFF7D56ABEF0004155550004154105D556AA",
INIT_22 => X"75FF08557DEBAA2FBEAAAA552E955EF5D0415410A2AE97545A2AE954BAF7FBD7",
INIT_23 => X"7DF55A2AEBDEAAFFFFC20AAFFFFFFFFFAAD5555FFFFAEAAB55A2D168B555D555",
INIT_24 => X"0000BAFFFBE8A00087FC20BA5D2A975EF5D0002010552E820AAFFD57FF55F7D1",
INIT_25 => X"8A38F45F7AA9217FA380AD400000000000000000000000000000000000000000",
INIT_26 => X"52E975EFFFDF68BFF557BEAA925551785D7BFD5EFE3F08002FA92EBA5FDE28FF",
INIT_27 => X"41017DE92BF8E3AA824924870BF5551555C7A28A821EFE3AABAE38005B575D75",
INIT_28 => X"8005A1041055716DB7DB6FBEFEA81C55D0A0516802AA28BEF5EDB7DAA8A15438",
INIT_29 => X"EF1C043FE28E3FBD55FFAADE2DAAAE3A5C51C71C042DF45A3D1D00281E8A1056",
INIT_2A => X"B45B47F6FB55A95555E90F78E17F52FEF5EDA82FD249057F080417492AAAFC7F",
INIT_2B => X"8AAAA95B7AF45FF8F7DFEDFFAFF8E005FAE92A3AE3DBFF57FA2DF555D257AAA8",
INIT_2C => X"000000000000000000000A8F571EAA150021C0092490E905FFFD0550BD75C5FF",
INIT_2D => X"43DE00A2C57DE08FFAAA8B55F7EE801F7F2849EE000000000000000000000000",
INIT_2E => X"AE29F067155543A15D2E955EFFFFBEABEF557FEAA10595169BED83D1EBCA8000",
INIT_2F => X"FD57DEEAAA15976EB0444BFEB086808A8E3082C954BA5D7DD6145AAAA821A6AA",
INIT_30 => X"FFD55D6107782001FF0812000A255D57FFBEF3B97EEAB2C40217B9778428ABAF",
INIT_31 => X"F003F17418AEE817B540D11CA80BAAFA825EFAABEBCA18FE803755D08079EB47",
INIT_32 => X"EBA2D757547D7862AF57ABFFCABE5553FD5FBEFE86353EFFFD03FE027500035F",
INIT_33 => X"1F70C6AA04537957D6FB4807FFFB45F7EFFDA58FF2AA88A0F3C5014018AC28BD",
INIT_34 => X"00000000000000000000000000000000000000B2DD7DEAA100069C14B25495A0",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000020",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(1),        -- Port A data input
DOA(0)   => data_read_a_lo_256(1),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(1),        -- Port B data input
DOB(0)   => data_read_b_lo_256(1),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_2_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10E44660018259B2843913100062C98004802322D3E030235201006009B2812",
INIT_01 => X"8005A188084900481C8024A542400340404000720885800802000906E4910204",
INIT_02 => X"5C010802020408040C640850AA055254090541A111240A104A0000000908B510",
INIT_03 => X"0C1101108800004481060A001204102802156020218808002440850008C80550",
INIT_04 => X"8840C08022050400482812C21C0804040968987810688899444090C10A124A69",
INIT_05 => X"4885109105400029210000010340086856B141212252142242A068A080106372",
INIT_06 => X"0082006020044004C240108005540A400440880000908281302852A6710AA420",
INIT_07 => X"08040860400008C022402502100AA00004404B5075460111044014002AAA2100",
INIT_08 => X"382A885244145048C860214020040505487C0800049000004220000110820204",
INIT_09 => X"88582833A24105145404D4694E710A832488C000002205C23600408C872A2A12",
INIT_0A => X"A211100D0828800A022025A81AE3048228002A7080012082C15C859D5073D520",
INIT_0B => X"3E00659A308809540009202A5820068019108A88B1D007285082002B10416820",
INIT_0C => X"1A0021A5021A1021A5021A1021A4021A0010C2010D010887470912171342A683",
INIT_0D => X"89180010084038220410042B2000715A0400200080623400380886086021A002",
INIT_0E => X"40000554015500481000300000C4480810000002040000000913000004C18402",
INIT_0F => X"00000001440002C052000400028000154052000400028000200501CCD28D206A",
INIT_10 => X"00000000048015405200040002800012C05200040002800014E0000100002000",
INIT_11 => X"00010008000000000002A0000D80060100004000000000180000294010240020",
INIT_12 => X"1011000000090000A310000881080102000A0000400000000000900002000684",
INIT_13 => X"204E008240000000483250000800000000000004E00007004120000000240A60",
INIT_14 => X"254000806000000000000560000942004110000000000000254C020220000001",
INIT_15 => X"00108840600002080200000000000020806000093000040000000000000B8000",
INIT_16 => X"008022200100000020A89068084D402120AAC005C00000000000000005408140",
INIT_17 => X"0802008020080601806018060180200802008020080601806018060180200802",
INIT_18 => X"8040080000800008000180401804018040080000800008060180601806018020",
INIT_19 => X"A2852F81F81F83F03F03F0018040180401804008000080000800018040180401",
INIT_1A => X"04609D21808205965965D64CC5B60040138D70C030B54284722B291C50C7D100",
INIT_1B => X"4A25128944A25041041041041041041041041041041041041041041041041041",
INIT_1C => X"44A25128944A25128944A25128944A25128944A25128944A25128944A2512894",
INIT_1D => X"055400000000000000000000000000000000000000000000001E1007FFE3F009",
INIT_1E => X"FF843DF45FFAEBDF55082A82155082AAAA10F7FFEAB455500175FF5D2A800100",
INIT_1F => X"F082ABDF455D7BD5545F7D5574BAFFD16AAAAA28428ABA000428AAA5D7FD7400",
INIT_20 => X"455D7BEAABA5D2A97545552E975FFFFD168AAA5D7BE8BFF5D557FFEFFFD16ABE",
INIT_21 => X"5555555555FFA2AE820BAFFFFEAABA5555554BA5D0417545F7D56AAAAAAFBEAB",
INIT_22 => X"AA00AAAEBDFFF08042AABA087BD54BA08043DEAAFF843FF5508517FF55552A95",
INIT_23 => X"82010AAD1401FF002EBFF45A2FBFDFEF00042AA00AAFBEAB5500003FF5500002",
INIT_24 => X"0000BA0004155550004154105D556AA00A2FBEAABA085542145082A800BA002A",
INIT_25 => X"00155FF552A87410007145400000000000000000000000000000000000000000",
INIT_26 => X"8002FABA4171D5400FF8A38F45F7AABA57D0000855FD1C2AAFA00EBA5E8B7D55",
INIT_27 => X"555178FD7BFD5FDFFA0020BFF78417BD5545F7F1554AAF7D16DABABFF57DE920",
INIT_28 => X"DFFDF6DAAAAAF1EFB6D417BEFA901C2E97F40552E975EFEBDF68ABA557BEAA92",
INIT_29 => X"7DA3FBD21C7492E9256D555B555C7A2ABC20AAE3AABAE38005B574AA49041756",
INIT_2A => X"B7D1E803AF6D400028E02AB8A3A012540E2AABABC75D043A00003FE10E3802DB",
INIT_2B => X"8B7D0AAA800AA147085000FFDA001C7B47BFABC7BFFF7AB4714042AA38BEF5ED",
INIT_2C => X"000000000000000000000821E8A10568005A1041055716DA38B6FBEFFEF1C0EB",
INIT_2D => X"EBDE00AAC16ABEF5500155EF552A954000855544000000000000000000000000",
INIT_2E => X"D57DE0AFAD1EBEB400043DEAA085555400FFAAAAB55F7AEA8BF77004147EF5D2",
INIT_2F => X"AFBEABAF557FEA8515951E8B4D83D1EBDFF082CBDFEF005756145FFD5574AAF7",
INIT_30 => X"5951550100004155EFF7FFFDE08AA557FFFF083FFCEB95104210405D2E955EFA",
INIT_31 => X"A002A3FE18AE803CBE7A3C014351082E951FF5D7FD6145AAAA820A2AAAD29E00",
INIT_32 => X"45550028ABAFFD17FFED01001FFEF5542ABEB2AA848AAA2552EA8ABA7551400A",
INIT_33 => X"EBAF3F95EEE95C00B7CF12AAA800BA551417105FFFFC21555556EAB4CD6D5EAD",
INIT_34 => X"00000000000000000000000000000000000000187782001FF0812000A255D57F",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000040",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(2),        -- Port A data input
DOA(0)   => data_read_a_lo_256(2),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(2),        -- Port B data input
DOB(0)   => data_read_b_lo_256(2),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_3_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"210C00A20020000108430020001600B815602110494074133520400E02B92206",
INIT_01 => X"A00C9BC048800168240442C99E004B61404040028804A0080A000D16A0990A08",
INIT_02 => X"4809A902031800444445089866E331352180D468B8200E600C0081110B80ACD0",
INIT_03 => X"6D0A60100C000142B1A30A040AC68428320006010A80881068A80D401C846330",
INIT_04 => X"482218076809C03B24841CD92CDD5A440209127847294C042640102107102D04",
INIT_05 => X"0583180353202129000104E40B04644B32A86D24014A0D204063297092000E34",
INIT_06 => X"0120D000808040181B5000A014CC662814442808805A52C03068280004629414",
INIT_07 => X"00444841428409C038B02523041994001C644C82732001190000B400E6640901",
INIT_08 => X"E8E64010248C4A5AA040308000440005487C285284B1D00BC22AC005B2820318",
INIT_09 => X"A8D588362040534C3B0E80A9DB742641620AC281826816925040408483008A10",
INIT_0A => X"040450A1439800840C32264119D004860110104004010001E732C0DF80F3B174",
INIT_0B => X"7C8575909088A4D010202422520090840B4028209AC1111954DA902230010002",
INIT_0C => X"032920329203692036920329203392036C900BC9019528100A0D30024BC8A283",
INIT_0D => X"446A101C05C0088A42D001032000333931001902010234888C68804808A03692",
INIT_0E => X"8601CCCC8B33004C0001004240140018380818040A0706009000028000903401",
INIT_0F => X"00000120000006000000000020004011000000000020004010072CC92416414C",
INIT_10 => X"0000001002001400000000002000401380000000002000401070000000000000",
INIT_11 => X"00000000000000000110000001A0000000000000000005002000244000000000",
INIT_12 => X"00000000010402049910000011000500000000000000000008000020000002C0",
INIT_13 => X"805500000000000820133000000000000000810000000C000000000004100B20",
INIT_14 => X"0530000000000000000180000011060000000000000001040154000000000020",
INIT_15 => X"0000820062000000000000000000040100000010700000000000000002400000",
INIT_16 => X"0680C2A05104100280A8D06C004044230B998021002004000001011000380000",
INIT_17 => X"280C0280C0280803808038080380803808038080380C0280C0280C0280C0280C",
INIT_18 => X"00C0280E0200C0280E030080380A030080380A030080380C0280C0280C0280C0",
INIT_19 => X"8A145D54AAB556AA9556AA830080380A030080380A030080380A0200C0280E02",
INIT_1A => X"04A20E858000049249240540430303C0C78C706428A141046016224C58629502",
INIT_1B => X"EA753A9D4EA75249249249249249249249249249249249249249041041041041",
INIT_1C => X"46A351A8D46A351A8D46A351A8D46A351A8D46A351A8D46A351A8D46A753A9D4",
INIT_1D => X"A8400000000000000000000000000000000000000000000000001007FEB6FECD",
INIT_1E => X"5500175FF5D2AA8A10005540155087BEABFF552ABDF45A2D16AAAAF7D540000A",
INIT_1F => X"000556AB55552ABDE00AAD140010F7D17FF45A2AA82155082AAAA10F7FFEAB45",
INIT_20 => X"55557FEAA10007FEAABA000428AAA557FD7400FF843DE00FFAEBFF55082A8201",
INIT_21 => X"A105D7BD5545F7D5574BAFF802AA00A2D168ABA085568BEFFFAE820000855421",
INIT_22 => X"FFEFF7D56ABEF557BD74BAFF8402145A2AEBFFEF552EAAABA5D0028BEF082AA8",
INIT_23 => X"3DEAAAAAA95410F7803FFFF55556AAAA552A975FFFFD16AAAA5D7BC01EF5D557",
INIT_24 => X"0000105D0417545F7D56AAAAAAFBEAB455D7BEAABA5D2A974005D55574005504",
INIT_25 => X"DF6FABAFFD547010AA8407400000000000000000000000000000000000000000",
INIT_26 => X"C2AAFA28EBF5E8B7D5500155FF552AAF0100071455451C75EABC74174BAF55B6",
INIT_27 => X"F7AABAF7D00009543D1C556AB6D4124BAE10BED542010FFD57AF55AAF5D756D1",
INIT_28 => X"FEBA0870281C5F4716D5D7FEDA3A0955FF48208002FABA4171D5400FF8A38F45",
INIT_29 => X"BA15203FFFF002AAFA384171D5545F7D0154AAF7D16DABABFF57DE92005F6ABF",
INIT_2A => X"ABA417BC01D7555178FD7BFD5FDF571575D24BA438E021D5B6A4BAFFF5D2EB8E",
INIT_2B => X"FE005D5B52428410E3AE92E3A490410EB843ABD71551FFE02552A975FFEBDF68",
INIT_2C => X"0000000000000000000003849041756DFFDF6DAAAAAF1EFB6D417BEFBD71C24B",
INIT_2D => X"56AB45081028B55FFFFFFEBAFFD557400A280144000000000000000000000000",
INIT_2E => X"D56ABF5AAD15455F5D2EBDEAAA2D16ABEF5500175EF552ABDE000855545455D5",
INIT_2F => X"85555400FFAAAAB14F7AE28BF77004146BA557DEABEF00002BE10FFD540000FF",
INIT_30 => X"F2D1EAEBA007FEABEFAA84174BA557FD55EF5D3BFEEB35055DEE1000043DEAA0",
INIT_31 => X"5FFAA28BF7592EABE0A0804ABFFB082EBDEAA005556145FFD5574AAF7D47DE0A",
INIT_32 => X"105D2E955EFAAFBE8AAA547FE21550853E8B4FABD5EBFF75D55420AA82AA8015",
INIT_33 => X"FFF087FFCEF90104B780A557FC20AA082AAAE10AA8000000A2AC2ABFD2151EB8",
INIT_34 => X"00000000000000000000000000000000000000AA0004155EFF7FFFDE08AA557F",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000020",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(3),        -- Port A data input
DOA(0)   => data_read_a_lo_256(3),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(3),        -- Port B data input
DOB(0)   => data_read_b_lo_256(3),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_4_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10804002061080A284201081034809800A00230350007833422C82904204006",
INIT_01 => X"204398001038084C0420050E12100368403008418984014902030906A0910204",
INIT_02 => X"480108A000000000446118E01E80F00A41043118680402000800000009882390",
INIT_03 => X"065140108C0000400026480000009120270072E03000000030808840888100F0",
INIT_04 => X"9100EB826A155C1AF0B81C160033B9440222BA281AE0D8B8E02010E81C22E821",
INIT_05 => X"5C0F20B36F08010924C084C501441C4CF21C48B133483C8042EAE1E0101074C4",
INIT_06 => X"010290102005118043508020543C1E480002820085D9C0C70000F2AA375A6071",
INIT_07 => X"00000860008008D200102502000786000C00C8025C00091B0400B00061F84020",
INIT_08 => X"991E02100C84C0480020010000004404087C8010009800004022800110000000",
INIT_09 => X"B83D6A2620418F7CF8084082425D01D123C2C040816A00708840408483000011",
INIT_0A => X"BB1B585C1304E002000064010E4007F7210010500400400800F0CC249C1401C1",
INIT_0B => X"7A04331814080458100134201A2086441B50A088078106C14540906D004068A0",
INIT_0C => X"186921829218692182921829218692182090D3490C352296CC60B11357088682",
INIT_0D => X"411050002500A9200A8014010001370F03080980912204883C28864860A18A92",
INIT_0E => X"C40903C1430F20025040102200441A040906008300418050501341208002A005",
INIT_0F => X"0000012004000BC01200000020004008C012000000200040000721CD86146108",
INIT_10 => X"0000001002000A40120000002000400DC01200000020004004D4400000000000",
INIT_11 => X"40000000000000000110200007600401000000000000050020005D4010040000",
INIT_12 => X"1010000001040004A3B000018008850200080000000000000800002002000650",
INIT_13 => X"80360082000000082034300000000000000081004000170041000000041005E0",
INIT_14 => X"2B200080400000000001804000192000401000000000010400F8020200000020",
INIT_15 => X"00114A00200002080000000000000401004000085C0000000000000002410000",
INIT_16 => X"459040281181004A8088986D045C24436C7840A6180300082001211304208140",
INIT_17 => X"1106409004110240904411024090040106419004010640900411064090440102",
INIT_18 => X"9024010041104409024190240104411004190240906411024190440102419004",
INIT_19 => X"021074B261934D964C3269C09064110040104409064190240104401004190640",
INIT_1A => X"8A74C1323433345145130282E6228A063807E05000143842130115063450454A",
INIT_1B => X"8D46A351A8D46AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA8A28A28A28A2",
INIT_1C => X"A0D068341A0D068341A0D068341A0D068341A0D068341A0D068341A0D46A351A",
INIT_1D => X"50015400000000000000000000000000000000000000000000001007FEA73FC1",
INIT_1E => X"A2D16AAAAF7D568A00AA8400000AAFFC21FFF7D542000FFAE821FF552EAAA105",
INIT_1F => X"0AAAE820BA550015400087FD74BAFFD540000F7D155555087BEABFF552ABDF45",
INIT_20 => X"AAF78015545FFD555555082AAAA10F7FFEAB455500175FF5D2AAAA1000554000",
INIT_21 => X"B45552ABDE00AAD140010F7D17FF45A2FBC2000A2FFC21555551554005D2EA8A",
INIT_22 => X"FF55082E82145A280001EFF78402145A2AE801555D2E95555552E9741000556A",
INIT_23 => X"7DF45557BD5410F7D555545F7AA97410000428AAA557FD5400FF843DE00FFAEB",
INIT_24 => X"0000AA085568BEFFFAE82000085542155557FEAA10007FEABEFAAD1400AA5D51",
INIT_25 => X"AA801EF4920AFA10490A17000000000000000000000000000000000000000000",
INIT_26 => X"C75EABEF4124BAF55B6DF6FABAFFD56F010AA8407428A2F1C01FFF7D142028EB",
INIT_27 => X"552AAFA10007155428A2AE850925D0010400087FD24AAE3DF47010E38E051451",
INIT_28 => X"55D51524004920ADA82EB8A12555EBFB4717D1C2AAFA28EBF5E8B7D5500155FF",
INIT_29 => X"55492A850381C5F6AB6D4124BAE10BED542010FFD57AF55AAF5D7410A2FBC015",
INIT_2A => X"400FF8A38E00F7AABAF7D0000955FDB684051D7F7840517DA2A4871554124925",
INIT_2B => X"75EFBED5400825D557FF55007BD7410EBDB5017DE38E8708008002FAAA4171D5",
INIT_2C => X"00000000000000000000082005F6ABFFEBA0870281C5F4716D5D7FEDB7D0955D",
INIT_2D => X"1401FFFFD5420BAA2AA821FF08043DE10002A964000000000000000000000000",
INIT_2E => X"FBD7410A2AE965555D556ABEF080028B55FFFFFDEBAFFD57FE00A280144BAAAD",
INIT_2F => X"2D16ABEF5500175EF552ABDE000855544AAAA82174105D0402000087FC00BAA2",
INIT_30 => X"AAD154400AAFBC015555554001008003FE00AAEA81154AAFFD65FF5D2EBDEAAA",
INIT_31 => X"FA2AA155550004021E5582A964BE557FEABEF00002BE10FFD540000FFD56ABF5",
INIT_32 => X"1000043DEAA085555400FFAAAAA10F7AC28BF558001454DF78017555F780175E",
INIT_33 => X"5EF5D7BFEEF35055487EFF7D1400105D517FF55087FD7410A2FBC01E7F2AE966",
INIT_34 => X"0000000000000000000000000000000000000010007FEABEFAA84174BA557FD5",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000040",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(4),        -- Port A data input
DOA(0)   => data_read_a_lo_256(4),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(4),        -- Port B data input
DOB(0)   => data_read_b_lo_256(4),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_5_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50DB4A0791B1B4B694369283C81F9996A091832102004AB37B20E07C0C1E006",
INIT_01 => X"285FBC448000804C446A00000034824841280A00084000C8C212892EE2953235",
INIT_02 => X"C809AD5CB118E640A4D118FC011FF0002080000082C8C66609DB7DDDCB1F2036",
INIT_03 => X"250907263A4C90D210A35C82484285720B20648A88800000B8E0F850A8C4500E",
INIT_04 => X"4005122126899100064D20001044429C78243A2C0436C887198AB916E0551A24",
INIT_05 => X"A370C14CA0E900004048002389CFE2F20F7D7A314CB5C20AE51437E044948912",
INIT_06 => X"90184D150505A1D84B7E2A285401412870B20A51842404C44437118630839B88",
INIT_07 => X"E640A94D1AB469D6300E2FFFAA7F8A4D23248130E259C903FBC403A9601A62E8",
INIT_08 => X"0A7E3016250D49CA3F83108186400000EBFD235488B9749BC1AAF325B35CB118",
INIT_09 => X"9B020B7E6AE46082032004904200C03DBC3BCA4860270BFA829968040B0800AC",
INIT_0A => X"22181A2B9203642840124098516CE0C3D825124111A79F802800F20DB4D6DA34",
INIT_0B => X"6824911331CA84D346A964F0125CD7AB1938A00AEFDD567DE480116848C9426A",
INIT_0C => X"01AD7016D701ED7012D701ED7016D701AAB8096B80F5A21828041846620F5AB8",
INIT_0D => X"847B053F48A8308A644A412BCA8470FF0209019081C706EABDAAC0DC0AF012D7",
INIT_0E => X"2194FFC044FF84B08FC862A2CD8F0A89014080A2425422151870500544991292",
INIT_0F => X"038ABBCBC7C7802F86FF87C002F87F002F86FF87C002F87F2000804821021004",
INIT_10 => X"0380230F2FFC002F94FF87C002F87F002F94FF87C002F87F2201BFFEBC2BA0C2",
INIT_11 => X"BFFE7C69E01804E1E7EABE3F000FF97D7C4BC0E008C7C3FE58FC029FEF5CD9A7",
INIT_12 => X"EC9C8120C4DFC802808B2EB22E777ADDE6F8A47CC0600C2683E0FFAAE3F1F001",
INIT_13 => X"FC14DFC5186104C6FE5037FFF00FC0000FC0FEE487A7066FA38C3082637F83BD",
INIT_14 => X"072FFF41C1C0C2038A7CED87A7D109FBBA5070380131CBFB2477BF919024189B",
INIT_15 => X"9F46DFBEB1B7F0380C4A80092E0FC1FDE607A7C077FFE828F0080AE1DFAA1E9F",
INIT_16 => X"5594254A10A03446128898494C09402081F83200A9442217159880640942320E",
INIT_17 => X"1940509465014251140519445094251142511445094451942511425014451940",
INIT_18 => X"9405094450944511425114650146501425194450944509405194250146501405",
INIT_19 => X"0A983124B2DA6924965B4D509445094051940501465014251142501465094451",
INIT_1A => X"BE5FDFF3F7F773CF3CF7D79FA8F5BB4E7F7B9DB7FF3A7E0FF4807F1B6DB7ED43",
INIT_1B => X"F77BBDDEEF77BBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEF",
INIT_1C => X"EF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEE",
INIT_1D => X"FFBFFE00000000000000000000000000000000000000000000001007FE1BFB5E",
INIT_1E => X"FFAE821FF552E820105500155555D2AA8A00AA843FFFFF78002155AAAE974AAF",
INIT_1F => X"0FFAE80000AAAE974BAFFAEAAB45AAAEBDEAAA2FFEAA00AAFFC21FFF7D542000",
INIT_20 => X"000055574BA557FFFF55087BEABFF552ABDF45A2D16AAAAF7D56AA00AA840000",
INIT_21 => X"0BA550015400087FD74BAFFD540000F780155555D7BE8B45085168BFFA2D17FE",
INIT_22 => X"AA10005140145FFFBC01EFAAFFD75FF002E97555A2AABDEAAAAAAAAA00AAAE82",
INIT_23 => X"174BA5D043FF45AAAA974AAF7AEBFF55082AAAA10F7FFEAB455500175FF5D2AA",
INIT_24 => X"000000A2FFC21555551554005D2EA8AAAF78015545FFD555410552EA8BEFAA84",
INIT_25 => X"8E0217DBEA4954AAE3FBFDE00000000000000000000000000000000000000000",
INIT_26 => X"2F1C01D7F7D142028EBAA801EF492087A10490A171455D2EADA28B6803FFFFFF",
INIT_27 => X"FFD56FA10AA8417428E3AE87010A2A4974AAE3AEAFB6DAAA4BDEAAA2F1EDA28A",
INIT_28 => X"D14516DBD7BEDB7DE381451554AA497FFFF451C75EABEF4124BAF55B6DF6FABA",
INIT_29 => X"AAAAA0AFA28A2A4850925D0010400087FD24AAE3DF47010E38E0516D5D7BE8B6",
INIT_2A => X"B7D5500155FF552AAFA10007155545F7F1C21D7AAF1D55FF082A9057DA2AABDE",
INIT_2B => X"70384124ADBFFBE84174AA55043FF6DBEAE950AAEB8ABDF7D1C2AAFA28EBF5E8",
INIT_2C => X"00000000000000000000010A2FBC01555D51524004920ADA82EB8A12410EBFB4",
INIT_2D => X"EBFEBAF7843DFEFF7AE801EFF780174AAAAFBFEE000000000000000000000000",
INIT_2E => X"803FEBAAAD17CEAAAAD140155FFD5420BAA2AA821FF080415410002A96555552",
INIT_2F => X"80028B55FFFFFDEBAFFD57FE00A280144AAA2AA97400A280174AAA2AEBDFEFA2",
INIT_30 => X"A2AE965FF557FE8BFF55557FF55FFFBFFEAA5D51554AA087BFEF555D556ABEF0",
INIT_31 => X"F0004821FFAAAEBDEAAAA843CEAAAA80174105D0402000087FC00BAA2FBD7410",
INIT_32 => X"FF5D2EBDEAAA2D16ABEF5500175EF552ABDE00005554545F7D140145A2D5555F",
INIT_33 => X"E00AAAA81114AAFFD64BA00043FFFFFF80174AA55043DFFFFFAE974BAA2AEBEF",
INIT_34 => X"0000000000000000000000000000000000000000AAFBC015555554001008003F",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000180",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(5),        -- Port A data input
DOA(0)   => data_read_a_lo_256(5),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(5),        -- Port B data input
DOB(0)   => data_read_b_lo_256(5),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_6_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10804B0061A010A2840012C030028180004003220200403302301C0381A0086",
INIT_01 => X"870041CA3839684D18A160000C52424841000000090800090210010008110204",
INIT_02 => X"080108200C1000004464480400C0080100000000010432400800800009882050",
INIT_03 => X"040001008C2340D0840208624210002182800584488000103080010E08C10000",
INIT_04 => X"00101611A029B08410044800000000040088102A440814040400900500001800",
INIT_05 => X"02800000400C820934E4A0002900404400820004000A00824004085011200A00",
INIT_06 => X"2210001A12100830434040870BFE004044420322C00812900308010000829400",
INIT_07 => X"00000860400108C22000A103090074120044800040001103005180911FE0C134",
INIT_08 => X"FD01C0120484C0580020C10000000000087C0800209100004228000110000C10",
INIT_09 => X"88FC08362240404100228080D200DFC1610200E40AA050000040D0C463008083",
INIT_0A => X"29561B22D77C720D2522400000400882091210008440005F8BF4C00002900004",
INIT_0B => X"7E25D11A200024541100342A5A2886285502A880C00107FD355E022005026BCA",
INIT_0C => X"D8282D8A82D8A82D8682D8682D8E82D8A016C1416C15A01D68209A127208A6B1",
INIT_0D => X"807888180A80910A1460150900013400410CB5C9D96236883460B60B602D8282",
INIT_0E => X"0062003C10002442006429124290034E85A742D1A368D0DA2004696884851806",
INIT_0F => X"000000157000604050000000028000D04050000000028000CE80004C00000000",
INIT_10 => X"000000000483D04042000000028000D04042000000028000C508000100000000",
INIT_11 => X"000100000000000000078000A40006000000000000000019A003080010200000",
INIT_12 => X"1001000000093490308001408000000200020000000000000000900518000508",
INIT_13 => X"23490002400000004993C000080000000000001FC000C8804020000000246800",
INIT_14 => X"C05000802000000000001740002256004100000000000000FD00000220000001",
INIT_15 => X"00A000404A000200020000000000002099C000330000040000000000001F0000",
INIT_16 => X"68DA308D09D0804880089A49461032040C07C1440C8190800020530865400540",
INIT_17 => X"9DA7695A1685A369DA7685A168DA369DA5685A168DA7695A5685A368DA7695A5",
INIT_18 => X"5A168DA7695A168DA1695A769DA1685A3695A569DA3685A169DA769DA1685A16",
INIT_19 => X"00046638C31C71C718638E68DA7695A568DA3685A769DA5685A368DA569DA368",
INIT_1A => X"8E76DDB3B7B377DF7DF7D7CEE7F78BCE7F8FF0F4FA957FC7F37F3F5F7CF7F108",
INIT_1B => X"7F3F9FCFE7F3F8E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E3",
INIT_1C => X"E7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE",
INIT_1D => X"AAABFE00000000000000000000000000000000000000000000181007FFDE534F",
INIT_1E => X"F78002155AAAE974AAFFFBFFE10F7FBE8BEF552E95555552EAABEF082E975EFA",
INIT_1F => X"0A2AAAAA10087FC01EF552EAAB45F7AE821550851555555D2AA8A00AA843FFFF",
INIT_20 => X"EFA2AEBDFFF552AAAA00AAFFC21FFF7D542000FFAE821FF552E8001055001541",
INIT_21 => X"000AAAE974BAFFAEAAB45AAAEBDEAAA2FFEAB45552E800AA555568A105D002AB",
INIT_22 => X"AA00AA8400000007BC21FFAA803FFEF5551420105D5568B45FF8400000FFAE80",
INIT_23 => X"C2155007FC20BAA2D5575FF087FFFF55087BEABFF552ABDF45A2D16AAAAF7D56",
INIT_24 => X"0001555D7BE8B45085168BFFA2D17FE000055574BA557FFFE10F7AAA8A00F7FB",
INIT_25 => X"24ADBD70820975FFA2A4BFE00000000000000000000000000000000000000000",
INIT_26 => X"D2EADA28B6803FFFFFF8E0217DBEA4954AAE3FBFDE38F7FFEABFF412A9056D49",
INIT_27 => X"492087010490A07038B6A0AFA38007BC51EF4920AFB55EBA4851450855555455",
INIT_28 => X"2555F68A3855002FBC7BEA4BFFFF492EADA28A2F1C01D7F7D142028EBAA801EF",
INIT_29 => X"45E38A07028E3AE87010A2A4974AAE3AEAFB6DAAA4BDEAAA2F1EDB55492A8508",
INIT_2A => X"F55B6DF6FABAFFD56FA10AA84174381C7FC01C7B68E3DFC75555400105D516DB",
INIT_2B => X"FE38F7A0AFA38E3FFC21450071C2092A2D5571FF0851FDF451C75EABEF4124BA",
INIT_2C => X"0000000000000000000016D5D7BE8B6D14516DBD7BEDB7DE381451554AA497FF",
INIT_2D => X"BEABEF002E801EF00003FF550800155FFA2803CE000000000000000000000000",
INIT_2E => X"8417555085154555552EBFEBAF7843DFEFF7AE801EFF780174AAAAFBFEEAAF7F",
INIT_2F => X"FD5420BAA2AA821FF080415410002A964AAFF803DEAA087FD55FF00043DF45A2",
INIT_30 => X"AAD17CF55002E95410557BEAABA55043DF55F7803FFEF002ABEEAAAAD140155F",
INIT_31 => X"55D51420105D517DF55AAAA964AAA2AA97400A280174AAA2AEBDFEFA2803FEBA",
INIT_32 => X"555D556ABEF080028B55FFFFFDEBAFFD57FE00A280144BA5D7FC2155FFAABDF4",
INIT_33 => X"EAA5D51554AA087BFEEAAF7803DEAAAAFBC0155085540000A2D5575FF08517CF",
INIT_34 => X"00000000000000000000000000000000000001FF557FE8BFF55557FF55FFFBFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000120",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(6),        -- Port A data input
DOA(0)   => data_read_a_lo_256(6),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(6),        -- Port B data input
DOB(0)   => data_read_b_lo_256(6),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_7_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10804B00482010A2842012C024500188000003000000003302300C018180002",
INIT_01 => X"0200084020084048040080000201024040000000080000080200010008110204",
INIT_02 => X"4801082248100000444008000080000041000000002222400800000009008010",
INIT_03 => X"0401008108A1444000020A400000002902006400088000003080040408C10000",
INIT_04 => X"0000100022418000000C80C00400000400201839040000050001140400201820",
INIT_05 => X"02000000400041092C80C0214144004400000000000800045004000020220800",
INIT_06 => X"0000300000000830435150020003004060000000080800801100000030829001",
INIT_07 => X"00000840000008C02000A503010002928040800062481919047140D40008C000",
INIT_08 => X"0A0002120484C0580850810000000000487C000000910000402A800110024810",
INIT_09 => X"8802083624504000022680A1DA20800164000400112284000004D404022A8800",
INIT_0A => X"30014050280040180020400011640CC72E029000084800503004C40100D21024",
INIT_0B => X"3801078228010454210028240082200081140800900220000000002011440009",
INIT_0C => X"40022400224002240822408224082240C1120211202008900800100242428280",
INIT_0D => X"807802988294900A00451109006230006E000800001280110050902901240022",
INIT_0E => X"0042C000C0002000000020020490000400020001020080401010813094801146",
INIT_0F => X"807144102420700052000003C00780B00052000003C007808450484C00000000",
INIT_10 => X"2C0E00E0D003300052000003C00780B00052000003C00780890800010000130C",
INIT_11 => X"000100000661801E18042100E000060100000B03803838012403800010240000",
INIT_12 => X"10111848322020512000414400000002000A1001058300C0741C005412080908",
INIT_13 => X"029F008240864231013BF00008000C3C003F00184040EF8041204321188053E0",
INIT_14 => X"F770008060130C8071821040403F5600411004C2600E3400C27C020223090644",
INIT_15 => X"00B8CA406A0002C812240B0201F038021140403F740004010472041E20110100",
INIT_16 => X"0080228011010042802890484040000008004945000100008844430060198941",
INIT_17 => X"0000000000000600802008020000400000000000080200802008000000000000",
INIT_18 => X"8020100000000008020080000000000020080200000000040080200802008060",
INIT_19 => X"0A14584104000208208000018020080200000010020080200800010000080200",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000442",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"82AAAA00000000000000000000000000000000000000000000001007FEBC3240",
INIT_1E => X"552EAABEF082E975EFAAAABFFEF002ABDF555D5157555F7FBC00AAAAD5400BA0",
INIT_1F => X"AAAAABDF55FFFBFDF55555568ABAAAD5401FF5D2AAAA10F7FBE8BEF552E95555",
INIT_20 => X"005D55554105D51401555D2AA8A00AA843FFFFF78002155AAAE974AAFFFBFFEA",
INIT_21 => X"A10087FC01EF552EAAB45F7AE821550851554AAF7FBFFEAA007BFFFEFF7D5400",
INIT_22 => X"00105500155EF5D2EBFF450000020AA5D7BC0000F7D555545A28000010A2AAAA",
INIT_23 => X"A8A10FFD568ABAA2D56AAAAF7AABFE00AAFFC21FFF7D542000FFAE821FF552E8",
INIT_24 => X"000145552E800AA555568A105D002ABEFA2AEBDFFF552AAAABAA2AE95555FFAA",
INIT_25 => X"F5C20BAAAD5420821C2EAAA00000000000000000000000000000000000000000",
INIT_26 => X"7FFEABFF412A9056D4924ADBD70820975FFA2A4BFFFF1C2EB8F45555550545E3",
INIT_27 => X"BEA4954AAE3FBFDE82B6AEBAF55E3FFFAF55555F6FA92BED5421C75D20AAA38F",
INIT_28 => X"20075FDFD7F7D5400385D51504385D55401455D2EADA28B6803FFFFFF8E0217D",
INIT_29 => X"7DB68E02038B6A0AFA38007BC51EF4920AFB55EBA485145085555492F7F5FFE9",
INIT_2A => X"028EBAA801EF492087010490A071EF4920B8F45140E07082417BC2000EBD5505",
INIT_2B => X"DA92A2A09257DE3A4AAA10F7D16FAAABED56AE82F780BAE28A2F1C01D7F7D142",
INIT_2C => X"00000000000000000000155492A85082555F68A3855002FBC7BEA4BFFFF492EA",
INIT_2D => X"EAAB455D5142155AAD1400AAA2D1420005D2EA9A000000000000000000000000",
INIT_2E => X"D1421555D042BAAAF7FBEABEF002E801EF00003FF550800155FFA2803CFFF552",
INIT_2F => X"7843DFEFF7AE801EFF780174AAAAFBFEE00F7AAAAB55AAFBEAB555D7BFDE00F7",
INIT_30 => X"085154400FFD17FE1000517FF55FFD5420BA5D55400BA555543155552EBFEBAF",
INIT_31 => X"0087BC0000A2D5421EFF7AE810AAFF803DEAA087FD55FF00043DF45A28417555",
INIT_32 => X"AAAAD140155FFD5420BAA2AA821FF080415410002A965FF080428B45552A9540",
INIT_33 => X"F55F7803FFEF002ABEE00A280001FFA28028A00FFD17DEAAF7D56AA10FF842BA",
INIT_34 => X"0000000000000000000000000000000000000155002E95410557BEAABA55043D",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"FFFFFFFE00000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000000000000000000001F",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(7),        -- Port A data input
DOA(0)   => data_read_a_lo_256(7),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(7),        -- Port B data input
DOB(0)   => data_read_b_lo_256(7),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_8_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10004B00000400E2840012C0000001800000070000000033022000000000082",
INIT_01 => X"000009C0183808481C0160000E02424040000000180800080200010048110204",
INIT_02 => X"080108000090000004400C000080000051000000000002400800000009000010",
INIT_03 => X"0000000004300840000200000000000002800504488000103080880008800000",
INIT_04 => X"00009410A028A084000440C00400000400001032040800150400008500221800",
INIT_05 => X"4280008040048A09302420202804400400800010200A00000204080011014A00",
INIT_06 => X"2B02000A32114192434010001FFC004240428122000800000008012000821400",
INIT_07 => X"00000840000008402001A50200000630404080006248381B000080837FF88114",
INIT_08 => X"0A000210040440480000090000000000087C0000009100000002000110000090",
INIT_09 => X"08020A322000400102260021DA2080114502002409A04400004282C4E1228800",
INIT_0A => X"904A4522920052012120400011641C4601005000041100002004800100C21024",
INIT_0B => X"78051792A8000454104020001280008845022000900000010444000000020009",
INIT_0C => X"000000000000000000000000000000000800040000452A9008001002424A8002",
INIT_0D => X"807880508202100A1000810B2020340041248548490004800400000008000800",
INIT_0E => X"20020000C000044214240932000001428CA14650A128508A2004284024840022",
INIT_0F => X"80000000001020404000783FC0000010404000783FC000000880084C01041008",
INIT_10 => X"FC7E0000000010404000783FC0000010404000783FC000000500000103D45F3D",
INIT_11 => X"000103961FE78000000000402400020003B43F1F800000002201080000202658",
INIT_12 => X"01617CD8000000803000804080000020090659833F9F03C00000000000040500",
INIT_13 => X"00400018639EC000000000000FE03FFC00000000400840000C31CF6000000800",
INIT_14 => X"4000001E2A3F3D80000000400802000401AA8FC7E00000000100002C2F5B0000",
INIT_15 => X"4020000104480DC372B47F060000000000400802000017570FF6000000010020",
INIT_16 => X"28CA30051851A0C0002890484600320408004444048090800022130864000540",
INIT_17 => X"84A1284A1284A328CA328CA328CA328CA328CA3284A1284A1284A1284A1284A1",
INIT_18 => X"CA328CA328CA3284A1284A1284A1284A328CA328CA328CA3284A1284A1284A12",
INIT_19 => X"080440000000000000000028CA328CA328CA328CA1284A1284A1284A128CA328",
INIT_1A => X"9EDFC8F33637D6CB6CB2900DA6128A0A543EBC57A10A244257C5051E75D64108",
INIT_1B => X"1F0F87C3E1F0F9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7",
INIT_1C => X"E1F4F87D3E1F4F87D3E1F4F87D3E1F4F87D3E1F4F87D3E1F4F87D3E1F0F87C3E",
INIT_1D => X"02ABFE00000000000000000000000000000000000000000000001007FE8A8913",
INIT_1E => X"F7FBC00AAAAD5400BA082AAAA10000000010F7D5421EF007BC01FF5D7FFFE100",
INIT_1F => X"A5551554AAFF80021EF002A820BAFF8428A00A2AAAABEF002ABDF555D5157555",
INIT_20 => X"EFFFFFEAB55002ABFE10F7FBE8BEF552E95555552EAABEF082E975EFAAAABFEA",
INIT_21 => X"F55FFFBFDF55555568ABAAAD5401FF5D2AAAB55FFD1400AA5D7FC01EFA2FFE8B",
INIT_22 => X"74AAFFFBFFEAA08001555555516ABEFA280020AA5D043DF55557BEAAAAAAAABD",
INIT_23 => X"2AB55005140145AAFFE8AAAF7D1401555D2AA8A00AA843FFFFF78002155AAAE9",
INIT_24 => X"0000AAF7FBFFEAA007BFFFEFF7D5400005D55554105D51400005551421EF0804",
INIT_25 => X"7FC21EF5D75FFE10142EBAE00000000000000000000000000000000000000000",
INIT_26 => X"C2EB8F45555550545E3F5C20BAAAD5420821C2EAAA101C0005000E3D1401D71C",
INIT_27 => X"0820975FFA2A4BFE925D51554AAE384001FF142E800AAFF802AA28AAAEAFBFF1",
INIT_28 => X"2557BC21D7BEF5EDBC7FFF1EFB6D1420BAE38F7FFEABFF412A9056D4924ADBD7",
INIT_29 => X"55417BEDA82B6AEBAF55E3FFFAF55555F6FA92BED5421C75D20AAB45F7D14709",
INIT_2A => X"FFFFF8E0217DBEA4954AAE3FBFDEAA1C001056D415F6ABEFA2840208249043AF",
INIT_2B => X"00385D51401EF00002FB45085F4016DAAF1EDAAAFFFB401455D2EADA28B6803F",
INIT_2C => X"00000000000000000000092F7F5FFE920075FDFD7F7D5400385D51504385D554",
INIT_2D => X"417410AAD540155557FC01EF5D557DE105D2AA8A000000000000000000000000",
INIT_2E => X"842AABAA2AEBDFFF552EAAB455D5142155AAD1400AAA2D1420005D2EA9A105D0",
INIT_2F => X"02E801EF00003FF550800155FFA2803CE105D55574BAA280021EF5D2E820BAF7",
INIT_30 => X"5D042BB45FFD157410557FC0155F7D57FF55F7D57FFEF550028AAAF7FBEABEF0",
INIT_31 => X"FAA8000000080428B55087FFFE00F7AAAAB55AAFBEAB555D7BFDE00F7D142155",
INIT_32 => X"55552EBFEBAF7843DFEFF7AE801EFF780174AAAAFBFEEBA5D04021EF087BE8BF",
INIT_33 => X"0BA5D55400BA5555430BA5555421EF00043FF45007BC21FFA2D57FEBAF7FBC21",
INIT_34 => X"0000000000000000000000000000000000000000FFD17FE1000517FF55FFD542",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000080",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(8),        -- Port A data input
DOA(0)   => data_read_a_lo_256(8),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(8),        -- Port B data input
DOB(0)   => data_read_b_lo_256(8),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_9_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10004B00018000A2840012C0000281800000030000000033022000000000006",
INIT_01 => X"000008000000004C0020000000100268413C0A61590001D90213C10008110204",
INIT_02 => X"680108200010000054400C000080000041000000010002400800800009082011",
INIT_03 => X"0004000000002040000200100000000042800584488000103081880008800000",
INIT_04 => X"00001610A00AB084000400C00600000400001030040010050020020400001880",
INIT_05 => X"02000200400C8A09206420000C00410400000000000800000804000000000800",
INIT_06 => X"2A10201A12104010435051000801004040000322980800000080000100821000",
INIT_07 => X"000018400000086020002502000002000040800062C8081B0000008000088034",
INIT_08 => X"0A000610040440480000010000000000187C0000009100002046000110000010",
INIT_09 => X"4802082220084001002400214A2080014400006400A000000000015421800800",
INIT_0A => X"4B505008020032032320400011640447000010040000000020048409004A9020",
INIT_0B => X"280005922000045400002001100000000D0000008000000041C48000002003EA",
INIT_0C => X"2080020000208002000020800200002080010000104100800000100202420142",
INIT_0D => X"C06800100240180A0010010921003400432C8CC8D80044000000080080020800",
INIT_0E => X"2002C000C000240004641932041403428DA146D0A36850DA3200684004800403",
INIT_0F => X"0000000144002000420000000280001000420000000280000000084C01041008",
INIT_10 => X"0000000004801000500000000280001000500000000280001100000100000000",
INIT_11 => X"00010000000000000002A0002000020100000000000000182001000000240000",
INIT_12 => X"00110000000900003000004000000000000A0000000000000000900002000100",
INIT_13 => X"205D0080400000004803F0000800000000000004E0004E800120000000240BA0",
INIT_14 => X"4770000060000000000005600013560001100000000000002574020020000001",
INIT_15 => X"0020CA406A0000080200000000000020806000137400040000000000000B8000",
INIT_16 => X"68DA320D19D1A0CA8028984D46543600080040440C8090800000130061400140",
INIT_17 => X"8DA368DA368DA1685A1685A1685A1685A1685A1685A1685A1685A1685A1685A1",
INIT_18 => X"5A1685A1685A1685A1685A1685A1685A368DA368DA368DA368DA368DA368DA36",
INIT_19 => X"801010000000000000000068DA368DA368DA368DA368DA368DA368DA3685A168",
INIT_1A => X"344A2D840100E492082405548817344CCCF48DE68A89004F98614C5C38E2540A",
INIT_1B => X"1A0D068341A0D14514514514514514514514514514514514514534D34D34D34D",
INIT_1C => X"41A4D268341A0D069349A0D069349A0D068341A4D268341A4D268341A0D06834",
INIT_1D => X"FD557400000000000000000000000000000000000000000000001FFFFE2CAD83",
INIT_1E => X"007BC01FF5D7FFFE10002ABFF55F7D168A00552E95555007BFFF55087BE8BFFF",
INIT_1F => X"0F7FBC0145F7AE801EFF7FBFFF455D7BC0155F7D557410000000010F7D5421EF",
INIT_20 => X"00AA803FFEF5D55421EF002ABDF555D5157555F7FBC00AAAAD5400BA082AAAA1",
INIT_21 => X"4AAFF80021EF002A820BAFF8428A00A2AAAAAAAF7D17DE00FFFBD5555A2AABDE",
INIT_22 => X"75EFAAAABFFEF002A954BA5551421EF552E954105D00021455555420AA555155",
INIT_23 => X"575EFA2FFD75455D7BE8A005D5557410F7FBE8BEF552E95555552EAABEF082E9",
INIT_24 => X"000155FFD1400AA5D7FC01EFA2FFE8BEFFFFFEAB55002ABFE10080028BFFF7D5",
INIT_25 => X"71F8F7D147BEFBEFEBD152400000000000000000000000000000000000000000",
INIT_26 => X"C0005000E3D1401D71C7FC21EF5D75FFE10142EBAF7DE3D16DA0041209056D1C",
INIT_27 => X"AAD5420821C2EAAA10E3FFC0145F7A0801FFEBFBF8F6D417BC716DEBD1524101",
INIT_28 => X"8F7F5D0545B6AAB8E38B68A3AFFF5551471FF1C2EB8F45555550545E3F5C20BA",
INIT_29 => X"455D5B470925D51554AAE384001FF142E800AAFF802AA28AAAEAFABAE3D17DE2",
INIT_2A => X"56D4924ADBD70820975FFA2A4BFFFF082E974BA4155401C7552097428550E021",
INIT_2B => X"AE0008002ABFFF7DB505FFAAFBD7555417FEFA00495B52438F7FFEABFF412A90",
INIT_2C => X"00000000000000000000145F7D147092557BC21D7BEF5EDBC7FFF1EFB6D1420B",
INIT_2D => X"17DE100804001EF55516ABFF557BFDFEFA2D5400000000000000000000000000",
INIT_2E => X"7FD55FFA2D5400105D0417410AAD540155557FC01EF5D557DE105D2AA8BEFAAD",
INIT_2F => X"D5142155AAD1400AAA2D1420005D2EA9A00A2FBC0145FF84001EFA2FFEABFF00",
INIT_30 => X"A2AEBDEAAAAD17DEBAFFD142155FFAAAAABAFFAAAABFF5551555FF552EAAB455",
INIT_31 => X"55D00154AA552E801455D7BD54105D55574BAA280021EF5D2E820BAF7842AABA",
INIT_32 => X"AAF7FBEABEF002E801EF00003FF550800155FFA2803CFFF002E954BA00514015",
INIT_33 => X"F55F7D57FFEF550028A10000428BEFF7FFC01FFA2FFD5545007BFDE10087FC00",
INIT_34 => X"0000000000000000000000000000000000000145FFD157410557FC0155F7D57F",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000100",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(9),        -- Port A data input
DOA(0)   => data_read_a_lo_256(9),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(9),        -- Port B data input
DOB(0)   => data_read_b_lo_256(9),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_10_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10040B0001824802840102C00002C18000202300500030B3132000400992006",
INIT_01 => X"A140098018300848180060000C00424040000000080000080200010008110200",
INIT_02 => X"0801080200100000046558040080000041000000002402400800000009008010",
INIT_03 => X"00010100840000D0842242024210810802006400088000003080054288C10000",
INIT_04 => X"0000100022008000000C08C00C00000400A83A3044200C840000800400101820",
INIT_05 => X"0200000040000000248080210044000402000025000800020004207010100800",
INIT_06 => X"0800200000004010435040A14001004844000800CC0812541020008230829000",
INIT_07 => X"00000860408108502000250208000600004080006248081B0040808000088000",
INIT_08 => X"0A000210040440480060010000000000087C0810209900000002000110020010",
INIT_09 => X"08020A2222004040000484214A2080110108C280022210020240000401080880",
INIT_0A => X"000000000200000C042040001164044609101000840000802004800100421020",
INIT_0B => X"782415809888A45010082408028010080110280800001001051A124810410800",
INIT_0C => X"0089000890000900009000890008900008800048004420910800120242488000",
INIT_0D => X"4110000006008820020010010001300040000100014000808C48004008800090",
INIT_0E => X"2002000040002000040020020490080400020001000482000010012080008005",
INIT_0F => X"0000010140002040100000000280401040100000000280400000204801041008",
INIT_10 => X"0000000006801040020000000280401040020000000280400500000000000000",
INIT_11 => X"0000000000000000010280002400040000000000000001182001080010000000",
INIT_12 => X"10000000000D0000808000408000000200000000000000000000902000000500",
INIT_13 => X"A000000200000000681000000000000000008004A00040004000000000340000",
INIT_14 => X"4000008000000000000085200002000040000000000001002400000200000001",
INIT_15 => X"00200000000002000000000000000021802000020000000000000000020A8000",
INIT_16 => X"040006E00100044200289048085D402008000040000100000000020065400000",
INIT_17 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_18 => X"0000000000000000000000000000000020080200802008020080200802008020",
INIT_19 => X"8290100000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"8A355950666151451453D5006F86890A940FE0D39712614261D20E4355520542",
INIT_1B => X"6532994CA65328A28A28A28A28A28A28A28A28A28A28A28A28A28A28A28A28A2",
INIT_1C => X"AE532994CA6532995CAE572B94CA6532994CA6572B95CAE532994CA6532994CA",
INIT_1D => X"FFBC2000000000000000000000000000000000000000000000001007FECF31DC",
INIT_1E => X"007BFFF55087BE8BFFFFD557400FF842ABEFA2AAA8B5500003DF55F7D568AAAF",
INIT_1F => X"008556ABFFA2D16AB550000021FFF7D17FFEF08042AB55F7D168A00552E95555",
INIT_20 => X"55A2D557400557BC2010000000010F7D5421EF007BC01FF5D7FFFE10002ABFE0",
INIT_21 => X"145F7AE801EFF7FBFFF455D7BC0155F7D557545FFAE820AA007BFDFEF55003FF",
INIT_22 => X"00BA082AAAA00FFAE820AAAAAABDFEFF78028BEF005140145A2842AA10F7FBC0",
INIT_23 => X"6AB55A2D157400552EBFFEF5D7BD75EF002ABDF555D5157555F7FBC00AAAAD54",
INIT_24 => X"0000AAF7D17DE00FFFBD5555A2AABDE00AA803FFEF5D55420BA08557FEBAAAD5",
INIT_25 => X"0E3AF55F7DF68ABAE3F1C0000000000000000000000000000000000000000000",
INIT_26 => X"3D16DA0041209056D1C71F8F7D147BEFBEFEBD152400F7842FBD7B6AAAAB551C",
INIT_27 => X"5D75FFE10142EBAE0008556FBD7B6DB6AB7D1C0A001D7FFD178FC71C0E28B7DE",
INIT_28 => X"2147BFAFEF49043AF45A2DF504285D71C00101C0005000E3D1401D71C7FC21EF",
INIT_29 => X"7DA28428A10E3FFC0145F7A0801FFEBFBF8F6D417BC716DEBD15256DF7AA8209",
INIT_2A => X"545E3F5C20BAAAD5420821C2EAAA00E3AA82092A2AABAFD7EB8A2ABC70855401",
INIT_2B => X"70821C557AE92A2DF6AB7DA2DF50410412ABDFC75D7BD55FF1C2EB8F45555550",
INIT_2C => X"000000000000000000000BAE3D17DE28F7F5D0545B6AAB8E38B68A3AFFF55514",
INIT_2D => X"03DF45FFAEA8B555D2EAAB45F7FBE8ABAAAD5400000000000000000000000000",
INIT_2E => X"D168B55552AA8BEFAAD17DE100804001EF55516ABFF557BFDFEFA2D540010FF8",
INIT_2F => X"AD540155557FC01EF5D557DE105D2AA8A0008557FF45FFFFE8BEF5D2E80155FF",
INIT_30 => X"A2D5401FFF7AA800105D7FE8BEF08002AB45AAFFC00AA5D51400105D0417410A",
INIT_31 => X"5AAAEAAB450055421FFAA8428A00A2FBC0145FF84001EFA2FFEABFF007FD55FF",
INIT_32 => X"FF552EAAB455D5142155AAD1400AAA2D1420005D2EA9A10A2AA82010AAAEAAB5",
INIT_33 => X"ABAFFAAAABFF555155400555568A10AAFBEABEFA2FFC0010082ABFF55557BD55",
INIT_34 => X"00000000000000000000000000000000000000AAAAD17DEBAFFD142155FFAAAA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"FFFFFFFE00000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000000000000000000011F",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(10),        -- Port A data input
DOA(0)   => data_read_a_lo_256(10),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(10),        -- Port B data input
DOB(0)   => data_read_b_lo_256(10),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_11_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10180B05A0010402840602C2D001019000000300000000330A20080EC180002",
INIT_01 => X"AB400986B830284D1820E0000C36424840000000080000088200080802512220",
INIT_02 => X"8801081438106400A4F55800008000004100000040CCE24208005000C9060032",
INIT_03 => X"000406A492E6E440842254D002108153432004800880000030C0315688C00006",
INIT_04 => X"00001201200090001205400000000094108C322644240C840008030440111800",
INIT_05 => X"222000444008010028404002A002009402400025080880000C04223000170900",
INIT_06 => X"01080C1020002810436532AB4003004864200A00540816544522008200821100",
INIT_07 => X"6400E96C488108502001295BA100022E4340800062D82819435143F20008C0A0",
INIT_08 => X"0A0012160585C1D809A3810000000000C8FD0B1420992419034A0221116C3810",
INIT_09 => X"4902083E2CB0400002020480C2008009000ACEC06B25500202988C84C0220028",
INIT_0A => X"004040000203600E06204000116C14474A36500499C49C802004C00800088000",
INIT_0B => X"6804110230CBA4576708201C0212100B492A2008000A1001C49A9348498B0808",
INIT_0C => X"410E5418E5410E5418E5418E5410E5418B2A0872A08428010000120202085000",
INIT_0D => X"41110244066C0820221480010AA7300042080980919580808C9A5002880A18E5",
INIT_0E => X"2022C000C0002020094030220C960A0409020481024482501A00401410088521",
INIT_0F => X"836090540355D86C046619A54052A5B86A046619694063168280004801041008",
INIT_10 => X"A2C60289802AB86A046619A54052A5B86C04661969406316AC018B0E2936DA02",
INIT_11 => X"CB0E1076D4A200B2AC611A3D0405886C6EB211550815A8A2686EC81E2A48B68A",
INIT_12 => X"8CE0C5E8F650E48000892B37885620C1E1A06D7016A90A4626D82B10F1B1FC09",
INIT_13 => X"4E02144D335546F28724001B030A56140A184483000C410A2699A2E32AC9C041",
INIT_14 => X"E8018A0A01B2990242E278056AAA203920E0BAE2012C08281808319C186F1E16",
INIT_15 => X"44F9051C049B18A12CB481042AD140C227002A0A02066954E7540CCDB58415AA",
INIT_16 => X"409024681181044080809A490C0964200800200108010003A02272400C19B80D",
INIT_17 => X"0902409024090240902409024090240902409024090240902409024090240902",
INIT_18 => X"1004010040100401004010040100401024090240902409024090240902409024",
INIT_19 => X"0284000000000000000000401004010040100401004010040100401004010040",
INIT_1A => X"20A069105251C0000001541148062608804180C0B10A04CA0900474210420140",
INIT_1B => X"0000000000000000000000000000000000000000000000000000208208208208",
INIT_1C => X"0000000000004020000000000000000000100800000000000000000000000000",
INIT_1D => X"00015400000000000000000000000000000000000000000000001007FE0FC1C0",
INIT_1E => X"00003DF55F7D568AAAFFFBC2010557BEAA10AAFBE8A00557BFFFEF007BC21550",
INIT_1F => X"55D7FE8BFF5D7FD540055003FFEFFFD142145000000000FF842ABEFA2AAA8B55",
INIT_20 => X"45557FC2010557FFDF55F7D168A00552E95555007BFFF55087BE8BFFFFD55754",
INIT_21 => X"BFFA2D16AB550000021FFF7D17FFEF08042AB55A2AAAAB4508517FE00557BC01",
INIT_22 => X"FE10002ABFE00AAFFE8AAAFF8402000550002145085555400F7FFE8A0008556A",
INIT_23 => X"3FEBA002A975EFF7D17DFFFAA8000010000000010F7D5421EF007BC01FF5D7FF",
INIT_24 => X"000145FFAE820AA007BFDFEF55003FF55A2D557400557BC2145A2D1421450804",
INIT_25 => X"7BF8FEF1C7FC516D080E15400000000000000000000000000000000000000000",
INIT_26 => X"7842FBD7B6AAAAB551C0E3AF55F7DF68ABAE3F1C00005D7BEDA00B6F1EFA2855",
INIT_27 => X"147BEFBEFEBD15257D5D7FEFBD7417BD5438550038FC7FFDF4216D080E07000F",
INIT_28 => X"514517FE105575C216D5571C50104171FDF7DE3D16DA0041209056D1C71F8F7D",
INIT_29 => X"00FFF1EFA0008556FBD7B6DB6AB7D1C0A001D7FFD178FC71C0E28B6DA2AEADB4",
INIT_2A => X"1D71C7FC21EF5D75FFE10142EBAE10A2FBEFA92F78A05028550E001451455524",
INIT_2B => X"016DB6D54514500003FEBA1420905FFFFDF78FC7BE84050101C0005000E3D140",
INIT_2C => X"0000000000000000000016DF7AA82092147BFAFEF49043AF45A2DF504285D71C",
INIT_2D => X"FFDE00F7D17FEBA557BEABEF557BD55EF082A974000000000000000000000000",
INIT_2E => X"FBC01FF082A97410FF803DF45FFAEA8B555D2EAAB45F7FBE8ABAAAD5400105D7",
INIT_2F => X"804001EF55516ABFF557BFDFEFA2D5401FF5D7FFDF55007BD74BA5D042AB45F7",
INIT_30 => X"552AA8BEFAAAABFF5555517FE005555401FF55515541000517FFEFAAD17DE100",
INIT_31 => X"A5D2A801455D5140000FFD57FE0008557FF45FFFFE8BEF5D2E80155FFD168B55",
INIT_32 => X"105D0417410AAD540155557FC01EF5D557DE105D2AA8A10AAFBFFE00F7AA974B",
INIT_33 => X"B45AAFFC00AA5D51401FFFFD15555500003FEBA5D04001EFFFFFE8B55FF84174",
INIT_34 => X"00000000000000000000000000000000000001FFF7AA800105D7FE8BEF08002A",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000100",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(11),        -- Port A data input
DOA(0)   => data_read_a_lo_256(11),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(11),        -- Port B data input
DOB(0)   => data_read_b_lo_256(11),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_12_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50080B01BC002006940202C0DE041196A83183000000023322287E0FC000006",
INIT_01 => X"0E000C048000C048400380000007026040000000080000088200002802153231",
INIT_02 => X"2809AD0E7D180040945008040090000061800000C0E2F66009DA3D11CB148015",
INIT_03 => X"210D050012F6F8D2108216E24842005B8A20640008800000B8E0141C28851006",
INIT_04 => X"0080100022408000060DE0000066630C70241827041000040800820480001AA4",
INIT_05 => X"0240000C400000003C808003E0C8001401000000040900020904004000070800",
INIT_06 => X"00006C00000008784B4D210E0001006050800000100804005784000130821200",
INIT_07 => X"A64019490A044860300FA3968B20028FC06080106249F819A19143FE00088200",
INIT_08 => X"0A002610240D494A0753D1810240000038FC234480B1709A81C67325B31EFD18",
INIT_09 => X"090209222EB84000010000104200802180210C007827C000009DBE040800008C",
INIT_0A => X"0000000002000030003040081164FC469227D20019F413503004900020000200",
INIT_0B => X"28200100004304D267C06CC500566003C13E0000000460000000000010CE0000",
INIT_0C => X"E1865E1065E1065E1865E1065E1065E1832F0C32F08000000004100202015940",
INIT_0D => X"0403CFE7E03E8080382FD0018FE670004000000000D5C023009278B7835E1065",
INIT_0E => X"01EA0000440000800A0040028108000000000000000000000A74812DF00E0BF4",
INIT_0F => X"8362F658A7E5F82CD23B6B0E403DBBE82C563B6A4E403DBB88C0E04820020004",
INIT_10 => X"BE5403AB992F282C563B6B0E403DBBE82CD23B6A4E403DBBB1084E4B25AC48DF",
INIT_11 => X"0E4B1D32BAB504BB74AD3F3FE04A8E0D0C319A7988B6F0C75CFD801A962454CF",
INIT_12 => X"18D994B866E2E8C3808B6B63040328E7A33AF99B0AC20DE634D06C437BF85100",
INIT_13 => X"5F6214CA5991C6A7177402C49CA354D808D358A927EAD10A652CC8E3538BEC41",
INIT_14 => X"E80083C3EAEB2003695430A7CDAA289553922990C11A4E494988231B32570CDC",
INIT_15 => X"D5B304AD05A946D81616970A225658940BA7CDAA0A312666BD600E5550B49F36",
INIT_16 => X"00000100000010420000904C0040000008003B81000000021CFEE02E2803BC0F",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"8020080200802008020080200802008000000000000000000000000000000000",
INIT_19 => X"0210100000000000000000008020080200802008020080200802008020080200",
INIT_1A => X"24481C040000B5145144015085C1B946088881360A95118D90215C090CB05442",
INIT_1B => X"32190C8643219041041041041041041041041041041041041041249249249249",
INIT_1C => X"4B2592C964B2592C964B2592C964B2592C964B2592C964B2592C964B2190C864",
INIT_1D => X"AFBC2000000000000000000000000000000000000000000000001007FEF001D6",
INIT_1E => X"557BFFFEF007BC2155000015555087FC0010AAFBFFE100004020BAAAFFD5400A",
INIT_1F => X"5AA8400000A2AABFF45550400000AAFBFFFEF550000010557BEAA10AAFBE8A00",
INIT_20 => X"10555155555FF8017400FF842ABEFA2AAA8B5500003DF55F7D568AAAFFFBC215",
INIT_21 => X"BFF5D7FD540055003FFEFFFD142145000000145A2AA821EFFFFFD7410007FC00",
INIT_22 => X"8BFFFFD5574000051420BA557FC2145557FC20AAA2D57DEBAA2FBD55455D7FE8",
INIT_23 => X"AAA00550415410AAFBFFFEF55042AB55F7D168A00552E95555007BFFF55087BE",
INIT_24 => X"000155A2AAAAB4508517FE00557BC0145557FC2010557FFDE10AA8400000082E",
INIT_25 => X"0A02092B6F5D2438A2FBC2000000000000000000000000000000000000000000",
INIT_26 => X"D7BEDA00B6F1EFA28557BF8FEF1C7FC516D080E1557D0075C7028B6F1FAE0000",
INIT_27 => X"F7DF68ABAE3F1C017DAA8E07028B6A0BFF6D490E00000BEF5FAFEF4904070005",
INIT_28 => X"FE3FBD0438007FC00385D555556DEB8410400F7842FBD7B6AAAAB551C0E3AF55",
INIT_29 => X"BAA2FBD557D5D7FEFBD7417BD5438550038FC7FFDF4216D080E0716DAAA0851F",
INIT_2A => X"56D1C71F8F7D147BEFBEFEBD152400005F450BA417BC51454971C20AAB6D17DE",
INIT_2B => X"DE10BE8E070280020AAA28410410400BEFBFAFEF49042AB7DE3D16DA00412090",
INIT_2C => X"0000000000000000000016DA2AEADB4514517FE105575C216D5571C50104171F",
INIT_2D => X"5574BAFFD568A10002A82000FFD5400AAA2FBC00000000000000000000000000",
INIT_2E => X"D568BEF0004174105D7FFDE00F7D17FEBA557BEABEF557BD55EF082A975EF005",
INIT_2F => X"FAEA8B555D2EAAB45F7FBE8ABAAAD5401EFA2AA974BAF7803FFFF002A82000FF",
INIT_30 => X"082A975EFA280175FFAAFFC00BA087FC20AA5D55555FFA28000010FF803DF45F",
INIT_31 => X"50851420BAFFD57DEAAAAFBD75FF5D7FFDF55007BD74BA5D042AB45F7FBC01FF",
INIT_32 => X"EFAAD17DE100804001EF55516ABFF557BFDFEFA2D540010007FD74AA007BD754",
INIT_33 => X"1FF55515541000517FE10F7AA954AA080428AAA000002010FFFFE8BEF080428B",
INIT_34 => X"00000000000000000000000000000000000001EFAAAABFF5555517FE00555540",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"FFFFFFFE00000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000000000000000000001F",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(12),        -- Port A data input
DOA(0)   => data_read_a_lo_256(12),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(12),        -- Port B data input
DOB(0)   => data_read_b_lo_256(12),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_13_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10110A0441812402840402822007818000E00700000000330A3000000008042",
INIT_01 => X"A1400984B830C848180260000C0042404001000008220008A200100802110200",
INIT_02 => X"88010C02801040002475580400800000410000000064024608134C0CC9018034",
INIT_03 => X"00010100926220D084234212421085084300648A0880000630C0654288C10000",
INIT_04 => X"0004122122029100100C00001200009C40A83A2044360C84190BAC04E0101820",
INIT_05 => X"027000004009050064C8C00104C10184034010250089C00EB004327064B60900",
INIT_06 => X"910000152500A050436A10A14003004864B00A50440812541027008230821380",
INIT_07 => X"640029605091495020002B8AAA000AF003408000E258081963F100C00008C2E8",
INIT_08 => X"0A001210040441C802E0010084000000AAFC09142899000B20020001105A0010",
INIT_09 => X"4A02096A62004000020004104200802D9838C2C80322100202020194408000A0",
INIT_0A => X"000000000203240E46204000516C04468C101005800E95802004B20020080200",
INIT_0B => X"28200101118BA4510008241D005211000910000A000A1000809A93485D610000",
INIT_0C => X"0000000800000000000000800000000000000400000000000000100202055040",
INIT_0D => X"0100000006C0802042501001C8017000C2190890904000508908000000000800",
INIT_0E => X"0010C000C00081A08BC832A209AB0A85094284A14254A2551010513080109404",
INIT_0F => X"01293C0F5012906A96DCD13042CE0C206E92DCD07042CE0C40D0204800000000",
INIT_10 => X"71CA2168ACB0E06E92DCD13042CE0C206A96DCD07042CE0C4408632C39530BA9",
INIT_11 => X"632C30D522CE80239CC2806AC44E954939AB299E000738F88296CA13B444CA42",
INIT_12 => X"D5306028F01990C080808494A64708B265CC4052B0F30302E060965EA0058408",
INIT_13 => X"28A2CA9722094650CCAC0629112BA89C04A228568547B1654B9104A32865145C",
INIT_14 => X"B80D4D8D48CB54012290470562EC29E44050B1DC60132282B68B9AA60C051E03",
INIT_15 => X"0A5C11B9008FE2FA38F87804251CB0FAD40562EC0B426149D17E0044B10A158B",
INIT_16 => X"5094246A10A10441010090480C0964201800044109012001A000726E45428000",
INIT_17 => X"0942509425094250942509425094250942509425094250942509425094250942",
INIT_18 => X"9425094250942509425094250942509425094250942509425094250942509425",
INIT_19 => X"02A8000000000000000000509425094250942509425094250942509425094250",
INIT_1A => X"BAFFD7F7F7F775555557DF9FE0FFBBEEFF3F7DF7FF3E7E2FF0087B9F7DF7E245",
INIT_1B => X"FD7EBF5FAFD7EBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAE",
INIT_1C => X"AFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FA",
INIT_1D => X"0557DE00000000000000000000000000000000000000000000001007FE0001DF",
INIT_1E => X"0004020BAAAFFD5400AAFBC2155AAAA97410FFFFEAAAAF7AA955EFF7803FF450",
INIT_1F => X"0F7AEBDE10FFFFFDEAAF7D568AAA5D002AB55005568B55087FC0010AAFBFFE10",
INIT_20 => X"FF5D04154BAAAAEAAA10557BEAA10AAFBE8A00557BFFFEF007BC215500001541",
INIT_21 => X"000A2AABFF45550400000AAFBFFFEF550000155A28415410F7AEAABFFA2D1555",
INIT_22 => X"8AAAFFFBC21555D517FF45F7AEA8BFFA2AEAAA10A280021EF5D557FF55AA8400",
INIT_23 => X"974AAF7D142145082A975FF555568A00FF842ABEFA2AAA8B5500003DF55F7D56",
INIT_24 => X"000145A2AA821EFFFFFD7410007FC0010555155555FF80174000055555EFAAAE",
INIT_25 => X"A0925C7E38E38F7D14557AE00000000000000000000000000000000000000000",
INIT_26 => X"075C7028B6F1FAE00000A02092B6F5D2438A2FBC2145B6A090428FFF5EAA92E3",
INIT_27 => X"1C7FC516D080E15438E3A4BAE00FFF5FAE92F7D16AAAA41042FB7D145568B7D0",
INIT_28 => X"8FFA4AFBFFAAD1505FF490E174AABEA0ADA005D7BEDA00B6F1EFA28557BF8FEF",
INIT_29 => X"FF555F7FF7DAA8E07028B6A0BFF6D490E00000BEF5FAFEF490407155BE8E1242",
INIT_2A => X"B551C0E3AF55F7DF68ABAE3F1C0145415B78F45FFA4AFBC7BEA4AAA10A284001",
INIT_2B => X"04380055525FFBEAE90482E3D54216D0024975FF555F68A00F7842FBD7B6AAAA",
INIT_2C => X"0000000000000000000016DAAA0851FFE3FBD0438007FC00385D555556DEB841",
INIT_2D => X"0020BAF7D16AA10A28402155A2AEA8BEF5D516AA000000000000000000000000",
INIT_2E => X"003DFEF55516ABEF0055574BAFFD568A10002A82000FFD5400AAA2FBC0145FF8",
INIT_2F => X"7D17FEBA557BEABEF557BD55EF082A974BAA28028A00F7D16AA10F7D56AABA08",
INIT_30 => X"000417545FFAA820BAFF843DFFFA2D5421FF002E954AAFF843DE105D7FFDE00F",
INIT_31 => X"5F7802AA10AA80001FF5D7FFDFEFA2AA974BAF7803FFFF002A82000FFD568BEF",
INIT_32 => X"10FF803DF45FFAEA8B555D2EAAB45F7FBE8ABAAAD540145007FE8B55FF843DF5",
INIT_33 => X"0AA5D55555FFA280000BA0855401EFF7AA82010AAD1421FF0004155FF557FEAA",
INIT_34 => X"00000000000000000000000000000000000001EFA280175FFAAFFC00BA087FC2",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"FFFFFFFE00000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000000000000000000019F",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(13),        -- Port A data input
DOA(0)   => data_read_a_lo_256(13),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(13),        -- Port B data input
DOB(0)   => data_read_b_lo_256(13),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_14_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10020A000180000284008280000281800000030000000033022000000580002",
INIT_01 => X"A140098018300848184860000C20C24040000000084000084200000000110200",
INIT_02 => X"88010C5A8010A600A4F558040080000041000000022C024008003CCCC9028030",
INIT_03 => X"000103A7A00904D0842242024210810803006480088000003081054288C10000",
INIT_04 => X"0000120122009000100C00000000000400A83A2044200C840000800400101820",
INIT_05 => X"020000004008010024C0C0010040000402000025000800020004207000100800",
INIT_06 => X"010000102000005043403AA14003004864000A00440812541020008230821000",
INIT_07 => X"2400A96850A16854200021DA2A0002000340800062C80819EBC402800008C020",
INIT_08 => X"0A0012140404414814E001000000000029FD0A10289924810182000110028010",
INIT_09 => X"080208222200400002000400420080010008C2C0032210020200008440000080",
INIT_0A => X"000000000203200E0620400011640446DA101004800005802004800000000000",
INIT_0B => X"282001001088A45000082408000010000910000800001000009A924810410000",
INIT_0C => X"0080000000000000080000000000000080000000000000000000100202000000",
INIT_0D => X"0100000004408020021010010001700042080880904000008808000000000800",
INIT_0E => X"00000000C00000000040302200800A0409020481024482501010413080008404",
INIT_0F => X"8090008142014840100002C38280000840100003838280000640204800000000",
INIT_10 => X"072C000444C00840020002C38280000840020003838280002C09D01086839746",
INIT_11 => X"D0104B01C57100440202900184414430534605E3804802180022480419183514",
INIT_12 => X"594C194000090450808802008830024F0E248C902AEF0024170CF18001003C09",
INIT_13 => X"20020E5A08E6000048200196264BCF1C030C0604800001076C04730000240049",
INIT_14 => X"2003DEDE82C78900902A0D0000080019FAAA32D9602490302409292B83280001",
INIT_15 => X"049100021171F6C34080240108AB292CA000000800AD1A19F6F000AA0C0A0000",
INIT_16 => X"4090246810810440000090480C0964200800000108010016000012004542800D",
INIT_17 => X"0902409024090240902409024090240902409024090240902409024090240902",
INIT_18 => X"9024090240902409024090240902409024090240902409024090240902409024",
INIT_19 => X"0280000000000000000000409024090240902409024090240902409024090240",
INIT_1A => X"9E7FDDF77777F3CF3CF7D54CEFD79B4E5C8FF0F7BE9D75C7F7B71F5F7DF65040",
INIT_1B => X"7F3F9FCFE7F3F9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7",
INIT_1C => X"E7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE",
INIT_1D => X"28417400000000000000000000000000000000000000000000001007FEFFFE0F",
INIT_1E => X"F7AA955EFF7803FF4500557DF45F7D16AB455D00001EFAAAAAAABA555557555A",
INIT_1F => X"555003FF450804001555D2AA8AAA002ABDE10082ABDF55AAAA97410FFFFEAAAA",
INIT_20 => X"EF5D5168A10082E80155087FC0010AAFBFFE100004020BAAAFFD5400AAFBC214",
INIT_21 => X"E10FFFFFDEAAF7D568AAA5D002AB55005568A00A2D5401455D00175FFFF84175",
INIT_22 => X"2155000015400AAD157545080402145087FD75FFF7AE82145A2D17FE10F7AEBD",
INIT_23 => X"000BAFFFBE8AAAA2FBFDE00087FD5410557BEAA10AAFBE8A00557BFFFEF007BC",
INIT_24 => X"000155A28415410F7AEAABFFA2D1555FF5D04154BAAAAEAAA005D002AB450000",
INIT_25 => X"A0AAA82555157555B68012400000000000000000000000000000000000000000",
INIT_26 => X"6A090428FFF5EAA92E3A0925C7E38E38F7D14557AF45FFDB6AB6D4100071C7B6",
INIT_27 => X"B6F5D2438A2FBC21455D0A3FF6D080407155552AAAA920020BFE10002EBAF45B",
INIT_28 => X"54100175C7E380125D7555B6DA1014248217D0075C7028B6F1FAE00000A02092",
INIT_29 => X"45AAD178E38E3A4BAE00FFF5FAE92F7D16AAAA41042FB7D145568A38AADF4014",
INIT_2A => X"A28557BF8FEF1C7FC516D080E15400A2DB5754508040716D007BD05EFEBAA821",
INIT_2B => X"DA0055002AB6D0000020BAFFF1E8ABABEF1FAE001C7FD54005D7BEDA00B6F1EF",
INIT_2C => X"00000000000000000000155BE8E12428FFA4AFBFFAAD1505FF490E174AABEA0A",
INIT_2D => X"FEABFF080015555F78028A00555155555FF84000000000000000000000000000",
INIT_2E => X"003DE10082EAAB45FF80020BAF7D16AA10A28402155A2AEA8BEF5D516AB45F7F",
INIT_2F => X"FD568A10002A82000FFD5400AAA2FBC0145552ABFFFF000417555552EA8A1000",
INIT_30 => X"55516AABAAAFFC0145000417555A280001455D7FFDE105504021EF0055574BAF",
INIT_31 => X"F007BC01FFAAAE80155AAD568ABAA28028A00F7D16AA10F7D56AABA08003DFEF",
INIT_32 => X"105D7FFDE00F7D17FEBA557BEABEF557BD55EF082A97410AAFFD55450800155F",
INIT_33 => X"1FF002E954AAFF843DE10550028BEF0004020BAF7D568AAAF7D168A105D7FD74",
INIT_34 => X"0000000000000000000000000000000000000145FFAA820BAFF843DFFFA2D542",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"FFFFFFFE00000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000000000000000000001F",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(14),        -- Port A data input
DOA(0)   => data_read_a_lo_256(14),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(14),        -- Port B data input
DOB(0)   => data_read_b_lo_256(14),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_15_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000A000000000284000280000001800020030000000033022000000180002",
INIT_01 => X"A140098018300848180060000C00424040000000080000080200000000110200",
INIT_02 => X"080108000010E60004E55800008000004100000000040240080000C009170016",
INIT_03 => X"0000000080000040842240000210810002000400888000003080014288C00000",
INIT_04 => X"0001100024A0800000440000000000040088322044200C840000011400151800",
INIT_05 => X"A200014C4000000020000000000B8094020000254C8800000514203000108800",
INIT_06 => X"000821000000A050434010A14001004844000801540812540020008600831000",
INIT_07 => X"C2000864489128502000210222000200034080006248081958C0008000088000",
INIT_08 => X"0A001214050540C800200101860000000B7C0910209900000002000110000010",
INIT_09 => X"0B0208222004400000000400420080010008C28002201002020001140800002C",
INIT_0A => X"000000000203000C04204000116404460810100080000F802004800000000000",
INIT_0B => X"280001001088A45000082008000010000100000800001000001A124800010000",
INIT_0C => X"0080000800008000000000000000000080000400004000000000100202000008",
INIT_0D => X"0100000004C00020025000018801600040000000000000008808000000000800",
INIT_0E => X"00108000C0000000000020020080080000000000000402000000000000009400",
INIT_0F => X"00000000000000404200000000000000404200000000000008C0004800000000",
INIT_10 => X"0000000000000040500000000000000040500000000000000400000100000000",
INIT_11 => X"0001000000000000000000000400020100000000000000000000080000240000",
INIT_12 => X"00110000000000C00080010180000000001A1024050000000000000000000400",
INIT_13 => X"0002008040000000002000000804002000000000000001000120000000000040",
INIT_14 => X"2000000061100280000000000008000001104422000000000008020020000000",
INIT_15 => X"00100000000009080E2E0A000000000000000008000004000000000000000000",
INIT_16 => X"0000046000000440000090480809402008000001000000000000000004188000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0280000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000040000000000040",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"8517DE00000000000000000000000000000000000000000000001007FE000000",
INIT_1E => X"AAAAAAABA555557555A284175FF000002010552A97400007BFDE10A2AA801EF0",
INIT_1F => X"F5D2AAAB45F7D17DF45087BC0155002A801FF08003DF45F7D16AB455D00001EF",
INIT_20 => X"45F7D568BEFAAD557555AAAA97410FFFFEAAAAF7AA955EFF7803FF4500557DFE",
INIT_21 => X"F450804001555D2AA8AAA002ABDE10082ABDFFFF7D17FE10002E954AAF7FBC21",
INIT_22 => X"5400AAFBC21EFA2AE95545A2D56ABFFAAD17DE10FFD1420AA007FC014555003F",
INIT_23 => X"801550055401555D00174BA002AA8B55087FC0010AAFBFFE100004020BAAAFFD",
INIT_24 => X"000000A2D5401455D00175FFFF84175EF5D5168A10082E801FFFF8428A10002A",
INIT_25 => X"71FAE00A2A0871EF145B7FE00000000000000000000000000000000000000000",
INIT_26 => X"FDB6AB6D4100071C7B6A0AAA82555157555B680125C71C0E0500049209543808",
INIT_27 => X"E38E38F7D14557AFC75524AFB45FFD178F7D1C71C2145002E801C7140A3FF45F",
INIT_28 => X"00024954AAFFFBC2145F7DB6DBEFA2D557545B6A090428FFF5EAA92E3A0925C7",
INIT_29 => X"820071C71455D0A3FF6D080407155552AAAA920020BFE10002EBAFC7FFDF7AE0",
INIT_2A => X"E00000A02092B6F5D2438A2FBC21FFBEA090545B6D568BFFAADB7AE10F7D5470",
INIT_2B => X"21FFE3802FA2808208017D1C5142155410A104AA1420AFB7D0075C7028B6F1FA",
INIT_2C => X"00000000000000000000038AADF401454100175C7E380125D7555B6DA1014248",
INIT_2D => X"E954100004174AA00516AA10AA80155EF5D7BFDE000000000000000000000000",
INIT_2E => X"2E801555D2EBDF45F7FFEABFF080015555F78028A00555155555FF8400155552",
INIT_2F => X"7D16AA10A28402155A2AEA8BEF5D516AB555D043DF55F7D56ABEF55514015508",
INIT_30 => X"082EAAB55FFFBE8A100804154AAF7FFC2145FFFFFDFEFAAD157545FF80020BAF",
INIT_31 => X"FA2FBE8A00FFD155410005555545552ABFFFF000417555552EA8A1000003DE10",
INIT_32 => X"EF0055574BAFFD568A10002A82000FFD5400AAA2FBC01FFF78400155F7D16ABE",
INIT_33 => X"1455D7FFDE105504021FFAA843DEBA0000021EF555142155002E800AA55003DF",
INIT_34 => X"00000000000000000000000000000000000000BAAAFFC0145000417555A28000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000180",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(15),        -- Port A data input
DOA(0)   => data_read_a_lo_256(15),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(15),        -- Port B data input
DOB(0)   => data_read_b_lo_256(15),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_16_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"DA22C618B1000482B688B186588884862A400438255FC38381441205BA803003",
INIT_01 => X"8645A80028404C211203A952A90341080B173340412000E1005D628000820484",
INIT_02 => X"A101A9006DC1084833011850AAC55001349B10881802821808B4110007005E11",
INIT_03 => X"010108A802BB00080080006020020001A61036202800000D2410104200404550",
INIT_04 => X"8BFA58800005C40A46240252145148B38248030356415A4E62B6FC660F287240",
INIT_05 => X"0F05EA11E570000D610000000710296E542B6E3A825C15FB30A643695BFC2D56",
INIT_06 => X"408003200040202B8584112645554B029006000140BCC0460050690A95C8383D",
INIT_07 => X"00480A2140040BE1480FA004342AA6F12000054004867415401DCDCF2AA10800",
INIT_08 => X"B32A8819064E48288012D45000005050247AA85220700009C06206C48080EDEA",
INIT_09 => X"445B2081340B6596594800400413CAC020894480000008C54C00311002000002",
INIT_0A => X"000000004B240028000342A00002FE00A3A1F06E491800AA29588181040A0020",
INIT_0B => X"2400848002912300200092BA80325A20000000000A8A5AA80018120E00066000",
INIT_0C => X"00220002200022000220002200022000210001100010000A40450100210072A0",
INIT_0D => X"002815014B90000205DA00880100095A648000000010006AC23000C7B69EC220",
INIT_0E => X"80922554515512174000000490009000000000000004010042A204A0C5817680",
INIT_0F => X"63EAA9C238B2D4C800632B266E828EE4C800632AAAB6830D0FC6B06C04102800",
INIT_10 => X"A149339E8FB964C800632B266E82B2E4C800632AAAB683310872800EDA52DA00",
INIT_11 => X"800EB090D4AAC91268FFCBE81397826C4A20D2B6C510E8624792A4A30A40839A",
INIT_12 => X"8849D5C532408DD6E004C90C06AC019D88B9795012CA96902C799912BC3C087A",
INIT_13 => X"531C74485BD42A30906057FADAA456218FD8E3ED83B60E3A242DC0F18983638E",
INIT_14 => X"A06FB555793057C444CF45C5C9E89543B8BC6E80193DC36F6C71D1093A478706",
INIT_15 => X"45DC02B331650CA8ACB4007E00D1C6A6A58395C917F7E74D936F650D69B51727",
INIT_16 => X"0000012000081500008A422150884081ACAAC0542054004FC588464050810DCD",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"147A7797E1E1A79E79E1560EEFBD11544C690DA64C1C69A9916D7E4F68A36040",
INIT_1B => X"7A7D1E9F47A7D345345345345345345345345345345345345345145145145145",
INIT_1C => X"4FA7D3E9F4FA3D1E8F47A3D1E8F47A3D1E9F4FA7D3E9F4FA7D3E9F4FA7D1E9F4",
INIT_1D => X"F8015400000000000000000000000000000000000000000000001007FE00001F",
INIT_1E => X"007BFDE10A2AA801EF08517DE10FFFFFDFEFA2D16AB55A2FFFFEAA5D7FC0000F",
INIT_1F => X"A5D2EBDFEFAAD17FFFF002EBDE000800174AA55043FFFF000002010552A97400",
INIT_20 => X"AAAA80000105D557FF45F7D16AB455D00001EFAAAAAAABA555557555A284174B",
INIT_21 => X"B45F7D17DF45087BC0155002A801FF08003DE000004154BA002A800BA087FE8A",
INIT_22 => X"FF4500557DEAAF7D57DEBA082A82010FFAE975555D7FFDEAAFF80155EF5D2AAA",
INIT_23 => X"7FFFF557FD55FF08003FE0055043FF55AAAA97410FFFFEAAAAF7AA955EFF7803",
INIT_24 => X"0001FFF7D17FE10002E954AAF7FBC2145F7D568BEFAAD557410552EA8BEFA2D5",
INIT_25 => X"FFFDEAA5571C7010FF8412400000000000000000000000000000000000000000",
INIT_26 => X"C0E050004920954380871FAE00A2A0871EF145B7FE10E3F1F8FC7AAD56DB7DB6",
INIT_27 => X"555157555B680124924124BDFEFA2D57FFC71C2EBDE280000174825D0E3FFC71",
INIT_28 => X"21424800AA007FEDAAAA284020385D5F7AF45FFDB6AB6D4100071C7B6A0AAA82",
INIT_29 => X"AAFF80175C75524AFB45FFD178F7D1C71C2145002E801C7140A3FE10080A1748",
INIT_2A => X"A92E3A0925C7E38E38F7D14557AE92EBDB78EAA1C2482010FFAE9556D557FF8E",
INIT_2B => X"7410492EADBEFA2D178FEF5575D55EF000A38E10490A3AF45B6A090428FFF5EA",
INIT_2C => X"000000000000000000001C7FFDF7AE000024954AAFFFBC2145F7DB6DBEFA2D55",
INIT_2D => X"56AB45A2D57DFFFF7FBFFEAA555555400F780000000000000000000000000000",
INIT_2E => X"0415400552ABDF55552E954100004174AA00516AA10AA80155EF5D7BFDE10A2D",
INIT_2F => X"80015555F78028A00555155555FF840000000043DFEFAAD17FF45552ABFEBA08",
INIT_30 => X"5D2EBDE10002E974005D04020BA007BFDEBAA284000BA557FE8B45F7FFEABFF0",
INIT_31 => X"0F7AE955EF5D7BE8ABAF784175555D043DF55F7D56ABEF555140155082E80155",
INIT_32 => X"45FF80020BAF7D16AA10A28402155A2AEA8BEF5D516AA00AAFBE8AAA55040000",
INIT_33 => X"145FFFFFDFEFAAD157410082ABFFEFAAD16ABFF5555575FF082AA8A00002AAAB",
INIT_34 => X"0000000000000000000000000000000000000155FFFBE8A100804154AAF7FFC2",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000080",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(16),        -- Port A data input
DOA(0)   => data_read_a_lo_256(16),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(16),        -- Port B data input
DOB(0)   => data_read_b_lo_256(16),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_17_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"5284CE4FB7BD2C8994A13392DBD02E14006B82AC7E800D44D3DD2FD5F9B961C0",
INIT_01 => X"F8ACD01F7E03FC6793F2199B39FC233C11D93AE6F3BB92B32091DBC339B24542",
INIT_02 => X"8F333007FD6808092A2AFA6667033DB50853379C10BFF70F1BD011110F205F18",
INIT_03 => X"294ADB4AFFCBF0DAD63ABF836B58EAFE060478202022234B2E0303FDC9E18339",
INIT_04 => X"DB7A40806FE4040840EBC563A0150A0926146FECB04196482236FC2005282AE1",
INIT_05 => X"0403DA0383200831C68206D7E6D0250834336D1E81500FDB306045255BFC2076",
INIT_06 => X"4470716040413D29AAC69F5FE33C072F06062C003670497AFF00291B3C0E2015",
INIT_07 => X"0849147160448EBB9537A0022DC67987042EE976ABEA77684653547819FF2000",
INIT_08 => X"E019C0C82A4E4820C15B089C380110002446045A31345000A84432409207F02D",
INIT_09 => X"983838A3BFF1030C397C060B4254064302042F803A69DB931FF4391C00002CC0",
INIT_0A => X"FB1F1F7BC81C003C001674BB55B5FBB4BB4F26A1BEE004F9D0DE08F7DE336DB2",
INIT_0B => X"28302F800633F1D0A7CC9AE74117FE01D34E82AC0CE8FCCC200A59BDD2FFE3E3",
INIT_0C => X"E9F79E9F79E9F79E9F79E9F79E9F79E9F7CF4FBCF4F000C2E225C8DE0BA05BB0",
INIT_0D => X"A5A99FD6D3FEF4BEB5FF994F0FEFFCCF8430000000D9D147E0D57AE7B79E9F79",
INIT_0E => X"0593F33FA0CF170F40006001B1A05C0000000000000008004BA78428C7AD7FE4",
INIT_0F => X"E46444357B3950A9BFBAC94CFA8581E0A9BFBAC8CCFA8580C7CAF51EF68B2976",
INIT_10 => X"B5DB54A09003E0A9BFBAC94CFA8581E0A9BFBAC8CCFA8580E46FBFCB0CBEDA57",
INIT_11 => X"BFCB1D5CFEB56A1A100D5345C1BFFE8FBDB892DB463034198E2881F3F787DF76",
INIT_12 => X"D39387F92B2935DFEAADDF38EBCFB9E3D636DCDF9B90F966BF92966D5D9E7467",
INIT_13 => X"27055EB6D555CB294981B7FB5B2954CD3013013FDF5E82AF5B6AAAE594A4E0AD",
INIT_14 => X"835C67E655BAA868610117575EA1C34BD6975D48B44A0405FC15BA7270FF2565",
INIT_15 => X"6CD2A47D0CBA96252756D7217E5E1C61DBDF5FA167F7AE5D3D21A414007F7D7E",
INIT_16 => X"000005F08000179C16DECF67F08BC02F9067ED55805600545DFE45A80E7BD07F",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"00C0000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"9A919261A1A6075D75D10DDF2F82003009EDCC4052E92E0826462117114F9818",
INIT_1B => X"8D068351A8D069A6BAE9A69A6BAE9A6BAE9A69A6BAE9A6BAE9A69A69A69A69A6",
INIT_1C => X"A8D46A351A8D46A351A8D46A351A8D46A341A0D068341A0D068341A0D068351A",
INIT_1D => X"AFFD5400000000000000000000000000000000000000000000001FFFFE000011",
INIT_1E => X"A2FFFFEAA5D7FC0000FF8015410FFFFFFFFFFFFFFDFEFF7D568A1008003DF55A",
INIT_1F => X"5A2D1400000804154BAF7D168A00A2803DE10FFAE95410FFFFFDFEFA2D16AB55",
INIT_20 => X"BAFFD56ABFF002EBDFFF000002010552A97400007BFDE10A2AA801EF08517DF5",
INIT_21 => X"FEFAAD17FFFF002EBDE000800174AA55043FEBA0004174AA5504000AA55042AA",
INIT_22 => X"7555A284175FFFFFBE8B55A2FFFFF55F7803DEBA002AAAAAAF7FBD74BA5D2EBD",
INIT_23 => X"17400FFD57DE00AAAAAAB45A2AA97545F7D16AB455D00001EFAAAAAAABA55555",
INIT_24 => X"0000000004154BA002A800BA087FE8AAAAA80000105D557FE00A2D5420AA5D04",
INIT_25 => X"D16AA00000E3DF6DBEF5D2400000000000000000000000000000000000000000",
INIT_26 => X"3F1F8FC7AAD56DB7DB6FFFDEAA5571C7010FF8412428FFFFFFFFFF7FBF8FD7EB",
INIT_27 => X"A2A0871EF145B7FF7DA2D547038140E10492FFDF6DA28A28E3DE00F7A092410E",
INIT_28 => X"2550A020BA55002AA82F7DF6DBD71C2EBFFC71C0E050004920954380871FAE00",
INIT_29 => X"BAF7F5D74924124BDFEFA2D57FFC71C2EBDE280000174825D0E3FEAA14001249",
INIT_2A => X"1C7B6A0AAA82555157555B680125FFEBFFEDB55BEFFFAF6DE38E3DEAA002EADA",
INIT_2B => X"AE28B6D545092490E10400FFDB7AE00A2AAADB45BEA092545FFDB6AB6D410007",
INIT_2C => X"00000000000000000000010080A174821424800AA007FEDAAAA284020385D5F7",
INIT_2D => X"BFDFEFF7FFEAB45A2D56AA00002EBDFFFF7D5400000000000000000000000000",
INIT_2E => X"AABDE10FF8400010A2D56AB45A2D57DFFFF7FBFFEAA555555400F780000AAFFF",
INIT_2F => X"004174AA00516AA10AA80155EF5D7BFDFEFAAD1554BA552E82000F7FFFFEAAA2",
INIT_30 => X"552ABDEBA5D0002000552A800BA55042AA10FFFFFDF55552EBDF55552E954100",
INIT_31 => X"FA2AEBFEAA082EBDEBAFFD55540000043DFEFAAD17FF45552ABFEBA080415400",
INIT_32 => X"45F7FFEABFF080015555F78028A00555155555FF84001FFAAFBFFF55FFFBEABF",
INIT_33 => X"EBAA284000BA557FE8AAAFFD155400082A82000F7FFE8A00A2AABDF45F780001",
INIT_34 => X"0000000000000000000000000000000000000010002E974005D04020BA007BFD",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"FFFFFFFE00000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000000000000000000019F",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(17),        -- Port A data input
DOA(0)   => data_read_a_lo_256(17),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(17),        -- Port B data input
DOB(0)   => data_read_b_lo_256(17),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_18_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"69844019080000A21A611406840014122A641074155FC28A2024001001801003",
INIT_01 => X"A643D920034004180005E9E3C90360C0041C0181002001602025800008440084",
INIT_02 => X"B7333980808408103F2000F81FC0FEDEAC2161B0B84D0002188011110C018041",
INIT_03 => X"0405D434003F2C020081587008020561E55116B0290000042B71240C800440F8",
INIT_04 => X"50805AC31007D6125724029216554A9847669903D640EC8E2001002604503004",
INIT_05 => X"07008000E0EA11803850C800010022660C1C0065003C0404002646DC20A02D40",
INIT_06 => X"0100001028040C093D0491A640FFC10028000280002C44D620F0228454C83810",
INIT_07 => X"08501620028007500CE801241021FE78E40486014006009044359DC707F55C20",
INIT_08 => X"9307CC082A0A4A6A01ECDCC40850001630080002A5CA500344040108120080AB",
INIT_09 => X"A0172083200B6186128040600C10C1C02009505081100088080BC6A052802001",
INIT_0A => X"002020000F0CA8428642430080438408A510185A40000008B83181C000141040",
INIT_0B => X"2E00C04C44C92A88DC42215C882E82240880000060D7030C30B885200D274404",
INIT_0C => X"10006100061000610006100061000610003080030800800C0540310130006E21",
INIT_0D => X"10202021000780004200408C1002003F66CA18A1B62622381B2B841840614006",
INIT_0E => X"806400FC503F08180050942E4200020C1B060D8306C182701404C19730108010",
INIT_0F => X"ABAF377DF1CA160820520EB3057E70E60820520F33057E72E915415900002900",
INIT_10 => X"5D48F37FAFEFE60820520EB3057E7CE60820520F33057E7EC658BF2DA7822AAB",
INIT_11 => X"BF2D4B2A80BF8FE39FD78EB0D882014A62C568FFAFC73FFDD9C2B30E0468A2AD",
INIT_12 => X"800DFC06F59F710107533C0C4E37619440FBFBAB2400AFC1600361D798F32658",
INIT_13 => X"EB9454005BAA36DEFF894823A3D1A88A2FE29D5FC6DCAA2A002DD51B6E7C728C",
INIT_14 => X"92A78606A28A5427AAB9FF4EDD251C7123E291660733EBF6FE519001BF40DEBB",
INIT_15 => X"AB58AFBFD5DE200A8EBE3A3EC110339E1DCEDC2590495BB2112E2BE4BF5F3B70",
INIT_16 => X"C1B06808348340000020301805002D008C1F92000A5F421B8000DB4910382202",
INIT_17 => X"1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06",
INIT_18 => X"B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C",
INIT_19 => X"000000000000000000000041B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1",
INIT_1A => X"8A244C16454170410412CA064A9BBECEB80EE173C2300FE3F1A3550F7DF16000",
INIT_1B => X"A552A944A2512AAA8A28A28A2AAAAAA8A28A28A2AAAAAA8A28A28A28A28A28A2",
INIT_1C => X"A25128944A25128944A25128944A25128944A25128944A25128944A25128954A",
INIT_1D => X"D2A80000000000000000000000000000000000000000000000001007FE000004",
INIT_1E => X"F7D568A1008003DF55AAFFD5410FFFFFFFFFFFFFFFFFFFFFBFDEBA552E974105",
INIT_1F => X"0FFFFFFFFFF7FBE8B55AAD16AA1000516AA005D0400010FFFFFFFFFFFFFFDFEF",
INIT_20 => X"00087BC2155087BC0010FFFFFDFEFA2D16AB55A2FFFFEAA5D7FC0000FF801541",
INIT_21 => X"0000804154BAF7D168A00A2803DE10FFAE95555FFFBE8B45A2D56ABEFFFFFFFE",
INIT_22 => X"01EF08517DF55000000010082A974AA08557DEBAFFAEBFF55AA8028B55A2D140",
INIT_23 => X"800105D2AAAA10A2D1420AAFFAEA8BFF000002010552A97400007BFDE10A2AA8",
INIT_24 => X"0000BA0004174AA5504000AA55042AABAFFD56ABFF002EBDEBA0004020BA552E",
INIT_25 => X"FBFFEBA552A95410552485000000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFF7FBF8FD7EBD16AA00000E3DF6DBEF5D2438FFFFFFFFFFFFFFFFEFF7",
INIT_27 => X"5571C7010FF8412410FFFBF8FC7E3F5EAB45BEDB6FA3800556FA00550405028F",
INIT_28 => X"5BEDB6FBC7EBF5F8E10007BC516D1C71C5010E3F1F8FC7AAD56DB7DB6FFFDEAA",
INIT_29 => X"55BE8A2DB7DA2D547038140E10492FFDF6DA28A28E3DE00F7A09256DE3F1EAB5",
INIT_2A => X"4380871FAE00A2A0871EF145B7FF45080E070280820924AA145578E92F7A4BFF",
INIT_2B => X"FEBA1C0A00092412E850005D2AAFA38A2DF45082F7AAA8BC71C0E05000492095",
INIT_2C => X"000000000000000000000AA140012492550A020BA55002AA82F7DF6DBD71C2EB",
INIT_2D => X"FFFFFFFFFBFDFEFF7FFFDEAA5D2E954105504154000000000000000000000000",
INIT_2E => X"557DE005500154AAFFFBFDFEFF7FFEAB45A2D56AA00002EBDFFFF7D5400AAFFF",
INIT_2F => X"2D57DFFFF7FBFFEAA555555400F78000010F7FBE8B55AAD16AB55F7FBFDEAA08",
INIT_30 => X"FF84001FFAAD568B45FFFBFFF55A2D568A00087BD55FF5D5555410A2D56AB45A",
INIT_31 => X"A555168A10FF803DF45FFAABDFEFAAD1554BA552E82000F7FFFFEAAA2AABDE10",
INIT_32 => X"55552E954100004174AA00516AA10AA80155EF5D7BFDF45002A974AA0800000A",
INIT_33 => X"A10FFFFFDF55552EBDEBA5D2E80010082A97410552EBDEBAA2FBD5400F7AAA8B",
INIT_34 => X"00000000000000000000000000000000000000BA5D0002000552A800BA55042A",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000080",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(18),        -- Port A data input
DOA(0)   => data_read_a_lo_256(18),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(18),        -- Port B data input
DOB(0)   => data_read_b_lo_256(18),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_19_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"042200000000000041088001001AA00000000000000000000000500802000003",
INIT_01 => X"200048000024000000000404000000000A22000800000800004A200000000001",
INIT_02 => X"032210008DEF00400060000001C008002489E0F0004037B00010101010000000",
INIT_03 => X"0000008128000000000000000000000024001620280000000000354200004008",
INIT_04 => X"000058800004C4024024001210001054B1C822009640000E2000002604003000",
INIT_05 => X"07008000E0200000000000000000200604000000001C04000026400000002C40",
INIT_06 => X"000000000000002600859AA1000D410000000000002C42010010200004C83810",
INIT_07 => X"0040380142810010564C41001140120024020280448088050008108100640000",
INIT_08 => X"83004C390242006200000868000040001020A850040AD0080426006933800DC4",
INIT_09 => X"0013200000016186100000000010C04002C00000000000707000000000000000",
INIT_0A => X"000000000B0C0000000101400040C0408100000000000008A810000000000000",
INIT_0B => X"00000000000400020000440000000000000000002F0001F00002024B20002000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"000210001D800000000000000002000964000000000000000000000000000000",
INIT_0E => X"0000000C50030008000000000000000000000000000000000000000000000000",
INIT_0F => X"101088A37034E156600D740022800EC156600D740022800D01E0412D06904000",
INIT_10 => X"0224081044914156600D7400228002C156600D7400228001098F00D0FB750500",
INIT_11 => X"00D0F2DD014010046037814EA63DBB31CE7605001008C41A061F0E7D693E6170",
INIT_12 => X"6D600000004089E12350C0E01FF23315422BABB46FEF5019146C0800380CC98F",
INIT_13 => X"130AA3592000000000629C03F3E60330C00C628908214551AC90000001036152",
INIT_14 => X"65C006070845039014460088235ACC3123E2A29148841008482A4DAC00000000",
INIT_15 => X"53A66BE7A5040018D8A8AD9090A1EC20A188235AC509FB50C2D0500B4094208D",
INIT_16 => X"000000000000000000000000000000008C01800270000061100084046086CD49",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"861A2882313054D34D301C862AA08BBA3F0C7010C6600A00200251C744192000",
INIT_1B => X"130984C261309861861861A69861861861861A69861861861861861861861861",
INIT_1C => X"6130984C26130984C26130984C26130984C26130984C26130984C261349A4C26",
INIT_1D => X"82E97400000000000000000000000000000000000000000000001007FE000002",
INIT_1E => X"FFFBFDEBA552E974105D2A801EFFFFFFFFFFFFFFFFFFFFFFFFFEAA552E954000",
INIT_1F => X"FFFFFFFFFFFFFFFFFEFF7FBFFEAA5D2E97545FFFFC2010FFFFFFFFFFFFFFFFFF",
INIT_20 => X"0008003DF555D5157410FFFFFFFFFFFFFFDFEFF7D568A1008003DF55AAFFD55E",
INIT_21 => X"FFFF7FBE8B55AAD16AA1000516AA005D04001EFFFFFFFFFFFFFBFDF45AAD16AA",
INIT_22 => X"0000FF80155EFFFFFFFFEFF7D16AB55A2D57DEBA557FEAA10080402010FFFFFF",
INIT_23 => X"6AB45FFFBFDEBA5D7FC0155FFFFD7410FFFFFDFEFA2D16AB55A2FFFFEAA5D7FC",
INIT_24 => X"000155FFFBE8B45A2D56ABEFFFFFFFE00087BC2155087BC00AAFFFBFDF45A2D5",
INIT_25 => X"FFFDEAA552E95400002095400000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFEFF7FBFFEBA552A954105524851C7FFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"000E3DF6DBEF5D25D7FFFFFFFFFFFFBFDFEFEBF5F8E92552E9556DEBF1C2038F",
INIT_28 => X"FE3F1FAF55A2D568A0000003FF7D495155428FFFFFFFFFF7FBF8FD7EBD16AA00",
INIT_29 => X"00000002010FFFBF8FC7E3F5EAB45BEDB6FA3800556FA005504051FFFFFFFDFE",
INIT_2A => X"B7DB6FFFDEAA5571C7010FF84125EFF7F1F8FC7EBD568B6DBEDF7DEBA5571EFA",
INIT_2B => X"5092E3F1F8F55AADB6DB7DEBF1FAE82557FC516DEBF1D0410E3F1F8FC7AAD56D",
INIT_2C => X"0000000000000000000016DE3F1EAB55BEDB6FBC7EBF5F8E10007BC516D1C71C",
INIT_2D => X"FFFFFFFFFFFFFFFFFFBFDEAA5D2A954000800154000000000000000000000000",
INIT_2E => X"2A955EFAAD1400AAFFFFFFFFFFFFBFDFEFF7FFFDEAA5D2E95410550415545FFF",
INIT_2F => X"7FFEAB45A2D56AA00002EBDFFFF7D540145FFFFFFFEFF7FBFFFFFAAD16AA0055",
INIT_30 => X"5500155EFF7FBFDFEFAAD568B55AAD568A0008003DFFF0855554AAFFFBFDFEFF",
INIT_31 => X"FFFFFFFEAA55517DE10080400010F7FBE8B55AAD16AB55F7FBFDEAA08557DE00",
INIT_32 => X"10A2D56AB45A2D57DFFFF7FBFFEAA555555400F780001FFF7D16AB55A2D16ABE",
INIT_33 => X"A00087BD55FF5D5555410AAD56AB45AAFFFFFEFAAD168A00557BD55FFA2D5400",
INIT_34 => X"00000000000000000000000000000000000001FFAAD568B45FFFBFFF55A2D568",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000100",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(19),        -- Port A data input
DOA(0)   => data_read_a_lo_256(19),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(19),        -- Port B data input
DOB(0)   => data_read_b_lo_256(19),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_20_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000003",
INIT_01 => X"A75FF80000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"14088080800008400F655001FFCFF80018FA8044000000000000011000000007",
INIT_03 => X"0000000000000000000000000000000024001660380000000000000000004FF8",
INIT_04 => X"000079800014CC02C034001600000000000000101EC0012EE0C0026E1E80F000",
INIT_05 => X"1F0FF433EFF0440C3902100002203F2EFC040388137C3E20C8EEC00284033CC0",
INIT_06 => X"4400080040440C000000000017FD5F239108000155FDC0000010E40087D8787A",
INIT_07 => X"08000EE00000000000000002101FF2002C00000004018001000030817FF50C00",
INIT_08 => X"FF7FCA302C0C00082148000008405550087C0000000000000002412489808000",
INIT_09 => X"44FF60000001EFBEF0040008023FDFC00000000040062A040001071004000013",
INIT_0A => X"000000002B7C0000008000000200000200A0C0040118400FABF9000000480002",
INIT_0B => X"0000000000000000000000000000004200310000000000000000200000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000400040",
INIT_0D => X"000000200000020000004000100203FF6C000000000000000000000000000000",
INIT_0E => X"00600FFC53FF001800000002004080000000000000040900005C848538000010",
INIT_0F => X"00009A9C300020080000800000003CC0080000800000003CC020007800000000",
INIT_10 => X"000000012963C0080000800000003CC0080000800000003CC100800000080000",
INIT_11 => X"800004000000000066C5000020020000000800000000C2E18001000200000800",
INIT_12 => X"000000000052B0200000014200040C2829000400000000000860F98798000100",
INIT_13 => X"4B00400000000002958000240400000000007E1B000040200000000001496004",
INIT_14 => X"4004181800000000005C5A00000200C40808000000000AF0D80080000000000A",
INIT_15 => X"0020141812737DC3020100400001C19C1D80000200400000000000015D140000",
INIT_16 => X"04010080800801810100000000000093EDFF8020000000000001001001000080",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0020000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0C8192608486879E79E681D903000030038200010089054D460400120104D204",
INIT_1B => X"86432190C86432CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB0C30C30C30C3",
INIT_1C => X"C86432190C86432190C86432190C86432190C86432190C86432190C86432190C",
INIT_1D => X"80402000000000000000000000000000000000000000000000001007FE000010",
INIT_1E => X"FFFFFFEAA552E95400082E975FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2A954100",
INIT_1F => X"0FFFFFFFFFFFFFFFFFFFFFFFDEAA5D2A954000800001EFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"BA5D2A97400FF8017410FFFFFFFFFFFFFFFFFFFFFBFDEBA552E974105D2A8000",
INIT_21 => X"FFFFFFFFFFEFF7FBFFEAA5D2E97545FFFFC21FFFFFFFFFFFFFFFFFFFFF7FBFFE",
INIT_22 => X"DF55AAFFD5400FFFFFFFFFFFFFFDFEFF7FFEAA10000417555AAD5555EFFFFFFF",
INIT_23 => X"FDFEFAAD568A0000043DF45AAFBC2010FFFFFFFFFFFFFFDFEFF7D568A1008003",
INIT_24 => X"0001EFFFFFFFFFFFFFBFDF45AAD16AA0008003DF555D51574BAFFFFFFFFFFFFB",
INIT_25 => X"FFFFEBA5D2A95410000A00000000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFDEAA552E954000020955FFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"552A95410552485010FFFFFFFFFFFFFFFFFFF7FBFDEBA5D2E95400140E001C7F",
INIT_28 => X"FFFFFFDFEFF7FFFFEAA5D2E95400E38A17438FFFFFFFFFFFFFFFFEFF7FBFFEBA",
INIT_29 => X"7DBEDF575D7FFFFFFFFFFFFBFDFEFEBF5F8E92552E9556DEBF1C21C7FFFFFFFF",
INIT_2A => X"FD7EBD16AA00000E3DF6DBEF5D2438FFFFFFFFFF7FBFDFC7EBF1E8A00080A155",
INIT_2B => X"5492FFFFFFFEFF7F1F8FD7A2D168A1008043FF6DAAFBC5028FFFFFFFFFF7FBF8",
INIT_2C => X"000000000000000000001FFFFFFFDFEFE3F1FAF55A2D568A0000003FF7D49515",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFEBA552A95410002E820000000000000000000000000",
INIT_2E => X"2E954005D2A82145FFFFFFFFFFFFFFFFFFFFFBFDEAA5D2A954000800155FFFFF",
INIT_2F => X"FFBFDFEFF7FFFDEAA5D2E95410550415410FFFFFFFFFFFFFFDFEFF7FBFFEBA55",
INIT_30 => X"AAD140155FFFFFFFFFF7FBFDFFFFFFBFDEBA5D2A95400A2AA974AAFFFFFFFFFF",
INIT_31 => X"5A2D568A10082E955FFFFFFD7545FFFFFFFEFF7FBFFFFFAAD16AA00552A955EF",
INIT_32 => X"AAFFFBFDFEFF7FFEAB45A2D56AA00002EBDFFFF7D5400BAFFFFFDFEFF7FBFFF5",
INIT_33 => X"A0008003DFFF085555410F7FBFDFEFFFD568B45AAD16AA1008003DFEFAAFBD74",
INIT_34 => X"00000000000000000000000000000000000001EFF7FBFDFEFAAD568B55AAD568",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"FFFFFFFE00000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000000000000000000001F",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(20),        -- Port A data input
DOA(0)   => data_read_a_lo_256(20),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(20),        -- Port B data input
DOB(0)   => data_read_b_lo_256(20),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_21_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"4A302428B824900A128C090A5C1800261500213C005FE812D10420054085A202",
INIT_01 => X"081FFE3440B609703B0427F801A40B8115BC4F655300340288A40D30040E4DD8",
INIT_02 => X"0109095C30C98809800000F9FFFFFFFF149FF1FCA4C0421B182E3490DF145FE4",
INIT_03 => X"084A76341244919000099486400026523C041660BA000100CC12701015007FF8",
INIT_04 => X"000079800014CC03C075161E001118653D2408041FC004AEF000816E1C11F541",
INIT_05 => X"3F0F807BFFE000240100004683103E7FFE02482553FC3C0204EFC25010143CC0",
INIT_06 => X"C42040304101118B84E4880817FD7F028000000101FFE4036450E08247F87870",
INIT_07 => X"0A09000D00204A855B000A08A61FF20C3D004D331D3400805984B7A1FFF00860",
INIT_08 => X"F7FFC08D234B4002030314D0001104500000034089902D0901A021E4015410EA",
INIT_09 => X"B4FFE10158E1FFBEF0440021083DFFCE22DC2880E24D1BFA7C98480802000023",
INIT_0A => X"A31514636FFC00080013029811240444A82422A85180778FAFF82A04B6356DD0",
INIT_0B => X"0600E20806520398C682157A49389667126880806FF917FC30010107688862A2",
INIT_0C => X"1B2451B2451B2451B2451B2451B2451B3228D9228D90800C6120881034003631",
INIT_0D => X"0403000A01282088624001201A8C43FF7C00100102A53208B2A246406081B245",
INIT_0E => X"C4053FFD5BFF00A04A00200602CA520011000880044402104803400400189000",
INIT_0F => X"63009140094D81A5040605800B506901A3040605401360562027218196506102",
INIT_10 => X"02811209062801A3040605800B506901A50406054013605604350B812822A002",
INIT_11 => X"0B811068C00049A0A5820A3C1725A8006C0A40404D058320496C2C9C600890A2",
INIT_12 => X"AC808127C454402483153A3A895BB3C1E2E820704020381702C1AAA2C4B3F435",
INIT_13 => X"CC1B154510413CC2A200501B400A40018A00C80400040D8AA288209AA2198361",
INIT_14 => X"0141AA00418080460678A4012288463B2050302019200B00206C35901024D910",
INIT_15 => X"2440470C8A9310280C0180302A01427D060022011606E800E00169C19A00048A",
INIT_16 => X"40100448008004000000E07008010003EFFFE0373056024B0111801198823314",
INIT_17 => X"0100401004010040100401004010040100401004010040100401004010040100",
INIT_18 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_19 => X"0000000000000000000000401004010040100401004010040100401004010040",
INIT_1A => X"BEFFFFF7F7FFF3CF3CFFFF9FE0FF9FEEFF7FFDF7FF3EFC2FF8107F3DFDF7E000",
INIT_1B => X"FF7FBFDFEFF7FBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEF",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FBFDFE",
INIT_1D => X"80002000000000000000000000000000000000000000000000001007FE00003F",
INIT_1E => X"FFFFFFEBA5D2A954100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974000",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFEBA552A97400082A975FFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"AA5D2E974100800155EFFFFFFFFFFFFFFFFFFFFFFFFFEAA552E95400082E975F",
INIT_21 => X"FFFFFFFFFFFFFFFFFDEAA5D2A95400080000000FFFFFFFFFFFFFFFFFFFFFFFDE",
INIT_22 => X"74105D2A80000FFFFFFFFFFFFFFFFFFFFFBFDEBA5D2E974005D2E80000FFFFFF",
INIT_23 => X"FFFFFF7FBFDEBA552A954005D2E97410FFFFFFFFFFFFFFFFFFFFFBFDEBA552E9",
INIT_24 => X"0001FFFFFFFFFFFFFFFFFFFFF7FBFFEBA5D2A97400FF80174BAFFFFFFFFFFFFF",
INIT_25 => X"FFFFEBA5D2E97400000400000000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFEBA5D2A95410000A001FFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"552E954000020955EFFFFFFFFFFFFFFFFFFFFFFFFFEAA552E97400002E955FFF",
INIT_28 => X"FFFFFFFFFFFFFBFDEAA5D2A974101400155C7FFFFFFFFFFFFFFFFFFFFFFFDEAA",
INIT_29 => X"00552A80010FFFFFFFFFFFFFFFFFFF7FBFDEBA5D2E95400140E00000FFFFFFFF",
INIT_2A => X"FEFF7FBFFEBA552A95410552485038FFFFFFFFFFFFFFFFFFF7FBFDEBA552E974",
INIT_2B => X"74AAFFFFFFFFFFFFFFFFEFF7FBFFEAA5D2E97400412497438FFFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000001C7FFFFFFFFFFFFFFDFEFF7FFFFEAA5D2E95400E38A1",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974000004000000000000000000000000000",
INIT_2E => X"2E97400002E975FFFFFFFFFFFFFFFFFFFFFFFFFFEBA552A95410002E821FFFFF",
INIT_2F => X"FFFFFFFFFFFBFDEAA5D2A954000800155EFFFFFFFFFFFFFFFFFFFFFFFFDEAA55",
INIT_30 => X"5D2A82010FFFFFFFFFFFFFFFFEFF7FBFDEBA552A974105D0015545FFFFFFFFFF",
INIT_31 => X"FF7FFFFEAA5D2A974005D2E82010FFFFFFFFFFFFFFDFEFF7FBFFEBA552E95400",
INIT_32 => X"AAFFFFFFFFFFFFBFDFEFF7FFFDEAA5D2E954105504154AAFFFFFFFFFFFFFFDFE",
INIT_33 => X"EBA5D2A95400A2AA974BAFFFFFFFFFF7FBFDFEFFFFFFDEBA552E974000004154",
INIT_34 => X"0000000000000000000000000000000000000155FFFFFFFFFF7FBFDFFFFFFBFD",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(21),        -- Port A data input
DOA(0)   => data_read_a_lo_256(21),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(21),        -- Port B data input
DOB(0)   => data_read_b_lo_256(21),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_22_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"5290F4CDE914905A14A43D33F488243E17122300F55FEB189B343A1140548380",
INIT_01 => X"A94007B259F6A975386262000C344BA9573C6FF57B18A5FB0ABFCD3C2C5F4F0C",
INIT_02 => X"877FE30EB378008D202551040030071869D0040180AC4B685F6E26FAA0810006",
INIT_03 => X"431965109E4481D6B5AAD6875AD6AB5A1815600802888808DEA83552954D3000",
INIT_04 => X"492C0020220001010E4916C884DCD607E5EC2A344103E48003D0800023D0072C",
INIT_05 => X"00107C441001100D620A06D683018001023D37E5088043620101179092540112",
INIT_06 => X"9108E1550544A451E0CE1AA94000206B541C08414402365774611E047020008E",
INIT_07 => X"809DA02F56A92FD7247E10305C40040D136E6A023F7FCF780C4C0528800C8028",
INIT_08 => X"00803A884B5B5206B7C3391F288551002401E993AF59012740A2E4F65586923D",
INIT_09 => X"040081C91AA010000560141801002028A83D2A08E06D0002FED9680A0E002A94",
INIT_0A => X"A71514E700838460402635019FBFE7FCA13520F8D580A08044081201206334A0",
INIT_0B => X"00A0220103D2A512C6A8C4F0011550070368000A0004D0000002126F30C902A2",
INIT_0C => X"0385503855038550385503855038550392A81C2A81C00280000C200006405A08",
INIT_0D => X"0D0E153941A8B1A262CA542A9A8D6C0010A1001002C500268ACA419412503855",
INIT_0E => X"089180008800143D83888281A2034A85014280A14050A01509E050854498B294",
INIT_0F => X"6706B3C189CD84ACD20B03001E387D04AC560B02401E387E1028AC0450080410",
INIT_10 => X"0201570B036C04AC560B03001E387D04ACD20B02401E387E24708E7E242000C2",
INIT_11 => X"8E7E1C20A0106EA167C84EBF052A8E010C0180606E86C3F459DC08DA90245887",
INIT_12 => X"189980254CDEC22A98032A22C50EAC462030A01800407C2700C2ACA2C0F04470",
INIT_13 => X"CC1154C258012D86F601A2E49003400138C0DA2443A208AA612C0096C3798225",
INIT_14 => X"025483C1E0C0006B085CEC03858958D15310201015504B512044A3133004A99B",
INIT_15 => X"9512C6FC01A1421006028038720640310643858162712020B001AA415F290E16",
INIT_16 => X"110445E22022365034A8EA754008004C0200323001182122548881649D16B046",
INIT_17 => X"1044110441104411044110441104411044110441104411044110441104411044",
INIT_18 => X"0401004010040100401004010040100401004010040100441104411044110441",
INIT_19 => X"22890000000003FFFFFFFF900401004010040100401004010040100401004010",
INIT_1A => X"9EFFDFF7F5F777DF7DF7DF5FEFBFBFDEFE8FF1F7DEBD6FEFF7EF6FDF7DF7D051",
INIT_1B => X"7F3F9FCFE7F3F9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7",
INIT_1C => X"E7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE",
INIT_1D => X"00000000000000000000000000000000000000000000000000001007FE00000F",
INIT_1E => X"FFFFFFEBA5D2E974000800021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E954000004001FFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"BA552A97400002A801FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2A954100804021F",
INIT_21 => X"FFFFFFFFFFFFFFFFFFEBA552A97400082A975FFFFFFFFFFFFFFFFFFFFFFFFFFE",
INIT_22 => X"5400082E975FFFFFFFFFFFFFFFFFFFFFFFFFFEAA552E95410002A955FFFFFFFF",
INIT_23 => X"FFFFFFFFFFFEAA552E95400002E975EFFFFFFFFFFFFFFFFFFFFFFFFFEAA552E9",
INIT_24 => X"000000FFFFFFFFFFFFFFFFFFFFFFFDEAA5D2E97410080015545FFFFFFFFFFFFF",
INIT_25 => X"FFFFEBA5D2E97410080002000000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974000004001FFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"5D2A95410000A001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2A954000804021FFF",
INIT_28 => X"FFFFFFFFFFFFFFFFEBA552A97400082E821FFFFFFFFFFFFFFFFFFFFFFFFFFEBA",
INIT_29 => X"10082A975EFFFFFFFFFFFFFFFFFFFFFFFFFEAA552E97400002E955FFFFFFFFFF",
INIT_2A => X"FFFFFFFFDEAA552E954000020955C7FFFFFFFFFFFFFFFFFFFFFFFFEAA552E954",
INIT_2B => X"5545FFFFFFFFFFFFFFFFFFFFFFFDEAA5D2A974001C24975C7FFFFFFFFFFFFFFF",
INIT_2C => X"00000000000000000000000FFFFFFFFFFFFFFFFFFFFFBFDEAA5D2A9741014001",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800020000000000000000000000000",
INIT_2E => X"2A954000800021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974000004001FFFFF",
INIT_2F => X"FFFFFFFFFFFFFFEBA552A95410002E821FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_30 => X"002E975EFFFFFFFFFFFFFFFFFFFFFFFFFEAA552A97400082A801FFFFFFFFFFFF",
INIT_31 => X"FFFFBFDEAA5D2E95410082E955EFFFFFFFFFFFFFFFFFFFFFFFFDEAA552E97400",
INIT_32 => X"45FFFFFFFFFFFFFFFFFFFFFBFDEAA5D2A95400080015545FFFFFFFFFFFFFFFFF",
INIT_33 => X"EBA552A974105D0015555FFFFFFFFFFFFFFFFFFF7FBFDEBA5D2A974005504175",
INIT_34 => X"0000000000000000000000000000000000000010FFFFFFFFFFFFFFFFEFF7FBFD",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"FFFFFFFE00000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000000000000000000001F",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(22),        -- Port A data input
DOA(0)   => data_read_a_lo_256(22),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(22),        -- Port B data input
DOB(0)   => data_read_b_lo_256(22),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_23_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"EF20906D902424807BC8241BC81801B97D38AD3C0800103362A6741C80A12A02",
INIT_01 => X"001FFF8409F089003B4422000D80C80106804A7951C5B9D1C828043EA28838F9",
INIT_02 => X"073B8858218C2C50801000F9FFEFF8E72CA7F5FC2E048026496834D84721DFE0",
INIT_03 => X"2C4360101A4001001005080400401420350016E0BB222341C312000014006FF8",
INIT_04 => X"00017B810015DC03D034201E14000036486008101FC0002EE006297E1C05F561",
INIT_05 => X"BF0F817FFFE80100004044800080BEFFFC0248005FFC3C18A5FFC2444484BCC0",
INIT_06 => X"00000070604191C93F02800017FF7F002000020001FFC0832050E00047F97870",
INIT_07 => X"AE4080091A0071070FA07A1CB23FFA403F0C4D23BF7C0EF85788B681FFFC6C20",
INIT_08 => X"F7FFD8880A034AC096620C46AC5055508401A24684227DB880000008B05001A3",
INIT_09 => X"21FFE0004047FFBEF2000000001DFFC612C0C04001000BF8000000804000003F",
INIT_0A => X"000000006FFEA002020626995FBE077430001E734020DF0FAFF5080496044B51",
INIT_0B => X"0600C48907120AC81083315A49388660180082A06FF907FC3081812048006000",
INIT_0C => X"182021820218202182021820218202182010C1010C10800C6120885430003631",
INIT_0D => X"80600020040030090000012A500003FF7E081881902233483828864860A18202",
INIT_0E => X"C7043FFD5FFF00A04BC010A7724B100008000400020000415003001000400002",
INIT_0F => X"290C2909080A872BC4FC8500054840072FC0FC8440054840200705F986106542",
INIT_10 => X"0180F1082E00072FC0FC8500054840072BC4FC84400548402214A380380B2080",
INIT_11 => X"A380344920080B21810240AB182EB37C380B40800707011001B43253EE50C822",
INIT_12 => X"E4000026C00C00042BD4149067465910640A0050C060A0028063672A00019214",
INIT_13 => X"800CCB050001344060211629580B80022480A444111706658280009A2030019C",
INIT_14 => X"232D6D0100C040250200845132C10BE200403018061101A220339C800004D801",
INIT_15 => X"2A5493B8E287E03808480060E40C83C1405132C90742E408D0082140820944CB",
INIT_16 => X"00802000100100000000000004002403EFFF8002385F03490101946500140210",
INIT_17 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_18 => X"8020080200802008020080200802008020080200802008020080200802008020",
INIT_19 => X"0000000000000000000000008020080200802008020080200802008020080200",
INIT_1A => X"0000000000000000000000000000000000000000000000000040000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"80400000000000000000000000000000000000000000000000001007FE000000",
INIT_1E => X"FFFFFFEBA5D2E974100000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100004021FFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"BA5D2E954000800001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974000800021F",
INIT_21 => X"FFFFFFFFFFFFFFFFFFEBA5D2E954000004001FFFFFFFFFFFFFFFFFFFFFFFFFFE",
INIT_22 => X"54100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2A954100000021FFFFFFFF",
INIT_23 => X"FFFFFFFFFFFEBA5D2A954100800021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2A9",
INIT_24 => X"0001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA552A97400002A801FFFFFFFFFFFFFFF",
INIT_25 => X"FFFFEBA5D2E97410080400000000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800021FFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"5D2E974000004001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100004021FFF",
INIT_28 => X"FFFFFFFFFFFFFFFFEBA5D2E954000800001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA",
INIT_29 => X"100004021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2A954000804021FFFFFFFFFF",
INIT_2A => X"FFFFFFFFFEBA5D2A95410000A001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2A954",
INIT_2B => X"21FFFFFFFFFFFFFFFFFFFFFFFFFFEBA552A97410080E001FFFFFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA552A97400082E8",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804000000000000000000000000000",
INIT_2E => X"2E974100000021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800021FFFFF",
INIT_2F => X"FFFFFFFFFFFFFFEBA5D2E974000004001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_30 => X"0800021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E954000804021FFFFFFFFFFFF",
INIT_31 => X"FFFFFFFEBA552A954100004001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2A95400",
INIT_32 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA552A95410002E821FFFFFFFFFFFFFFFFFFF",
INIT_33 => X"EAA552A97400082A801EFFFFFFFFFFFFFFFFFFFFFFFFFEAA552A97410002A821",
INIT_34 => X"00000000000000000000000000000000000001EFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"FFFFFFFE00000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000000000000000000001F",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(23),        -- Port A data input
DOA(0)   => data_read_a_lo_256(23),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(23),        -- Port B data input
DOB(0)   => data_read_b_lo_256(23),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_24_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100600007FFF000080108004000800020000840041000080808",
INIT_02 => X"172A00D000EF8210000000F9FFEFF8E7240FF1FC224087B1000639401D005FC0",
INIT_03 => X"00003A2E200811000000000400000000340016603A0000004860400014006FFF",
INIT_04 => X"000079800014CC03C034001E04010850300000101FC0002EE000006E1C00F500",
INIT_05 => X"1F0F8033FFE000000000000000003E2FFC024800137C3C0000EFC00000003CC0",
INIT_06 => X"00000040004111CE08AA800017FD7F000000000001FFC0000010E00007F87870",
INIT_07 => X"001080040814210254000A00B21FF2003F2A80D5000006E461803081FFF40000",
INIT_08 => X"F7FFD88D2B4A02C0940018EB0A1000058400810205E2D8030900004D925821CC",
INIT_09 => X"20FFE0000001FFBEF0000000001DFFC002C0000000000BF80000000000000003",
INIT_0A => X"000000006FFE80000015406A80000338800002500000470FAFF0080496044950",
INIT_0B => X"0600C008140800080000100248288660100080806FD107FC3000000000006000",
INIT_0C => X"182001820018200182001820018200182000C1000C10800C6020881030002431",
INIT_0D => X"000900160000000000000000000003FF7C001001002032083020060060018200",
INIT_0E => X"C4043FFD5BFF0000410000000041100000000000000000004003000000000000",
INIT_0F => X"1080012302010049400086C02200420049400087802200412027059996516100",
INIT_10 => X"0300081406100049400086C0220042004940008780220041248190818403A042",
INIT_11 => X"90814C09C01010400132100106836001504240E01040051200200D06410C1924",
INIT_12 => X"680C0100010408240BD80008983596CD86EA84104060503C0B00002025023481",
INIT_13 => X"90164F40086000082062C1B6600BC000C300818044000B27A0043000041202CD",
INIT_14 => X"2577FE4080C08010842180C40018545BBA00301808A0810C0059AD0180200020",
INIT_15 => X"04100852B931F00800010081980B042D2044001850ED8808F00050A002C11000",
INIT_16 => X"00000000000000000000000000000003EFFF80037046031E0110001100A4820C",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"BEC99E61848655D75D7FCB598CC0AEEAF6E7CC1132CD73C8261273B444199000",
INIT_1B => X"0F0783C1E0F07BEFBEFBEF9E79E79E79E79E7BEFBEFBEFBEFBEFBE7BE7BE7BE7",
INIT_1C => X"E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E",
INIT_1D => X"80402000000000000000000000000000000000000000000000001007FE000001",
INIT_1E => X"FFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800021FFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"BA5D2E974100000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100000001F",
INIT_21 => X"FFFFFFFFFFFFFFFFFFEBA5D2E974100004021FFFFFFFFFFFFFFFFFFFFFFFFFFE",
INIT_22 => X"74000800021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974000004001FFFFFFFF",
INIT_23 => X"FFFFFFFFFFFEBA5D2E974000800001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9",
INIT_24 => X"0001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E954000800001FFFFFFFFFFFFFFF",
INIT_25 => X"FFFFEBA5D2E97410080402000000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"5D2E974100800021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800021FFF",
INIT_28 => X"FFFFFFFFFFFFFFFFEBA5D2E974100000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA",
INIT_29 => X"000004001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100004021FFFFFFFFFF",
INIT_2A => X"FFFFFFFFFEBA5D2E974000004001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_2B => X"01FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E954000800021FFFFFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9540008000",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804020000000000000000000000000",
INIT_2E => X"2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFF",
INIT_2F => X"FFFFFFFFFFFFFFEBA5D2E974100800021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_30 => X"0000021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100000001FFFFFFFFFFFF",
INIT_31 => X"FFFFFFFEBA5D2E974000004021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E97410",
INIT_32 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974000004001FFFFFFFFFFFFFFFFFFF",
INIT_33 => X"EBA5D2E954000804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E954000004021",
INIT_34 => X"00000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(24),        -- Port A data input
DOA(0)   => data_read_a_lo_256(24),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(24),        -- Port B data input
DOB(0)   => data_read_b_lo_256(24),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_25_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100200002000000080100004000000020000800041000080808",
INIT_02 => X"1000218000000800000000F9FFEFF8E738FFF1FC20400400000004455A375FE0",
INIT_03 => X"00002000000001000000000400000000340016623A0000004000000014006FFF",
INIT_04 => X"924279824C94CC1BE0B4001F20000000020380401FE0082EF000106E1C00F500",
INIT_05 => X"1F0F8033FFF048202582800100523E2FFE024820137C3C0040EFE02000003CE4",
INIT_06 => X"D4A00671414191800000800017FD7F038100201101FFC0000010E08A07FC7870",
INIT_07 => X"080000000000000000000A00B21FF2003E0000000000066041803081FFFC2C60",
INIT_08 => X"F7FFFA0008000200A0400002280000050400800204000000000201202B800000",
INIT_09 => X"B4FFF0008001FFBEF80C40630C7DFFEEBAF0008002021BF80000400A02000003",
INIT_0A => X"000000006FFF800C0400000000000330080000500006470FAFFD29F7DE565971",
INIT_0B => X"0600C008040000080000100248688760101080806FD107FC3018000000006000",
INIT_0C => X"182001820018200182001820018200182000C1000C10800EE6618911398524B1",
INIT_0D => X"000000000000000000000002500003FF7C001001002032083120060060018200",
INIT_0E => X"C6043FFD5BFF00A04B80608003CB120C11060883044582114013412080000000",
INIT_0F => X"000000200200000900000400200000000900000400200000200701E186106140",
INIT_10 => X"0000001000000009000004002000000009000004002000000000808000002000",
INIT_11 => X"8080000800000000001010000002200000004000000004000000000240000020",
INIT_12 => X"2000000001000004031802000004100000100024400000000800800001000000",
INIT_13 => X"0000410000000008000000204004000000000100040000208000000004000004",
INIT_14 => X"0004200001000200000100040000004200004020000000040000840000000020",
INIT_15 => X"00000010800000000C0A00000000040000040000004080000000000000401000",
INIT_16 => X"451044C82082068C0200000008014023EFFFC006304602080100000100000308",
INIT_17 => X"1104411044110441104411044110441104411044110441104411044110441104",
INIT_18 => X"1044110441104411044110441104411044110441104411044110441104411044",
INIT_19 => X"00002FFFFFFFFFFFFFFFFFC11044110441104411044110441104411044110441",
INIT_1A => X"042824014C48569A69AFEE9E50B2894A196A8C5A2932F7C8086034EC15DA0808",
INIT_1B => X"6231188C46231249249249249249249249249041041041041041041249041249",
INIT_1C => X"562B158AC562B158AC562B158AC562B158AC562B158AC562B158AC56231188C4",
INIT_1D => X"80400000000000000000000000000000000000000000000000001FFFFE00002C",
INIT_1E => X"FFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"BA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001F",
INIT_21 => X"FFFFFFFFFFFFFFFFFFEBA5D2E974100800021FFFFFFFFFFFFFFFFFFFFFFFFFFE",
INIT_22 => X"74100000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800001FFFFFFFF",
INIT_23 => X"FFFFFFFFFFFEBA5D2E974100000021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9",
INIT_24 => X"0001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100000001FFFFFFFFFFFFFFF",
INIT_25 => X"FFFFEBA5D2E97410080400000000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFF",
INIT_28 => X"FFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA",
INIT_29 => X"100800001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800021FFFFFFFFFF",
INIT_2A => X"FFFFFFFFFEBA5D2E974100800021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_2B => X"01FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100000021FFFFFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741000000",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804000000000000000000000000000",
INIT_2E => X"2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFF",
INIT_2F => X"FFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_30 => X"0804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFF",
INIT_31 => X"FFFFFFFEBA5D2E974100800001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E97410",
INIT_32 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800021FFFFFFFFFFFFFFFFFFF",
INIT_33 => X"EBA5D2E974100000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800021",
INIT_34 => X"00000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"FFFFFFFE00000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000000000000000000001F",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(25),        -- Port A data input
DOA(0)   => data_read_a_lo_256(25),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(25),        -- Port B data input
DOB(0)   => data_read_b_lo_256(25),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_26_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"E9264EAB20190CA3BA4997AA9002AE9C001006B0778015CFA17E0811039879C7",
INIT_01 => X"F1FFF9BB1F773C7F9BB07DFFFDD863FC5FFF3FEFFBBF9FFB22FFFBC7B9F30686",
INIT_02 => X"1B33188302E708180F6FFBFFFFCFFFFF9C7FF7FC24350B99082400001D00DFD8",
INIT_03 => X"4A53D958C50000DCE7366303739CD98C27C57EF57980014F271807E3C9E9CFF8",
INIT_04 => X"DBFAFBD7FB1CDEBEF1BE17F7AC88042787FBFFF8FEE9FF7EE6F4C0EE1FFAF869",
INIT_05 => X"5F0FFEB3EFFEFFBDA7F7FED508707E2EFEBF6FFEB37C3FF302EEEDFF9B487CF6",
INIT_06 => X"67F2B27AFAD11587B7C094F1FFFFDF0FAF4E8FAA67FDDB7FB870FF30FFDEF87F",
INIT_07 => X"08180EF060C18E5BEFB051225CDFF7002C4EEDE77F6E0EFD044ABC817FFFDD35",
INIT_08 => X"FF7FC8790E46426CE06C2C7E381041460C7E8C1A35DF80000C0084C9188302E7",
INIT_09 => X"2CFF7A27B303EFBEFAFCC2E35E7FDFD147CCF3F583FA3FFF7D6000EC75088ED3",
INIT_0A => X"5A3A3B5AFF7CFACFAFE776F39FF7077E29D83CFAE601602FEBFFCDF7DEE77DF7",
INIT_0B => X"3EB1EDDCDEBCFF589807B70AD9A99EE41FD18884FFF19FFC71FEFED7B251E747",
INIT_0C => X"1AF181AF181AF181AF181AF181AF181AF4C0D78C0D718ADEEE61D99B7BE2A433",
INIT_0D => X"B9EC20181CC1F73F87501DED3409BFFFEFFEBCEBFE68370CFA6D07407481EF18",
INIT_0E => X"CE04FFFFF3FF1F5F5475BD7F72E4D75EBFAF5FD7AFEFDFFAF59B6FF28FE1D406",
INIT_0F => X"7C040101480807D17B0004001F804007D17B0004001F8040212F35FFC6D86D70",
INIT_10 => X"0001DC00068007D17B0004001F804007D17B0004001F804006F6008140002000",
INIT_11 => X"0081800800007B000102C0801FB02683800040007700011801003DE050A70020",
INIT_12 => X"32130207080D012CEFF41008D188D502100B02004000F01900039020040206F6",
INIT_13 => X"A01F21A2C40039006823F80048100003F0008004D8100F90D162001C803403E2",
INIT_14 => X"27F020A07400007C040085581019D602451500001EC00100247C46426080E101",
INIT_15 => X"2010EA40EA00020C830100F0D000022180581019F40084800001F100020B6040",
INIT_16 => X"EFFBFEFDFDDFE7DD87FEFF7FF796FFFFFDFFC017FEFFD7E841001D8197DCC3F0",
INIT_17 => X"BFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAF",
INIT_18 => X"FAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFE",
INIT_19 => X"88646FFFFFFFFFFFFFFFFFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEB",
INIT_1A => X"86EBCAF55357E1C71C751D53C44B15BCF491E166CC853E8117696853F86EDB5C",
INIT_1B => X"130984C261309861861861861861861861861861861861861861861A69A69861",
INIT_1C => X"6130984C26130984C26130984C26130984C26130984C26130984C26130984C26",
INIT_1D => X"80400000000000000000000000000000000000000000000000001007FE000002",
INIT_1E => X"FFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"BA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021F",
INIT_21 => X"FFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFE",
INIT_22 => X"74100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFF",
INIT_23 => X"FFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9",
INIT_24 => X"0001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFF",
INIT_25 => X"FFFFEBA5D2E97410080400000000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFF",
INIT_28 => X"FFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA",
INIT_29 => X"100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFF",
INIT_2A => X"FFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_2B => X"21FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008040",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804000000000000000000000000000",
INIT_2E => X"2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFF",
INIT_2F => X"FFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_30 => X"0804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFF",
INIT_31 => X"FFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E97410",
INIT_32 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFF",
INIT_33 => X"EBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001",
INIT_34 => X"00000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(26),        -- Port A data input
DOA(0)   => data_read_a_lo_256(26),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(26),        -- Port B data input
DOB(0)   => data_read_b_lo_256(26),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_27_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"00080A40000A41248002029000050A088000008242A0004404480002000A1155",
INIT_01 => X"F1FFF1C11F781C129C107DFFFE0860941E81258CA2B71C2220EC1B86E1A00002",
INIT_02 => X"4000002100000014400FF6FFFF0FFFFF8007F1FC211100014200800000887FC0",
INIT_03 => X"0842D85841000098C63061026318C18404C459757000015F00088BE3C0618FF8",
INIT_04 => X"DBEAE5D6D91C2EBCE1B21EA72C00000007FBE7C8F8E9EF79E6D440E91FDAE061",
INIT_05 => X"5C8FFCB38FF6B68984B5BCE408347E28FEBF6FEEB3723F7102E8EDBF8A4872F6",
INIT_06 => X"6E62106ADAD14180035044F1FFFC9F0C0E4C8DAAEFF1DB7FA868FE30EF1CE47E",
INIT_07 => X"0014401060C180190310540118DFF1000C0849673F6C06FE000A38007FF13115",
INIT_08 => X"F47FC80208808210880C00020814000044008C1A340C00000A08000000210000",
INIT_09 => X"04FC721491038F7DF8BEC2E39C5F1FD047CEF1B582D83FF779200062B12A8EC3",
INIT_0A => X"02606042787C5AC5ADC424B39FB6073D00D8048A6201002F83F04DFFDE83FDD6",
INIT_0B => X"56B5F0DEFABC705488069302DBA98EAC16C1A884FFE18FFD757E7ED7A211EC0C",
INIT_0C => X"186881868818688186881868818688187840C3440C35A8DFEE61CB9979AAA433",
INIT_0D => X"D1F820101441DA3A8310198C34089BFF8DD6B56B6F28378C7E2D07007801C688",
INIT_0E => X"E4047FFD23FF315D54358D593474955AB6AD5B56ADAB5FAAE58B2F628EA0C407",
INIT_0F => X"7C0400004C080791290004001D80001791290004001D8000210F15879715710A",
INIT_10 => X"0001DC0000801791290004001D80001791290004001D800012F6008040002000",
INIT_11 => X"0080800800007B000000E0801BB020828000400077000008210035E040830020",
INIT_12 => X"220202070801010C6F1410085188D500100102004000F01900031000060202F6",
INIT_13 => X"205D2120840039000813F80040100003F0000000F8100E909042001C80040BA2",
INIT_14 => X"07F020201400007C040001781011D602040500001EC00000057444404080E100",
INIT_15 => X"2000EA40EA000004810100F0D000020080781011F40080800001F1000003E040",
INIT_16 => X"AB6BDE75ED5EC71385FC2512E3565BBBF1FFC00636EED7E841000D81924C43F0",
INIT_17 => X"B6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6AD",
INIT_18 => X"6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADA",
INIT_19 => X"88747FFFFFFFFFFFFFFFFFAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB",
INIT_1A => X"00780401CBC8400000052412F84E2168100481CA8604368008402F02104A4716",
INIT_1B => X"4020100804020000000000000000000000000000000000000000208000000000",
INIT_1C => X"140A05028140A05028140A05028140A05028140A05028140A050281402010080",
INIT_1D => X"80400000000000000000000000000000000000000000000000001007FE000028",
INIT_1E => X"FFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"BA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001F",
INIT_21 => X"FFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFE",
INIT_22 => X"74100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFF",
INIT_23 => X"FFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9",
INIT_24 => X"0001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFF",
INIT_25 => X"FFFFEBA5D2E97410080400000000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFF",
INIT_28 => X"FFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA",
INIT_29 => X"100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFF",
INIT_2A => X"FFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_2B => X"21FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008040",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804000000000000000000000000000",
INIT_2E => X"2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFF",
INIT_2F => X"FFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_30 => X"0804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFF",
INIT_31 => X"FFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E97410",
INIT_32 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFF",
INIT_33 => X"EBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021",
INIT_34 => X"00000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"FFFFFFFE00000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000000000000000000001F",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(27),        -- Port A data input
DOA(0)   => data_read_a_lo_256(27),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(27),        -- Port B data input
DOB(0)   => data_read_b_lo_256(27),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_28_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"02200AA400180030808802A900002A08001280A08A801044104A1000001818C3",
INIT_01 => X"50A00011460214428114180000882214413D0A71592A01D92213D28005210202",
INIT_02 => X"1444428102100884000AA30200000000C1000401041108404400022220800000",
INIT_03 => X"461080404900000C6314A900318C52A40051081000888806108802A141288001",
INIT_04 => X"00800040110102000902002000888400081045A8A00003C00000500000080008",
INIT_05 => X"0000000000024CA0A0101800032000400000000B800000014000000B08180000",
INIT_06 => X"0040B0000804001040000450A00080444A002480220009A88800009A88000000",
INIT_07 => X"088400122448908A204020004080010000408200000001000002080000099000",
INIT_08 => X"0000028040101004200C21002084555500004489120509244022801244810210",
INIT_09 => X"9000008101400000049016080102000220001110001020058320402A16002650",
INIT_0A => X"A53534A50000080080E041000000008000C81000220020A00004000000300003",
INIT_0B => X"0090024440245400082D0220800008000081022C0000080000206CB0821086A6",
INIT_0C => X"02C0A02C0A02C0A02C0A02C0A02C0A02C050160501600240010860CC04200280",
INIT_0D => X"1884200810C1631181500CA60400B40080720020240A00004005800800206C0A",
INIT_0E => X"0A00C000200005000010040A0020CC000200010000800920040804020A605400",
INIT_0F => X"0000000140000010290000000280000010290000000280000100180210410442",
INIT_10 => X"0000000004800010290000000280000010290000000280000002000040000000",
INIT_11 => X"0000800000000000000280000010008280000000000000180000002000830000",
INIT_12 => X"0202020000090100548000000080000010010200000000000000900000000002",
INIT_13 => X"2000202084000000480008000010000000000004880000101042000000240002",
INIT_14 => X"0080002014000000000005080000800004050000000000002400404040800001",
INIT_15 => X"00002000000000048100000000000020800800008000008000000000000A2000",
INIT_16 => X"80210810840861CD33548542A10209D4100000010200400000000880035840A0",
INIT_17 => X"0200802008020080200802008020080200802008020080200802008020080200",
INIT_18 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_19 => X"22E1000000000000000000002008020080200802008020080200802008020080",
INIT_1A => X"200360D4141D630C30C7788C0211102C110A00246972C0C19D0154BD89A40A0C",
INIT_1B => X"6030180C06030208208208208208208208208208208208208208208208208208",
INIT_1C => X"160B0582C160B0582C160B0582C160B0582C160B0582C160B0582C16030180C0",
INIT_1D => X"80400000000000000000000000000000000000000000000000001007FE00002C",
INIT_1E => X"FFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"BA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001F",
INIT_21 => X"FFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFE",
INIT_22 => X"74100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFF",
INIT_23 => X"FFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9",
INIT_24 => X"0001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFF",
INIT_25 => X"FFFFEBA5D2E97410080400000000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFF",
INIT_28 => X"FFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA",
INIT_29 => X"100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFF",
INIT_2A => X"FFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_2B => X"01FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008040",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804000000000000000000000000000",
INIT_2E => X"2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFF",
INIT_2F => X"FFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_30 => X"0804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFF",
INIT_31 => X"FFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E97410",
INIT_32 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFF",
INIT_33 => X"EBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001",
INIT_34 => X"00000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"FFFFFFFE00000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000000000000000000001F",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(28),        -- Port A data input
DOA(0)   => data_read_a_lo_256(28),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(28),        -- Port B data input
DOB(0)   => data_read_b_lo_256(28),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_29_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"79964E4BA01DACAB9E659792D00AAE160002829C7FDFEFCEE97C2815039D70C3",
INIT_01 => X"50BFF9AB0775343F9AB01DF80D5821FC0FFF3FEFD1AF9FF1207FFBC7B9720586",
INIT_02 => X"0B33180300E700080F6AAA7BFFC007189C7FF2FC003503980A0000001D00DFD8",
INIT_03 => X"0401D940CD0000C8421A2B03210868AC23403E903900010E271006A148A0C000",
INIT_04 => X"49B87A417315D20A313E17F1800000058013DDF8BE21F36E02F0D06E03E8F800",
INIT_05 => X"1F007E33E01A4D9C87525E5101603E6E023D27DA937C03E340EE25CB9B483C12",
INIT_06 => X"4570301028001487B7809450B7FFC007AB0E068023FC3BFC98101F109FC6780F",
INIT_07 => X"00080EF020408EC8CFA01122149FF700200665A35D260B250442BC8100177C20",
INIT_08 => X"FF00007906464068406C0C7E100000020C7E840A15D6800044200049180300E7",
INIT_09 => X"A8FF18222341E0820AD40201423FC00122C4935001722BFD056040A452000443",
INIT_0A => X"5A2A2B5AAF00A80A82C332D18ED301D229C82C7AA600402FE80B8813485534A2",
INIT_0B => X"28102D445624DB481806A628810018400B9100042FF0180000ABFEF892508545",
INIT_0C => X"00D1A00D1A00D1A00D1A00D1A00D1A00D4D0068D006000428200508A0A600280",
INIT_0D => X"B0E8201018C1561E855008C50401B7FFE27A08A0B64A0100CA45814814A04D1A",
INIT_0E => X"4400DFFFF0001F1F0050342D42A086040B02058102C48970541944B20FA15402",
INIT_0F => X"00000101480000507B00000002804000507B000000028040212034FAD2892832",
INIT_10 => X"00000000068000507B00000002804000507B0000000280400402000140000000",
INIT_11 => X"00018000000000000102C0000410068380000000000001180000082010A70000",
INIT_12 => X"12130200000D0120ED64000080800002100B0200000000000000902004000402",
INIT_13 => X"A00220A2C4000000682008000810000000008004D80001105162000000340042",
INIT_14 => X"208000A074000000000085580008800045150000000001002408424260800001",
INIT_15 => X"001020000000020C8300000000000021805800088000048000000000020B6000",
INIT_16 => X"C4B12C989489418D13FE7F3FFD8BADB7FC004012CA5141600000198087D8C0F0",
INIT_17 => X"0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02",
INIT_18 => X"B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C",
INIT_19 => X"00602FFFFFFFFFFFFFFFFFC0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0",
INIT_1A => X"AEFFFFF7E7EFBFFFFFFAEF1DE1EF9F96EE7FFDF7FE78FC2FE8847F3FFDFFEA0C",
INIT_1B => X"F7FBFDFEFF7FBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBAEBAEBAEBAEB",
INIT_1C => X"FF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEF",
INIT_1D => X"80400000000000000000000000000000000000000000000000001007FE00003E",
INIT_1E => X"FFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"BA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001F",
INIT_21 => X"FFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFE",
INIT_22 => X"74100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFF",
INIT_23 => X"FFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9",
INIT_24 => X"0001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFF",
INIT_25 => X"FFFFEBA5D2E97410080400000000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFF",
INIT_28 => X"FFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA",
INIT_29 => X"100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFF",
INIT_2A => X"FFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_2B => X"01FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008040",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804000000000000000000000000000",
INIT_2E => X"2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFF",
INIT_2F => X"FFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_30 => X"0804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFF",
INIT_31 => X"FFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E97410",
INIT_32 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFF",
INIT_33 => X"EBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001",
INIT_34 => X"00000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(29),        -- Port A data input
DOA(0)   => data_read_a_lo_256(29),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(29),        -- Port B data input
DOB(0)   => data_read_b_lo_256(29),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_30_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"9EEBFEF5D7D7F7DF7DFFDFDFCEFFBFFEFF9FE1F7FFBFEFC9B77B7FFFFDFFD000",
INIT_1B => X"7F3F9FCFE7F3F9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7",
INIT_1C => X"E7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE",
INIT_1D => X"80400000000000000000000000000000000000000000000000001007FE00000F",
INIT_1E => X"FFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"BA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001F",
INIT_21 => X"FFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFE",
INIT_22 => X"74100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFF",
INIT_23 => X"FFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9",
INIT_24 => X"0001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFF",
INIT_25 => X"FFFFEBA5D2E97410080400000000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFF",
INIT_28 => X"FFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA",
INIT_29 => X"100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFF",
INIT_2A => X"FFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_2B => X"01FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008040",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804000000000000000000000000000",
INIT_2E => X"2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFF",
INIT_2F => X"FFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_30 => X"0804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFF",
INIT_31 => X"FFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E97410",
INIT_32 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFF",
INIT_33 => X"EBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001",
INIT_34 => X"00000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(30),        -- Port A data input
DOA(0)   => data_read_a_lo_256(30),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(30),        -- Port B data input
DOB(0)   => data_read_b_lo_256(30),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_31_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"129000008004A00804A40000400800020000000C005FEA005800200400050100",
INIT_01 => X"A15FF18019700810180065FFFC0040801E80258CA2951C2200EC0906A0804140",
INIT_02 => X"0000000000000011000550FDFF0FFFFF0007F1FC200000011000000000205FC0",
INIT_03 => X"08425818000000908428C0024210A30004045060302223490002014280410FF8",
INIT_04 => X"DB6A618248140C18E0B016872400000007EBA24058E1ECA8E2D400681FD0E061",
INIT_05 => X"1C0FFC338FF01009048084C400103E28FE3F6FE513703F7000E8E5B4825030F6",
INIT_06 => X"4420006040410180034000A157FC1F08040C080045F1F2572060FE82671C607E",
INIT_07 => X"001100004081001103107000185FF0000C0849673F6C06FC000830007FF00000",
INIT_08 => X"F47FC80008000200800000020811000004008812240800000800000000000000",
INIT_09 => X"04FC700090038F3CF82C44630C5D1FC002CCE08082481BF27A00000000000883",
INIT_0A => X"00000000687C0044040424B39FB6073C0010048A4000008F83F009F7DE037DD0",
INIT_0B => X"0620E08812982050800A910249298624124080886FE187FC301B124F20016000",
INIT_0C => X"182001820018200182001820018200183000C1000C10808EE661891139802431",
INIT_0D => X"816800100400902A0200110810080BFF0C8010010220330C3A28070070018200",
INIT_0E => X"C4043FFD03FF101D400080013040180810040802040102004183012084808006",
INIT_0F => X"7C04000008080781000004001D00000781000004001D0000200F018586106100",
INIT_10 => X"0001DC0000000781000004001D00000781000004001D000002F4008000002000",
INIT_11 => X"0080000800007B00000040801BA020000000400077000000010035C040000020",
INIT_12 => X"200000070800000C231410085108D500000000004000F01900030000040202F4",
INIT_13 => X"001D0100000039000003F00040000003F000000050100E808000001C800003A0",
INIT_14 => X"077020000000007C0400005010115602000000001EC00000007404000000E100",
INIT_15 => X"2000CA40EA000000000100F0D000020000501011740080000001F10000014040",
INIT_16 => X"010044602002061004A820104809402BE1FFC006304E03684100050190040350",
INIT_17 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_18 => X"0040100401004010040100401004010040100401004010040100401004010040",
INIT_19 => X"00802FFFFFFFFFFFFFFFFF810040100401004010040100401004010040100401",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000010",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"80400000000000000000000000000000000000000000000000001007FE000000",
INIT_1E => X"FFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"BA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001F",
INIT_21 => X"FFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFE",
INIT_22 => X"74100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFF",
INIT_23 => X"FFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9",
INIT_24 => X"0001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFF",
INIT_25 => X"FFFFEBA5D2E97410080400000000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFF",
INIT_28 => X"FFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA",
INIT_29 => X"100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFF",
INIT_2A => X"FFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_2B => X"01FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008040",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804000000000000000000000000000",
INIT_2E => X"2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFF",
INIT_2F => X"FFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_30 => X"0804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFF",
INIT_31 => X"FFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E97410",
INIT_32 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFF",
INIT_33 => X"EBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001",
INIT_34 => X"00000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(31),        -- Port A data input
DOA(0)   => data_read_a_lo_256(31),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(31),        -- Port B data input
DOB(0)   => data_read_b_lo_256(31),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_0_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"ED39BA795990D275FB4A6E96ACC4731DEA4598B0AFB54867F6EE4618C3749807",
INIT_01 => X"58A0047D8607944AC7DA180001ECA2544042106208408208C20022E9173734B3",
INIT_02 => X"9F775E7CB273E6CCA7DAAF00001000000478020113C9C38E09FB7CCCDD9F203E",
INIT_03 => X"441406267B4CB04443163C91110C58F24A31000B8028A810A3D0F8B169A01006",
INIT_04 => X"0005802424830120024121209088809DF81454ACA01E03501D0A3B91E00F0A00",
INIT_05 => X"E0F001CC00012034C20B0232838F80D001C0100AEC83C008EF101A034C8CC300",
INIT_06 => X"908A0D058584A45164BE6E58A000000583F08459A2000DA8C40F003C80030780",
INIT_07 => X"E6CCAFDC3870EEEEC44E2BDFE220094D03022210C011C103FB860B28000007C9",
INIT_08 => X"080032BF07C7C1FC3F87253D96C45557ABFF070C19D62C9065EAF36919FCB273",
INIT_09 => X"DB0009EF68EC0000045082984202002DB93119096025040581B9691E8A88262C",
INIT_0A => X"8014546E000344A0488111084048E082D0ED020133A6BF200005F60820B88206",
INIT_0B => X"28000947E16656074EA560F08054490B01280A26900C4800814069B0C8888008",
INIT_0C => X"03DCF03CCF03DCF03CCF03DCF03CCF038E780C6781C008500804708A42255A88",
INIT_0D => X"7095352BD2A90515A1CA44E7EA84B00001010012008700624187C09C0E707CCF",
INIT_0E => X"0B92800224008AE09F8942C48D1BC49120489024481225058860128543287291",
INIT_0F => X"038ABACB83C7E03EA5FF83C002783F103EA5FF83C002783F0120847A70470C7E",
INIT_10 => X"0380230F2D7C103EACFF83C002783F103EACFF83C002783F310BBF7EFC2B80C2",
INIT_11 => X"BF7EFC61E01804E1E6EA1E3FA01FD97EFC4B80E008C7C2F678FF023FAF5BD987",
INIT_12 => X"CC8E8320C4DAC9220C6B2FF22EF72ADDE6F1A67C80600C2683E0EF8AE1F1F10B",
INIT_13 => X"5C00FE651C6104C6D6400FFFB01FC0000FC07EE42FA7C07F22CE3082636B801F",
INIT_14 => X"C08FDF4195C0C2038A7C6CAFA7E289F9BA4570380131CAFB2003F9D190A4189B",
INIT_15 => X"9FE635BE11B7F0308D4A80092E0FC1FC662FA7E283FF68A8F0080AE1DDA8BE9F",
INIT_16 => X"12058312C1241140A056954AB0D680D000003350013024179498C2EC6B9270AE",
INIT_17 => X"2048120481204812048120481204812048120481204812048120481204812048",
INIT_18 => X"0481204812048120481204812048120481204812048120481204812048120481",
INIT_19 => X"2859400000000000000000120481204812048120481204812048120481204812",
INIT_1A => X"082218821390771C71C557C449F3898E09B56C74DAB16787E0760E5D1CF13043",
INIT_1B => X"7C3E1F0F87C3E082082082082082082082082082082082082082082082082082",
INIT_1C => X"87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F8",
INIT_1D => X"D7BD7400000000000000000000000000000000000000000000061007FE00000F",
INIT_1E => X"A2D1574005D0428A10A2AAA8BEF552EBDFFF557BC01FF5D7BFFEBA5D55555EF5",
INIT_1F => X"AFFFFC2000AA8428AAAFFAAA8BFF00002AA10FF802ABEFA2D16AA00F7FBE8A10",
INIT_20 => X"EFFF8002010002EAAAAAAAD1555FFFFAEA8B550051401450055575FF00517DEB",
INIT_21 => X"5FF0855575455D2AA8BFFA2D1575EF5D5555545FFFBE8A00087FC20BA5D2A975",
INIT_22 => X"8A00FFAE800AA082A820005D2E974BAA2D140145A2842AA00A284021FF5D0415",
INIT_23 => X"7FFEF000017400FFD1555FF007FFFEBA55042AA00000017400FFAABFEBAFF802",
INIT_24 => X"000155F7D540000F7FBFFE105D7BE8ABAA284000105D0428BFFA2FBFDFFFA2D1",
INIT_25 => X"7BFAEBA5551501D51C5FC7E00000000000000000000000000000000000000000",
INIT_26 => X"6D16AA28EBF5EDA38AADE1543849557D492BF8E2DE00552EBFFC7552BC01D75D",
INIT_27 => X"A85400E00E38A175FDE3F5C002DAAD42DAAAF784AFA82BC042DF47E3D1F8028B",
INIT_28 => X"50021C0092490E904BAFFD550A90FFA495FC7A05B555C257AAA8B45007540000",
INIT_29 => X"02402ABD4AD1D0E175D7140B455D516A1EAB45E2A000B4748717A095F571EAA1",
INIT_2A => X"4A8BC0ABFF7D03A17D1D5147540B454AA080038E9748542AE3D0051C7B6F02DA",
INIT_2B => X"D4B8FC7BFFFD2168B68F57492F505FF5FA550490BFA482B420B8428A3DA85400",
INIT_2C => X"0000000000000000000016ABD554201543A1EDE9016D4AAB454AF400547ABFB6",
INIT_2D => X"EBDF55556BC35E7557FE8AB25D11415FD0151614000000000000000000000000",
INIT_2E => X"6CBEA41D7D3DECFAF7D43FABAAAD57DEBAAAFFD74AA04547EE18D680BE9A55D2",
INIT_2F => X"78228E5000EA422E10439C1FBCD282351BDAAF9C20AAAABCBEB1DFF803FC5959",
INIT_30 => X"284683ABBDD7DEAA100069C14B25495A00F38EBAC0E198B9760501805357547D",
INIT_31 => X"8FE6A755ED8EFEFE41B2D17EAF02552BC0545556BD61E501001DF5DD3EBA31E6",
INIT_32 => X"F922ACA8AB8283C8310FAB1588916D3861C0422C44082B52A81550A828141440",
INIT_33 => X"DBCD7D262E5AFAC4B6AADDD562AF57D7C369AF25495A23068A8301BA7FB95556",
INIT_34 => X"FE0000003FE0000003FE0000003FE0000003FE03D5789700282E9FEFB501EA5F",
INIT_35 => X"3FE0000003FE0000003FE0000003FE0000003FE0000003FE0000003FE0000003",
INIT_36 => X"00000000000000000000000000000000000000000000000000000003FE000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000020",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(0),        -- Port A data input
DOA(0)   => data_read_a_hi_256(0),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(0),        -- Port B data input
DOB(0)   => data_read_b_hi_256(0),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_1_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"212C001411984004084D000508C53810A03D1450E839B003342114428A000807",
INIT_01 => X"08000010400A0008010600000084004000400002000000000000000000140000",
INIT_02 => X"484DEBA0111800C004400D000000000028800001CC404E6008B4933336880010",
INIT_03 => X"650C00000848A0423183089008C604224200000100A200002C280810098C0001",
INIT_04 => X"00000004208B00200E010800006667BE7000102C00080000040012010000080C",
INIT_05 => X"0080000000002020600100208D04414000800000000200004800080000800200",
INIT_06 => X"0000CB008084001C481040080000006050402008080000800488000000020400",
INIT_07 => X"00C00843060C19E2300221036000004400208000400041034001042000000101",
INIT_08 => X"08000290248CC84E0801318000C45555087C60C182B1592FE26AD7B7F7A01118",
INIT_09 => X"D8000AA220480040050080085200001161020001202100008008611687A28000",
INIT_0A => X"2640440000000080081040000040208300041000008004104006840000B80004",
INIT_0B => X"78051112A80000840200202112800001010828008000000105400020082800A8",
INIT_0C => X"2358323483234832358323583234832340190AC191A52801000C1002020883C2",
INIT_0D => X"4417882F82C00181707044212080300001002102010244800400C80C80323183",
INIT_0E => X"0B92C000000000400001004200004010200810040802040080200284401C1C11",
INIT_0F => X"00000043C2016000000F03C00280030000000F03C00280030000004860C60C0C",
INIT_10 => X"03800000049C0000000F03C00280030000000F03C002800321080000BC2380C2",
INIT_11 => X"00007861E0180000002A9001A00000007C4380E00000001E002300000008D187",
INIT_12 => X"4C0C81200009480010280340000008082430A07C80600C000000900861001108",
INIT_13 => X"34400241186100004A500007B00FC000000000E4A402C001208C308000268800",
INIT_14 => X"C0001E0181C0C200000025A400A200812A4070380000000B2500098190240001",
INIT_15 => X"04A0002410A170300C4A800800000020E22400A200096828F008000000AA9002",
INIT_16 => X"0200820040041002000010080014000000002340002004118010C22861400008",
INIT_17 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_18 => X"0080200802008020080200802008020080200802008020080200802008020080",
INIT_19 => X"0A04000000000000000000020080200802008020080200802008020080200802",
INIT_1A => X"8AB2048634B03249249604C061028A46BABEFC54A08170062002340C7452B500",
INIT_1B => X"DD6EB75BADD6EAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA8A28A28A28A2",
INIT_1C => X"A5D2E974BA5D2E974BA5D2E974BA5D2E974BA5D2E974BA5D2E974BA5D6EB75BA",
INIT_1D => X"AAAAAA00000000000000000000000000000000000000000000181FFFFF00000B",
INIT_1E => X"5D7BE8ABA5D557DFEFFFD17FEBA00042AAAAFFFFFFE00FF843DF45FFAE95555A",
INIT_1F => X"F552A800AA5555575FFA2AE820BAFFAEBFF555500155EF552E975FFF7D168BEF",
INIT_20 => X"00A2FBEAABA5D55420AA00002AA00AAFBE8B55A280175455D002AA00A2AABDFE",
INIT_21 => X"5FFAA802AAAAFFAA801EF00517FFFFF7D56ABEF0004155550004154105D556AA",
INIT_22 => X"75FF08557DEBAA2FBEAAAA552E955EF5D0415410A2AE97545A2AE954BAF7FBD7",
INIT_23 => X"7DF55A2AEBDEAAFFFFC20AAFFFFFFFFFAAD5555FFFFAEAAB55A2D168B555D555",
INIT_24 => X"0000BAFFFBE8A00087FC20BA5D2A975EF5D0002010552E820AAFFD57FF55F7D1",
INIT_25 => X"8A38F45F7AA9217FA380AD400000000000000000000000000000000000000000",
INIT_26 => X"52E975EFFFDF68BFF557BEAA925551785D7BFD5EFE3F08002FA92EBA5FDE28FF",
INIT_27 => X"41017DE92BF8E3AA824924870BF5551555C7A28A821EFE3AABAE38005B575D75",
INIT_28 => X"8005A1041055716DB7DB6FBEFEA81C55D0A0516802AA28BEF5EDB7DAA8A15438",
INIT_29 => X"EF1C043FE28E3FBD55FFAADE2DAAAE3A5C51C71C042DF45A3D1D00281E8A1056",
INIT_2A => X"B45B47F6FB55A95555E90F78E17F52FEF5EDA82FD249057F080417492AAAFC7F",
INIT_2B => X"8AAAA95B7AF45FF8F7DFEDFFAFF8E005FAE92A3AE3DBFF57FA2DF555D257AAA8",
INIT_2C => X"000000000000000000000A8F571EAA150021C0092490E905FFFD0550BD75C5FF",
INIT_2D => X"43DE00A2C57DE08FFAAA8B55F7EE801F7F2849EE000000000000000000000000",
INIT_2E => X"AE29F067155543A15D2E955EFFFFBEABEF557FEAA10595169BED83D1EBCA8000",
INIT_2F => X"FD57DEEAAA15976EB0444BFEB086808A8E3082C954BA5D7DD6145AAAA821A6AA",
INIT_30 => X"FFD55D6107782001FF0812000A255D57FFBEF3B97EEAB2C40217B9778428ABAF",
INIT_31 => X"F003F17418AEE817B540D11CA80BAAFA825EFAABEBCA18FE803755D08079EB47",
INIT_32 => X"EBA2D757547D7862AF57ABFFCABE5553FD5FBEFE86353EFFFD03FE027500035F",
INIT_33 => X"1F70C6AA04537957D6FB4807FFFB45F7EFFDA58FF2AA88A0F3C5014018AC28BD",
INIT_34 => X"00000000000000000000000000000000000000B2DD7DEAA100069C14B25495A0",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000020",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(1),        -- Port A data input
DOA(0)   => data_read_a_hi_256(1),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(1),        -- Port B data input
DOB(0)   => data_read_b_hi_256(1),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_2_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10E44660018259B2843913100062C98004802322D3E030235201006009B2812",
INIT_01 => X"8005A188084900481C8024A542400340404000720885800802000906E4910204",
INIT_02 => X"5C010802020408040C640850AA055254090541A111240A104A0000000908B510",
INIT_03 => X"0C1101108800004481060A001204102802156020218808002440850008C80550",
INIT_04 => X"8840C08022050400482812C21C0804040968987810688899444090C10A124A69",
INIT_05 => X"4885109105400029210000010340086856B141212252142242A068A080106372",
INIT_06 => X"0082006020044004C240108005540A400440880000908281302852A6710AA420",
INIT_07 => X"08040860400008C022402502100AA00004404B5075460111044014002AAA2100",
INIT_08 => X"382A885244145048C860214020040505487C0800049000004220000110820204",
INIT_09 => X"88582833A24105145404D4694E710A832488C000002205C23600408C872A2A12",
INIT_0A => X"A211100D0828800A022025A81AE3048228002A7080012082C15C859D5073D520",
INIT_0B => X"3E00659A308809540009202A5820068019108A88B1D007285082002B10416820",
INIT_0C => X"1A0021A5021A1021A5021A1021A4021A0010C2010D010887470912171342A683",
INIT_0D => X"89180010084038220410042B2000715A0400200080623400380886086021A002",
INIT_0E => X"40000554015500481000300000C4480810000002040000000913000004C18402",
INIT_0F => X"00000001440002C052000400028000154052000400028000200501CCD28D206A",
INIT_10 => X"00000000048015405200040002800012C05200040002800014E0000100002000",
INIT_11 => X"00010008000000000002A0000D80060100004000000000180000294010240020",
INIT_12 => X"1011000000090000A310000881080102000A0000400000000000900002000684",
INIT_13 => X"204E008240000000483250000800000000000004E00007004120000000240A60",
INIT_14 => X"254000806000000000000560000942004110000000000000254C020220000001",
INIT_15 => X"00108840600002080200000000000020806000093000040000000000000B8000",
INIT_16 => X"008022200100000020A89068084D402120AAC005C00000000000000005408140",
INIT_17 => X"0802008020080601806018060180200802008020080601806018060180200802",
INIT_18 => X"8040080000800008000180401804018040080000800008060180601806018020",
INIT_19 => X"A2852F81F81F83F03F03F0018040180401804008000080000800018040180401",
INIT_1A => X"04609D21808205965965D64CC5B60040138D70C030B54284722B291C50C7D100",
INIT_1B => X"4A25128944A25041041041041041041041041041041041041041041041041041",
INIT_1C => X"44A25128944A25128944A25128944A25128944A25128944A25128944A2512894",
INIT_1D => X"055400000000000000000000000000000000000000000000001E1007FFE3F009",
INIT_1E => X"FF843DF45FFAEBDF55082A82155082AAAA10F7FFEAB455500175FF5D2A800100",
INIT_1F => X"F082ABDF455D7BD5545F7D5574BAFFD16AAAAA28428ABA000428AAA5D7FD7400",
INIT_20 => X"455D7BEAABA5D2A97545552E975FFFFD168AAA5D7BE8BFF5D557FFEFFFD16ABE",
INIT_21 => X"5555555555FFA2AE820BAFFFFEAABA5555554BA5D0417545F7D56AAAAAAFBEAB",
INIT_22 => X"AA00AAAEBDFFF08042AABA087BD54BA08043DEAAFF843FF5508517FF55552A95",
INIT_23 => X"82010AAD1401FF002EBFF45A2FBFDFEF00042AA00AAFBEAB5500003FF5500002",
INIT_24 => X"0000BA0004155550004154105D556AA00A2FBEAABA085542145082A800BA002A",
INIT_25 => X"00155FF552A87410007145400000000000000000000000000000000000000000",
INIT_26 => X"8002FABA4171D5400FF8A38F45F7AABA57D0000855FD1C2AAFA00EBA5E8B7D55",
INIT_27 => X"555178FD7BFD5FDFFA0020BFF78417BD5545F7F1554AAF7D16DABABFF57DE920",
INIT_28 => X"DFFDF6DAAAAAF1EFB6D417BEFA901C2E97F40552E975EFEBDF68ABA557BEAA92",
INIT_29 => X"7DA3FBD21C7492E9256D555B555C7A2ABC20AAE3AABAE38005B574AA49041756",
INIT_2A => X"B7D1E803AF6D400028E02AB8A3A012540E2AABABC75D043A00003FE10E3802DB",
INIT_2B => X"8B7D0AAA800AA147085000FFDA001C7B47BFABC7BFFF7AB4714042AA38BEF5ED",
INIT_2C => X"000000000000000000000821E8A10568005A1041055716DA38B6FBEFFEF1C0EB",
INIT_2D => X"EBDE00AAC16ABEF5500155EF552A954000855544000000000000000000000000",
INIT_2E => X"D57DE0AFAD1EBEB400043DEAA085555400FFAAAAB55F7AEA8BF77004147EF5D2",
INIT_2F => X"AFBEABAF557FEA8515951E8B4D83D1EBDFF082CBDFEF005756145FFD5574AAF7",
INIT_30 => X"5951550100004155EFF7FFFDE08AA557FFFF083FFCEB95104210405D2E955EFA",
INIT_31 => X"A002A3FE18AE803CBE7A3C014351082E951FF5D7FD6145AAAA820A2AAAD29E00",
INIT_32 => X"45550028ABAFFD17FFED01001FFEF5542ABEB2AA848AAA2552EA8ABA7551400A",
INIT_33 => X"EBAF3F95EEE95C00B7CF12AAA800BA551417105FFFFC21555556EAB4CD6D5EAD",
INIT_34 => X"00000000000000000000000000000000000000187782001FF0812000A255D57F",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000040",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(2),        -- Port A data input
DOA(0)   => data_read_a_hi_256(2),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(2),        -- Port B data input
DOB(0)   => data_read_b_hi_256(2),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_3_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"210C00A20020000108430020001600B815602110494074133520400E02B92206",
INIT_01 => X"A00C9BC048800168240442C99E004B61404040028804A0080A000D16A0990A08",
INIT_02 => X"4809A902031800444445089866E331352180D468B8200E600C0081110B80ACD0",
INIT_03 => X"6D0A60100C000142B1A30A040AC68428320006010A80881068A80D401C846330",
INIT_04 => X"482218076809C03B24841CD92CDD5A440209127847294C042640102107102D04",
INIT_05 => X"0583180353202129000104E40B04644B32A86D24014A0D204063297092000E34",
INIT_06 => X"0120D000808040181B5000A014CC662814442808805A52C03068280004629414",
INIT_07 => X"00444841428409C038B02523041994001C644C82732001190000B400E6640901",
INIT_08 => X"E8E64010248C4A5AA040308000440005487C285284B1D00BC22AC005B2820318",
INIT_09 => X"A8D588362040534C3B0E80A9DB742641620AC281826816925040408483008A10",
INIT_0A => X"040450A1439800840C32264119D004860110104004010001E732C0DF80F3B174",
INIT_0B => X"7C8575909088A4D010202422520090840B4028209AC1111954DA902230010002",
INIT_0C => X"032920329203692036920329203392036C900BC9019528100A0D30024BC8A283",
INIT_0D => X"446A101C05C0088A42D001032000333931001902010234888C68804808A03692",
INIT_0E => X"8601CCCC8B33004C0001004240140018380818040A0706009000028000903401",
INIT_0F => X"00000120000006000000000020004011000000000020004010072CC92416414C",
INIT_10 => X"0000001002001400000000002000401380000000002000401070000000000000",
INIT_11 => X"00000000000000000110000001A0000000000000000005002000244000000000",
INIT_12 => X"00000000010402049910000011000500000000000000000008000020000002C0",
INIT_13 => X"805500000000000820133000000000000000810000000C000000000004100B20",
INIT_14 => X"0530000000000000000180000011060000000000000001040154000000000020",
INIT_15 => X"0000820062000000000000000000040100000010700000000000000002400000",
INIT_16 => X"0680C2A05104100280A8D06C004044230B998021002004000001011000380000",
INIT_17 => X"280C0280C0280803808038080380803808038080380C0280C0280C0280C0280C",
INIT_18 => X"00C0280E0200C0280E030080380A030080380A030080380C0280C0280C0280C0",
INIT_19 => X"8A145D54AAB556AA9556AA830080380A030080380A030080380A0200C0280E02",
INIT_1A => X"04A20E858000049249240540430303C0C78C706428A141046016224C58629502",
INIT_1B => X"EA753A9D4EA75249249249249249249249249249249249249249041041041041",
INIT_1C => X"46A351A8D46A351A8D46A351A8D46A351A8D46A351A8D46A351A8D46A753A9D4",
INIT_1D => X"A8400000000000000000000000000000000000000000000000001007FEB6FECD",
INIT_1E => X"5500175FF5D2AA8A10005540155087BEABFF552ABDF45A2D16AAAAF7D540000A",
INIT_1F => X"000556AB55552ABDE00AAD140010F7D17FF45A2AA82155082AAAA10F7FFEAB45",
INIT_20 => X"55557FEAA10007FEAABA000428AAA557FD7400FF843DE00FFAEBFF55082A8201",
INIT_21 => X"A105D7BD5545F7D5574BAFF802AA00A2D168ABA085568BEFFFAE820000855421",
INIT_22 => X"FFEFF7D56ABEF557BD74BAFF8402145A2AEBFFEF552EAAABA5D0028BEF082AA8",
INIT_23 => X"3DEAAAAAA95410F7803FFFF55556AAAA552A975FFFFD16AAAA5D7BC01EF5D557",
INIT_24 => X"0000105D0417545F7D56AAAAAAFBEAB455D7BEAABA5D2A974005D55574005504",
INIT_25 => X"DF6FABAFFD547010AA8407400000000000000000000000000000000000000000",
INIT_26 => X"C2AAFA28EBF5E8B7D5500155FF552AAF0100071455451C75EABC74174BAF55B6",
INIT_27 => X"F7AABAF7D00009543D1C556AB6D4124BAE10BED542010FFD57AF55AAF5D756D1",
INIT_28 => X"FEBA0870281C5F4716D5D7FEDA3A0955FF48208002FABA4171D5400FF8A38F45",
INIT_29 => X"BA15203FFFF002AAFA384171D5545F7D0154AAF7D16DABABFF57DE92005F6ABF",
INIT_2A => X"ABA417BC01D7555178FD7BFD5FDF571575D24BA438E021D5B6A4BAFFF5D2EB8E",
INIT_2B => X"FE005D5B52428410E3AE92E3A490410EB843ABD71551FFE02552A975FFEBDF68",
INIT_2C => X"0000000000000000000003849041756DFFDF6DAAAAAF1EFB6D417BEFBD71C24B",
INIT_2D => X"56AB45081028B55FFFFFFEBAFFD557400A280144000000000000000000000000",
INIT_2E => X"D56ABF5AAD15455F5D2EBDEAAA2D16ABEF5500175EF552ABDE000855545455D5",
INIT_2F => X"85555400FFAAAAB14F7AE28BF77004146BA557DEABEF00002BE10FFD540000FF",
INIT_30 => X"F2D1EAEBA007FEABEFAA84174BA557FD55EF5D3BFEEB35055DEE1000043DEAA0",
INIT_31 => X"5FFAA28BF7592EABE0A0804ABFFB082EBDEAA005556145FFD5574AAF7D47DE0A",
INIT_32 => X"105D2E955EFAAFBE8AAA547FE21550853E8B4FABD5EBFF75D55420AA82AA8015",
INIT_33 => X"FFF087FFCEF90104B780A557FC20AA082AAAE10AA8000000A2AC2ABFD2151EB8",
INIT_34 => X"00000000000000000000000000000000000000AA0004155EFF7FFFDE08AA557F",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000020",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(3),        -- Port A data input
DOA(0)   => data_read_a_hi_256(3),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(3),        -- Port B data input
DOB(0)   => data_read_b_hi_256(3),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_4_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10804002061080A284201081034809800A00230350007833422C82904204006",
INIT_01 => X"204398001038084C0420050E12100368403008418984014902030906A0910204",
INIT_02 => X"480108A000000000446118E01E80F00A41043118680402000800000009882390",
INIT_03 => X"065140108C0000400026480000009120270072E03000000030808840888100F0",
INIT_04 => X"9100EB826A155C1AF0B81C160033B9440222BA281AE0D8B8E02010E81C22E821",
INIT_05 => X"5C0F20B36F08010924C084C501441C4CF21C48B133483C8042EAE1E0101074C4",
INIT_06 => X"010290102005118043508020543C1E480002820085D9C0C70000F2AA375A6071",
INIT_07 => X"00000860008008D200102502000786000C00C8025C00091B0400B00061F84020",
INIT_08 => X"991E02100C84C0480020010000004404087C8010009800004022800110000000",
INIT_09 => X"B83D6A2620418F7CF8084082425D01D123C2C040816A00708840408483000011",
INIT_0A => X"BB1B585C1304E002000064010E4007F7210010500400400800F0CC249C1401C1",
INIT_0B => X"7A04331814080458100134201A2086441B50A088078106C14540906D004068A0",
INIT_0C => X"186921829218692182921829218692182090D3490C352296CC60B11357088682",
INIT_0D => X"411050002500A9200A8014010001370F03080980912204883C28864860A18A92",
INIT_0E => X"C40903C1430F20025040102200441A040906008300418050501341208002A005",
INIT_0F => X"0000012004000BC01200000020004008C012000000200040000721CD86146108",
INIT_10 => X"0000001002000A40120000002000400DC01200000020004004D4400000000000",
INIT_11 => X"40000000000000000110200007600401000000000000050020005D4010040000",
INIT_12 => X"1010000001040004A3B000018008850200080000000000000800002002000650",
INIT_13 => X"80360082000000082034300000000000000081004000170041000000041005E0",
INIT_14 => X"2B200080400000000001804000192000401000000000010400F8020200000020",
INIT_15 => X"00114A00200002080000000000000401004000085C0000000000000002410000",
INIT_16 => X"459040281181004A8088986D045C24436C7840A6180300082001211304208140",
INIT_17 => X"1106409004110240904411024090040106419004010640900411064090440102",
INIT_18 => X"9024010041104409024190240104411004190240906411024190440102419004",
INIT_19 => X"021074B261934D964C3269C09064110040104409064190240104401004190640",
INIT_1A => X"8A74C1323433345145130282E6228A063807E05000143842130115063450454A",
INIT_1B => X"8D46A351A8D46AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA8A28A28A28A2",
INIT_1C => X"A0D068341A0D068341A0D068341A0D068341A0D068341A0D068341A0D46A351A",
INIT_1D => X"50015400000000000000000000000000000000000000000000001007FEA73FC1",
INIT_1E => X"A2D16AAAAF7D568A00AA8400000AAFFC21FFF7D542000FFAE821FF552EAAA105",
INIT_1F => X"0AAAE820BA550015400087FD74BAFFD540000F7D155555087BEABFF552ABDF45",
INIT_20 => X"AAF78015545FFD555555082AAAA10F7FFEAB455500175FF5D2AAAA1000554000",
INIT_21 => X"B45552ABDE00AAD140010F7D17FF45A2FBC2000A2FFC21555551554005D2EA8A",
INIT_22 => X"FF55082E82145A280001EFF78402145A2AE801555D2E95555552E9741000556A",
INIT_23 => X"7DF45557BD5410F7D555545F7AA97410000428AAA557FD5400FF843DE00FFAEB",
INIT_24 => X"0000AA085568BEFFFAE82000085542155557FEAA10007FEABEFAAD1400AA5D51",
INIT_25 => X"AA801EF4920AFA10490A17000000000000000000000000000000000000000000",
INIT_26 => X"C75EABEF4124BAF55B6DF6FABAFFD56F010AA8407428A2F1C01FFF7D142028EB",
INIT_27 => X"552AAFA10007155428A2AE850925D0010400087FD24AAE3DF47010E38E051451",
INIT_28 => X"55D51524004920ADA82EB8A12555EBFB4717D1C2AAFA28EBF5E8B7D5500155FF",
INIT_29 => X"55492A850381C5F6AB6D4124BAE10BED542010FFD57AF55AAF5D7410A2FBC015",
INIT_2A => X"400FF8A38E00F7AABAF7D0000955FDB684051D7F7840517DA2A4871554124925",
INIT_2B => X"75EFBED5400825D557FF55007BD7410EBDB5017DE38E8708008002FAAA4171D5",
INIT_2C => X"00000000000000000000082005F6ABFFEBA0870281C5F4716D5D7FEDB7D0955D",
INIT_2D => X"1401FFFFD5420BAA2AA821FF08043DE10002A964000000000000000000000000",
INIT_2E => X"FBD7410A2AE965555D556ABEF080028B55FFFFFDEBAFFD57FE00A280144BAAAD",
INIT_2F => X"2D16ABEF5500175EF552ABDE000855544AAAA82174105D0402000087FC00BAA2",
INIT_30 => X"AAD154400AAFBC015555554001008003FE00AAEA81154AAFFD65FF5D2EBDEAAA",
INIT_31 => X"FA2AA155550004021E5582A964BE557FEABEF00002BE10FFD540000FFD56ABF5",
INIT_32 => X"1000043DEAA085555400FFAAAAA10F7AC28BF558001454DF78017555F780175E",
INIT_33 => X"5EF5D7BFEEF35055487EFF7D1400105D517FF55087FD7410A2FBC01E7F2AE966",
INIT_34 => X"0000000000000000000000000000000000000010007FEABEFAA84174BA557FD5",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000040",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(4),        -- Port A data input
DOA(0)   => data_read_a_hi_256(4),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(4),        -- Port B data input
DOB(0)   => data_read_b_hi_256(4),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_5_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50DB4A0791B1B4B694369283C81F9996A091832102004AB37B20E07C0C1E006",
INIT_01 => X"285FBC448000804C446A00000034824841280A00084000C8C212892EE2953235",
INIT_02 => X"C809AD5CB118E640A4D118FC011FF0002080000082C8C66609DB7DDDCB1F2036",
INIT_03 => X"250907263A4C90D210A35C82484285720B20648A88800000B8E0F850A8C4500E",
INIT_04 => X"4005122126899100064D20001044429C78243A2C0436C887198AB916E0551A24",
INIT_05 => X"A370C14CA0E900004048002389CFE2F20F7D7A314CB5C20AE51437E044948912",
INIT_06 => X"90184D150505A1D84B7E2A285401412870B20A51842404C44437118630839B88",
INIT_07 => X"E640A94D1AB469D6300E2FFFAA7F8A4D23248130E259C903FBC403A9601A62E8",
INIT_08 => X"0A7E3016250D49CA3F83108186400000EBFD235488B9749BC1AAF325B35CB118",
INIT_09 => X"9B020B7E6AE46082032004904200C03DBC3BCA4860270BFA829968040B0800AC",
INIT_0A => X"22181A2B9203642840124098516CE0C3D825124111A79F802800F20DB4D6DA34",
INIT_0B => X"6824911331CA84D346A964F0125CD7AB1938A00AEFDD567DE480116848C9426A",
INIT_0C => X"01AD7016D701ED7012D701ED7016D701AAB8096B80F5A21828041846620F5AB8",
INIT_0D => X"847B053F48A8308A644A412BCA8470FF0209019081C706EABDAAC0DC0AF012D7",
INIT_0E => X"2194FFC044FF84B08FC862A2CD8F0A89014080A2425422151870500544991292",
INIT_0F => X"038ABBCBC7C7802F86FF87C002F87F002F86FF87C002F87F2000804821021004",
INIT_10 => X"0380230F2FFC002F94FF87C002F87F002F94FF87C002F87F2201BFFEBC2BA0C2",
INIT_11 => X"BFFE7C69E01804E1E7EABE3F000FF97D7C4BC0E008C7C3FE58FC029FEF5CD9A7",
INIT_12 => X"EC9C8120C4DFC802808B2EB22E777ADDE6F8A47CC0600C2683E0FFAAE3F1F001",
INIT_13 => X"FC14DFC5186104C6FE5037FFF00FC0000FC0FEE487A7066FA38C3082637F83BD",
INIT_14 => X"072FFF41C1C0C2038A7CED87A7D109FBBA5070380131CBFB2477BF919024189B",
INIT_15 => X"9F46DFBEB1B7F0380C4A80092E0FC1FDE607A7C077FFE828F0080AE1DFAA1E9F",
INIT_16 => X"5594254A10A03446128898494C09402081F83200A9442217159880640942320E",
INIT_17 => X"1940509465014251140519445094251142511445094451942511425014451940",
INIT_18 => X"9405094450944511425114650146501425194450944509405194250146501405",
INIT_19 => X"0A983124B2DA6924965B4D509445094051940501465014251142501465094451",
INIT_1A => X"BE5FDFF3F7F773CF3CF7D79FA8F5BB4E7F7B9DB7FF3A7E0FF4807F1B6DB7ED43",
INIT_1B => X"F77BBDDEEF77BBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEF",
INIT_1C => X"EF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEE",
INIT_1D => X"FFBFFE00000000000000000000000000000000000000000000001007FE1BFB5E",
INIT_1E => X"FFAE821FF552E820105500155555D2AA8A00AA843FFFFF78002155AAAE974AAF",
INIT_1F => X"0FFAE80000AAAE974BAFFAEAAB45AAAEBDEAAA2FFEAA00AAFFC21FFF7D542000",
INIT_20 => X"000055574BA557FFFF55087BEABFF552ABDF45A2D16AAAAF7D56AA00AA840000",
INIT_21 => X"0BA550015400087FD74BAFFD540000F780155555D7BE8B45085168BFFA2D17FE",
INIT_22 => X"AA10005140145FFFBC01EFAAFFD75FF002E97555A2AABDEAAAAAAAAA00AAAE82",
INIT_23 => X"174BA5D043FF45AAAA974AAF7AEBFF55082AAAA10F7FFEAB455500175FF5D2AA",
INIT_24 => X"000000A2FFC21555551554005D2EA8AAAF78015545FFD555410552EA8BEFAA84",
INIT_25 => X"8E0217DBEA4954AAE3FBFDE00000000000000000000000000000000000000000",
INIT_26 => X"2F1C01D7F7D142028EBAA801EF492087A10490A171455D2EADA28B6803FFFFFF",
INIT_27 => X"FFD56FA10AA8417428E3AE87010A2A4974AAE3AEAFB6DAAA4BDEAAA2F1EDA28A",
INIT_28 => X"D14516DBD7BEDB7DE381451554AA497FFFF451C75EABEF4124BAF55B6DF6FABA",
INIT_29 => X"AAAAA0AFA28A2A4850925D0010400087FD24AAE3DF47010E38E0516D5D7BE8B6",
INIT_2A => X"B7D5500155FF552AAFA10007155545F7F1C21D7AAF1D55FF082A9057DA2AABDE",
INIT_2B => X"70384124ADBFFBE84174AA55043FF6DBEAE950AAEB8ABDF7D1C2AAFA28EBF5E8",
INIT_2C => X"00000000000000000000010A2FBC01555D51524004920ADA82EB8A12410EBFB4",
INIT_2D => X"EBFEBAF7843DFEFF7AE801EFF780174AAAAFBFEE000000000000000000000000",
INIT_2E => X"803FEBAAAD17CEAAAAD140155FFD5420BAA2AA821FF080415410002A96555552",
INIT_2F => X"80028B55FFFFFDEBAFFD57FE00A280144AAA2AA97400A280174AAA2AEBDFEFA2",
INIT_30 => X"A2AE965FF557FE8BFF55557FF55FFFBFFEAA5D51554AA087BFEF555D556ABEF0",
INIT_31 => X"F0004821FFAAAEBDEAAAA843CEAAAA80174105D0402000087FC00BAA2FBD7410",
INIT_32 => X"FF5D2EBDEAAA2D16ABEF5500175EF552ABDE00005554545F7D140145A2D5555F",
INIT_33 => X"E00AAAA81114AAFFD64BA00043FFFFFF80174AA55043DFFFFFAE974BAA2AEBEF",
INIT_34 => X"0000000000000000000000000000000000000000AAFBC015555554001008003F",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000180",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(5),        -- Port A data input
DOA(0)   => data_read_a_hi_256(5),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(5),        -- Port B data input
DOB(0)   => data_read_b_hi_256(5),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_6_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10804B0061A010A2840012C030028180004003220200403302301C0381A0086",
INIT_01 => X"870041CA3839684D18A160000C52424841000000090800090210010008110204",
INIT_02 => X"080108200C1000004464480400C0080100000000010432400800800009882050",
INIT_03 => X"040001008C2340D0840208624210002182800584488000103080010E08C10000",
INIT_04 => X"00101611A029B08410044800000000040088102A440814040400900500001800",
INIT_05 => X"02800000400C820934E4A0002900404400820004000A00824004085011200A00",
INIT_06 => X"2210001A12100830434040870BFE004044420322C00812900308010000829400",
INIT_07 => X"00000860400108C22000A103090074120044800040001103005180911FE0C134",
INIT_08 => X"FD01C0120484C0580020C10000000000087C0800209100004228000110000C10",
INIT_09 => X"88FC08362240404100228080D200DFC1610200E40AA050000040D0C463008083",
INIT_0A => X"29561B22D77C720D2522400000400882091210008440005F8BF4C00002900004",
INIT_0B => X"7E25D11A200024541100342A5A2886285502A880C00107FD355E022005026BCA",
INIT_0C => X"D8282D8A82D8A82D8682D8682D8E82D8A016C1416C15A01D68209A127208A6B1",
INIT_0D => X"807888180A80910A1460150900013400410CB5C9D96236883460B60B602D8282",
INIT_0E => X"0062003C10002442006429124290034E85A742D1A368D0DA2004696884851806",
INIT_0F => X"000000157000604050000000028000D04050000000028000CE80004C00000000",
INIT_10 => X"000000000483D04042000000028000D04042000000028000C508000100000000",
INIT_11 => X"000100000000000000078000A40006000000000000000019A003080010200000",
INIT_12 => X"1001000000093490308001408000000200020000000000000000900518000508",
INIT_13 => X"23490002400000004993C000080000000000001FC000C8804020000000246800",
INIT_14 => X"C05000802000000000001740002256004100000000000000FD00000220000001",
INIT_15 => X"00A000404A000200020000000000002099C000330000040000000000001F0000",
INIT_16 => X"68DA308D09D0804880089A49461032040C07C1440C8190800020530865400540",
INIT_17 => X"9DA7695A1685A369DA7685A168DA369DA5685A168DA7695A5685A368DA7695A5",
INIT_18 => X"5A168DA7695A168DA1695A769DA1685A3695A569DA3685A169DA769DA1685A16",
INIT_19 => X"00046638C31C71C718638E68DA7695A568DA3685A769DA5685A368DA569DA368",
INIT_1A => X"8E76DDB3B7B377DF7DF7D7CEE7F78BCE7F8FF0F4FA957FC7F37F3F5F7CF7F108",
INIT_1B => X"7F3F9FCFE7F3F8E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E3",
INIT_1C => X"E7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE",
INIT_1D => X"AAABFE00000000000000000000000000000000000000000000181007FFDE534F",
INIT_1E => X"F78002155AAAE974AAFFFBFFE10F7FBE8BEF552E95555552EAABEF082E975EFA",
INIT_1F => X"0A2AAAAA10087FC01EF552EAAB45F7AE821550851555555D2AA8A00AA843FFFF",
INIT_20 => X"EFA2AEBDFFF552AAAA00AAFFC21FFF7D542000FFAE821FF552E8001055001541",
INIT_21 => X"000AAAE974BAFFAEAAB45AAAEBDEAAA2FFEAB45552E800AA555568A105D002AB",
INIT_22 => X"AA00AA8400000007BC21FFAA803FFEF5551420105D5568B45FF8400000FFAE80",
INIT_23 => X"C2155007FC20BAA2D5575FF087FFFF55087BEABFF552ABDF45A2D16AAAAF7D56",
INIT_24 => X"0001555D7BE8B45085168BFFA2D17FE000055574BA557FFFE10F7AAA8A00F7FB",
INIT_25 => X"24ADBD70820975FFA2A4BFE00000000000000000000000000000000000000000",
INIT_26 => X"D2EADA28B6803FFFFFF8E0217DBEA4954AAE3FBFDE38F7FFEABFF412A9056D49",
INIT_27 => X"492087010490A07038B6A0AFA38007BC51EF4920AFB55EBA4851450855555455",
INIT_28 => X"2555F68A3855002FBC7BEA4BFFFF492EADA28A2F1C01D7F7D142028EBAA801EF",
INIT_29 => X"45E38A07028E3AE87010A2A4974AAE3AEAFB6DAAA4BDEAAA2F1EDB55492A8508",
INIT_2A => X"F55B6DF6FABAFFD56FA10AA84174381C7FC01C7B68E3DFC75555400105D516DB",
INIT_2B => X"FE38F7A0AFA38E3FFC21450071C2092A2D5571FF0851FDF451C75EABEF4124BA",
INIT_2C => X"0000000000000000000016D5D7BE8B6D14516DBD7BEDB7DE381451554AA497FF",
INIT_2D => X"BEABEF002E801EF00003FF550800155FFA2803CE000000000000000000000000",
INIT_2E => X"8417555085154555552EBFEBAF7843DFEFF7AE801EFF780174AAAAFBFEEAAF7F",
INIT_2F => X"FD5420BAA2AA821FF080415410002A964AAFF803DEAA087FD55FF00043DF45A2",
INIT_30 => X"AAD17CF55002E95410557BEAABA55043DF55F7803FFEF002ABEEAAAAD140155F",
INIT_31 => X"55D51420105D517DF55AAAA964AAA2AA97400A280174AAA2AEBDFEFA2803FEBA",
INIT_32 => X"555D556ABEF080028B55FFFFFDEBAFFD57FE00A280144BA5D7FC2155FFAABDF4",
INIT_33 => X"EAA5D51554AA087BFEEAAF7803DEAAAAFBC0155085540000A2D5575FF08517CF",
INIT_34 => X"00000000000000000000000000000000000001FF557FE8BFF55557FF55FFFBFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000120",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(6),        -- Port A data input
DOA(0)   => data_read_a_hi_256(6),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(6),        -- Port B data input
DOB(0)   => data_read_b_hi_256(6),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_7_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10804B00482010A2842012C024500188000003000000003302300C018180002",
INIT_01 => X"0200084020084048040080000201024040000000080000080200010008110204",
INIT_02 => X"4801082248100000444008000080000041000000002222400800000009008010",
INIT_03 => X"0401008108A1444000020A400000002902006400088000003080040408C10000",
INIT_04 => X"0000100022418000000C80C00400000400201839040000050001140400201820",
INIT_05 => X"02000000400041092C80C0214144004400000000000800045004000020220800",
INIT_06 => X"0000300000000830435150020003004060000000080800801100000030829001",
INIT_07 => X"00000840000008C02000A503010002928040800062481919047140D40008C000",
INIT_08 => X"0A0002120484C0580850810000000000487C000000910000402A800110024810",
INIT_09 => X"8802083624504000022680A1DA20800164000400112284000004D404022A8800",
INIT_0A => X"30014050280040180020400011640CC72E029000084800503004C40100D21024",
INIT_0B => X"3801078228010454210028240082200081140800900220000000002011440009",
INIT_0C => X"40022400224002240822408224082240C1120211202008900800100242428280",
INIT_0D => X"807802988294900A00451109006230006E000800001280110050902901240022",
INIT_0E => X"0042C000C0002000000020020490000400020001020080401010813094801146",
INIT_0F => X"807144102420700052000003C00780B00052000003C007808450484C00000000",
INIT_10 => X"2C0E00E0D003300052000003C00780B00052000003C00780890800010000130C",
INIT_11 => X"000100000661801E18042100E000060100000B03803838012403800010240000",
INIT_12 => X"10111848322020512000414400000002000A1001058300C0741C005412080908",
INIT_13 => X"029F008240864231013BF00008000C3C003F00184040EF8041204321188053E0",
INIT_14 => X"F770008060130C8071821040403F5600411004C2600E3400C27C020223090644",
INIT_15 => X"00B8CA406A0002C812240B0201F038021140403F740004010472041E20110100",
INIT_16 => X"0080228011010042802890484040000008004945000100008844430060198941",
INIT_17 => X"0000000000000600802008020000400000000000080200802008000000000000",
INIT_18 => X"8020100000000008020080000000000020080200000000040080200802008060",
INIT_19 => X"0A14584104000208208000018020080200000010020080200800010000080200",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000442",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"82AAAA00000000000000000000000000000000000000000000001007FEBC3240",
INIT_1E => X"552EAABEF082E975EFAAAABFFEF002ABDF555D5157555F7FBC00AAAAD5400BA0",
INIT_1F => X"AAAAABDF55FFFBFDF55555568ABAAAD5401FF5D2AAAA10F7FBE8BEF552E95555",
INIT_20 => X"005D55554105D51401555D2AA8A00AA843FFFFF78002155AAAE974AAFFFBFFEA",
INIT_21 => X"A10087FC01EF552EAAB45F7AE821550851554AAF7FBFFEAA007BFFFEFF7D5400",
INIT_22 => X"00105500155EF5D2EBFF450000020AA5D7BC0000F7D555545A28000010A2AAAA",
INIT_23 => X"A8A10FFD568ABAA2D56AAAAF7AABFE00AAFFC21FFF7D542000FFAE821FF552E8",
INIT_24 => X"000145552E800AA555568A105D002ABEFA2AEBDFFF552AAAABAA2AE95555FFAA",
INIT_25 => X"F5C20BAAAD5420821C2EAAA00000000000000000000000000000000000000000",
INIT_26 => X"7FFEABFF412A9056D4924ADBD70820975FFA2A4BFFFF1C2EB8F45555550545E3",
INIT_27 => X"BEA4954AAE3FBFDE82B6AEBAF55E3FFFAF55555F6FA92BED5421C75D20AAA38F",
INIT_28 => X"20075FDFD7F7D5400385D51504385D55401455D2EADA28B6803FFFFFF8E0217D",
INIT_29 => X"7DB68E02038B6A0AFA38007BC51EF4920AFB55EBA485145085555492F7F5FFE9",
INIT_2A => X"028EBAA801EF492087010490A071EF4920B8F45140E07082417BC2000EBD5505",
INIT_2B => X"DA92A2A09257DE3A4AAA10F7D16FAAABED56AE82F780BAE28A2F1C01D7F7D142",
INIT_2C => X"00000000000000000000155492A85082555F68A3855002FBC7BEA4BFFFF492EA",
INIT_2D => X"EAAB455D5142155AAD1400AAA2D1420005D2EA9A000000000000000000000000",
INIT_2E => X"D1421555D042BAAAF7FBEABEF002E801EF00003FF550800155FFA2803CFFF552",
INIT_2F => X"7843DFEFF7AE801EFF780174AAAAFBFEE00F7AAAAB55AAFBEAB555D7BFDE00F7",
INIT_30 => X"085154400FFD17FE1000517FF55FFD5420BA5D55400BA555543155552EBFEBAF",
INIT_31 => X"0087BC0000A2D5421EFF7AE810AAFF803DEAA087FD55FF00043DF45A28417555",
INIT_32 => X"AAAAD140155FFD5420BAA2AA821FF080415410002A965FF080428B45552A9540",
INIT_33 => X"F55F7803FFEF002ABEE00A280001FFA28028A00FFD17DEAAF7D56AA10FF842BA",
INIT_34 => X"0000000000000000000000000000000000000155002E95410557BEAABA55043D",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"FFFFFFFE00000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000000000000000000001F",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(7),        -- Port A data input
DOA(0)   => data_read_a_hi_256(7),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(7),        -- Port B data input
DOB(0)   => data_read_b_hi_256(7),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_8_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10004B00000400E2840012C0000001800000070000000033022000000000082",
INIT_01 => X"000009C0183808481C0160000E02424040000000180800080200010048110204",
INIT_02 => X"080108000090000004400C000080000051000000000002400800000009000010",
INIT_03 => X"0000000004300840000200000000000002800504488000103080880008800000",
INIT_04 => X"00009410A028A084000440C00400000400001032040800150400008500221800",
INIT_05 => X"4280008040048A09302420202804400400800010200A00000204080011014A00",
INIT_06 => X"2B02000A32114192434010001FFC004240428122000800000008012000821400",
INIT_07 => X"00000840000008402001A50200000630404080006248381B000080837FF88114",
INIT_08 => X"0A000210040440480000090000000000087C0000009100000002000110000090",
INIT_09 => X"08020A322000400102260021DA2080114502002409A04400004282C4E1228800",
INIT_0A => X"904A4522920052012120400011641C4601005000041100002004800100C21024",
INIT_0B => X"78051792A8000454104020001280008845022000900000010444000000020009",
INIT_0C => X"000000000000000000000000000000000800040000452A9008001002424A8002",
INIT_0D => X"807880508202100A1000810B2020340041248548490004800400000008000800",
INIT_0E => X"20020000C000044214240932000001428CA14650A128508A2004284024840022",
INIT_0F => X"80000000001020404000783FC0000010404000783FC000000880084C01041008",
INIT_10 => X"FC7E0000000010404000783FC0000010404000783FC000000500000103D45F3D",
INIT_11 => X"000103961FE78000000000402400020003B43F1F800000002201080000202658",
INIT_12 => X"01617CD8000000803000804080000020090659833F9F03C00000000000040500",
INIT_13 => X"00400018639EC000000000000FE03FFC00000000400840000C31CF6000000800",
INIT_14 => X"4000001E2A3F3D80000000400802000401AA8FC7E00000000100002C2F5B0000",
INIT_15 => X"4020000104480DC372B47F060000000000400802000017570FF6000000010020",
INIT_16 => X"28CA30051851A0C0002890484600320408004444048090800022130864000540",
INIT_17 => X"84A1284A1284A328CA328CA328CA328CA328CA3284A1284A1284A1284A1284A1",
INIT_18 => X"CA328CA328CA3284A1284A1284A1284A328CA328CA328CA3284A1284A1284A12",
INIT_19 => X"080440000000000000000028CA328CA328CA328CA1284A1284A1284A128CA328",
INIT_1A => X"9EDFC8F33637D6CB6CB2900DA6128A0A543EBC57A10A244257C5051E75D64108",
INIT_1B => X"1F0F87C3E1F0F9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7",
INIT_1C => X"E1F4F87D3E1F4F87D3E1F4F87D3E1F4F87D3E1F4F87D3E1F4F87D3E1F0F87C3E",
INIT_1D => X"02ABFE00000000000000000000000000000000000000000000001007FE8A8913",
INIT_1E => X"F7FBC00AAAAD5400BA082AAAA10000000010F7D5421EF007BC01FF5D7FFFE100",
INIT_1F => X"A5551554AAFF80021EF002A820BAFF8428A00A2AAAABEF002ABDF555D5157555",
INIT_20 => X"EFFFFFEAB55002ABFE10F7FBE8BEF552E95555552EAABEF082E975EFAAAABFEA",
INIT_21 => X"F55FFFBFDF55555568ABAAAD5401FF5D2AAAB55FFD1400AA5D7FC01EFA2FFE8B",
INIT_22 => X"74AAFFFBFFEAA08001555555516ABEFA280020AA5D043DF55557BEAAAAAAAABD",
INIT_23 => X"2AB55005140145AAFFE8AAAF7D1401555D2AA8A00AA843FFFFF78002155AAAE9",
INIT_24 => X"0000AAF7FBFFEAA007BFFFEFF7D5400005D55554105D51400005551421EF0804",
INIT_25 => X"7FC21EF5D75FFE10142EBAE00000000000000000000000000000000000000000",
INIT_26 => X"C2EB8F45555550545E3F5C20BAAAD5420821C2EAAA101C0005000E3D1401D71C",
INIT_27 => X"0820975FFA2A4BFE925D51554AAE384001FF142E800AAFF802AA28AAAEAFBFF1",
INIT_28 => X"2557BC21D7BEF5EDBC7FFF1EFB6D1420BAE38F7FFEABFF412A9056D4924ADBD7",
INIT_29 => X"55417BEDA82B6AEBAF55E3FFFAF55555F6FA92BED5421C75D20AAB45F7D14709",
INIT_2A => X"FFFFF8E0217DBEA4954AAE3FBFDEAA1C001056D415F6ABEFA2840208249043AF",
INIT_2B => X"00385D51401EF00002FB45085F4016DAAF1EDAAAFFFB401455D2EADA28B6803F",
INIT_2C => X"00000000000000000000092F7F5FFE920075FDFD7F7D5400385D51504385D554",
INIT_2D => X"417410AAD540155557FC01EF5D557DE105D2AA8A000000000000000000000000",
INIT_2E => X"842AABAA2AEBDFFF552EAAB455D5142155AAD1400AAA2D1420005D2EA9A105D0",
INIT_2F => X"02E801EF00003FF550800155FFA2803CE105D55574BAA280021EF5D2E820BAF7",
INIT_30 => X"5D042BB45FFD157410557FC0155F7D57FF55F7D57FFEF550028AAAF7FBEABEF0",
INIT_31 => X"FAA8000000080428B55087FFFE00F7AAAAB55AAFBEAB555D7BFDE00F7D142155",
INIT_32 => X"55552EBFEBAF7843DFEFF7AE801EFF780174AAAAFBFEEBA5D04021EF087BE8BF",
INIT_33 => X"0BA5D55400BA5555430BA5555421EF00043FF45007BC21FFA2D57FEBAF7FBC21",
INIT_34 => X"0000000000000000000000000000000000000000FFD17FE1000517FF55FFD542",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000080",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(8),        -- Port A data input
DOA(0)   => data_read_a_hi_256(8),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(8),        -- Port B data input
DOB(0)   => data_read_b_hi_256(8),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_9_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10004B00018000A2840012C0000281800000030000000033022000000000006",
INIT_01 => X"000008000000004C0020000000100268413C0A61590001D90213C10008110204",
INIT_02 => X"680108200010000054400C000080000041000000010002400800800009082011",
INIT_03 => X"0004000000002040000200100000000042800584488000103081880008800000",
INIT_04 => X"00001610A00AB084000400C00600000400001030040010050020020400001880",
INIT_05 => X"02000200400C8A09206420000C00410400000000000800000804000000000800",
INIT_06 => X"2A10201A12104010435051000801004040000322980800000080000100821000",
INIT_07 => X"000018400000086020002502000002000040800062C8081B0000008000088034",
INIT_08 => X"0A000610040440480000010000000000187C0000009100002046000110000010",
INIT_09 => X"4802082220084001002400214A2080014400006400A000000000015421800800",
INIT_0A => X"4B505008020032032320400011640447000010040000000020048409004A9020",
INIT_0B => X"280005922000045400002001100000000D0000008000000041C48000002003EA",
INIT_0C => X"2080020000208002000020800200002080010000104100800000100202420142",
INIT_0D => X"C06800100240180A0010010921003400432C8CC8D80044000000080080020800",
INIT_0E => X"2002C000C000240004641932041403428DA146D0A36850DA3200684004800403",
INIT_0F => X"0000000144002000420000000280001000420000000280000000084C01041008",
INIT_10 => X"0000000004801000500000000280001000500000000280001100000100000000",
INIT_11 => X"00010000000000000002A0002000020100000000000000182001000000240000",
INIT_12 => X"00110000000900003000004000000000000A0000000000000000900002000100",
INIT_13 => X"205D0080400000004803F0000800000000000004E0004E800120000000240BA0",
INIT_14 => X"4770000060000000000005600013560001100000000000002574020020000001",
INIT_15 => X"0020CA406A0000080200000000000020806000137400040000000000000B8000",
INIT_16 => X"68DA320D19D1A0CA8028984D46543600080040440C8090800000130061400140",
INIT_17 => X"8DA368DA368DA1685A1685A1685A1685A1685A1685A1685A1685A1685A1685A1",
INIT_18 => X"5A1685A1685A1685A1685A1685A1685A368DA368DA368DA368DA368DA368DA36",
INIT_19 => X"801010000000000000000068DA368DA368DA368DA368DA368DA368DA3685A168",
INIT_1A => X"344A2D840100E492082405548817344CCCF48DE68A89004F98614C5C38E2540A",
INIT_1B => X"1A0D068341A0D14514514514514514514514514514514514514534D34D34D34D",
INIT_1C => X"41A4D268341A0D069349A0D069349A0D068341A4D268341A4D268341A0D06834",
INIT_1D => X"FD557400000000000000000000000000000000000000000000001FFFFE2CAD83",
INIT_1E => X"007BC01FF5D7FFFE10002ABFF55F7D168A00552E95555007BFFF55087BE8BFFF",
INIT_1F => X"0F7FBC0145F7AE801EFF7FBFFF455D7BC0155F7D557410000000010F7D5421EF",
INIT_20 => X"00AA803FFEF5D55421EF002ABDF555D5157555F7FBC00AAAAD5400BA082AAAA1",
INIT_21 => X"4AAFF80021EF002A820BAFF8428A00A2AAAAAAAF7D17DE00FFFBD5555A2AABDE",
INIT_22 => X"75EFAAAABFFEF002A954BA5551421EF552E954105D00021455555420AA555155",
INIT_23 => X"575EFA2FFD75455D7BE8A005D5557410F7FBE8BEF552E95555552EAABEF082E9",
INIT_24 => X"000155FFD1400AA5D7FC01EFA2FFE8BEFFFFFEAB55002ABFE10080028BFFF7D5",
INIT_25 => X"71F8F7D147BEFBEFEBD152400000000000000000000000000000000000000000",
INIT_26 => X"C0005000E3D1401D71C7FC21EF5D75FFE10142EBAF7DE3D16DA0041209056D1C",
INIT_27 => X"AAD5420821C2EAAA10E3FFC0145F7A0801FFEBFBF8F6D417BC716DEBD1524101",
INIT_28 => X"8F7F5D0545B6AAB8E38B68A3AFFF5551471FF1C2EB8F45555550545E3F5C20BA",
INIT_29 => X"455D5B470925D51554AAE384001FF142E800AAFF802AA28AAAEAFABAE3D17DE2",
INIT_2A => X"56D4924ADBD70820975FFA2A4BFFFF082E974BA4155401C7552097428550E021",
INIT_2B => X"AE0008002ABFFF7DB505FFAAFBD7555417FEFA00495B52438F7FFEABFF412A90",
INIT_2C => X"00000000000000000000145F7D147092557BC21D7BEF5EDBC7FFF1EFB6D1420B",
INIT_2D => X"17DE100804001EF55516ABFF557BFDFEFA2D5400000000000000000000000000",
INIT_2E => X"7FD55FFA2D5400105D0417410AAD540155557FC01EF5D557DE105D2AA8BEFAAD",
INIT_2F => X"D5142155AAD1400AAA2D1420005D2EA9A00A2FBC0145FF84001EFA2FFEABFF00",
INIT_30 => X"A2AEBDEAAAAD17DEBAFFD142155FFAAAAABAFFAAAABFF5551555FF552EAAB455",
INIT_31 => X"55D00154AA552E801455D7BD54105D55574BAA280021EF5D2E820BAF7842AABA",
INIT_32 => X"AAF7FBEABEF002E801EF00003FF550800155FFA2803CFFF002E954BA00514015",
INIT_33 => X"F55F7D57FFEF550028A10000428BEFF7FFC01FFA2FFD5545007BFDE10087FC00",
INIT_34 => X"0000000000000000000000000000000000000145FFD157410557FC0155F7D57F",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000100",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(9),        -- Port A data input
DOA(0)   => data_read_a_hi_256(9),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(9),        -- Port B data input
DOB(0)   => data_read_b_hi_256(9),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_10_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10040B0001824802840102C00002C18000202300500030B3132000400992006",
INIT_01 => X"A140098018300848180060000C00424040000000080000080200010008110200",
INIT_02 => X"0801080200100000046558040080000041000000002402400800000009008010",
INIT_03 => X"00010100840000D0842242024210810802006400088000003080054288C10000",
INIT_04 => X"0000100022008000000C08C00C00000400A83A3044200C840000800400101820",
INIT_05 => X"0200000040000000248080210044000402000025000800020004207010100800",
INIT_06 => X"0800200000004010435040A14001004844000800CC0812541020008230829000",
INIT_07 => X"00000860408108502000250208000600004080006248081B0040808000088000",
INIT_08 => X"0A000210040440480060010000000000087C0810209900000002000110020010",
INIT_09 => X"08020A2222004040000484214A2080110108C280022210020240000401080880",
INIT_0A => X"000000000200000C042040001164044609101000840000802004800100421020",
INIT_0B => X"782415809888A45010082408028010080110280800001001051A124810410800",
INIT_0C => X"0089000890000900009000890008900008800048004420910800120242488000",
INIT_0D => X"4110000006008820020010010001300040000100014000808C48004008800090",
INIT_0E => X"2002000040002000040020020490080400020001000482000010012080008005",
INIT_0F => X"0000010140002040100000000280401040100000000280400000204801041008",
INIT_10 => X"0000000006801040020000000280401040020000000280400500000000000000",
INIT_11 => X"0000000000000000010280002400040000000000000001182001080010000000",
INIT_12 => X"10000000000D0000808000408000000200000000000000000000902000000500",
INIT_13 => X"A000000200000000681000000000000000008004A00040004000000000340000",
INIT_14 => X"4000008000000000000085200002000040000000000001002400000200000001",
INIT_15 => X"00200000000002000000000000000021802000020000000000000000020A8000",
INIT_16 => X"040006E00100044200289048085D402008000040000100000000020065400000",
INIT_17 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_18 => X"0000000000000000000000000000000020080200802008020080200802008020",
INIT_19 => X"8290100000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"8A355950666151451453D5006F86890A940FE0D39712614261D20E4355520542",
INIT_1B => X"6532994CA65328A28A28A28A28A28A28A28A28A28A28A28A28A28A28A28A28A2",
INIT_1C => X"AE532994CA6532995CAE572B94CA6532994CA6572B95CAE532994CA6532994CA",
INIT_1D => X"FFBC2000000000000000000000000000000000000000000000001007FECF31DC",
INIT_1E => X"007BFFF55087BE8BFFFFD557400FF842ABEFA2AAA8B5500003DF55F7D568AAAF",
INIT_1F => X"008556ABFFA2D16AB550000021FFF7D17FFEF08042AB55F7D168A00552E95555",
INIT_20 => X"55A2D557400557BC2010000000010F7D5421EF007BC01FF5D7FFFE10002ABFE0",
INIT_21 => X"145F7AE801EFF7FBFFF455D7BC0155F7D557545FFAE820AA007BFDFEF55003FF",
INIT_22 => X"00BA082AAAA00FFAE820AAAAAABDFEFF78028BEF005140145A2842AA10F7FBC0",
INIT_23 => X"6AB55A2D157400552EBFFEF5D7BD75EF002ABDF555D5157555F7FBC00AAAAD54",
INIT_24 => X"0000AAF7D17DE00FFFBD5555A2AABDE00AA803FFEF5D55420BA08557FEBAAAD5",
INIT_25 => X"0E3AF55F7DF68ABAE3F1C0000000000000000000000000000000000000000000",
INIT_26 => X"3D16DA0041209056D1C71F8F7D147BEFBEFEBD152400F7842FBD7B6AAAAB551C",
INIT_27 => X"5D75FFE10142EBAE0008556FBD7B6DB6AB7D1C0A001D7FFD178FC71C0E28B7DE",
INIT_28 => X"2147BFAFEF49043AF45A2DF504285D71C00101C0005000E3D1401D71C7FC21EF",
INIT_29 => X"7DA28428A10E3FFC0145F7A0801FFEBFBF8F6D417BC716DEBD15256DF7AA8209",
INIT_2A => X"545E3F5C20BAAAD5420821C2EAAA00E3AA82092A2AABAFD7EB8A2ABC70855401",
INIT_2B => X"70821C557AE92A2DF6AB7DA2DF50410412ABDFC75D7BD55FF1C2EB8F45555550",
INIT_2C => X"000000000000000000000BAE3D17DE28F7F5D0545B6AAB8E38B68A3AFFF55514",
INIT_2D => X"03DF45FFAEA8B555D2EAAB45F7FBE8ABAAAD5400000000000000000000000000",
INIT_2E => X"D168B55552AA8BEFAAD17DE100804001EF55516ABFF557BFDFEFA2D540010FF8",
INIT_2F => X"AD540155557FC01EF5D557DE105D2AA8A0008557FF45FFFFE8BEF5D2E80155FF",
INIT_30 => X"A2D5401FFF7AA800105D7FE8BEF08002AB45AAFFC00AA5D51400105D0417410A",
INIT_31 => X"5AAAEAAB450055421FFAA8428A00A2FBC0145FF84001EFA2FFEABFF007FD55FF",
INIT_32 => X"FF552EAAB455D5142155AAD1400AAA2D1420005D2EA9A10A2AA82010AAAEAAB5",
INIT_33 => X"ABAFFAAAABFF555155400555568A10AAFBEABEFA2FFC0010082ABFF55557BD55",
INIT_34 => X"00000000000000000000000000000000000000AAAAD17DEBAFFD142155FFAAAA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"FFFFFFFE00000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000000000000000000011F",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(10),        -- Port A data input
DOA(0)   => data_read_a_hi_256(10),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(10),        -- Port B data input
DOB(0)   => data_read_b_hi_256(10),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_11_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10180B05A0010402840602C2D001019000000300000000330A20080EC180002",
INIT_01 => X"AB400986B830284D1820E0000C36424840000000080000088200080802512220",
INIT_02 => X"8801081438106400A4F55800008000004100000040CCE24208005000C9060032",
INIT_03 => X"000406A492E6E440842254D002108153432004800880000030C0315688C00006",
INIT_04 => X"00001201200090001205400000000094108C322644240C840008030440111800",
INIT_05 => X"222000444008010028404002A002009402400025080880000C04223000170900",
INIT_06 => X"01080C1020002810436532AB4003004864200A00540816544522008200821100",
INIT_07 => X"6400E96C488108502001295BA100022E4340800062D82819435143F20008C0A0",
INIT_08 => X"0A0012160585C1D809A3810000000000C8FD0B1420992419034A0221116C3810",
INIT_09 => X"4902083E2CB0400002020480C2008009000ACEC06B25500202988C84C0220028",
INIT_0A => X"004040000203600E06204000116C14474A36500499C49C802004C00800088000",
INIT_0B => X"6804110230CBA4576708201C0212100B492A2008000A1001C49A9348498B0808",
INIT_0C => X"410E5418E5410E5418E5418E5410E5418B2A0872A08428010000120202085000",
INIT_0D => X"41110244066C0820221480010AA7300042080980919580808C9A5002880A18E5",
INIT_0E => X"2022C000C0002020094030220C960A0409020481024482501A00401410088521",
INIT_0F => X"836090540355D86C046619A54052A5B86A046619694063168280004801041008",
INIT_10 => X"A2C60289802AB86A046619A54052A5B86C04661969406316AC018B0E2936DA02",
INIT_11 => X"CB0E1076D4A200B2AC611A3D0405886C6EB211550815A8A2686EC81E2A48B68A",
INIT_12 => X"8CE0C5E8F650E48000892B37885620C1E1A06D7016A90A4626D82B10F1B1FC09",
INIT_13 => X"4E02144D335546F28724001B030A56140A184483000C410A2699A2E32AC9C041",
INIT_14 => X"E8018A0A01B2990242E278056AAA203920E0BAE2012C08281808319C186F1E16",
INIT_15 => X"44F9051C049B18A12CB481042AD140C227002A0A02066954E7540CCDB58415AA",
INIT_16 => X"409024681181044080809A490C0964200800200108010003A02272400C19B80D",
INIT_17 => X"0902409024090240902409024090240902409024090240902409024090240902",
INIT_18 => X"1004010040100401004010040100401024090240902409024090240902409024",
INIT_19 => X"0284000000000000000000401004010040100401004010040100401004010040",
INIT_1A => X"20A069105251C0000001541148062608804180C0B10A04CA0900474210420140",
INIT_1B => X"0000000000000000000000000000000000000000000000000000208208208208",
INIT_1C => X"0000000000004020000000000000000000100800000000000000000000000000",
INIT_1D => X"00015400000000000000000000000000000000000000000000001007FE0FC1C0",
INIT_1E => X"00003DF55F7D568AAAFFFBC2010557BEAA10AAFBE8A00557BFFFEF007BC21550",
INIT_1F => X"55D7FE8BFF5D7FD540055003FFEFFFD142145000000000FF842ABEFA2AAA8B55",
INIT_20 => X"45557FC2010557FFDF55F7D168A00552E95555007BFFF55087BE8BFFFFD55754",
INIT_21 => X"BFFA2D16AB550000021FFF7D17FFEF08042AB55A2AAAAB4508517FE00557BC01",
INIT_22 => X"FE10002ABFE00AAFFE8AAAFF8402000550002145085555400F7FFE8A0008556A",
INIT_23 => X"3FEBA002A975EFF7D17DFFFAA8000010000000010F7D5421EF007BC01FF5D7FF",
INIT_24 => X"000145FFAE820AA007BFDFEF55003FF55A2D557400557BC2145A2D1421450804",
INIT_25 => X"7BF8FEF1C7FC516D080E15400000000000000000000000000000000000000000",
INIT_26 => X"7842FBD7B6AAAAB551C0E3AF55F7DF68ABAE3F1C00005D7BEDA00B6F1EFA2855",
INIT_27 => X"147BEFBEFEBD15257D5D7FEFBD7417BD5438550038FC7FFDF4216D080E07000F",
INIT_28 => X"514517FE105575C216D5571C50104171FDF7DE3D16DA0041209056D1C71F8F7D",
INIT_29 => X"00FFF1EFA0008556FBD7B6DB6AB7D1C0A001D7FFD178FC71C0E28B6DA2AEADB4",
INIT_2A => X"1D71C7FC21EF5D75FFE10142EBAE10A2FBEFA92F78A05028550E001451455524",
INIT_2B => X"016DB6D54514500003FEBA1420905FFFFDF78FC7BE84050101C0005000E3D140",
INIT_2C => X"0000000000000000000016DF7AA82092147BFAFEF49043AF45A2DF504285D71C",
INIT_2D => X"FFDE00F7D17FEBA557BEABEF557BD55EF082A974000000000000000000000000",
INIT_2E => X"FBC01FF082A97410FF803DF45FFAEA8B555D2EAAB45F7FBE8ABAAAD5400105D7",
INIT_2F => X"804001EF55516ABFF557BFDFEFA2D5401FF5D7FFDF55007BD74BA5D042AB45F7",
INIT_30 => X"552AA8BEFAAAABFF5555517FE005555401FF55515541000517FFEFAAD17DE100",
INIT_31 => X"A5D2A801455D5140000FFD57FE0008557FF45FFFFE8BEF5D2E80155FFD168B55",
INIT_32 => X"105D0417410AAD540155557FC01EF5D557DE105D2AA8A10AAFBFFE00F7AA974B",
INIT_33 => X"B45AAFFC00AA5D51401FFFFD15555500003FEBA5D04001EFFFFFE8B55FF84174",
INIT_34 => X"00000000000000000000000000000000000001FFF7AA800105D7FE8BEF08002A",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000100",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(11),        -- Port A data input
DOA(0)   => data_read_a_hi_256(11),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(11),        -- Port B data input
DOB(0)   => data_read_b_hi_256(11),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_12_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50080B01BC002006940202C0DE041196A83183000000023322287E0FC000006",
INIT_01 => X"0E000C048000C048400380000007026040000000080000088200002802153231",
INIT_02 => X"2809AD0E7D180040945008040090000061800000C0E2F66009DA3D11CB148015",
INIT_03 => X"210D050012F6F8D2108216E24842005B8A20640008800000B8E0141C28851006",
INIT_04 => X"0080100022408000060DE0000066630C70241827041000040800820480001AA4",
INIT_05 => X"0240000C400000003C808003E0C8001401000000040900020904004000070800",
INIT_06 => X"00006C00000008784B4D210E0001006050800000100804005784000130821200",
INIT_07 => X"A64019490A044860300FA3968B20028FC06080106249F819A19143FE00088200",
INIT_08 => X"0A002610240D494A0753D1810240000038FC234480B1709A81C67325B31EFD18",
INIT_09 => X"090209222EB84000010000104200802180210C007827C000009DBE040800008C",
INIT_0A => X"0000000002000030003040081164FC469227D20019F413503004900020000200",
INIT_0B => X"28200100004304D267C06CC500566003C13E0000000460000000000010CE0000",
INIT_0C => X"E1865E1065E1065E1865E1065E1065E1832F0C32F08000000004100202015940",
INIT_0D => X"0403CFE7E03E8080382FD0018FE670004000000000D5C023009278B7835E1065",
INIT_0E => X"01EA0000440000800A0040028108000000000000000000000A74812DF00E0BF4",
INIT_0F => X"8362F658A7E5F82CD23B6B0E403DBBE82C563B6A4E403DBB88C0E04820020004",
INIT_10 => X"BE5403AB992F282C563B6B0E403DBBE82CD23B6A4E403DBBB1084E4B25AC48DF",
INIT_11 => X"0E4B1D32BAB504BB74AD3F3FE04A8E0D0C319A7988B6F0C75CFD801A962454CF",
INIT_12 => X"18D994B866E2E8C3808B6B63040328E7A33AF99B0AC20DE634D06C437BF85100",
INIT_13 => X"5F6214CA5991C6A7177402C49CA354D808D358A927EAD10A652CC8E3538BEC41",
INIT_14 => X"E80083C3EAEB2003695430A7CDAA289553922990C11A4E494988231B32570CDC",
INIT_15 => X"D5B304AD05A946D81616970A225658940BA7CDAA0A312666BD600E5550B49F36",
INIT_16 => X"00000100000010420000904C0040000008003B81000000021CFEE02E2803BC0F",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"8020080200802008020080200802008000000000000000000000000000000000",
INIT_19 => X"0210100000000000000000008020080200802008020080200802008020080200",
INIT_1A => X"24481C040000B5145144015085C1B946088881360A95118D90215C090CB05442",
INIT_1B => X"32190C8643219041041041041041041041041041041041041041249249249249",
INIT_1C => X"4B2592C964B2592C964B2592C964B2592C964B2592C964B2592C964B2190C864",
INIT_1D => X"AFBC2000000000000000000000000000000000000000000000001007FEF001D6",
INIT_1E => X"557BFFFEF007BC2155000015555087FC0010AAFBFFE100004020BAAAFFD5400A",
INIT_1F => X"5AA8400000A2AABFF45550400000AAFBFFFEF550000010557BEAA10AAFBE8A00",
INIT_20 => X"10555155555FF8017400FF842ABEFA2AAA8B5500003DF55F7D568AAAFFFBC215",
INIT_21 => X"BFF5D7FD540055003FFEFFFD142145000000145A2AA821EFFFFFD7410007FC00",
INIT_22 => X"8BFFFFD5574000051420BA557FC2145557FC20AAA2D57DEBAA2FBD55455D7FE8",
INIT_23 => X"AAA00550415410AAFBFFFEF55042AB55F7D168A00552E95555007BFFF55087BE",
INIT_24 => X"000155A2AAAAB4508517FE00557BC0145557FC2010557FFDE10AA8400000082E",
INIT_25 => X"0A02092B6F5D2438A2FBC2000000000000000000000000000000000000000000",
INIT_26 => X"D7BEDA00B6F1EFA28557BF8FEF1C7FC516D080E1557D0075C7028B6F1FAE0000",
INIT_27 => X"F7DF68ABAE3F1C017DAA8E07028B6A0BFF6D490E00000BEF5FAFEF4904070005",
INIT_28 => X"FE3FBD0438007FC00385D555556DEB8410400F7842FBD7B6AAAAB551C0E3AF55",
INIT_29 => X"BAA2FBD557D5D7FEFBD7417BD5438550038FC7FFDF4216D080E0716DAAA0851F",
INIT_2A => X"56D1C71F8F7D147BEFBEFEBD152400005F450BA417BC51454971C20AAB6D17DE",
INIT_2B => X"DE10BE8E070280020AAA28410410400BEFBFAFEF49042AB7DE3D16DA00412090",
INIT_2C => X"0000000000000000000016DA2AEADB4514517FE105575C216D5571C50104171F",
INIT_2D => X"5574BAFFD568A10002A82000FFD5400AAA2FBC00000000000000000000000000",
INIT_2E => X"D568BEF0004174105D7FFDE00F7D17FEBA557BEABEF557BD55EF082A975EF005",
INIT_2F => X"FAEA8B555D2EAAB45F7FBE8ABAAAD5401EFA2AA974BAF7803FFFF002A82000FF",
INIT_30 => X"082A975EFA280175FFAAFFC00BA087FC20AA5D55555FFA28000010FF803DF45F",
INIT_31 => X"50851420BAFFD57DEAAAAFBD75FF5D7FFDF55007BD74BA5D042AB45F7FBC01FF",
INIT_32 => X"EFAAD17DE100804001EF55516ABFF557BFDFEFA2D540010007FD74AA007BD754",
INIT_33 => X"1FF55515541000517FE10F7AA954AA080428AAA000002010FFFFE8BEF080428B",
INIT_34 => X"00000000000000000000000000000000000001EFAAAABFF5555517FE00555540",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"FFFFFFFE00000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000000000000000000001F",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(12),        -- Port A data input
DOA(0)   => data_read_a_hi_256(12),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(12),        -- Port B data input
DOB(0)   => data_read_b_hi_256(12),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_13_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10110A0441812402840402822007818000E00700000000330A3000000008042",
INIT_01 => X"A1400984B830C848180260000C0042404001000008220008A200100802110200",
INIT_02 => X"88010C02801040002475580400800000410000000064024608134C0CC9018034",
INIT_03 => X"00010100926220D084234212421085084300648A0880000630C0654288C10000",
INIT_04 => X"0004122122029100100C00001200009C40A83A2044360C84190BAC04E0101820",
INIT_05 => X"027000004009050064C8C00104C10184034010250089C00EB004327064B60900",
INIT_06 => X"910000152500A050436A10A14003004864B00A50440812541027008230821380",
INIT_07 => X"640029605091495020002B8AAA000AF003408000E258081963F100C00008C2E8",
INIT_08 => X"0A001210040441C802E0010084000000AAFC09142899000B20020001105A0010",
INIT_09 => X"4A02096A62004000020004104200802D9838C2C80322100202020194408000A0",
INIT_0A => X"000000000203240E46204000516C04468C101005800E95802004B20020080200",
INIT_0B => X"28200101118BA4510008241D005211000910000A000A1000809A93485D610000",
INIT_0C => X"0000000800000000000000800000000000000400000000000000100202055040",
INIT_0D => X"0100000006C0802042501001C8017000C2190890904000508908000000000800",
INIT_0E => X"0010C000C00081A08BC832A209AB0A85094284A14254A2551010513080109404",
INIT_0F => X"01293C0F5012906A96DCD13042CE0C206E92DCD07042CE0C40D0204800000000",
INIT_10 => X"71CA2168ACB0E06E92DCD13042CE0C206A96DCD07042CE0C4408632C39530BA9",
INIT_11 => X"632C30D522CE80239CC2806AC44E954939AB299E000738F88296CA13B444CA42",
INIT_12 => X"D5306028F01990C080808494A64708B265CC4052B0F30302E060965EA0058408",
INIT_13 => X"28A2CA9722094650CCAC0629112BA89C04A228568547B1654B9104A32865145C",
INIT_14 => X"B80D4D8D48CB54012290470562EC29E44050B1DC60132282B68B9AA60C051E03",
INIT_15 => X"0A5C11B9008FE2FA38F87804251CB0FAD40562EC0B426149D17E0044B10A158B",
INIT_16 => X"5094246A10A10441010090480C0964201800044109012001A000726E45428000",
INIT_17 => X"0942509425094250942509425094250942509425094250942509425094250942",
INIT_18 => X"9425094250942509425094250942509425094250942509425094250942509425",
INIT_19 => X"02A8000000000000000000509425094250942509425094250942509425094250",
INIT_1A => X"BAFFD7F7F7F775555557DF9FE0FFBBEEFF3F7DF7FF3E7E2FF0087B9F7DF7E245",
INIT_1B => X"FD7EBF5FAFD7EBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAE",
INIT_1C => X"AFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FA",
INIT_1D => X"0557DE00000000000000000000000000000000000000000000001007FE0001DF",
INIT_1E => X"0004020BAAAFFD5400AAFBC2155AAAA97410FFFFEAAAAF7AA955EFF7803FF450",
INIT_1F => X"0F7AEBDE10FFFFFDEAAF7D568AAA5D002AB55005568B55087FC0010AAFBFFE10",
INIT_20 => X"FF5D04154BAAAAEAAA10557BEAA10AAFBE8A00557BFFFEF007BC215500001541",
INIT_21 => X"000A2AABFF45550400000AAFBFFFEF550000155A28415410F7AEAABFFA2D1555",
INIT_22 => X"8AAAFFFBC21555D517FF45F7AEA8BFFA2AEAAA10A280021EF5D557FF55AA8400",
INIT_23 => X"974AAF7D142145082A975FF555568A00FF842ABEFA2AAA8B5500003DF55F7D56",
INIT_24 => X"000145A2AA821EFFFFFD7410007FC0010555155555FF80174000055555EFAAAE",
INIT_25 => X"A0925C7E38E38F7D14557AE00000000000000000000000000000000000000000",
INIT_26 => X"075C7028B6F1FAE00000A02092B6F5D2438A2FBC2145B6A090428FFF5EAA92E3",
INIT_27 => X"1C7FC516D080E15438E3A4BAE00FFF5FAE92F7D16AAAA41042FB7D145568B7D0",
INIT_28 => X"8FFA4AFBFFAAD1505FF490E174AABEA0ADA005D7BEDA00B6F1EFA28557BF8FEF",
INIT_29 => X"FF555F7FF7DAA8E07028B6A0BFF6D490E00000BEF5FAFEF490407155BE8E1242",
INIT_2A => X"B551C0E3AF55F7DF68ABAE3F1C0145415B78F45FFA4AFBC7BEA4AAA10A284001",
INIT_2B => X"04380055525FFBEAE90482E3D54216D0024975FF555F68A00F7842FBD7B6AAAA",
INIT_2C => X"0000000000000000000016DAAA0851FFE3FBD0438007FC00385D555556DEB841",
INIT_2D => X"0020BAF7D16AA10A28402155A2AEA8BEF5D516AA000000000000000000000000",
INIT_2E => X"003DFEF55516ABEF0055574BAFFD568A10002A82000FFD5400AAA2FBC0145FF8",
INIT_2F => X"7D17FEBA557BEABEF557BD55EF082A974BAA28028A00F7D16AA10F7D56AABA08",
INIT_30 => X"000417545FFAA820BAFF843DFFFA2D5421FF002E954AAFF843DE105D7FFDE00F",
INIT_31 => X"5F7802AA10AA80001FF5D7FFDFEFA2AA974BAF7803FFFF002A82000FFD568BEF",
INIT_32 => X"10FF803DF45FFAEA8B555D2EAAB45F7FBE8ABAAAD540145007FE8B55FF843DF5",
INIT_33 => X"0AA5D55555FFA280000BA0855401EFF7AA82010AAD1421FF0004155FF557FEAA",
INIT_34 => X"00000000000000000000000000000000000001EFA280175FFAAFFC00BA087FC2",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"FFFFFFFE00000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000000000000000000019F",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(13),        -- Port A data input
DOA(0)   => data_read_a_hi_256(13),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(13),        -- Port B data input
DOB(0)   => data_read_b_hi_256(13),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_14_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10020A000180000284008280000281800000030000000033022000000580002",
INIT_01 => X"A140098018300848184860000C20C24040000000084000084200000000110200",
INIT_02 => X"88010C5A8010A600A4F558040080000041000000022C024008003CCCC9028030",
INIT_03 => X"000103A7A00904D0842242024210810803006480088000003081054288C10000",
INIT_04 => X"0000120122009000100C00000000000400A83A2044200C840000800400101820",
INIT_05 => X"020000004008010024C0C0010040000402000025000800020004207000100800",
INIT_06 => X"010000102000005043403AA14003004864000A00440812541020008230821000",
INIT_07 => X"2400A96850A16854200021DA2A0002000340800062C80819EBC402800008C020",
INIT_08 => X"0A0012140404414814E001000000000029FD0A10289924810182000110028010",
INIT_09 => X"080208222200400002000400420080010008C2C0032210020200008440000080",
INIT_0A => X"000000000203200E0620400011640446DA101004800005802004800000000000",
INIT_0B => X"282001001088A45000082408000010000910000800001000009A924810410000",
INIT_0C => X"0080000000000000080000000000000080000000000000000000100202000000",
INIT_0D => X"0100000004408020021010010001700042080880904000008808000000000800",
INIT_0E => X"00000000C00000000040302200800A0409020481024482501010413080008404",
INIT_0F => X"8090008142014840100002C38280000840100003838280000640204800000000",
INIT_10 => X"072C000444C00840020002C38280000840020003838280002C09D01086839746",
INIT_11 => X"D0104B01C57100440202900184414430534605E3804802180022480419183514",
INIT_12 => X"594C194000090450808802008830024F0E248C902AEF0024170CF18001003C09",
INIT_13 => X"20020E5A08E6000048200196264BCF1C030C0604800001076C04730000240049",
INIT_14 => X"2003DEDE82C78900902A0D0000080019FAAA32D9602490302409292B83280001",
INIT_15 => X"049100021171F6C34080240108AB292CA000000800AD1A19F6F000AA0C0A0000",
INIT_16 => X"4090246810810440000090480C0964200800000108010016000012004542800D",
INIT_17 => X"0902409024090240902409024090240902409024090240902409024090240902",
INIT_18 => X"9024090240902409024090240902409024090240902409024090240902409024",
INIT_19 => X"0280000000000000000000409024090240902409024090240902409024090240",
INIT_1A => X"9E7FDDF77777F3CF3CF7D54CEFD79B4E5C8FF0F7BE9D75C7F7B71F5F7DF65040",
INIT_1B => X"7F3F9FCFE7F3F9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7",
INIT_1C => X"E7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE",
INIT_1D => X"28417400000000000000000000000000000000000000000000001007FEFFFE0F",
INIT_1E => X"F7AA955EFF7803FF4500557DF45F7D16AB455D00001EFAAAAAAABA555557555A",
INIT_1F => X"555003FF450804001555D2AA8AAA002ABDE10082ABDF55AAAA97410FFFFEAAAA",
INIT_20 => X"EF5D5168A10082E80155087FC0010AAFBFFE100004020BAAAFFD5400AAFBC214",
INIT_21 => X"E10FFFFFDEAAF7D568AAA5D002AB55005568A00A2D5401455D00175FFFF84175",
INIT_22 => X"2155000015400AAD157545080402145087FD75FFF7AE82145A2D17FE10F7AEBD",
INIT_23 => X"000BAFFFBE8AAAA2FBFDE00087FD5410557BEAA10AAFBE8A00557BFFFEF007BC",
INIT_24 => X"000155A28415410F7AEAABFFA2D1555FF5D04154BAAAAEAAA005D002AB450000",
INIT_25 => X"A0AAA82555157555B68012400000000000000000000000000000000000000000",
INIT_26 => X"6A090428FFF5EAA92E3A0925C7E38E38F7D14557AF45FFDB6AB6D4100071C7B6",
INIT_27 => X"B6F5D2438A2FBC21455D0A3FF6D080407155552AAAA920020BFE10002EBAF45B",
INIT_28 => X"54100175C7E380125D7555B6DA1014248217D0075C7028B6F1FAE00000A02092",
INIT_29 => X"45AAD178E38E3A4BAE00FFF5FAE92F7D16AAAA41042FB7D145568A38AADF4014",
INIT_2A => X"A28557BF8FEF1C7FC516D080E15400A2DB5754508040716D007BD05EFEBAA821",
INIT_2B => X"DA0055002AB6D0000020BAFFF1E8ABABEF1FAE001C7FD54005D7BEDA00B6F1EF",
INIT_2C => X"00000000000000000000155BE8E12428FFA4AFBFFAAD1505FF490E174AABEA0A",
INIT_2D => X"FEABFF080015555F78028A00555155555FF84000000000000000000000000000",
INIT_2E => X"003DE10082EAAB45FF80020BAF7D16AA10A28402155A2AEA8BEF5D516AB45F7F",
INIT_2F => X"FD568A10002A82000FFD5400AAA2FBC0145552ABFFFF000417555552EA8A1000",
INIT_30 => X"55516AABAAAFFC0145000417555A280001455D7FFDE105504021EF0055574BAF",
INIT_31 => X"F007BC01FFAAAE80155AAD568ABAA28028A00F7D16AA10F7D56AABA08003DFEF",
INIT_32 => X"105D7FFDE00F7D17FEBA557BEABEF557BD55EF082A97410AAFFD55450800155F",
INIT_33 => X"1FF002E954AAFF843DE10550028BEF0004020BAF7D568AAAF7D168A105D7FD74",
INIT_34 => X"0000000000000000000000000000000000000145FFAA820BAFF843DFFFA2D542",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"FFFFFFFE00000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000000000000000000001F",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(14),        -- Port A data input
DOA(0)   => data_read_a_hi_256(14),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(14),        -- Port B data input
DOB(0)   => data_read_b_hi_256(14),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_15_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000A000000000284000280000001800020030000000033022000000180002",
INIT_01 => X"A140098018300848180060000C00424040000000080000080200000000110200",
INIT_02 => X"080108000010E60004E55800008000004100000000040240080000C009170016",
INIT_03 => X"0000000080000040842240000210810002000400888000003080014288C00000",
INIT_04 => X"0001100024A0800000440000000000040088322044200C840000011400151800",
INIT_05 => X"A200014C4000000020000000000B8094020000254C8800000514203000108800",
INIT_06 => X"000821000000A050434010A14001004844000801540812540020008600831000",
INIT_07 => X"C2000864489128502000210222000200034080006248081958C0008000088000",
INIT_08 => X"0A001214050540C800200101860000000B7C0910209900000002000110000010",
INIT_09 => X"0B0208222004400000000400420080010008C28002201002020001140800002C",
INIT_0A => X"000000000203000C04204000116404460810100080000F802004800000000000",
INIT_0B => X"280001001088A45000082008000010000100000800001000001A124800010000",
INIT_0C => X"0080000800008000000000000000000080000400004000000000100202000008",
INIT_0D => X"0100000004C00020025000018801600040000000000000008808000000000800",
INIT_0E => X"00108000C0000000000020020080080000000000000402000000000000009400",
INIT_0F => X"00000000000000404200000000000000404200000000000008C0004800000000",
INIT_10 => X"0000000000000040500000000000000040500000000000000400000100000000",
INIT_11 => X"0001000000000000000000000400020100000000000000000000080000240000",
INIT_12 => X"00110000000000C00080010180000000001A1024050000000000000000000400",
INIT_13 => X"0002008040000000002000000804002000000000000001000120000000000040",
INIT_14 => X"2000000061100280000000000008000001104422000000000008020020000000",
INIT_15 => X"00100000000009080E2E0A000000000000000008000004000000000000000000",
INIT_16 => X"0000046000000440000090480809402008000001000000000000000004188000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0280000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000040000000000040",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"8517DE00000000000000000000000000000000000000000000001007FE000000",
INIT_1E => X"AAAAAAABA555557555A284175FF000002010552A97400007BFDE10A2AA801EF0",
INIT_1F => X"F5D2AAAB45F7D17DF45087BC0155002A801FF08003DF45F7D16AB455D00001EF",
INIT_20 => X"45F7D568BEFAAD557555AAAA97410FFFFEAAAAF7AA955EFF7803FF4500557DFE",
INIT_21 => X"F450804001555D2AA8AAA002ABDE10082ABDFFFF7D17FE10002E954AAF7FBC21",
INIT_22 => X"5400AAFBC21EFA2AE95545A2D56ABFFAAD17DE10FFD1420AA007FC014555003F",
INIT_23 => X"801550055401555D00174BA002AA8B55087FC0010AAFBFFE100004020BAAAFFD",
INIT_24 => X"000000A2D5401455D00175FFFF84175EF5D5168A10082E801FFFF8428A10002A",
INIT_25 => X"71FAE00A2A0871EF145B7FE00000000000000000000000000000000000000000",
INIT_26 => X"FDB6AB6D4100071C7B6A0AAA82555157555B680125C71C0E0500049209543808",
INIT_27 => X"E38E38F7D14557AFC75524AFB45FFD178F7D1C71C2145002E801C7140A3FF45F",
INIT_28 => X"00024954AAFFFBC2145F7DB6DBEFA2D557545B6A090428FFF5EAA92E3A0925C7",
INIT_29 => X"820071C71455D0A3FF6D080407155552AAAA920020BFE10002EBAFC7FFDF7AE0",
INIT_2A => X"E00000A02092B6F5D2438A2FBC21FFBEA090545B6D568BFFAADB7AE10F7D5470",
INIT_2B => X"21FFE3802FA2808208017D1C5142155410A104AA1420AFB7D0075C7028B6F1FA",
INIT_2C => X"00000000000000000000038AADF401454100175C7E380125D7555B6DA1014248",
INIT_2D => X"E954100004174AA00516AA10AA80155EF5D7BFDE000000000000000000000000",
INIT_2E => X"2E801555D2EBDF45F7FFEABFF080015555F78028A00555155555FF8400155552",
INIT_2F => X"7D16AA10A28402155A2AEA8BEF5D516AB555D043DF55F7D56ABEF55514015508",
INIT_30 => X"082EAAB55FFFBE8A100804154AAF7FFC2145FFFFFDFEFAAD157545FF80020BAF",
INIT_31 => X"FA2FBE8A00FFD155410005555545552ABFFFF000417555552EA8A1000003DE10",
INIT_32 => X"EF0055574BAFFD568A10002A82000FFD5400AAA2FBC01FFF78400155F7D16ABE",
INIT_33 => X"1455D7FFDE105504021FFAA843DEBA0000021EF555142155002E800AA55003DF",
INIT_34 => X"00000000000000000000000000000000000000BAAAFFC0145000417555A28000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000180",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(15),        -- Port A data input
DOA(0)   => data_read_a_hi_256(15),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(15),        -- Port B data input
DOB(0)   => data_read_b_hi_256(15),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_16_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"DA22C618B1000482B688B186588884862A400438255FC38381441205BA803003",
INIT_01 => X"8645A80028404C211203A952A90341080B173340412000E1005D628000820484",
INIT_02 => X"A101A9006DC1084833011850AAC55001349B10881802821808B4110007005E11",
INIT_03 => X"010108A802BB00080080006020020001A61036202800000D2410104200404550",
INIT_04 => X"8BFA58800005C40A46240252145148B38248030356415A4E62B6FC660F287240",
INIT_05 => X"0F05EA11E570000D610000000710296E542B6E3A825C15FB30A643695BFC2D56",
INIT_06 => X"408003200040202B8584112645554B029006000140BCC0460050690A95C8383D",
INIT_07 => X"00480A2140040BE1480FA004342AA6F12000054004867415401DCDCF2AA10800",
INIT_08 => X"B32A8819064E48288012D45000005050247AA85220700009C06206C48080EDEA",
INIT_09 => X"445B2081340B6596594800400413CAC020894480000008C54C00311002000002",
INIT_0A => X"000000004B240028000342A00002FE00A3A1F06E491800AA29588181040A0020",
INIT_0B => X"2400848002912300200092BA80325A20000000000A8A5AA80018120E00066000",
INIT_0C => X"00220002200022000220002200022000210001100010000A40450100210072A0",
INIT_0D => X"002815014B90000205DA00880100095A648000000010006AC23000C7B69EC220",
INIT_0E => X"80922554515512174000000490009000000000000004010042A204A0C5817680",
INIT_0F => X"63EAA9C238B2D4C800632B266E828EE4C800632AAAB6830D0FC6B06C04102800",
INIT_10 => X"A149339E8FB964C800632B266E82B2E4C800632AAAB683310872800EDA52DA00",
INIT_11 => X"800EB090D4AAC91268FFCBE81397826C4A20D2B6C510E8624792A4A30A40839A",
INIT_12 => X"8849D5C532408DD6E004C90C06AC019D88B9795012CA96902C799912BC3C087A",
INIT_13 => X"531C74485BD42A30906057FADAA456218FD8E3ED83B60E3A242DC0F18983638E",
INIT_14 => X"A06FB555793057C444CF45C5C9E89543B8BC6E80193DC36F6C71D1093A478706",
INIT_15 => X"45DC02B331650CA8ACB4007E00D1C6A6A58395C917F7E74D936F650D69B51727",
INIT_16 => X"0000012000081500008A422150884081ACAAC0542054004FC588464050810DCD",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"147A7797E1E1A79E79E1560EEFBD11544C690DA64C1C69A9916D7E4F68A36040",
INIT_1B => X"7A7D1E9F47A7D345345345345345345345345345345345345345145145145145",
INIT_1C => X"4FA7D3E9F4FA3D1E8F47A3D1E8F47A3D1E9F4FA7D3E9F4FA7D3E9F4FA7D1E9F4",
INIT_1D => X"F8015400000000000000000000000000000000000000000000001007FE00001F",
INIT_1E => X"007BFDE10A2AA801EF08517DE10FFFFFDFEFA2D16AB55A2FFFFEAA5D7FC0000F",
INIT_1F => X"A5D2EBDFEFAAD17FFFF002EBDE000800174AA55043FFFF000002010552A97400",
INIT_20 => X"AAAA80000105D557FF45F7D16AB455D00001EFAAAAAAABA555557555A284174B",
INIT_21 => X"B45F7D17DF45087BC0155002A801FF08003DE000004154BA002A800BA087FE8A",
INIT_22 => X"FF4500557DEAAF7D57DEBA082A82010FFAE975555D7FFDEAAFF80155EF5D2AAA",
INIT_23 => X"7FFFF557FD55FF08003FE0055043FF55AAAA97410FFFFEAAAAF7AA955EFF7803",
INIT_24 => X"0001FFF7D17FE10002E954AAF7FBC2145F7D568BEFAAD557410552EA8BEFA2D5",
INIT_25 => X"FFFDEAA5571C7010FF8412400000000000000000000000000000000000000000",
INIT_26 => X"C0E050004920954380871FAE00A2A0871EF145B7FE10E3F1F8FC7AAD56DB7DB6",
INIT_27 => X"555157555B680124924124BDFEFA2D57FFC71C2EBDE280000174825D0E3FFC71",
INIT_28 => X"21424800AA007FEDAAAA284020385D5F7AF45FFDB6AB6D4100071C7B6A0AAA82",
INIT_29 => X"AAFF80175C75524AFB45FFD178F7D1C71C2145002E801C7140A3FE10080A1748",
INIT_2A => X"A92E3A0925C7E38E38F7D14557AE92EBDB78EAA1C2482010FFAE9556D557FF8E",
INIT_2B => X"7410492EADBEFA2D178FEF5575D55EF000A38E10490A3AF45B6A090428FFF5EA",
INIT_2C => X"000000000000000000001C7FFDF7AE000024954AAFFFBC2145F7DB6DBEFA2D55",
INIT_2D => X"56AB45A2D57DFFFF7FBFFEAA555555400F780000000000000000000000000000",
INIT_2E => X"0415400552ABDF55552E954100004174AA00516AA10AA80155EF5D7BFDE10A2D",
INIT_2F => X"80015555F78028A00555155555FF840000000043DFEFAAD17FF45552ABFEBA08",
INIT_30 => X"5D2EBDE10002E974005D04020BA007BFDEBAA284000BA557FE8B45F7FFEABFF0",
INIT_31 => X"0F7AE955EF5D7BE8ABAF784175555D043DF55F7D56ABEF555140155082E80155",
INIT_32 => X"45FF80020BAF7D16AA10A28402155A2AEA8BEF5D516AA00AAFBE8AAA55040000",
INIT_33 => X"145FFFFFDFEFAAD157410082ABFFEFAAD16ABFF5555575FF082AA8A00002AAAB",
INIT_34 => X"0000000000000000000000000000000000000155FFFBE8A100804154AAF7FFC2",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000080",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(16),        -- Port A data input
DOA(0)   => data_read_a_hi_256(16),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(16),        -- Port B data input
DOB(0)   => data_read_b_hi_256(16),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_17_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"5284CE4FB7BD2C8994A13392DBD02E14006B82AC7E800D44D3DD2FD5F9B961C0",
INIT_01 => X"F8ACD01F7E03FC6793F2199B39FC233C11D93AE6F3BB92B32091DBC339B24542",
INIT_02 => X"8F333007FD6808092A2AFA6667033DB50853379C10BFF70F1BD011110F205F18",
INIT_03 => X"294ADB4AFFCBF0DAD63ABF836B58EAFE060478202022234B2E0303FDC9E18339",
INIT_04 => X"DB7A40806FE4040840EBC563A0150A0926146FECB04196482236FC2005282AE1",
INIT_05 => X"0403DA0383200831C68206D7E6D0250834336D1E81500FDB306045255BFC2076",
INIT_06 => X"4470716040413D29AAC69F5FE33C072F06062C003670497AFF00291B3C0E2015",
INIT_07 => X"0849147160448EBB9537A0022DC67987042EE976ABEA77684653547819FF2000",
INIT_08 => X"E019C0C82A4E4820C15B089C380110002446045A31345000A84432409207F02D",
INIT_09 => X"983838A3BFF1030C397C060B4254064302042F803A69DB931FF4391C00002CC0",
INIT_0A => X"FB1F1F7BC81C003C001674BB55B5FBB4BB4F26A1BEE004F9D0DE08F7DE336DB2",
INIT_0B => X"28302F800633F1D0A7CC9AE74117FE01D34E82AC0CE8FCCC200A59BDD2FFE3E3",
INIT_0C => X"E9F79E9F79E9F79E9F79E9F79E9F79E9F7CF4FBCF4F000C2E225C8DE0BA05BB0",
INIT_0D => X"A5A99FD6D3FEF4BEB5FF994F0FEFFCCF8430000000D9D147E0D57AE7B79E9F79",
INIT_0E => X"0593F33FA0CF170F40006001B1A05C0000000000000008004BA78428C7AD7FE4",
INIT_0F => X"E46444357B3950A9BFBAC94CFA8581E0A9BFBAC8CCFA8580C7CAF51EF68B2976",
INIT_10 => X"B5DB54A09003E0A9BFBAC94CFA8581E0A9BFBAC8CCFA8580E46FBFCB0CBEDA57",
INIT_11 => X"BFCB1D5CFEB56A1A100D5345C1BFFE8FBDB892DB463034198E2881F3F787DF76",
INIT_12 => X"D39387F92B2935DFEAADDF38EBCFB9E3D636DCDF9B90F966BF92966D5D9E7467",
INIT_13 => X"27055EB6D555CB294981B7FB5B2954CD3013013FDF5E82AF5B6AAAE594A4E0AD",
INIT_14 => X"835C67E655BAA868610117575EA1C34BD6975D48B44A0405FC15BA7270FF2565",
INIT_15 => X"6CD2A47D0CBA96252756D7217E5E1C61DBDF5FA167F7AE5D3D21A414007F7D7E",
INIT_16 => X"000005F08000179C16DECF67F08BC02F9067ED55805600545DFE45A80E7BD07F",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"00C0000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"9A919261A1A6075D75D10DDF2F82003009EDCC4052E92E0826462117114F9818",
INIT_1B => X"8D068351A8D069A6BAE9A69A6BAE9A6BAE9A69A6BAE9A6BAE9A69A69A69A69A6",
INIT_1C => X"A8D46A351A8D46A351A8D46A351A8D46A341A0D068341A0D068341A0D068351A",
INIT_1D => X"AFFD5400000000000000000000000000000000000000000000001FFFFE000011",
INIT_1E => X"A2FFFFEAA5D7FC0000FF8015410FFFFFFFFFFFFFFDFEFF7D568A1008003DF55A",
INIT_1F => X"5A2D1400000804154BAF7D168A00A2803DE10FFAE95410FFFFFDFEFA2D16AB55",
INIT_20 => X"BAFFD56ABFF002EBDFFF000002010552A97400007BFDE10A2AA801EF08517DF5",
INIT_21 => X"FEFAAD17FFFF002EBDE000800174AA55043FEBA0004174AA5504000AA55042AA",
INIT_22 => X"7555A284175FFFFFBE8B55A2FFFFF55F7803DEBA002AAAAAAF7FBD74BA5D2EBD",
INIT_23 => X"17400FFD57DE00AAAAAAB45A2AA97545F7D16AB455D00001EFAAAAAAABA55555",
INIT_24 => X"0000000004154BA002A800BA087FE8AAAAA80000105D557FE00A2D5420AA5D04",
INIT_25 => X"D16AA00000E3DF6DBEF5D2400000000000000000000000000000000000000000",
INIT_26 => X"3F1F8FC7AAD56DB7DB6FFFDEAA5571C7010FF8412428FFFFFFFFFF7FBF8FD7EB",
INIT_27 => X"A2A0871EF145B7FF7DA2D547038140E10492FFDF6DA28A28E3DE00F7A092410E",
INIT_28 => X"2550A020BA55002AA82F7DF6DBD71C2EBFFC71C0E050004920954380871FAE00",
INIT_29 => X"BAF7F5D74924124BDFEFA2D57FFC71C2EBDE280000174825D0E3FEAA14001249",
INIT_2A => X"1C7B6A0AAA82555157555B680125FFEBFFEDB55BEFFFAF6DE38E3DEAA002EADA",
INIT_2B => X"AE28B6D545092490E10400FFDB7AE00A2AAADB45BEA092545FFDB6AB6D410007",
INIT_2C => X"00000000000000000000010080A174821424800AA007FEDAAAA284020385D5F7",
INIT_2D => X"BFDFEFF7FFEAB45A2D56AA00002EBDFFFF7D5400000000000000000000000000",
INIT_2E => X"AABDE10FF8400010A2D56AB45A2D57DFFFF7FBFFEAA555555400F780000AAFFF",
INIT_2F => X"004174AA00516AA10AA80155EF5D7BFDFEFAAD1554BA552E82000F7FFFFEAAA2",
INIT_30 => X"552ABDEBA5D0002000552A800BA55042AA10FFFFFDF55552EBDF55552E954100",
INIT_31 => X"FA2AEBFEAA082EBDEBAFFD55540000043DFEFAAD17FF45552ABFEBA080415400",
INIT_32 => X"45F7FFEABFF080015555F78028A00555155555FF84001FFAAFBFFF55FFFBEABF",
INIT_33 => X"EBAA284000BA557FE8AAAFFD155400082A82000F7FFE8A00A2AABDF45F780001",
INIT_34 => X"0000000000000000000000000000000000000010002E974005D04020BA007BFD",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"FFFFFFFE00000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000000000000000000019F",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(17),        -- Port A data input
DOA(0)   => data_read_a_hi_256(17),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(17),        -- Port B data input
DOB(0)   => data_read_b_hi_256(17),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_18_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"69844019080000A21A611406840014122A641074155FC28A2024001001801003",
INIT_01 => X"A643D920034004180005E9E3C90360C0041C0181002001602025800008440084",
INIT_02 => X"B7333980808408103F2000F81FC0FEDEAC2161B0B84D0002188011110C018041",
INIT_03 => X"0405D434003F2C020081587008020561E55116B0290000042B71240C800440F8",
INIT_04 => X"50805AC31007D6125724029216554A9847669903D640EC8E2001002604503004",
INIT_05 => X"07008000E0EA11803850C800010022660C1C0065003C0404002646DC20A02D40",
INIT_06 => X"0100001028040C093D0491A640FFC10028000280002C44D620F0228454C83810",
INIT_07 => X"08501620028007500CE801241021FE78E40486014006009044359DC707F55C20",
INIT_08 => X"9307CC082A0A4A6A01ECDCC40850001630080002A5CA500344040108120080AB",
INIT_09 => X"A0172083200B6186128040600C10C1C02009505081100088080BC6A052802001",
INIT_0A => X"002020000F0CA8428642430080438408A510185A40000008B83181C000141040",
INIT_0B => X"2E00C04C44C92A88DC42215C882E82240880000060D7030C30B885200D274404",
INIT_0C => X"10006100061000610006100061000610003080030800800C0540310130006E21",
INIT_0D => X"10202021000780004200408C1002003F66CA18A1B62622381B2B841840614006",
INIT_0E => X"806400FC503F08180050942E4200020C1B060D8306C182701404C19730108010",
INIT_0F => X"ABAF377DF1CA160820520EB3057E70E60820520F33057E72E915415900002900",
INIT_10 => X"5D48F37FAFEFE60820520EB3057E7CE60820520F33057E7EC658BF2DA7822AAB",
INIT_11 => X"BF2D4B2A80BF8FE39FD78EB0D882014A62C568FFAFC73FFDD9C2B30E0468A2AD",
INIT_12 => X"800DFC06F59F710107533C0C4E37619440FBFBAB2400AFC1600361D798F32658",
INIT_13 => X"EB9454005BAA36DEFF894823A3D1A88A2FE29D5FC6DCAA2A002DD51B6E7C728C",
INIT_14 => X"92A78606A28A5427AAB9FF4EDD251C7123E291660733EBF6FE519001BF40DEBB",
INIT_15 => X"AB58AFBFD5DE200A8EBE3A3EC110339E1DCEDC2590495BB2112E2BE4BF5F3B70",
INIT_16 => X"C1B06808348340000020301805002D008C1F92000A5F421B8000DB4910382202",
INIT_17 => X"1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06",
INIT_18 => X"B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C",
INIT_19 => X"000000000000000000000041B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1",
INIT_1A => X"8A244C16454170410412CA064A9BBECEB80EE173C2300FE3F1A3550F7DF16000",
INIT_1B => X"A552A944A2512AAA8A28A28A2AAAAAA8A28A28A2AAAAAA8A28A28A28A28A28A2",
INIT_1C => X"A25128944A25128944A25128944A25128944A25128944A25128944A25128954A",
INIT_1D => X"D2A80000000000000000000000000000000000000000000000001007FE000004",
INIT_1E => X"F7D568A1008003DF55AAFFD5410FFFFFFFFFFFFFFFFFFFFFBFDEBA552E974105",
INIT_1F => X"0FFFFFFFFFF7FBE8B55AAD16AA1000516AA005D0400010FFFFFFFFFFFFFFDFEF",
INIT_20 => X"00087BC2155087BC0010FFFFFDFEFA2D16AB55A2FFFFEAA5D7FC0000FF801541",
INIT_21 => X"0000804154BAF7D168A00A2803DE10FFAE95555FFFBE8B45A2D56ABEFFFFFFFE",
INIT_22 => X"01EF08517DF55000000010082A974AA08557DEBAFFAEBFF55AA8028B55A2D140",
INIT_23 => X"800105D2AAAA10A2D1420AAFFAEA8BFF000002010552A97400007BFDE10A2AA8",
INIT_24 => X"0000BA0004174AA5504000AA55042AABAFFD56ABFF002EBDEBA0004020BA552E",
INIT_25 => X"FBFFEBA552A95410552485000000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFF7FBF8FD7EBD16AA00000E3DF6DBEF5D2438FFFFFFFFFFFFFFFFEFF7",
INIT_27 => X"5571C7010FF8412410FFFBF8FC7E3F5EAB45BEDB6FA3800556FA00550405028F",
INIT_28 => X"5BEDB6FBC7EBF5F8E10007BC516D1C71C5010E3F1F8FC7AAD56DB7DB6FFFDEAA",
INIT_29 => X"55BE8A2DB7DA2D547038140E10492FFDF6DA28A28E3DE00F7A09256DE3F1EAB5",
INIT_2A => X"4380871FAE00A2A0871EF145B7FF45080E070280820924AA145578E92F7A4BFF",
INIT_2B => X"FEBA1C0A00092412E850005D2AAFA38A2DF45082F7AAA8BC71C0E05000492095",
INIT_2C => X"000000000000000000000AA140012492550A020BA55002AA82F7DF6DBD71C2EB",
INIT_2D => X"FFFFFFFFFBFDFEFF7FFFDEAA5D2E954105504154000000000000000000000000",
INIT_2E => X"557DE005500154AAFFFBFDFEFF7FFEAB45A2D56AA00002EBDFFFF7D5400AAFFF",
INIT_2F => X"2D57DFFFF7FBFFEAA555555400F78000010F7FBE8B55AAD16AB55F7FBFDEAA08",
INIT_30 => X"FF84001FFAAD568B45FFFBFFF55A2D568A00087BD55FF5D5555410A2D56AB45A",
INIT_31 => X"A555168A10FF803DF45FFAABDFEFAAD1554BA552E82000F7FFFFEAAA2AABDE10",
INIT_32 => X"55552E954100004174AA00516AA10AA80155EF5D7BFDF45002A974AA0800000A",
INIT_33 => X"A10FFFFFDF55552EBDEBA5D2E80010082A97410552EBDEBAA2FBD5400F7AAA8B",
INIT_34 => X"00000000000000000000000000000000000000BA5D0002000552A800BA55042A",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000080",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(18),        -- Port A data input
DOA(0)   => data_read_a_hi_256(18),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(18),        -- Port B data input
DOB(0)   => data_read_b_hi_256(18),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_19_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"042200000000000041088001001AA00000000000000000000000500802000003",
INIT_01 => X"200048000024000000000404000000000A22000800000800004A200000000001",
INIT_02 => X"032210008DEF00400060000001C008002489E0F0004037B00010101010000000",
INIT_03 => X"0000008128000000000000000000000024001620280000000000354200004008",
INIT_04 => X"000058800004C4024024001210001054B1C822009640000E2000002604003000",
INIT_05 => X"07008000E0200000000000000000200604000000001C04000026400000002C40",
INIT_06 => X"000000000000002600859AA1000D410000000000002C42010010200004C83810",
INIT_07 => X"0040380142810010564C41001140120024020280448088050008108100640000",
INIT_08 => X"83004C390242006200000868000040001020A850040AD0080426006933800DC4",
INIT_09 => X"0013200000016186100000000010C04002C00000000000707000000000000000",
INIT_0A => X"000000000B0C0000000101400040C0408100000000000008A810000000000000",
INIT_0B => X"00000000000400020000440000000000000000002F0001F00002024B20002000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"000210001D800000000000000002000964000000000000000000000000000000",
INIT_0E => X"0000000C50030008000000000000000000000000000000000000000000000000",
INIT_0F => X"101088A37034E156600D740022800EC156600D740022800D01E0412D06904000",
INIT_10 => X"0224081044914156600D7400228002C156600D7400228001098F00D0FB750500",
INIT_11 => X"00D0F2DD014010046037814EA63DBB31CE7605001008C41A061F0E7D693E6170",
INIT_12 => X"6D600000004089E12350C0E01FF23315422BABB46FEF5019146C0800380CC98F",
INIT_13 => X"130AA3592000000000629C03F3E60330C00C628908214551AC90000001036152",
INIT_14 => X"65C006070845039014460088235ACC3123E2A29148841008482A4DAC00000000",
INIT_15 => X"53A66BE7A5040018D8A8AD9090A1EC20A188235AC509FB50C2D0500B4094208D",
INIT_16 => X"000000000000000000000000000000008C01800270000061100084046086CD49",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"861A2882313054D34D301C862AA08BBA3F0C7010C6600A00200251C744192000",
INIT_1B => X"130984C261309861861861A69861861861861A69861861861861861861861861",
INIT_1C => X"6130984C26130984C26130984C26130984C26130984C26130984C261349A4C26",
INIT_1D => X"82E97400000000000000000000000000000000000000000000001007FE000002",
INIT_1E => X"FFFBFDEBA552E974105D2A801EFFFFFFFFFFFFFFFFFFFFFFFFFEAA552E954000",
INIT_1F => X"FFFFFFFFFFFFFFFFFEFF7FBFFEAA5D2E97545FFFFC2010FFFFFFFFFFFFFFFFFF",
INIT_20 => X"0008003DF555D5157410FFFFFFFFFFFFFFDFEFF7D568A1008003DF55AAFFD55E",
INIT_21 => X"FFFF7FBE8B55AAD16AA1000516AA005D04001EFFFFFFFFFFFFFBFDF45AAD16AA",
INIT_22 => X"0000FF80155EFFFFFFFFEFF7D16AB55A2D57DEBA557FEAA10080402010FFFFFF",
INIT_23 => X"6AB45FFFBFDEBA5D7FC0155FFFFD7410FFFFFDFEFA2D16AB55A2FFFFEAA5D7FC",
INIT_24 => X"000155FFFBE8B45A2D56ABEFFFFFFFE00087BC2155087BC00AAFFFBFDF45A2D5",
INIT_25 => X"FFFDEAA552E95400002095400000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFEFF7FBFFEBA552A954105524851C7FFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"000E3DF6DBEF5D25D7FFFFFFFFFFFFBFDFEFEBF5F8E92552E9556DEBF1C2038F",
INIT_28 => X"FE3F1FAF55A2D568A0000003FF7D495155428FFFFFFFFFF7FBF8FD7EBD16AA00",
INIT_29 => X"00000002010FFFBF8FC7E3F5EAB45BEDB6FA3800556FA005504051FFFFFFFDFE",
INIT_2A => X"B7DB6FFFDEAA5571C7010FF84125EFF7F1F8FC7EBD568B6DBEDF7DEBA5571EFA",
INIT_2B => X"5092E3F1F8F55AADB6DB7DEBF1FAE82557FC516DEBF1D0410E3F1F8FC7AAD56D",
INIT_2C => X"0000000000000000000016DE3F1EAB55BEDB6FBC7EBF5F8E10007BC516D1C71C",
INIT_2D => X"FFFFFFFFFFFFFFFFFFBFDEAA5D2A954000800154000000000000000000000000",
INIT_2E => X"2A955EFAAD1400AAFFFFFFFFFFFFBFDFEFF7FFFDEAA5D2E95410550415545FFF",
INIT_2F => X"7FFEAB45A2D56AA00002EBDFFFF7D540145FFFFFFFEFF7FBFFFFFAAD16AA0055",
INIT_30 => X"5500155EFF7FBFDFEFAAD568B55AAD568A0008003DFFF0855554AAFFFBFDFEFF",
INIT_31 => X"FFFFFFFEAA55517DE10080400010F7FBE8B55AAD16AB55F7FBFDEAA08557DE00",
INIT_32 => X"10A2D56AB45A2D57DFFFF7FBFFEAA555555400F780001FFF7D16AB55A2D16ABE",
INIT_33 => X"A00087BD55FF5D5555410AAD56AB45AAFFFFFEFAAD168A00557BD55FFA2D5400",
INIT_34 => X"00000000000000000000000000000000000001FFAAD568B45FFFBFFF55A2D568",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000100",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(19),        -- Port A data input
DOA(0)   => data_read_a_hi_256(19),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(19),        -- Port B data input
DOB(0)   => data_read_b_hi_256(19),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_20_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000003",
INIT_01 => X"A75FF80000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"14088080800008400F655001FFCFF80018FA8044000000000000011000000007",
INIT_03 => X"0000000000000000000000000000000024001660380000000000000000004FF8",
INIT_04 => X"000079800014CC02C034001600000000000000101EC0012EE0C0026E1E80F000",
INIT_05 => X"1F0FF433EFF0440C3902100002203F2EFC040388137C3E20C8EEC00284033CC0",
INIT_06 => X"4400080040440C000000000017FD5F239108000155FDC0000010E40087D8787A",
INIT_07 => X"08000EE00000000000000002101FF2002C00000004018001000030817FF50C00",
INIT_08 => X"FF7FCA302C0C00082148000008405550087C0000000000000002412489808000",
INIT_09 => X"44FF60000001EFBEF0040008023FDFC00000000040062A040001071004000013",
INIT_0A => X"000000002B7C0000008000000200000200A0C0040118400FABF9000000480002",
INIT_0B => X"0000000000000000000000000000004200310000000000000000200000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000400040",
INIT_0D => X"000000200000020000004000100203FF6C000000000000000000000000000000",
INIT_0E => X"00600FFC53FF001800000002004080000000000000040900005C848538000010",
INIT_0F => X"00009A9C300020080000800000003CC0080000800000003CC020007800000000",
INIT_10 => X"000000012963C0080000800000003CC0080000800000003CC100800000080000",
INIT_11 => X"800004000000000066C5000020020000000800000000C2E18001000200000800",
INIT_12 => X"000000000052B0200000014200040C2829000400000000000860F98798000100",
INIT_13 => X"4B00400000000002958000240400000000007E1B000040200000000001496004",
INIT_14 => X"4004181800000000005C5A00000200C40808000000000AF0D80080000000000A",
INIT_15 => X"0020141812737DC3020100400001C19C1D80000200400000000000015D140000",
INIT_16 => X"04010080800801810100000000000093EDFF8020000000000001001001000080",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0020000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0C8192608486879E79E681D903000030038200010089054D460400120104D204",
INIT_1B => X"86432190C86432CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB0C30C30C30C3",
INIT_1C => X"C86432190C86432190C86432190C86432190C86432190C86432190C86432190C",
INIT_1D => X"80402000000000000000000000000000000000000000000000001007FE000010",
INIT_1E => X"FFFFFFEAA552E95400082E975FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2A954100",
INIT_1F => X"0FFFFFFFFFFFFFFFFFFFFFFFDEAA5D2A954000800001EFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"BA5D2A97400FF8017410FFFFFFFFFFFFFFFFFFFFFBFDEBA552E974105D2A8000",
INIT_21 => X"FFFFFFFFFFEFF7FBFFEAA5D2E97545FFFFC21FFFFFFFFFFFFFFFFFFFFF7FBFFE",
INIT_22 => X"DF55AAFFD5400FFFFFFFFFFFFFFDFEFF7FFEAA10000417555AAD5555EFFFFFFF",
INIT_23 => X"FDFEFAAD568A0000043DF45AAFBC2010FFFFFFFFFFFFFFDFEFF7D568A1008003",
INIT_24 => X"0001EFFFFFFFFFFFFFBFDF45AAD16AA0008003DF555D51574BAFFFFFFFFFFFFB",
INIT_25 => X"FFFFEBA5D2A95410000A00000000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFDEAA552E954000020955FFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"552A95410552485010FFFFFFFFFFFFFFFFFFF7FBFDEBA5D2E95400140E001C7F",
INIT_28 => X"FFFFFFDFEFF7FFFFEAA5D2E95400E38A17438FFFFFFFFFFFFFFFFEFF7FBFFEBA",
INIT_29 => X"7DBEDF575D7FFFFFFFFFFFFBFDFEFEBF5F8E92552E9556DEBF1C21C7FFFFFFFF",
INIT_2A => X"FD7EBD16AA00000E3DF6DBEF5D2438FFFFFFFFFF7FBFDFC7EBF1E8A00080A155",
INIT_2B => X"5492FFFFFFFEFF7F1F8FD7A2D168A1008043FF6DAAFBC5028FFFFFFFFFF7FBF8",
INIT_2C => X"000000000000000000001FFFFFFFDFEFE3F1FAF55A2D568A0000003FF7D49515",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFEBA552A95410002E820000000000000000000000000",
INIT_2E => X"2E954005D2A82145FFFFFFFFFFFFFFFFFFFFFBFDEAA5D2A954000800155FFFFF",
INIT_2F => X"FFBFDFEFF7FFFDEAA5D2E95410550415410FFFFFFFFFFFFFFDFEFF7FBFFEBA55",
INIT_30 => X"AAD140155FFFFFFFFFF7FBFDFFFFFFBFDEBA5D2A95400A2AA974AAFFFFFFFFFF",
INIT_31 => X"5A2D568A10082E955FFFFFFD7545FFFFFFFEFF7FBFFFFFAAD16AA00552A955EF",
INIT_32 => X"AAFFFBFDFEFF7FFEAB45A2D56AA00002EBDFFFF7D5400BAFFFFFDFEFF7FBFFF5",
INIT_33 => X"A0008003DFFF085555410F7FBFDFEFFFD568B45AAD16AA1008003DFEFAAFBD74",
INIT_34 => X"00000000000000000000000000000000000001EFF7FBFDFEFAAD568B55AAD568",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"FFFFFFFE00000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000000000000000000001F",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(20),        -- Port A data input
DOA(0)   => data_read_a_hi_256(20),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(20),        -- Port B data input
DOB(0)   => data_read_b_hi_256(20),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_21_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"4A302428B824900A128C090A5C1800261500213C005FE812D10420054085A202",
INIT_01 => X"081FFE3440B609703B0427F801A40B8115BC4F655300340288A40D30040E4DD8",
INIT_02 => X"0109095C30C98809800000F9FFFFFFFF149FF1FCA4C0421B182E3490DF145FE4",
INIT_03 => X"084A76341244919000099486400026523C041660BA000100CC12701015007FF8",
INIT_04 => X"000079800014CC03C075161E001118653D2408041FC004AEF000816E1C11F541",
INIT_05 => X"3F0F807BFFE000240100004683103E7FFE02482553FC3C0204EFC25010143CC0",
INIT_06 => X"C42040304101118B84E4880817FD7F028000000101FFE4036450E08247F87870",
INIT_07 => X"0A09000D00204A855B000A08A61FF20C3D004D331D3400805984B7A1FFF00860",
INIT_08 => X"F7FFC08D234B4002030314D0001104500000034089902D0901A021E4015410EA",
INIT_09 => X"B4FFE10158E1FFBEF0440021083DFFCE22DC2880E24D1BFA7C98480802000023",
INIT_0A => X"A31514636FFC00080013029811240444A82422A85180778FAFF82A04B6356DD0",
INIT_0B => X"0600E20806520398C682157A49389667126880806FF917FC30010107688862A2",
INIT_0C => X"1B2451B2451B2451B2451B2451B2451B3228D9228D90800C6120881034003631",
INIT_0D => X"0403000A01282088624001201A8C43FF7C00100102A53208B2A246406081B245",
INIT_0E => X"C4053FFD5BFF00A04A00200602CA520011000880044402104803400400189000",
INIT_0F => X"63009140094D81A5040605800B506901A3040605401360562027218196506102",
INIT_10 => X"02811209062801A3040605800B506901A50406054013605604350B812822A002",
INIT_11 => X"0B811068C00049A0A5820A3C1725A8006C0A40404D058320496C2C9C600890A2",
INIT_12 => X"AC808127C454402483153A3A895BB3C1E2E820704020381702C1AAA2C4B3F435",
INIT_13 => X"CC1B154510413CC2A200501B400A40018A00C80400040D8AA288209AA2198361",
INIT_14 => X"0141AA00418080460678A4012288463B2050302019200B00206C35901024D910",
INIT_15 => X"2440470C8A9310280C0180302A01427D060022011606E800E00169C19A00048A",
INIT_16 => X"40100448008004000000E07008010003EFFFE0373056024B0111801198823314",
INIT_17 => X"0100401004010040100401004010040100401004010040100401004010040100",
INIT_18 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_19 => X"0000000000000000000000401004010040100401004010040100401004010040",
INIT_1A => X"BEFFFFF7F7FFF3CF3CFFFF9FE0FF9FEEFF7FFDF7FF3EFC2FF8107F3DFDF7E000",
INIT_1B => X"FF7FBFDFEFF7FBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEF",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FBFDFE",
INIT_1D => X"80002000000000000000000000000000000000000000000000001007FE00003F",
INIT_1E => X"FFFFFFEBA5D2A954100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974000",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFEBA552A97400082A975FFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"AA5D2E974100800155EFFFFFFFFFFFFFFFFFFFFFFFFFEAA552E95400082E975F",
INIT_21 => X"FFFFFFFFFFFFFFFFFDEAA5D2A95400080000000FFFFFFFFFFFFFFFFFFFFFFFDE",
INIT_22 => X"74105D2A80000FFFFFFFFFFFFFFFFFFFFFBFDEBA5D2E974005D2E80000FFFFFF",
INIT_23 => X"FFFFFF7FBFDEBA552A954005D2E97410FFFFFFFFFFFFFFFFFFFFFBFDEBA552E9",
INIT_24 => X"0001FFFFFFFFFFFFFFFFFFFFF7FBFFEBA5D2A97400FF80174BAFFFFFFFFFFFFF",
INIT_25 => X"FFFFEBA5D2E97400000400000000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFEBA5D2A95410000A001FFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"552E954000020955EFFFFFFFFFFFFFFFFFFFFFFFFFEAA552E97400002E955FFF",
INIT_28 => X"FFFFFFFFFFFFFBFDEAA5D2A974101400155C7FFFFFFFFFFFFFFFFFFFFFFFDEAA",
INIT_29 => X"00552A80010FFFFFFFFFFFFFFFFFFF7FBFDEBA5D2E95400140E00000FFFFFFFF",
INIT_2A => X"FEFF7FBFFEBA552A95410552485038FFFFFFFFFFFFFFFFFFF7FBFDEBA552E974",
INIT_2B => X"74AAFFFFFFFFFFFFFFFFEFF7FBFFEAA5D2E97400412497438FFFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000001C7FFFFFFFFFFFFFFDFEFF7FFFFEAA5D2E95400E38A1",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974000004000000000000000000000000000",
INIT_2E => X"2E97400002E975FFFFFFFFFFFFFFFFFFFFFFFFFFEBA552A95410002E821FFFFF",
INIT_2F => X"FFFFFFFFFFFBFDEAA5D2A954000800155EFFFFFFFFFFFFFFFFFFFFFFFFDEAA55",
INIT_30 => X"5D2A82010FFFFFFFFFFFFFFFFEFF7FBFDEBA552A974105D0015545FFFFFFFFFF",
INIT_31 => X"FF7FFFFEAA5D2A974005D2E82010FFFFFFFFFFFFFFDFEFF7FBFFEBA552E95400",
INIT_32 => X"AAFFFFFFFFFFFFBFDFEFF7FFFDEAA5D2E954105504154AAFFFFFFFFFFFFFFDFE",
INIT_33 => X"EBA5D2A95400A2AA974BAFFFFFFFFFF7FBFDFEFFFFFFDEBA552E974000004154",
INIT_34 => X"0000000000000000000000000000000000000155FFFFFFFFFF7FBFDFFFFFFBFD",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(21),        -- Port A data input
DOA(0)   => data_read_a_hi_256(21),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(21),        -- Port B data input
DOB(0)   => data_read_b_hi_256(21),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_22_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"5290F4CDE914905A14A43D33F488243E17122300F55FEB189B343A1140548380",
INIT_01 => X"A94007B259F6A975386262000C344BA9573C6FF57B18A5FB0ABFCD3C2C5F4F0C",
INIT_02 => X"877FE30EB378008D202551040030071869D0040180AC4B685F6E26FAA0810006",
INIT_03 => X"431965109E4481D6B5AAD6875AD6AB5A1815600802888808DEA83552954D3000",
INIT_04 => X"492C0020220001010E4916C884DCD607E5EC2A344103E48003D0800023D0072C",
INIT_05 => X"00107C441001100D620A06D683018001023D37E5088043620101179092540112",
INIT_06 => X"9108E1550544A451E0CE1AA94000206B541C08414402365774611E047020008E",
INIT_07 => X"809DA02F56A92FD7247E10305C40040D136E6A023F7FCF780C4C0528800C8028",
INIT_08 => X"00803A884B5B5206B7C3391F288551002401E993AF59012740A2E4F65586923D",
INIT_09 => X"040081C91AA010000560141801002028A83D2A08E06D0002FED9680A0E002A94",
INIT_0A => X"A71514E700838460402635019FBFE7FCA13520F8D580A08044081201206334A0",
INIT_0B => X"00A0220103D2A512C6A8C4F0011550070368000A0004D0000002126F30C902A2",
INIT_0C => X"0385503855038550385503855038550392A81C2A81C00280000C200006405A08",
INIT_0D => X"0D0E153941A8B1A262CA542A9A8D6C0010A1001002C500268ACA419412503855",
INIT_0E => X"089180008800143D83888281A2034A85014280A14050A01509E050854498B294",
INIT_0F => X"6706B3C189CD84ACD20B03001E387D04AC560B02401E387E1028AC0450080410",
INIT_10 => X"0201570B036C04AC560B03001E387D04ACD20B02401E387E24708E7E242000C2",
INIT_11 => X"8E7E1C20A0106EA167C84EBF052A8E010C0180606E86C3F459DC08DA90245887",
INIT_12 => X"189980254CDEC22A98032A22C50EAC462030A01800407C2700C2ACA2C0F04470",
INIT_13 => X"CC1154C258012D86F601A2E49003400138C0DA2443A208AA612C0096C3798225",
INIT_14 => X"025483C1E0C0006B085CEC03858958D15310201015504B512044A3133004A99B",
INIT_15 => X"9512C6FC01A1421006028038720640310643858162712020B001AA415F290E16",
INIT_16 => X"110445E22022365034A8EA754008004C0200323001182122548881649D16B046",
INIT_17 => X"1044110441104411044110441104411044110441104411044110441104411044",
INIT_18 => X"0401004010040100401004010040100401004010040100441104411044110441",
INIT_19 => X"22890000000003FFFFFFFF900401004010040100401004010040100401004010",
INIT_1A => X"9EFFDFF7F5F777DF7DF7DF5FEFBFBFDEFE8FF1F7DEBD6FEFF7EF6FDF7DF7D051",
INIT_1B => X"7F3F9FCFE7F3F9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7",
INIT_1C => X"E7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE",
INIT_1D => X"00000000000000000000000000000000000000000000000000001007FE00000F",
INIT_1E => X"FFFFFFEBA5D2E974000800021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E954000004001FFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"BA552A97400002A801FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2A954100804021F",
INIT_21 => X"FFFFFFFFFFFFFFFFFFEBA552A97400082A975FFFFFFFFFFFFFFFFFFFFFFFFFFE",
INIT_22 => X"5400082E975FFFFFFFFFFFFFFFFFFFFFFFFFFEAA552E95410002A955FFFFFFFF",
INIT_23 => X"FFFFFFFFFFFEAA552E95400002E975EFFFFFFFFFFFFFFFFFFFFFFFFFEAA552E9",
INIT_24 => X"000000FFFFFFFFFFFFFFFFFFFFFFFDEAA5D2E97410080015545FFFFFFFFFFFFF",
INIT_25 => X"FFFFEBA5D2E97410080002000000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974000004001FFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"5D2A95410000A001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2A954000804021FFF",
INIT_28 => X"FFFFFFFFFFFFFFFFEBA552A97400082E821FFFFFFFFFFFFFFFFFFFFFFFFFFEBA",
INIT_29 => X"10082A975EFFFFFFFFFFFFFFFFFFFFFFFFFEAA552E97400002E955FFFFFFFFFF",
INIT_2A => X"FFFFFFFFDEAA552E954000020955C7FFFFFFFFFFFFFFFFFFFFFFFFEAA552E954",
INIT_2B => X"5545FFFFFFFFFFFFFFFFFFFFFFFDEAA5D2A974001C24975C7FFFFFFFFFFFFFFF",
INIT_2C => X"00000000000000000000000FFFFFFFFFFFFFFFFFFFFFBFDEAA5D2A9741014001",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800020000000000000000000000000",
INIT_2E => X"2A954000800021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974000004001FFFFF",
INIT_2F => X"FFFFFFFFFFFFFFEBA552A95410002E821FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_30 => X"002E975EFFFFFFFFFFFFFFFFFFFFFFFFFEAA552A97400082A801FFFFFFFFFFFF",
INIT_31 => X"FFFFBFDEAA5D2E95410082E955EFFFFFFFFFFFFFFFFFFFFFFFFDEAA552E97400",
INIT_32 => X"45FFFFFFFFFFFFFFFFFFFFFBFDEAA5D2A95400080015545FFFFFFFFFFFFFFFFF",
INIT_33 => X"EBA552A974105D0015555FFFFFFFFFFFFFFFFFFF7FBFDEBA5D2A974005504175",
INIT_34 => X"0000000000000000000000000000000000000010FFFFFFFFFFFFFFFFEFF7FBFD",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"FFFFFFFE00000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000000000000000000001F",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(22),        -- Port A data input
DOA(0)   => data_read_a_hi_256(22),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(22),        -- Port B data input
DOB(0)   => data_read_b_hi_256(22),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_23_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"EF20906D902424807BC8241BC81801B97D38AD3C0800103362A6741C80A12A02",
INIT_01 => X"001FFF8409F089003B4422000D80C80106804A7951C5B9D1C828043EA28838F9",
INIT_02 => X"073B8858218C2C50801000F9FFEFF8E72CA7F5FC2E048026496834D84721DFE0",
INIT_03 => X"2C4360101A4001001005080400401420350016E0BB222341C312000014006FF8",
INIT_04 => X"00017B810015DC03D034201E14000036486008101FC0002EE006297E1C05F561",
INIT_05 => X"BF0F817FFFE80100004044800080BEFFFC0248005FFC3C18A5FFC2444484BCC0",
INIT_06 => X"00000070604191C93F02800017FF7F002000020001FFC0832050E00047F97870",
INIT_07 => X"AE4080091A0071070FA07A1CB23FFA403F0C4D23BF7C0EF85788B681FFFC6C20",
INIT_08 => X"F7FFD8880A034AC096620C46AC5055508401A24684227DB880000008B05001A3",
INIT_09 => X"21FFE0004047FFBEF2000000001DFFC612C0C04001000BF8000000804000003F",
INIT_0A => X"000000006FFEA002020626995FBE077430001E734020DF0FAFF5080496044B51",
INIT_0B => X"0600C48907120AC81083315A49388660180082A06FF907FC3081812048006000",
INIT_0C => X"182021820218202182021820218202182010C1010C10800C6120885430003631",
INIT_0D => X"80600020040030090000012A500003FF7E081881902233483828864860A18202",
INIT_0E => X"C7043FFD5FFF00A04BC010A7724B100008000400020000415003001000400002",
INIT_0F => X"290C2909080A872BC4FC8500054840072FC0FC8440054840200705F986106542",
INIT_10 => X"0180F1082E00072FC0FC8500054840072BC4FC84400548402214A380380B2080",
INIT_11 => X"A380344920080B21810240AB182EB37C380B40800707011001B43253EE50C822",
INIT_12 => X"E4000026C00C00042BD4149067465910640A0050C060A0028063672A00019214",
INIT_13 => X"800CCB050001344060211629580B80022480A444111706658280009A2030019C",
INIT_14 => X"232D6D0100C040250200845132C10BE200403018061101A220339C800004D801",
INIT_15 => X"2A5493B8E287E03808480060E40C83C1405132C90742E408D0082140820944CB",
INIT_16 => X"00802000100100000000000004002403EFFF8002385F03490101946500140210",
INIT_17 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_18 => X"8020080200802008020080200802008020080200802008020080200802008020",
INIT_19 => X"0000000000000000000000008020080200802008020080200802008020080200",
INIT_1A => X"0000000000000000000000000000000000000000000000000040000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"80400000000000000000000000000000000000000000000000001007FE000000",
INIT_1E => X"FFFFFFEBA5D2E974100000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100004021FFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"BA5D2E954000800001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974000800021F",
INIT_21 => X"FFFFFFFFFFFFFFFFFFEBA5D2E954000004001FFFFFFFFFFFFFFFFFFFFFFFFFFE",
INIT_22 => X"54100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2A954100000021FFFFFFFF",
INIT_23 => X"FFFFFFFFFFFEBA5D2A954100800021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2A9",
INIT_24 => X"0001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA552A97400002A801FFFFFFFFFFFFFFF",
INIT_25 => X"FFFFEBA5D2E97410080400000000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800021FFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"5D2E974000004001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100004021FFF",
INIT_28 => X"FFFFFFFFFFFFFFFFEBA5D2E954000800001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA",
INIT_29 => X"100004021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2A954000804021FFFFFFFFFF",
INIT_2A => X"FFFFFFFFFEBA5D2A95410000A001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2A954",
INIT_2B => X"21FFFFFFFFFFFFFFFFFFFFFFFFFFEBA552A97410080E001FFFFFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA552A97400082E8",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804000000000000000000000000000",
INIT_2E => X"2E974100000021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800021FFFFF",
INIT_2F => X"FFFFFFFFFFFFFFEBA5D2E974000004001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_30 => X"0800021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E954000804021FFFFFFFFFFFF",
INIT_31 => X"FFFFFFFEBA552A954100004001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2A95400",
INIT_32 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA552A95410002E821FFFFFFFFFFFFFFFFFFF",
INIT_33 => X"EAA552A97400082A801EFFFFFFFFFFFFFFFFFFFFFFFFFEAA552A97410002A821",
INIT_34 => X"00000000000000000000000000000000000001EFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"FFFFFFFE00000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000000000000000000001F",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(23),        -- Port A data input
DOA(0)   => data_read_a_hi_256(23),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(23),        -- Port B data input
DOB(0)   => data_read_b_hi_256(23),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_24_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100600007FFF000080108004000800020000840041000080808",
INIT_02 => X"172A00D000EF8210000000F9FFEFF8E7240FF1FC224087B1000639401D005FC0",
INIT_03 => X"00003A2E200811000000000400000000340016603A0000004860400014006FFF",
INIT_04 => X"000079800014CC03C034001E04010850300000101FC0002EE000006E1C00F500",
INIT_05 => X"1F0F8033FFE000000000000000003E2FFC024800137C3C0000EFC00000003CC0",
INIT_06 => X"00000040004111CE08AA800017FD7F000000000001FFC0000010E00007F87870",
INIT_07 => X"001080040814210254000A00B21FF2003F2A80D5000006E461803081FFF40000",
INIT_08 => X"F7FFD88D2B4A02C0940018EB0A1000058400810205E2D8030900004D925821CC",
INIT_09 => X"20FFE0000001FFBEF0000000001DFFC002C0000000000BF80000000000000003",
INIT_0A => X"000000006FFE80000015406A80000338800002500000470FAFF0080496044950",
INIT_0B => X"0600C008140800080000100248288660100080806FD107FC3000000000006000",
INIT_0C => X"182001820018200182001820018200182000C1000C10800C6020881030002431",
INIT_0D => X"000900160000000000000000000003FF7C001001002032083020060060018200",
INIT_0E => X"C4043FFD5BFF0000410000000041100000000000000000004003000000000000",
INIT_0F => X"1080012302010049400086C02200420049400087802200412027059996516100",
INIT_10 => X"0300081406100049400086C0220042004940008780220041248190818403A042",
INIT_11 => X"90814C09C01010400132100106836001504240E01040051200200D06410C1924",
INIT_12 => X"680C0100010408240BD80008983596CD86EA84104060503C0B00002025023481",
INIT_13 => X"90164F40086000082062C1B6600BC000C300818044000B27A0043000041202CD",
INIT_14 => X"2577FE4080C08010842180C40018545BBA00301808A0810C0059AD0180200020",
INIT_15 => X"04100852B931F00800010081980B042D2044001850ED8808F00050A002C11000",
INIT_16 => X"00000000000000000000000000000003EFFF80037046031E0110001100A4820C",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"BEC99E61848655D75D7FCB598CC0AEEAF6E7CC1132CD73C8261273B444199000",
INIT_1B => X"0F0783C1E0F07BEFBEFBEF9E79E79E79E79E7BEFBEFBEFBEFBEFBE7BE7BE7BE7",
INIT_1C => X"E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E",
INIT_1D => X"80402000000000000000000000000000000000000000000000001007FE000001",
INIT_1E => X"FFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800021FFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"BA5D2E974100000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100000001F",
INIT_21 => X"FFFFFFFFFFFFFFFFFFEBA5D2E974100004021FFFFFFFFFFFFFFFFFFFFFFFFFFE",
INIT_22 => X"74000800021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974000004001FFFFFFFF",
INIT_23 => X"FFFFFFFFFFFEBA5D2E974000800001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9",
INIT_24 => X"0001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E954000800001FFFFFFFFFFFFFFF",
INIT_25 => X"FFFFEBA5D2E97410080402000000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"5D2E974100800021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800021FFF",
INIT_28 => X"FFFFFFFFFFFFFFFFEBA5D2E974100000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA",
INIT_29 => X"000004001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100004021FFFFFFFFFF",
INIT_2A => X"FFFFFFFFFEBA5D2E974000004001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_2B => X"01FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E954000800021FFFFFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9540008000",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804020000000000000000000000000",
INIT_2E => X"2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFF",
INIT_2F => X"FFFFFFFFFFFFFFEBA5D2E974100800021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_30 => X"0000021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100000001FFFFFFFFFFFF",
INIT_31 => X"FFFFFFFEBA5D2E974000004021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E97410",
INIT_32 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974000004001FFFFFFFFFFFFFFFFFFF",
INIT_33 => X"EBA5D2E954000804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E954000004021",
INIT_34 => X"00000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(24),        -- Port A data input
DOA(0)   => data_read_a_hi_256(24),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(24),        -- Port B data input
DOB(0)   => data_read_b_hi_256(24),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_25_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100200002000000080100004000000020000800041000080808",
INIT_02 => X"1000218000000800000000F9FFEFF8E738FFF1FC20400400000004455A375FE0",
INIT_03 => X"00002000000001000000000400000000340016623A0000004000000014006FFF",
INIT_04 => X"924279824C94CC1BE0B4001F20000000020380401FE0082EF000106E1C00F500",
INIT_05 => X"1F0F8033FFF048202582800100523E2FFE024820137C3C0040EFE02000003CE4",
INIT_06 => X"D4A00671414191800000800017FD7F038100201101FFC0000010E08A07FC7870",
INIT_07 => X"080000000000000000000A00B21FF2003E0000000000066041803081FFFC2C60",
INIT_08 => X"F7FFFA0008000200A0400002280000050400800204000000000201202B800000",
INIT_09 => X"B4FFF0008001FFBEF80C40630C7DFFEEBAF0008002021BF80000400A02000003",
INIT_0A => X"000000006FFF800C0400000000000330080000500006470FAFFD29F7DE565971",
INIT_0B => X"0600C008040000080000100248688760101080806FD107FC3018000000006000",
INIT_0C => X"182001820018200182001820018200182000C1000C10800EE6618911398524B1",
INIT_0D => X"000000000000000000000002500003FF7C001001002032083120060060018200",
INIT_0E => X"C6043FFD5BFF00A04B80608003CB120C11060883044582114013412080000000",
INIT_0F => X"000000200200000900000400200000000900000400200000200701E186106140",
INIT_10 => X"0000001000000009000004002000000009000004002000000000808000002000",
INIT_11 => X"8080000800000000001010000002200000004000000004000000000240000020",
INIT_12 => X"2000000001000004031802000004100000100024400000000800800001000000",
INIT_13 => X"0000410000000008000000204004000000000100040000208000000004000004",
INIT_14 => X"0004200001000200000100040000004200004020000000040000840000000020",
INIT_15 => X"00000010800000000C0A00000000040000040000004080000000000000401000",
INIT_16 => X"451044C82082068C0200000008014023EFFFC006304602080100000100000308",
INIT_17 => X"1104411044110441104411044110441104411044110441104411044110441104",
INIT_18 => X"1044110441104411044110441104411044110441104411044110441104411044",
INIT_19 => X"00002FFFFFFFFFFFFFFFFFC11044110441104411044110441104411044110441",
INIT_1A => X"042824014C48569A69AFEE9E50B2894A196A8C5A2932F7C8086034EC15DA0808",
INIT_1B => X"6231188C46231249249249249249249249249041041041041041041249041249",
INIT_1C => X"562B158AC562B158AC562B158AC562B158AC562B158AC562B158AC56231188C4",
INIT_1D => X"80400000000000000000000000000000000000000000000000001FFFFE00002C",
INIT_1E => X"FFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"BA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001F",
INIT_21 => X"FFFFFFFFFFFFFFFFFFEBA5D2E974100800021FFFFFFFFFFFFFFFFFFFFFFFFFFE",
INIT_22 => X"74100000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800001FFFFFFFF",
INIT_23 => X"FFFFFFFFFFFEBA5D2E974100000021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9",
INIT_24 => X"0001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100000001FFFFFFFFFFFFFFF",
INIT_25 => X"FFFFEBA5D2E97410080400000000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFF",
INIT_28 => X"FFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA",
INIT_29 => X"100800001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800021FFFFFFFFFF",
INIT_2A => X"FFFFFFFFFEBA5D2E974100800021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_2B => X"01FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100000021FFFFFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741000000",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804000000000000000000000000000",
INIT_2E => X"2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFF",
INIT_2F => X"FFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_30 => X"0804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFF",
INIT_31 => X"FFFFFFFEBA5D2E974100800001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E97410",
INIT_32 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800021FFFFFFFFFFFFFFFFFFF",
INIT_33 => X"EBA5D2E974100000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100800021",
INIT_34 => X"00000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"FFFFFFFE00000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000000000000000000001F",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(25),        -- Port A data input
DOA(0)   => data_read_a_hi_256(25),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(25),        -- Port B data input
DOB(0)   => data_read_b_hi_256(25),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_26_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"E9264EAB20190CA3BA4997AA9002AE9C001006B0778015CFA17E0811039879C7",
INIT_01 => X"F1FFF9BB1F773C7F9BB07DFFFDD863FC5FFF3FEFFBBF9FFB22FFFBC7B9F30686",
INIT_02 => X"1B33188302E708180F6FFBFFFFCFFFFF9C7FF7FC24350B99082400001D00DFD8",
INIT_03 => X"4A53D958C50000DCE7366303739CD98C27C57EF57980014F271807E3C9E9CFF8",
INIT_04 => X"DBFAFBD7FB1CDEBEF1BE17F7AC88042787FBFFF8FEE9FF7EE6F4C0EE1FFAF869",
INIT_05 => X"5F0FFEB3EFFEFFBDA7F7FED508707E2EFEBF6FFEB37C3FF302EEEDFF9B487CF6",
INIT_06 => X"67F2B27AFAD11587B7C094F1FFFFDF0FAF4E8FAA67FDDB7FB870FF30FFDEF87F",
INIT_07 => X"08180EF060C18E5BEFB051225CDFF7002C4EEDE77F6E0EFD044ABC817FFFDD35",
INIT_08 => X"FF7FC8790E46426CE06C2C7E381041460C7E8C1A35DF80000C0084C9188302E7",
INIT_09 => X"2CFF7A27B303EFBEFAFCC2E35E7FDFD147CCF3F583FA3FFF7D6000EC75088ED3",
INIT_0A => X"5A3A3B5AFF7CFACFAFE776F39FF7077E29D83CFAE601602FEBFFCDF7DEE77DF7",
INIT_0B => X"3EB1EDDCDEBCFF589807B70AD9A99EE41FD18884FFF19FFC71FEFED7B251E747",
INIT_0C => X"1AF181AF181AF181AF181AF181AF181AF4C0D78C0D718ADEEE61D99B7BE2A433",
INIT_0D => X"B9EC20181CC1F73F87501DED3409BFFFEFFEBCEBFE68370CFA6D07407481EF18",
INIT_0E => X"CE04FFFFF3FF1F5F5475BD7F72E4D75EBFAF5FD7AFEFDFFAF59B6FF28FE1D406",
INIT_0F => X"7C040101480807D17B0004001F804007D17B0004001F8040212F35FFC6D86D70",
INIT_10 => X"0001DC00068007D17B0004001F804007D17B0004001F804006F6008140002000",
INIT_11 => X"0081800800007B000102C0801FB02683800040007700011801003DE050A70020",
INIT_12 => X"32130207080D012CEFF41008D188D502100B02004000F01900039020040206F6",
INIT_13 => X"A01F21A2C40039006823F80048100003F0008004D8100F90D162001C803403E2",
INIT_14 => X"27F020A07400007C040085581019D602451500001EC00100247C46426080E101",
INIT_15 => X"2010EA40EA00020C830100F0D000022180581019F40084800001F100020B6040",
INIT_16 => X"EFFBFEFDFDDFE7DD87FEFF7FF796FFFFFDFFC017FEFFD7E841001D8197DCC3F0",
INIT_17 => X"BFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAF",
INIT_18 => X"FAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFE",
INIT_19 => X"88646FFFFFFFFFFFFFFFFFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEB",
INIT_1A => X"86EBCAF55357E1C71C751D53C44B15BCF491E166CC853E8117696853F86EDB5C",
INIT_1B => X"130984C261309861861861861861861861861861861861861861861A69A69861",
INIT_1C => X"6130984C26130984C26130984C26130984C26130984C26130984C26130984C26",
INIT_1D => X"80400000000000000000000000000000000000000000000000001007FE000002",
INIT_1E => X"FFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"BA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021F",
INIT_21 => X"FFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFE",
INIT_22 => X"74100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFF",
INIT_23 => X"FFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9",
INIT_24 => X"0001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFF",
INIT_25 => X"FFFFEBA5D2E97410080400000000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFF",
INIT_28 => X"FFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA",
INIT_29 => X"100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFF",
INIT_2A => X"FFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_2B => X"21FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008040",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804000000000000000000000000000",
INIT_2E => X"2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFF",
INIT_2F => X"FFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_30 => X"0804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFF",
INIT_31 => X"FFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E97410",
INIT_32 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFF",
INIT_33 => X"EBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001",
INIT_34 => X"00000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(26),        -- Port A data input
DOA(0)   => data_read_a_hi_256(26),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(26),        -- Port B data input
DOB(0)   => data_read_b_hi_256(26),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_27_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"00080A40000A41248002029000050A088000008242A0004404480002000A1155",
INIT_01 => X"F1FFF1C11F781C129C107DFFFE0860941E81258CA2B71C2220EC1B86E1A00002",
INIT_02 => X"4000002100000014400FF6FFFF0FFFFF8007F1FC211100014200800000887FC0",
INIT_03 => X"0842D85841000098C63061026318C18404C459757000015F00088BE3C0618FF8",
INIT_04 => X"DBEAE5D6D91C2EBCE1B21EA72C00000007FBE7C8F8E9EF79E6D440E91FDAE061",
INIT_05 => X"5C8FFCB38FF6B68984B5BCE408347E28FEBF6FEEB3723F7102E8EDBF8A4872F6",
INIT_06 => X"6E62106ADAD14180035044F1FFFC9F0C0E4C8DAAEFF1DB7FA868FE30EF1CE47E",
INIT_07 => X"0014401060C180190310540118DFF1000C0849673F6C06FE000A38007FF13115",
INIT_08 => X"F47FC80208808210880C00020814000044008C1A340C00000A08000000210000",
INIT_09 => X"04FC721491038F7DF8BEC2E39C5F1FD047CEF1B582D83FF779200062B12A8EC3",
INIT_0A => X"02606042787C5AC5ADC424B39FB6073D00D8048A6201002F83F04DFFDE83FDD6",
INIT_0B => X"56B5F0DEFABC705488069302DBA98EAC16C1A884FFE18FFD757E7ED7A211EC0C",
INIT_0C => X"186881868818688186881868818688187840C3440C35A8DFEE61CB9979AAA433",
INIT_0D => X"D1F820101441DA3A8310198C34089BFF8DD6B56B6F28378C7E2D07007801C688",
INIT_0E => X"E4047FFD23FF315D54358D593474955AB6AD5B56ADAB5FAAE58B2F628EA0C407",
INIT_0F => X"7C0400004C080791290004001D80001791290004001D8000210F15879715710A",
INIT_10 => X"0001DC0000801791290004001D80001791290004001D800012F6008040002000",
INIT_11 => X"0080800800007B000000E0801BB020828000400077000008210035E040830020",
INIT_12 => X"220202070801010C6F1410085188D500100102004000F01900031000060202F6",
INIT_13 => X"205D2120840039000813F80040100003F0000000F8100E909042001C80040BA2",
INIT_14 => X"07F020201400007C040001781011D602040500001EC00000057444404080E100",
INIT_15 => X"2000EA40EA000004810100F0D000020080781011F40080800001F1000003E040",
INIT_16 => X"AB6BDE75ED5EC71385FC2512E3565BBBF1FFC00636EED7E841000D81924C43F0",
INIT_17 => X"B6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6AD",
INIT_18 => X"6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADA",
INIT_19 => X"88747FFFFFFFFFFFFFFFFFAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB",
INIT_1A => X"00780401CBC8400000052412F84E2168100481CA8604368008402F02104A4716",
INIT_1B => X"4020100804020000000000000000000000000000000000000000208000000000",
INIT_1C => X"140A05028140A05028140A05028140A05028140A05028140A050281402010080",
INIT_1D => X"80400000000000000000000000000000000000000000000000001007FE000028",
INIT_1E => X"FFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"BA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001F",
INIT_21 => X"FFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFE",
INIT_22 => X"74100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFF",
INIT_23 => X"FFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9",
INIT_24 => X"0001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFF",
INIT_25 => X"FFFFEBA5D2E97410080400000000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFF",
INIT_28 => X"FFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA",
INIT_29 => X"100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFF",
INIT_2A => X"FFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_2B => X"21FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008040",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804000000000000000000000000000",
INIT_2E => X"2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFF",
INIT_2F => X"FFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_30 => X"0804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFF",
INIT_31 => X"FFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E97410",
INIT_32 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021FFFFFFFFFFFFFFFFFFF",
INIT_33 => X"EBA5D2E974100804021FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804021",
INIT_34 => X"00000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"FFFFFFFE00000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000000000000000000001F",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(27),        -- Port A data input
DOA(0)   => data_read_a_hi_256(27),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(27),        -- Port B data input
DOB(0)   => data_read_b_hi_256(27),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_28_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"02200AA400180030808802A900002A08001280A08A801044104A1000001818C3",
INIT_01 => X"50A00011460214428114180000882214413D0A71592A01D92213D28005210202",
INIT_02 => X"1444428102100884000AA30200000000C1000401041108404400022220800000",
INIT_03 => X"461080404900000C6314A900318C52A40051081000888806108802A141288001",
INIT_04 => X"00800040110102000902002000888400081045A8A00003C00000500000080008",
INIT_05 => X"0000000000024CA0A0101800032000400000000B800000014000000B08180000",
INIT_06 => X"0040B0000804001040000450A00080444A002480220009A88800009A88000000",
INIT_07 => X"088400122448908A204020004080010000408200000001000002080000099000",
INIT_08 => X"0000028040101004200C21002084555500004489120509244022801244810210",
INIT_09 => X"9000008101400000049016080102000220001110001020058320402A16002650",
INIT_0A => X"A53534A50000080080E041000000008000C81000220020A00004000000300003",
INIT_0B => X"0090024440245400082D0220800008000081022C0000080000206CB0821086A6",
INIT_0C => X"02C0A02C0A02C0A02C0A02C0A02C0A02C050160501600240010860CC04200280",
INIT_0D => X"1884200810C1631181500CA60400B40080720020240A00004005800800206C0A",
INIT_0E => X"0A00C000200005000010040A0020CC000200010000800920040804020A605400",
INIT_0F => X"0000000140000010290000000280000010290000000280000100180210410442",
INIT_10 => X"0000000004800010290000000280000010290000000280000002000040000000",
INIT_11 => X"0000800000000000000280000010008280000000000000180000002000830000",
INIT_12 => X"0202020000090100548000000080000010010200000000000000900000000002",
INIT_13 => X"2000202084000000480008000010000000000004880000101042000000240002",
INIT_14 => X"0080002014000000000005080000800004050000000000002400404040800001",
INIT_15 => X"00002000000000048100000000000020800800008000008000000000000A2000",
INIT_16 => X"80210810840861CD33548542A10209D4100000010200400000000880035840A0",
INIT_17 => X"0200802008020080200802008020080200802008020080200802008020080200",
INIT_18 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_19 => X"22E1000000000000000000002008020080200802008020080200802008020080",
INIT_1A => X"200360D4141D630C30C7788C0211102C110A00246972C0C19D0154BD89A40A0C",
INIT_1B => X"6030180C06030208208208208208208208208208208208208208208208208208",
INIT_1C => X"160B0582C160B0582C160B0582C160B0582C160B0582C160B0582C16030180C0",
INIT_1D => X"80400000000000000000000000000000000000000000000000001007FE00002C",
INIT_1E => X"FFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"BA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001F",
INIT_21 => X"FFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFE",
INIT_22 => X"74100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFF",
INIT_23 => X"FFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9",
INIT_24 => X"0001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFF",
INIT_25 => X"FFFFEBA5D2E97410080400000000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFF",
INIT_28 => X"FFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA",
INIT_29 => X"100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFF",
INIT_2A => X"FFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_2B => X"01FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008040",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804000000000000000000000000000",
INIT_2E => X"2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFF",
INIT_2F => X"FFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_30 => X"0804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFF",
INIT_31 => X"FFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E97410",
INIT_32 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFF",
INIT_33 => X"EBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001",
INIT_34 => X"00000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"FFFFFFFE00000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000000000000000000001F",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(28),        -- Port A data input
DOA(0)   => data_read_a_hi_256(28),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(28),        -- Port B data input
DOB(0)   => data_read_b_hi_256(28),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_29_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"79964E4BA01DACAB9E659792D00AAE160002829C7FDFEFCEE97C2815039D70C3",
INIT_01 => X"50BFF9AB0775343F9AB01DF80D5821FC0FFF3FEFD1AF9FF1207FFBC7B9720586",
INIT_02 => X"0B33180300E700080F6AAA7BFFC007189C7FF2FC003503980A0000001D00DFD8",
INIT_03 => X"0401D940CD0000C8421A2B03210868AC23403E903900010E271006A148A0C000",
INIT_04 => X"49B87A417315D20A313E17F1800000058013DDF8BE21F36E02F0D06E03E8F800",
INIT_05 => X"1F007E33E01A4D9C87525E5101603E6E023D27DA937C03E340EE25CB9B483C12",
INIT_06 => X"4570301028001487B7809450B7FFC007AB0E068023FC3BFC98101F109FC6780F",
INIT_07 => X"00080EF020408EC8CFA01122149FF700200665A35D260B250442BC8100177C20",
INIT_08 => X"FF00007906464068406C0C7E100000020C7E840A15D6800044200049180300E7",
INIT_09 => X"A8FF18222341E0820AD40201423FC00122C4935001722BFD056040A452000443",
INIT_0A => X"5A2A2B5AAF00A80A82C332D18ED301D229C82C7AA600402FE80B8813485534A2",
INIT_0B => X"28102D445624DB481806A628810018400B9100042FF0180000ABFEF892508545",
INIT_0C => X"00D1A00D1A00D1A00D1A00D1A00D1A00D4D0068D006000428200508A0A600280",
INIT_0D => X"B0E8201018C1561E855008C50401B7FFE27A08A0B64A0100CA45814814A04D1A",
INIT_0E => X"4400DFFFF0001F1F0050342D42A086040B02058102C48970541944B20FA15402",
INIT_0F => X"00000101480000507B00000002804000507B000000028040212034FAD2892832",
INIT_10 => X"00000000068000507B00000002804000507B0000000280400402000140000000",
INIT_11 => X"00018000000000000102C0000410068380000000000001180000082010A70000",
INIT_12 => X"12130200000D0120ED64000080800002100B0200000000000000902004000402",
INIT_13 => X"A00220A2C4000000682008000810000000008004D80001105162000000340042",
INIT_14 => X"208000A074000000000085580008800045150000000001002408424260800001",
INIT_15 => X"001020000000020C8300000000000021805800088000048000000000020B6000",
INIT_16 => X"C4B12C989489418D13FE7F3FFD8BADB7FC004012CA5141600000198087D8C0F0",
INIT_17 => X"0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02",
INIT_18 => X"B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C",
INIT_19 => X"00602FFFFFFFFFFFFFFFFFC0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0",
INIT_1A => X"AEFFFFF7E7EFBFFFFFFAEF1DE1EF9F96EE7FFDF7FE78FC2FE8847F3FFDFFEA0C",
INIT_1B => X"F7FBFDFEFF7FBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBAEBAEBAEBAEB",
INIT_1C => X"FF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEF",
INIT_1D => X"80400000000000000000000000000000000000000000000000001007FE00003E",
INIT_1E => X"FFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"BA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001F",
INIT_21 => X"FFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFE",
INIT_22 => X"74100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFF",
INIT_23 => X"FFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9",
INIT_24 => X"0001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFF",
INIT_25 => X"FFFFEBA5D2E97410080400000000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFF",
INIT_28 => X"FFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA",
INIT_29 => X"100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFF",
INIT_2A => X"FFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_2B => X"01FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008040",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804000000000000000000000000000",
INIT_2E => X"2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFF",
INIT_2F => X"FFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_30 => X"0804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFF",
INIT_31 => X"FFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E97410",
INIT_32 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFF",
INIT_33 => X"EBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001",
INIT_34 => X"00000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(29),        -- Port A data input
DOA(0)   => data_read_a_hi_256(29),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(29),        -- Port B data input
DOB(0)   => data_read_b_hi_256(29),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_30_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"9EEBFEF5D7D7F7DF7DFFDFDFCEFFBFFEFF9FE1F7FFBFEFC9B77B7FFFFDFFD000",
INIT_1B => X"7F3F9FCFE7F3F9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7",
INIT_1C => X"E7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE",
INIT_1D => X"80400000000000000000000000000000000000000000000000001007FE00000F",
INIT_1E => X"FFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"BA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001F",
INIT_21 => X"FFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFE",
INIT_22 => X"74100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFF",
INIT_23 => X"FFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9",
INIT_24 => X"0001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFF",
INIT_25 => X"FFFFEBA5D2E97410080400000000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFF",
INIT_28 => X"FFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA",
INIT_29 => X"100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFF",
INIT_2A => X"FFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_2B => X"01FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008040",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804000000000000000000000000000",
INIT_2E => X"2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFF",
INIT_2F => X"FFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_30 => X"0804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFF",
INIT_31 => X"FFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E97410",
INIT_32 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFF",
INIT_33 => X"EBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001",
INIT_34 => X"00000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(30),        -- Port A data input
DOA(0)   => data_read_a_hi_256(30),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(30),        -- Port B data input
DOB(0)   => data_read_b_hi_256(30),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_31_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"129000008004A00804A40000400800020000000C005FEA005800200400050100",
INIT_01 => X"A15FF18019700810180065FFFC0040801E80258CA2951C2200EC0906A0804140",
INIT_02 => X"0000000000000011000550FDFF0FFFFF0007F1FC200000011000000000205FC0",
INIT_03 => X"08425818000000908428C0024210A30004045060302223490002014280410FF8",
INIT_04 => X"DB6A618248140C18E0B016872400000007EBA24058E1ECA8E2D400681FD0E061",
INIT_05 => X"1C0FFC338FF01009048084C400103E28FE3F6FE513703F7000E8E5B4825030F6",
INIT_06 => X"4420006040410180034000A157FC1F08040C080045F1F2572060FE82671C607E",
INIT_07 => X"001100004081001103107000185FF0000C0849673F6C06FC000830007FF00000",
INIT_08 => X"F47FC80008000200800000020811000004008812240800000800000000000000",
INIT_09 => X"04FC700090038F3CF82C44630C5D1FC002CCE08082481BF27A00000000000883",
INIT_0A => X"00000000687C0044040424B39FB6073C0010048A4000008F83F009F7DE037DD0",
INIT_0B => X"0620E08812982050800A910249298624124080886FE187FC301B124F20016000",
INIT_0C => X"182001820018200182001820018200183000C1000C10808EE661891139802431",
INIT_0D => X"816800100400902A0200110810080BFF0C8010010220330C3A28070070018200",
INIT_0E => X"C4043FFD03FF101D400080013040180810040802040102004183012084808006",
INIT_0F => X"7C04000008080781000004001D00000781000004001D0000200F018586106100",
INIT_10 => X"0001DC0000000781000004001D00000781000004001D000002F4008000002000",
INIT_11 => X"0080000800007B00000040801BA020000000400077000000010035C040000020",
INIT_12 => X"200000070800000C231410085108D500000000004000F01900030000040202F4",
INIT_13 => X"001D0100000039000003F00040000003F000000050100E808000001C800003A0",
INIT_14 => X"077020000000007C0400005010115602000000001EC00000007404000000E100",
INIT_15 => X"2000CA40EA000000000100F0D000020000501011740080000001F10000014040",
INIT_16 => X"010044602002061004A820104809402BE1FFC006304E03684100050190040350",
INIT_17 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_18 => X"0040100401004010040100401004010040100401004010040100401004010040",
INIT_19 => X"00802FFFFFFFFFFFFFFFFF810040100401004010040100401004010040100401",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000010",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"80400000000000000000000000000000000000000000000000001007FE000000",
INIT_1E => X"FFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"BA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001F",
INIT_21 => X"FFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFE",
INIT_22 => X"74100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFF",
INIT_23 => X"FFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9",
INIT_24 => X"0001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFF",
INIT_25 => X"FFFFEBA5D2E97410080400000000000000000000000000000000000000000000",
INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFF",
INIT_28 => X"FFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA",
INIT_29 => X"100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFF",
INIT_2A => X"FFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974",
INIT_2B => X"01FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFF",
INIT_2C => X"000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E9741008040",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804000000000000000000000000000",
INIT_2E => X"2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFF",
INIT_2F => X"FFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D",
INIT_30 => X"0804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFF",
INIT_31 => X"FFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E97410",
INIT_32 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001FFFFFFFFFFFFFFFFFFF",
INIT_33 => X"EBA5D2E974100804001FFFFFFFFFFFFFFFFFFFFFFFFFFEBA5D2E974100804001",
INIT_34 => X"00000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(31),        -- Port A data input
DOA(0)   => data_read_a_hi_256(31),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(31),        -- Port B data input
DOB(0)   => data_read_b_hi_256(31),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


end;