library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_misc.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library UNISIM;
use UNISIM.vcomponents.all;

entity ram_master is
	port(clk             : in  std_logic;
        address_a       : in  std_logic_vector(31 downto 2);
        enable_a        : in  std_logic;
        wbe_a           : in  std_logic_vector(3 downto 0);
        data_write_a    : in  std_logic_vector(31 downto 0);
        data_read_a     : out std_logic_vector(31 downto 0);

        address_b       : in  std_logic_vector(31 downto 2);
        enable_b        : in  std_logic;
        wbe_b           : in  std_logic_vector(3 downto 0);
        data_write_b    : in  std_logic_vector(31 downto 0);
        data_read_b     : out std_logic_vector(31 downto 0));
end; --entity ram     

architecture ram_master of ram_master is
signal enable_a_lo       : std_logic;
signal wbe_a_lo          : std_logic_vector(3 downto 0);
signal data_write_a_lo   : std_logic_vector(31 downto 0);
signal data_read_a_lo    : std_logic_vector(31 downto 0);
signal enable_b_lo       : std_logic;
signal wbe_b_lo          : std_logic_vector(3 downto 0);
signal data_read_b_lo    : std_logic_vector(31 downto 0);
signal enable_a_hi       : std_logic;
signal wbe_a_hi          : std_logic_vector(3 downto 0);
signal data_read_a_hi   : std_logic_vector(31 downto 0);
signal enable_b_hi       : std_logic;
signal wbe_b_hi          : std_logic_vector(3 downto 0);
signal data_read_b_hi    : std_logic_vector(31 downto 0);
signal address_a_reg     : std_logic_vector(31 downto 2);
signal address_b_reg     : std_logic_vector(31 downto 2);
signal enable_a_lo_256       : std_logic;
signal wbe_a_lo_256          : std_logic_vector(3 downto 0);
signal data_write_a_lo_256   : std_logic_vector(31 downto 0);
signal data_read_a_lo_256    : std_logic_vector(31 downto 0);
signal enable_b_lo_256       : std_logic;
signal wbe_b_lo_256          : std_logic_vector(3 downto 0);
signal data_read_b_lo_256    : std_logic_vector(31 downto 0);
signal enable_a_hi_256       : std_logic;
signal wbe_a_hi_256          : std_logic_vector(3 downto 0);
signal data_read_a_hi_256   : std_logic_vector(31 downto 0);
signal enable_b_hi_256       : std_logic;
signal wbe_b_hi_256          : std_logic_vector(3 downto 0);
signal data_read_b_hi_256    : std_logic_vector(31 downto 0);
begin
process(clk)
begin
if rising_edge(clk) then
	address_a_reg <= address_a;
	address_b_reg <= address_b;
	end if;
end process;
data_read_a <= data_read_a_lo when (address_a_reg < x"0001000"&"00") else
data_read_a_hi when ((address_a_reg >= x"0001000"&"00") and (address_a_reg < x"0002000"&"00")) else 
data_read_a_lo_256 when ((address_a_reg >= x"0002000"&"00") and (address_a_reg < x"0003000"&"00")) else 
data_read_a_hi_256 when ((address_a_reg >= x"0003000"&"00") and (address_a_reg < x"0004000"&"00"));
data_read_b <= data_read_b_lo when (address_b_reg < x"0001000"&"00") else
data_read_b_hi when ((address_b_reg >= x"0001000"&"00") and (address_b_reg < x"0002000"&"00")) else
data_read_b_lo_256 when ((address_b_reg >= x"0002000"&"00") and (address_a_reg < x"0003000"&"00")) else 
data_read_b_hi_256 when ((address_b_reg >= x"0003000"&"00") and (address_b_reg< x"0004000"&"00"));
enable_a_lo <= enable_a when (address_a < x"0001000"&"00") else '0';
enable_b_lo <= enable_b when (address_b < x"0001000"&"00") else '0';
enable_a_hi <= enable_a when ((address_a >= x"0001000"&"00") and (address_a < x"0002000"&"00")) else '0';
enable_b_hi <= enable_b when ((address_b >= x"0001000"&"00") and (address_b < x"0002000"&"00")) else '0';
enable_a_lo_256 <= enable_a when ((address_a >= x"0002000"&"00") and (address_a < x"0003000"&"00")) else '0';
enable_b_lo_256 <= enable_b when ((address_b >= x"0002000"&"00") and (address_b < x"0003000"&"00")) else '0';
enable_a_hi_256 <= enable_a when ((address_a >= x"0003000"&"00") and (address_a < x"0004000"&"00")) else '0';
enable_b_hi_256 <= enable_b when ((address_b >= x"0003000"&"00") and (address_b < x"0004000"&"00")) else '0';
wbe_a_lo <= wbe_a when  enable_a_lo='1' else x"0";
wbe_a_hi <= wbe_a when  enable_a_hi='1' else x"0";
wbe_b_lo <= wbe_b when  enable_b_lo='1' else x"0";
wbe_b_hi <= wbe_b when  enable_b_hi='1' else x"0";
wbe_a_lo_256 <= wbe_a when  enable_a_lo_256='1' else x"0";
wbe_a_hi_256 <= wbe_a when  enable_a_hi_256='1' else x"0";
wbe_b_lo_256 <= wbe_b when  enable_b_lo_256='1' else x"0";
wbe_b_hi_256 <= wbe_b when  enable_b_hi_256='1' else x"0";



ram_bit_0_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"ED39BA795990D275FB4A6E96ACC4731DEA4598B0AFB54867F6EE4618C3749803",
INIT_01 => X"58A0047D8607944AC7DA180001ECA2544042106208408208C20022E9173734B3",
INIT_02 => X"9F775E7CB273E6CCA7DAAF00001000000478020113C9C38E09FB7CCCDD9F203E",
INIT_03 => X"441406267B4CB04443163C91110C58F24A31000B8028A810A3D0F8B169A01006",
INIT_04 => X"0005802424830120024121209088809DF81454ACA01E03501D0A3B91E00F0A00",
INIT_05 => X"E0F001CC00012034C20B0232838F80D001C0100AEC83C008EF101A034C8CC300",
INIT_06 => X"582541A028D584E40CB0583CCA0100000161F84322000DA8C40F003C80030780",
INIT_07 => X"2BF70E1C3BBBB1138AF7F888025340C0888430047040FEE182CA00044BC5827C",
INIT_08 => X"0CAFC1F1F07F0FE1C94F65B11555EAFFC1C306758B24197ABCDA467F2C9CF9B3",
INIT_09 => X"027BDA3B0000011420A61080800B6E4C464258094101606E5A47A2A2098B0200",
INIT_0A => X"40198000D1281220444210123820B43B40804CE9AFC800017D82082E2081B6C0",
INIT_0B => X"CA2E0B32B01A752B078412A24844B01302A26900C4801854069B0C888890A081",
INIT_0C => X"C0F33C0F73C0F33C0F73C0F33C0E39E0319E0710A9402011C22908B56A21A020",
INIT_0D => X"8429A95E954868AD0E52273F542580000808061C0389161F027039C1F33C0F73",
INIT_0E => X"5C94001120055704FC4A1624485E2489024481224091282C4300942A19439481",
INIT_0F => X"1C55D65C3E3F01F52FFC1E0013C1F801F52FFC1E0013C1F8090423D38A18E3B1",
INIT_10 => X"1C0118796BE001F567FC1E0013C1F801F567FC1E0013C1F9085DFBF7E15C0610",
INIT_11 => X"FBF7E30F00C0270F3751F1FD00FECBF7E25C0700463E17B2C7F811FD7ADECC38",
INIT_12 => X"6474190626D6491063597F9177B956EF378D33E4030061341F077C571F8F885D",
INIT_13 => X"E207F328E3082636B2807FFD80FE00007E03F7207D3E03F9167184131B5C40FE",
INIT_14 => X"047EFA0CAE06101C53E3647D3F144FCDD22B81C0098E57D9081FCE8C8520C4DA",
INIT_15 => X"FF31ADF08DBF81846A540049707E0FE3307D3F141FFB45478040570EED41F4FE",
INIT_16 => X"902C189601208A1502B4AA5584B4068000019A80098120BCA4C617635C938574",
INIT_17 => X"0240902409024090240902409024090240902409024090240902409024090240",
INIT_18 => X"2409024090240902409024090240902409024090240902409024090240902409",
INIT_19 => X"424A800000000000000000902409024090240902409024090240902409024090",
INIT_1A => X"08208208208831042720EE38E38AAF9C4C704DAB63A6D58B3C10BAE8E789AA09",
INIT_1B => X"0F87C3E1F0F87C3E1F0F82082082082082082082082082082082082082082082",
INIT_1C => X"F800003E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F",
INIT_1D => X"55557BD75EF5D00000000000000000000000000000000000000000000018401F",
INIT_1E => X"FEFA28428B455D0017410A28428AAAA2FBD54BAF7FFD55EF007FD75EFFFAE975",
INIT_1F => X"0145F7AEBFFFF08002AA10A2AABFEAAA2FFC0000AA843FE00AAFBE8B45AA803D",
INIT_20 => X"974AA5D7BFFE000804000BAAAAAAAB45557FFFEBAA2D5401450051401555D7FC",
INIT_21 => X"FD7410557FC21555D51574AAA2FFE8B455D7BD755555517FFEFA280021FF082E",
INIT_22 => X"AEBFE00A2803FEBA002A820AA0800174BA5D2EA8B45005168A10AA8028A10087",
INIT_23 => X"7FFE8B45FFFBC00005D003FF45557FC01FFFFAE95410AA80000005D003FEAAFF",
INIT_24 => X"00000000000557DF5500003DFEFFF84175EFA2AEA8A10000417410A2FFE8BEFF",
INIT_25 => X"F0075D75EFEBAE9554540754717F1F8000000000000000000000000000000000",
INIT_26 => X"47E00A2DB45AA8A3AFD7B68E2AB78550E12555F524AFE38B780154BAFFF1D54A",
INIT_27 => X"1D500002A150038038E285D7F78FD7000B6AB50B6AABDE12BEA0AF010B7D1F8F",
INIT_28 => X"D5C7AA854008700249243A412EBFF5542A43FE9257F1E816D557095EAAA2D140",
INIT_29 => X"EDBC0B680900AAF52B474385D75C502D157545A87AAD178A8002D1D21C5E8257",
INIT_2A => X"F6A150012A2F02AFFDF40E85F475451D502D152A82000E3A5D2150AB8F401471",
INIT_2B => X"51EAFEDB52E3F1EFFFF485A2DA3D5D24BD417FD7E9541242FE920AD082E10A28",
INIT_2C => X"00000000000000000000000000005AAF555080550E87B7A405B52AAD152BD001",
INIT_2D => X"FA69574BAF7D5555AF0D79D55FFA2AC97445057F405458500000000000000000",
INIT_2E => X"0FF16565B2FA9075F4F7B3EBDF50FEAEAAB55F7AEAABFF5D2A81151FB8635A02",
INIT_2F => X"4D5D51F5E08A394003A908B8410E707EF34A08D46F6ABE7082AAAAF2FAC77FE0",
INIT_30 => X"FAE8C798A11A0EAEF75F7AA84001A7052C95256803CE3AEB038662E5D8140601",
INIT_31 => X"A05051023F9A9D57B63BFBF906CB45FABC0954AF0151555AF58794040077D774",
INIT_32 => X"FEE5555BE48AB2A2AE0A0F20C43EAC562245B4E1870108B11020AD4AA05542A0",
INIT_33 => X"D407A97F6F35F498B96BEB12DAAB77558ABD5F5F0DA6BC9525688C1A2A0C06E9",
INIT_34 => X"8000000FF8000000FF8000000FF8000000FF8000000FF80F55E25C00A0BA7FBE",
INIT_35 => X"F8000000FF8000000FF8000000FF8000000FF8000000FF8000000FF8000000FF",
INIT_36 => X"000000000000000000000000000000000000000000000000000000000000000F",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000008000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(0),        -- Port A data input
DOA(0)   => data_read_a_lo(0),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(0),        -- Port B data input
DOB(0)   => data_read_b_lo(0),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_1_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"212C001411984004084D000508C53810A03D1450E839B003342114428A000807",
INIT_01 => X"08000010400A0008010600000084004000400002000000000000000000140000",
INIT_02 => X"484DEBA0111800C004400D000000000028800001CC404E6008B4933336880010",
INIT_03 => X"650C00000848A0423183089008C604224200000100A200002C280810098C0001",
INIT_04 => X"00000004208B00200E010800006667BE7000102C00080000040012010000080C",
INIT_05 => X"0080000000002020600100208D04414000800000000200004800080000800200",
INIT_06 => X"0820196100006044401008100208000008082010000000800488000000020400",
INIT_07 => X"1210C18306788C00894098000011000820001000104050004108000001008250",
INIT_08 => X"00A48903121780004C6000311555521F183060AC564BF818B5EDFDE004460030",
INIT_09 => X"02AD881200100140A0223480000458400000480840002002184581A020000200",
INIT_0A => X"140040001020020410000010082080010400002001041001B102002E20013600",
INIT_0B => X"0895400004201001010884000000901100800800000004140002008280A8A815",
INIT_0C => X"C8D00C8D00C8D40C8D40C8D00C8D20642A06468400000030480808020F08E008",
INIT_0D => X"20BC417C16004C0B83822109040180000801000910000003203220C8C40C8D40",
INIT_0E => X"5C96000000010200200802100022008100408020401020040100142200E0E08A",
INIT_0F => X"0000021E300B000000781E00140018000000781E00140018000002430E30E061",
INIT_10 => X"1C00000024E0000000781E00140018000000781E0014001908400005E11C0610",
INIT_11 => X"0003C30F00C000000155800D00000003E21C0700000000F00118000000468C38",
INIT_12 => X"60640900004A400081401A0000004041218503E4030060000004804318008840",
INIT_13 => X"A0001208C30800025200003D807E000000000725201600090461840001340002",
INIT_14 => X"0000F00C0E06100000012D2005100409520381C00000005920004C0C81200009",
INIT_15 => X"25000120850B8180625400400000010711200510004B41478040000005548016",
INIT_16 => X"10040002002080040000804000A0000000011A000100208C008611430A000040",
INIT_17 => X"0040100401004010040100401004010040100401004010040100401004010040",
INIT_18 => X"0401004010040100401004010040100401004010040100401004010040100401",
INIT_19 => X"5000800000000000000000100401004010040100401004010040100401004010",
INIT_1A => X"8A28A28A2AC8090C69606492492C09945235D5F7E2A5040B80E1C863A2958000",
INIT_1B => X"5BADD6EB75BADD6EB75BAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA28A2",
INIT_1C => X"FC00002E974BA5D2E974BA5D2E974BA5D2E974BA5D2E974BA5D2E974BA5D2E97",
INIT_1D => X"BA55556AAAAAA800000000000000000000000000000000000000000000607FFF",
INIT_1E => X"F45A2FBD75EFA2AE97555F7FBFFF45FFAE80010AAAABFFFFFF803FE10F7D17FE",
INIT_1F => X"8AAAF7FBD54AA002A955555D7FE8ABA082EBFEBAFFD555400557BD54BA5D7FFD",
INIT_20 => X"17555AA8028BEFAAAE97555082A80000AA802ABEFA2D568A005D5157400AA802",
INIT_21 => X"EBDFEF5D7FEAA00AAAABFEAA007BC0145FFFFFDF55AAFBC00105555400105504",
INIT_22 => X"D5575555D7FC2155F7AEA8BEFAAAA954BA557BD7410550428ABA5D5168ABA552",
INIT_23 => X"FD57DF45F7D568ABAF7AABFFFF082ABFFFFFFFFEAB55557FFFEBAAAD568B45A2",
INIT_24 => X"000000000002EBFFEFA280021FF082E974AA5D7BD74000804154BA082ABFF55F",
INIT_25 => X"7F78A3FE28E3D17DEAA485FE8E02B50000000000000000000000000000000000",
INIT_26 => X"6D5D75D54BA5D7BFFF7DA2FFD55EFAAA495545E175EFF57BF8FC2000BEA4BAE9",
INIT_27 => X"A28550E10405F7A4AFE38EAA0924921C2FD55455571E8A2A087BF8EAAEB8E001",
INIT_28 => X"7A28415A001684104155C5B6DF6DBEFBFAA07157428145A00AA8A2FBD7B6DF6A",
INIT_29 => X"AAABF1FFBC7010FF8A38FEF557FEAB78B6AAB8E971471C7010B7D168F47400A0",
INIT_2A => X"495EAAA2D16D1FDBED56A55557A43DE385FD4BFBD7B6A0BF492415FC20105D24",
INIT_2B => X"F5D717FE2AAAA56DEBD17FE3DF7FB7FEBFE38017EBA4A8EB8F6FFD5FE8B7D557",
INIT_2C => X"00000000000000000000000000002A3D5C7AA854008700249243A417FFF41542",
INIT_2D => X"AF2A00010F78028B15F7823FEAAA2D57DFBA007DFCA127B80000000000000000",
INIT_2E => X"A0869AAAB8A7C19C55550E8574BA557BFFFEFAAFBD55FFAA8416545A6FB60F47",
INIT_2F => X"10A2AEBFF55F7BAAA8565DBAC1112FFAC21A022A38C20B2552E975F758516AAA",
INIT_30 => X"01E7AD1FFF5575841DE08007FC2048002895755FFEFBCEE5FBAACB10085EE5DE",
INIT_31 => X"D4000D7FC00FC5D062BBA05ED5034472A02EABEA097BEAAFAF2863FA00DD5742",
INIT_32 => X"62B0A2F7AE8B5D5D51F5E18ABD5EAFFF2AF9554FF57EFBFA18D4FBFFF40FF809",
INIT_33 => X"C95256807DC31AA8114DE55F5BED201FFFED17DFBFF6963FCAAA2283CF140500",
INIT_34 => X"0000000000000000000000000000000000000000000002CB75F7AA84001A7052",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000008000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(1),        -- Port A data input
DOA(0)   => data_read_a_lo(1),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(1),        -- Port B data input
DOB(0)   => data_read_b_lo(1),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_2_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10E44660018259B2843913100062C98004802322D3E030235201006009B2816",
INIT_01 => X"8005A188084900481C8024A542400340404000720885800802000906E4910204",
INIT_02 => X"5C010802020408040C640850AA055254090541A111240A104A0000000908B510",
INIT_03 => X"0C1101108800004481060A001204102803156020218808002440850008C80550",
INIT_04 => X"8840C08122050400582812C21C0804040968987810688899444090C10A124A69",
INIT_05 => X"4885109105400129210040010340086856B141212252142242A068A080106372",
INIT_06 => X"047450004062400090000202000054C28012204400908281302852A6710AA420",
INIT_07 => X"121810000230089008408402A800011012D41D518044411005000AA8A5004390",
INIT_08 => X"A214110514163218085008010141421F02000124000010880000442080810201",
INIT_09 => X"0A09E89041451581B53A739C42A0C9223000004881708D80100331CA8A848E0A",
INIT_0A => X"1009020A30020008096A06B8C1208A000A9C20004820B0573165541CD5482216",
INIT_0B => X"ACC084404A8000490152D100344001108AA88B1D007291402802B1041632A011",
INIT_0C => X"8696086860869608686086920868004309043414A2191C24485C4D2A9A0DF823",
INIT_0D => X"484000804201C1102080215900038AD030014588D200F0221821808682086820",
INIT_0E => X"00002AA00AA80240A001010026824040C000201030000200C8980080260C201E",
INIT_0F => X"0000000A20001602900020001400002A029000200014000100280E6694490312",
INIT_10 => X"0000000024002A02900020001400001602900020001400002700000800010000",
INIT_11 => X"0008004000000000001500006C00300800020000000000C100014A0081200100",
INIT_12 => X"8088000000480005188000440840081000500002000000000004800010003420",
INIT_13 => X"0070041200000002411280004000000000000026000038020900000001201300",
INIT_14 => X"2A0004030000000000002A00004A100208800000000000012260101100000009",
INIT_15 => X"0084420300001040100000000000010402000049800020000000000000580001",
INIT_16 => X"040111000008001505448340606B21090556002E00000000000080002A040A00",
INIT_17 => X"401004010040300C0300C0300C0100401004010040300C0300C0300C01004010",
INIT_18 => X"0200400004000040000C0200C0200C0200400004000040300C0300C0300C0100",
INIT_19 => X"14A97C0FC0FC1F81F81F800C0200C0200C0200400004000040000C0200C0200C",
INIT_1A => X"0410410411823A4301040B2CB2CBACB002009C6B860185AA1491B0E2863EA015",
INIT_1B => X"8944A25128944A25128941041041041041041041041041041041041041041041",
INIT_1C => X"FC703F25128944A25128944A25128944A25128944A25128944A25128944A2512",
INIT_1D => X"AA0004001550000000000000000000000000000000000000000000000078401F",
INIT_1E => X"5FF5D003FE10F7D17FEBAF7D5420AA0855420AAAA843DFFFAAD1554005D7FD74",
INIT_1F => X"FF45AAFBC20AAF7D1575EF55517DF555D2EBFF45AAAAA8A10A2AE80010A2AA97",
INIT_20 => X"AABEFAAD1575EFAAAE974AA5D51554BA5D7FFFF45A2AA975EFA2FFD7555FFFBF",
INIT_21 => X"5554AA555555555557FE8ABA082EBFFFFAAAE95555552E974105D517DF55AAAA",
INIT_22 => X"D540000AA802AABAF7FFC2010AAAE821EF552E82010F7AABFE10FFD542145FFD",
INIT_23 => X"02E800AA08042AB45007FC00BAFFD168BEFF7FBC0010AA802ABEFAAD540000FF",
INIT_24 => X"000000000002E80010555540010550417555AA8028BEFAAAE821550851420AA0",
INIT_25 => X"7A2DF55400557FD54AA1D04001C5150000000000000000000000000000000000",
INIT_26 => X"D5F7A482000BEAE905C755003FE28E3D17DEAAE95F40002157F470AABE803AE9",
INIT_27 => X"5EFAAA495545E3F5EFF57F7FE80082FFDE105EF55517DFC5552ABDF45B6AEAFF",
INIT_28 => X"24105D5B7FF7DB6AAAABC7BEDB505EFBEA4070BA5FD0154BA5D7BFAF7DA2AE95",
INIT_29 => X"38E00B6DF68FEF4871D24BA495B5556D5571E8AAF082AB8EAAEB8E0016D5D2A9",
INIT_2A => X"E2FBD7B6DF47A00EBDB50000A380AAE28E80495038AAAEAF1D7410E80000FF84",
INIT_2B => X"FBC703AE2DF42AAA002A851C214003FF680071ED1EFEAF1EFFFDEAD1C5010AA8",
INIT_2C => X"00000000000000000000000000002087A28415A001684104155C5B68E2DBEFBF",
INIT_2D => X"51FBD74BAF7802AB05AAFBD5400557BD54AA5500021555100000000000000000",
INIT_2E => X"55D2ABDF55F782BEB47AFAD00010F7AA8215555003FEAAAAD57DEBAA2FDDC010",
INIT_2F => X"BA557BEABEFAAEBD55FFAA1456547A2D360F47AF7FC20B2F7FBC015D58517FF5",
INIT_30 => X"AB4A78016545540400010557BFDFFFF7822A955FFFFC20FFF3AE544108410174",
INIT_31 => X"D545002A800A8FF862BA00F2F9E8F0050D4420BA547FD75FF58516AAAA0828AA",
INIT_32 => X"35B57AB5155400A2AEBFF45FFFB404007FFBD550AAFACAAA122AA8954BAA2AE9",
INIT_33 => X"895755FFAEBCFE57BBA57002DF3C4AAAA002E954505C417FFFF08555555BAAD3",
INIT_34 => X"000000000000000000000000000000000000000000000061DE08007FC2048002",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000010000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(2),        -- Port A data input
DOA(0)   => data_read_a_lo(2),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(2),        -- Port B data input
DOB(0)   => data_read_b_lo(2),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_3_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"210C44A20020248B08431120001604B8156023104C40771B3430400A02380206",
INIT_01 => X"014C9A4250B0296D3C2422C992100B49404040028804A0080A000416A8D90A0C",
INIT_02 => X"4809A900031800444460589C66E331352180D468B8040E600C0081110B802CD0",
INIT_03 => X"6D0B6110880001D23583480648D60520330066810A80881068A808029CC56330",
INIT_04 => X"48221A066A09D03B348C1C1928DD5A4402A13868070940842640902107002D24",
INIT_05 => X"058318035328202004C1C4E50B44644B30A86D01014A0D224063090082100E34",
INIT_06 => X"08381A010040200AC2190ED2002ACD99881822104C5A40942048288234629414",
INIT_07 => X"0218408142740E2C0948C3066400071913209CC8004640100D003999552083D2",
INIT_08 => X"900409231292A8080C2000110001521F0810A92E7402F08AB0016CA000C60011",
INIT_09 => X"620C889014D30E4A210214D5099058808010605A81A41480102130C020A43A39",
INIT_0A => X"512850E61822020C899046740121820004102000402079CCA037A02C68552A35",
INIT_0B => X"8895000026A00141015290040460C0B4828289AC1011954C0026A20400882914",
INIT_0C => X"80CA080DA080DA080CA080CE080DB0402F040654A2442834C0092E228A0DF2AB",
INIT_0D => X"289080600E04C50206808059000999C98840C508D220108200202080DA080CA0",
INIT_0E => X"300E6660599802602209021204A050E1C850C428521C208480821D842085A03E",
INIT_0F => X"0000010000003202900000010000000A02900000010000008038666920920A24",
INIT_10 => X"0000008000002202900000010000001E02900000010000002380000800000000",
INIT_11 => X"0008000000000000008000002D00300800000000000020010001620081200000",
INIT_12 => X"8088000008001021C88000048800281000500000000000004000000000003600",
INIT_13 => X"00B8041200000040011980004000000000000803000068020900000020001B00",
INIT_14 => X"29800403000000000008030000C83002088000000000002002E0101100000100",
INIT_15 => X"00841003100010401000000000002000030000C38000200000000000020C0001",
INIT_16 => X"108722420420A0100006D34A404800185CCE0128410820000008008021C40A00",
INIT_17 => X"0872108721085218852188521885218852188521887210872108721087210872",
INIT_18 => X"8721086214872108621C852188421C852188421C852188721087210872108721",
INIT_19 => X"54A2EAA555AAB554AAB5561C852188421C852188421C85218842148721086214",
INIT_1A => X"0410410412881D0B0000092492480A981E063C638321450A08899A62C314A014",
INIT_1B => X"9D4EA753A9D4EA753A9D49249249249249249249249249249249249249241041",
INIT_1C => X"FAABC4351A8D46A351A8D46A351A8D46A351A8D46A351A8D46A351A8D46A351A",
INIT_1D => X"5500002AA100000000000000000000000000000000000000000000000000401F",
INIT_1E => X"FFFAAD1554005D7FD74AAA284001550055421EFAAFFD54AAF7D168B45AAAABDF",
INIT_1F => X"20AA080400155AAD5554AAF7802AB4500043DF45FFD168AAA0855420AAAA843D",
INIT_20 => X"021550855555FFAA84001FFAAAE80010A2AA955FF5D003FE10F7803FEBAFFD54",
INIT_21 => X"BC20AAA284175EF55517DF555D2EBFE00AA8028B45A2AE82155A2FBFFEBA0800",
INIT_22 => X"7BD7555FFFBFDF55AAFBD55EF5D2EBFE10085168ABAFFFBD54BAAAAE97400A2F",
INIT_23 => X"D0015410F7AAAAAAA55043DE00FFFFD5555AAAA954AA5D7FFFF45AAAA975EF00",
INIT_24 => X"0000000000004174105D517DF55AAAAAABEFAAD1575EFAAAE974AA5D00175555",
INIT_25 => X"2EBD56DB7DBEAEBFF551C042AA101D0000000000000000000000000000000000",
INIT_26 => X"D75D5B470AABE8A3AFD7A2DF55400557FD54AABC04001C51551471D7AAF1D05D",
INIT_27 => X"E28E3D17DEAAEBDF40002550F47155AADB50492EB842FB5508043FF55EBD56AB",
INIT_28 => X"017DAAFFFAE821C0A0717D1C5B575FFB68E82557FD2082000BEAE905C755003F",
INIT_29 => X"D74BAE3AE85480FFFFC00AABE8E105C755517DF40552ABDF45B6AEAFFD5F7A48",
INIT_2A => X"FFAF7DA2AE905EF0075D5545E3F5EFF57F7D5C55D7492E90E3808756DA92EBFF",
INIT_2B => X"F5C7092FF801756D490A10438EBA4B8E9241043AE10EAF5C5547FF80954AA5D7",
INIT_2C => X"00000000000000000000000000000E124105D5B7FF7DB6AAAABC7BEDB505EFBE",
INIT_2D => X"515157555AAD142040A2D57FFFFFFAEBFF555D0028A005100000000000000000",
INIT_2E => X"500003FF55AAFD6AB455157D74BAF7AAA8B45AAFBD54005D7BD54AAF78002155",
INIT_2F => X"10F7AA8215555003FEAAAAC53DEB8A2FDDC01051AE955F7AAFBC0000AF843FF5",
INIT_30 => X"F51F782BCB47ABAE801FFAAFBEAA105D2E955FF557BD74EFFBACD41577B84000",
INIT_31 => X"0AAA00557FEA8A2FDD64BAAF8282012AFFEC20BAF7AA8015558517FF555D2ABD",
INIT_32 => X"48547AE04174BA557BEABEFA2AA951FF88554214FA2D3EAF57AFFDD7555082AA",
INIT_33 => X"22A955FFFFC21FFF3BE40412DE02955FF082A820AAAB842AA00000028AB0AAFF",
INIT_34 => X"0000000000000000000000000000000000000000000002A80010557BFDFFFF78",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000008000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(3),        -- Port A data input
DOA(0)   => data_read_a_lo(3),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(3),        -- Port B data input
DOB(0)   => data_read_b_lo(3),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_4_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10804002061080A284201081034809800A00230340007833522C82D04A16006",
INIT_01 => X"804399801838084C0420450E1E104348403008418984014902030006A0910204",
INIT_02 => X"480108A200000000446418E01E80F00A4104311868240200080000000988A390",
INIT_03 => X"065140108800004080064A0002001128270072E03000000030808D00888100F0",
INIT_04 => X"9100EB836A155C1AF0B81CD60433B944022AB8385AC0D4B8E02010E81C32E821",
INIT_05 => X"5C0F20B36F08000024C084C501441C4CF01C489533483C8042EAC190001074C4",
INIT_06 => X"0034420151620118120106902406C3C7800201448DD9D2871020F2AA375A6071",
INIT_07 => X"12181000023480040840C001E080030032009700024641000C00187A442007C2",
INIT_08 => X"8084830110160218004000001101121F220000260000108AA000440880000000",
INIT_09 => X"5A8C881063DF3E839008F29F407448F200B020DA841CA2001001008882046647",
INIT_0A => X"C61504C1380101801900439001FD8804041400001002003C230B6715A4786E0F",
INIT_0B => X"ACD1240522E000098100D104B26041348A088078116C105DA006D10416BE3002",
INIT_0C => X"8608086180860808608086180860A0434C0430D4A25F3182CC4D5D221A09E821",
INIT_0D => X"0BC28081080549504400A8080009B878184044881222D1821821A08628086180",
INIT_0E => X"20481E0E18790012820001100200D02048300418022C1282809A09040415002A",
INIT_0F => X"0000010020005E0090000001000000C6009000000100000000380E6C30830806",
INIT_10 => X"000000800000D20090000001000000EE0090000001000000A6A2000000000000",
INIT_11 => X"0000000000000000008100003B00200800000000000020010002EA0080200000",
INIT_12 => X"80800000080000211D80000C0044281000400000000000004000000010003282",
INIT_13 => X"03B00410000000400121800000000000000008020000B8020800000020006F00",
INIT_14 => X"59000402000000000008020000C9000200800000000000200FC0101000000100",
INIT_15 => X"008A500100001040000000000000200002000042E00000000000000002080001",
INIT_16 => X"08820440040802500104C34820E3031B63C20530C01800410009009821040A00",
INIT_17 => X"C832008020C812008220C81200802048320880204832008020C8320082204812",
INIT_18 => X"8120481208822008020C812048320880208802048320C8120882204812088020",
INIT_19 => X"10A3A5930C9A6CB261934E048320C81200822008220C81204832008020882204",
INIT_1A => X"8A28A28A2BD30264686668A28A2605145031C03F028000A1C2ED7831A2822250",
INIT_1B => X"51A8D46A351A8D46A351AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA28A2",
INIT_1C => X"F94304068341A0D068341A0D068341A0D068341A0D068341A0D068341A0D0683",
INIT_1D => X"BAAA84154005500000000000000000000000000000000000000000000000401F",
INIT_1E => X"4AAF7D168B45AAAABDF55A2802AA1000002ABFF087FFDF5508003FEBA087FD54",
INIT_1F => X"015500002AABA082E954005500021FF5D2EBFF5500003DF455555421EFAAFFD5",
INIT_20 => X"174BAA2AABDE0055517FF555555420AAAA843DFFFAAD1554005D7FD74AAAA840",
INIT_21 => X"400155AAD1554AAF7802AB4500043DF45FFD168BEF080028BFF0855555455500",
INIT_22 => X"803FEBAFFD5420BA085168A00007BFDE10085168ABA0055574BA5555554BA5D0",
INIT_23 => X"02A97545F7D1555EF55043DF5555517DEAA5D0400010A2AA955FF55003FE10F7",
INIT_24 => X"000000000002A82155A2FBFFEBA0800021550855555FFAA84001FFAAFBEAB450",
INIT_25 => X"5080A3AEAA007BD2482BE84124285C0000000000000000000000000000000000",
INIT_26 => X"381451471D7AAFBD0492EBD56DB7DBEAEBFF55BC042AA101D0A28BC7007FFDF4",
INIT_27 => X"400557FD54AABE84001C5550A28ABA1424974004100021FF492AB8F7D1C0438E",
INIT_28 => X"8BEF005557545490012482B6A0BAE2849557AFED1C5F470AABE8A3AFD7A2DF55",
INIT_29 => X"504924955524AA140E0717DAADB50492EB842FB5508043FF55EBD56ABD75D042",
INIT_2A => X"A905C755003FE28E3803DEAAEBDF40002557F6DA101475FDE10145F68A921C55",
INIT_2B => X"DF425575D7BEFB55002097555FFD5401EF5D043AF6D405F78E3A1C2002000BEA",
INIT_2C => X"0000000000000000000000000000208017DAAFFFAE821C0A0717D1C5B575FFB6",
INIT_2D => X"512EAAB45007FFFF55082EA8AAA087FC2010F784000AA5900000000000000000",
INIT_2E => X"F002EA8BEF5D0428ABA595557555AAFBC2000A2D57FFFFF7AEBFF55FF8028A00",
INIT_2F => X"BAF7AAA8B45AAFBD54005D7BD54AAF78002155512AAAA085D04174100800021F",
INIT_30 => X"F55AAFD6AB4551002ABEF005555555000402000FF802ABAA04552ABFF597FD74",
INIT_31 => X"DE005D7BE8AA85555400100879560AA592F955FFAAFBC0000AF843FF5500003F",
INIT_32 => X"FCABA598400010F7AA8215555003FEAAAA843DEB0A2FD5600051537DE005D557",
INIT_33 => X"E955FF557BD75EFFBBCD415521FBFDF45000417545FFD5421FF5D0428BEF0079",
INIT_34 => X"00000000000000000000000000000000000000000000004001FFAAFBEAA105D2",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000010000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(4),        -- Port A data input
DOA(0)   => data_read_a_lo(4),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(4),        -- Port B data input
DOB(0)   => data_read_b_lo(4),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_5_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50DB4A0791B1B4B694369283C81F9996A091832112004AB37B20E07C0C1E006",
INIT_01 => X"085FBC448000804C446A00000034826841280A00084000C8C212802EE2953235",
INIT_02 => X"C809AD5CB118E640A4D018FC011FF0002080000082C8C66609DB7DDDCB1F2036",
INIT_03 => X"250907263E4C90D210835C82484205720B20640A88800000B8E0F810A8C4500E",
INIT_04 => X"4005102126898100064D20001044429C7824382C0416C087198AB916E0551A24",
INIT_05 => X"A370C14CA0E101094008002389CFE2F20D7D7A114CB5C20AE514178054948912",
INIT_06 => X"547319A1499121D4C0A046FC4E06C030581859058C2404844437118630839B88",
INIT_07 => X"2A53468D1A758C038AFFEA9FE39348C9204C389672407EF120EA5806E6C543AC",
INIT_08 => X"8C05896372728FE0C420619000003AFF48D1222E5D26F06ABCC96CD72C463990",
INIT_09 => X"82DE9AB9182080C801041080300F6F0E42821809C2FEA0B65A212282002B029F",
INIT_0A => X"1688E480D10A90049026145B3830B64944904569E7E00A002C836D35B68D26C0",
INIT_0B => X"88990E14269AB54B078092E6BD4431138A00AEFDD567DA480816848C94180846",
INIT_0C => X"C0591C0791C0491C0791C0591C06A8E0248E03D68860A0106119883D6AE1A0A4",
INIT_0D => X"23D829FA654184533252095E542387F81008071C1BAAD68B027029C0491C0691",
INIT_0E => X"0CA7FE0227FC25847C4395166C5844480204011210A11028C380802A24C89494",
INIT_0F => X"1C55D65E3E3C017C37FC3E0017C1F8017C37FC3E0017C1F90005024108308061",
INIT_10 => X"1C0118796FE0017CA7FC3E0017C1F8017CA7FC3E0017C1F9100DFFF5E15D0610",
INIT_11 => X"FFF3E34F00C0270F3755F1F8007FCBEBE25E0700463E17F2C7E014FF7AE6CD38",
INIT_12 => X"64E4090626DE40100459759173BBD6EF37C523E6030061341F07FC571F8F800D",
INIT_13 => X"E0A6FE28C3082636F201BFFF807E00007E03F7243D38337D1C6184131B7C1DEF",
INIT_14 => X"397FFA0E0E06101C53E36C3D3E884FDDD28381C0098E57D923BDFC8C8120C4DB",
INIT_15 => X"FA36FDF58DBF81C062540049707E0FE7303D3E03BFFF41478040570EED50F4F8",
INIT_16 => X"88212B100901A2349004C26A624A21040FC190050A2110B8ACC40B204A119074",
INIT_17 => X"C20080230802108C2008C22080210882108C220842208821088210842208C200",
INIT_18 => X"20084220842208C2008823080230802108823084220842008821080230842008",
INIT_19 => X"54C1892596D34924B2DA6884220842008C20084220802108821080230802308C",
INIT_1A => X"BEFBEFBEFB7F7FE7EFEEE79E79EFAF2DDA73FBDCEDBFF9D3F0FDE0DB6DBF6218",
INIT_1B => X"DEEF77BBDDEEF77BBDDEEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEF",
INIT_1C => X"FAF3167BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBD",
INIT_1D => X"BA5D2ABFFEFFF80000000000000000000000000000000000000000000000401F",
INIT_1E => X"F5508003FEBA087FD54BA0804154005555574AAA2802AA10FFFFFDE0008556AA",
INIT_1F => X"AA1000003FEBA00002AABA5D2EBFEBAAAD16AABAF7AAA8BFFAA802ABFF087FFD",
INIT_20 => X"E8B45FF80001555D2E955FFFFD5421EFAAFFD54AAF7D168B45AAAABDF55AA802",
INIT_21 => X"02AABA082E954005500021FF5D2EBFF5500003DE005555575EFA2D142145A2FF",
INIT_22 => X"7FD74AAAA840014500517FFEF007BEABFF5D7FC00BA5D5568AAAF7AAAAAAAAA8",
INIT_23 => X"2FBEAA105D2E97410FFD16AAAA5D2ABDEBAFFD5420AAAA843DFFFAAD1554005D",
INIT_24 => X"000000000000028BFF0855555455500174BAA2AABDE0055517FF555504154BAA",
INIT_25 => X"0FFFFFFE38085F6FA92552AB8FEFF78000000000000000000000000000000000",
INIT_26 => X"C7B68A28BC70075FDF45080A3AEAA007BD24821E84124285C51574BAB68A2DA0",
INIT_27 => X"B7DBEAEBFF55BE842AA105D0A38EBA1C0428A925D2AB8EBABEDB6AA92F7AAA8B",
INIT_28 => X"75EFA2DB45145B6F5EFB6DF78E05145552A925FFFFD1471D7AAFBD0492EBD56D",
INIT_29 => X"68AAAF7AAAAA82BE8A28A921424974004100021FF492AB8F7D1C0438E38145B5",
INIT_2A => X"A3AFD7A2DF55400557FD54AABE84001C555517DFC70875EABC7557FC20AA415F",
INIT_2B => X"043AFED1C0E10492B6FFEFA105D2A95410FFDB6FABA542ABAE2AF7DF470AABE8",
INIT_2C => X"00000000000000000000000000000428BEF005557545490012482B6A0BAE2849",
INIT_2D => X"5955554BAFFAEBDE10F7FBFDEBA007BFDE005D2AAABEFFB80000000000000000",
INIT_2E => X"AF7FBE8A00FFAEAAB45F3AAAAB4500557FF55082EA8AAA087FC20105504000AA",
INIT_2F => X"55AAFBC2000A2D57FFFFF7AEBFF55FF8028A00512AA8AAA5D0028A005D2AA8AB",
INIT_30 => X"BEF5D0428ABA597FD55FFA2FFD5555FFD57FFEFFFAA97545552A821EFFBD5575",
INIT_31 => X"8B55557FC0012087FEAABAF7AAAAA10F3AAAAA005D04174100800021FF002EA8",
INIT_32 => X"A8ABAFBFFD74BAF7AAA8B45AAFBD54005D7BD54AAF7800015551517DF4500516",
INIT_33 => X"402000FF802AAAA04452ABFF592E80010FFFFFFE005D2A95410F7FFFFEBA5D2E",
INIT_34 => X"000000000000000000000000000000000000000000000002ABEF005555555000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000060000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(5),        -- Port A data input
DOA(0)   => data_read_a_lo(5),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(5),        -- Port B data input
DOB(0)   => data_read_b_lo(5),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_6_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10804B0061A010A2840012C030028180004003220200403302301C0381A0086",
INIT_01 => X"A70041CA3839684D18A160000C52424841000000090800090210080008110204",
INIT_02 => X"080108200C1000004465480400C0080100000000010432400800800009882050",
INIT_03 => X"040001008C2340D0842208624210802182800584488000103080014E08C10000",
INIT_04 => X"00101611A029B08410044800000000040088122A44281C040400900500001800",
INIT_05 => X"02800000400C820934E4A0002900404402820024000A00824004283011200A00",
INIT_06 => X"2632000004084804134DA7C011A83FC012122100C80812D00308010000829400",
INIT_07 => X"02181020423088002940C2401D0480112000100004404014602447F805326393",
INIT_08 => X"7004812130160008304000000000021F020408244000108A0000440003040000",
INIT_09 => X"020C889010104088A000348037F05840303902E814000010341108802020FF40",
INIT_0A => X"86C8B5DF1C83C9C8900000100220C244840021100017E2FD200000A40001223F",
INIT_0B => X"88D1804122A088018152D144317205502A880C00107FD75DE922005026A62A15",
INIT_0C => X"B6284B6284B6184B6184B6384B62825B0425B0568075A0826849C8229AC5F8AE",
INIT_0D => X"03C440C054048850A300A8480009A0020865A588DA20F1A2D92D82B6084B6084",
INIT_0E => X"031001E0800122100321C89214A01A742D3A168D1B4686D100234B442428C034",
INIT_0F => X"000008AB80030202800000001402068202800000001402067400026000000000",
INIT_10 => X"00000000341E8202100000001402068202100000001402062840000800000000",
INIT_11 => X"0008000000000000083C00052000300000000000000008CD0018400081000000",
INIT_12 => X"800800000069A48584000A0400000010001000000000000000048128C0002840",
INIT_13 => X"1A480012000000034C1E000040000000000400FE000644020100000001A34000",
INIT_14 => X"02800401000000000004BA000112B0020800000000000807E80000110000000D",
INIT_15 => X"0500020250001000100000000000010CCE000198000020000000000010F80006",
INIT_16 => X"62D18468CE8402440404D24A3081B020603E0A20640C8400010298432A002A00",
INIT_17 => X"ED3B4ED0B42D1B4ED3B42D0B42D1B4ED2B42D0B46D3B4ED2B42D1B46D3B4AD2B",
INIT_18 => X"D0B46D3B4AD0B46D1B4AD3B4ED0B42D1B4ED2B4ED1B42D0B4AD3B4ED0B42D0B4",
INIT_19 => X"002331C618E38E38C31C7346D3B4AD2B46D1B42D2B4ED2B42D1B46D2B4AD1B42",
INIT_1A => X"8E38E38E39DB3B676F66EFBEFBEFAFBC5E73FC7F87A7D4ABFE7CFAFBE7BF8040",
INIT_1B => X"CFE7F3F9FCFE7F3F9FCFE38E38E38E38E38E38E38E38E38E38E38E38E38E38E3",
INIT_1C => X"FF75A43F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9F",
INIT_1D => X"BA5D7BEAAAAFF80000000000000000000000000000000000000000000060401F",
INIT_1E => X"A10FFFFFDE0008556AABA5D2ABFFEFFF843DFEFA2FBD54BA5555554BAAAFBC20",
INIT_1F => X"5400550428AAAAA84021FF007BD54BAAAD17DEBA0855421455555574AAA2802A",
INIT_20 => X"17400AAFBE8ABAF7FFD54AAAA802ABFF087FFDF5508003FEBA087FD54BA00041",
INIT_21 => X"03FEBA00002AABA5D2EBFEBAAAD16AABAF7AAA8BFFAAD1554BA002A95555A284",
INIT_22 => X"AABDF55AA802AA100000001EF087FEAA00FFFBD5545080417555A2D17FE10000",
INIT_23 => X"2803DFEF0855401FF082EA8B555D7FC21FFFFD5421EFAAFFD54AAF7D168B45AA",
INIT_24 => X"0000000000055575EFA2D142145A2FFE8B45FF80001555D2E955FFFF843DEAAA",
INIT_25 => X"A415B52492B6F5C20825D7FE8A92FF8000000000000000000000000000000000",
INIT_26 => X"555551574BAB68A2DA00FFFFFFE38085F6FA92552AB8FEFF78E3DFFFAAFFD04A",
INIT_27 => X"EAA007BD24821C04124281C0E2DA82BE8E001EF147BD2482BED57AE921451421",
INIT_28 => X"24AA14209557DA28E15400BEF1EFA92FFFFD24BAB68A28BC70075FDF45080A3A",
INIT_29 => X"17545B6D178E281C0A38EBA1C0428A925D2AB8EBABEDB6AA92F7AAA8BC7B6D55",
INIT_2A => X"BD0492EBD56DB7DBEAEBFF55BE842AA105D0E071FF0071EDA38F7F1D55550004",
INIT_2B => X"2A925FFFF8E3DE82BE8E38FFF0851401C70824A8B555C7FC2147F7D1471D7AAF",
INIT_2C => X"00000000000000000000000000005B575EFA2DB45145B6F5EFB6DF78E0514555",
INIT_2D => X"FBAABDFEFAAFBC00BA007BC0000FFD542000557FE8A00F380000000000000000",
INIT_2E => X"0F7D168A105D55421455155554BAFFAEBDE10F7FBFDEBA007BFDE005D2AAABEF",
INIT_2F => X"4500557FF55082EA8AAA087FC20105504000AA592ABFE00F7AA821FF557FC001",
INIT_30 => X"A00FFAEAAB45F3D5400BA5504155EFAAAE95410F7D57DE00FFFBC00AAFBAAAAB",
INIT_31 => X"FEAAF7D157545080417545F7D56AAAA592AA8AAA5D0028A005D2AA8ABAF7FBE8",
INIT_32 => X"C2145F3D557555AAFBC2000A2D57FFFFF7AEBFF55FF8028A00512E975FF08557",
INIT_33 => X"57FFEFFFAA97545552A821EFFBAABDE00F7AAAABEF005542155000028B555D7F",
INIT_34 => X"0000000000000000000000000000000000000000000007FD55FFA2FFD5555FFD",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000048000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(6),        -- Port A data input
DOA(0)   => data_read_a_lo(6),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(6),        -- Port B data input
DOB(0)   => data_read_b_lo(6),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_7_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10840B0048225802842102C02450418800002300500030B313300C418992002",
INIT_01 => X"A34009C23838684D1C20E0000E11426840000000080000080200090000510200",
INIT_02 => X"4801082048100000446558040080000041000000000622400800000009000010",
INIT_03 => X"040001818CA144D0842248424210812102000400088000003080014688800000",
INIT_04 => X"000010002041800000048000000000040088322944200C850001940400301800",
INIT_05 => X"0200000040004100280040204104004402000025000800065004203030320800",
INIT_06 => X"0430060044084804900806D1112A002012120004440812D40120008200829001",
INIT_07 => X"02181020423408002940C24001A4A010200018920646C10C7035000244004380",
INIT_08 => X"008481213016020C204000000000121F020408264000100AA000440012040000",
INIT_09 => X"820C899410000000A100348020005902B1A0048825008091350100CAA0200280",
INIT_0A => X"50140A0010058188100004590331C9C4A400231200340C012100002400012200",
INIT_0B => X"1811C44D22A1884141600411800008104080890023000009A926801050001C00",
INIT_0C => X"9002C9002C9022C9022C9022C903064809648080204020004009080A0A00E088",
INIT_0D => X"0880144434A0010012280008031980036000014A0046206241A4069002C9002C",
INIT_0E => X"0216000200010000000081102080400040002000002010000004008080048A00",
INIT_0F => X"038A2881210382000000001E003E0582000000001E003E042283424000000000",
INIT_10 => X"60700706901982000000001E003E0582000000001E003E046840000000009864",
INIT_11 => X"00000000330C00F0C8210807200000000000581C01C1C809201C400000000001",
INIT_12 => X"0000C2419121028C00020A2400000000000080082C180603A0E003A090406840",
INIT_13 => X"14E8000004321189085F8000000061E001FC00C00207740000021908C4829D00",
INIT_14 => X"BB800000009864038C14800201BAB000000026130071A80613A0000018483224",
INIT_15 => X"0546520350000600812058100F81C018880201BBA0000008239020F110800806",
INIT_16 => X"24003300080022140444D268624B210040004A08000000044222900320C84008",
INIT_17 => X"4010040100402000000000000003004010040100000000000000100401004010",
INIT_18 => X"0000C01004010000000001004010040000000004010040300400000000000200",
INIT_19 => X"54A2C208200010410400000800000000040100C01000000000100C0100400000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000002A10",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FAF8800000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"55002E820AAAA80000000000000000000000000000000000000000000000401F",
INIT_1E => X"4BA5555554BAAAFBC20BA5D7BEAAAAFFFBC00AAF7D5575455D557DFEF002AAAB",
INIT_1F => X"FFEFFFAAAAAAAF7D57FFEFF7D555555A2AEAAB55007FD74AAAA843DFEFA2FBD5",
INIT_20 => X"FDF550000175555504175450055574AAA2802AA10FFFFFDE0008556AABA5D2AB",
INIT_21 => X"428AAAAA84021FF007BD54BAAAD17DEBA085542145552ABDFEFFFAA801EFFFFB",
INIT_22 => X"7FD54BA000415400557BD74BAFFD140000082A975EF00003DF55555168A00000",
INIT_23 => X"5557FEAAA2843FF55A2AEA8B55AAAABDEAAFF802ABFF087FFDF5508003FEBA08",
INIT_24 => X"0000000000051554BA002A95555A28417400AAFBE8ABAF7FFD54AAAAAEA8ABA5",
INIT_25 => X"5415178FD7082EAAB550820870BAAA8000000000000000000000000000000000",
INIT_26 => X"82AA8E3DFFFAAFFD04AA415B52492B6F5C20825D7FE8A92FFFFC70BAE3D15555",
INIT_27 => X"E38085F6FA92552AB8FEFF7A0ADABAEBD578FFFEBD55557DBEA4AFB550871D74",
INIT_28 => X"DFD7FFA4801D7F7F5FDF55000E17545410E175550051574BAB68A2DA00FFFFFF",
INIT_29 => X"3AF55415F6DA38080E2DA82BE8E001EF147BD2482BED57AE921451421555524B",
INIT_2A => X"5FDF45080A3AEAA007BD24821C04124281C7BD2482E3D1450381C20905EF0800",
INIT_2B => X"FFD24BAB6A4A8A82495F78E92AA843DF45BEAAAFB55ABA0BDE02EB8A28BC7007",
INIT_2C => X"000000000000000000000000000055524AA14209557DA28E15400BEF1EFA92FF",
INIT_2D => X"F3FFD54BAAAD15754508556AB45002AA8B450800174BAA680000000000000000",
INIT_2E => X"FF7803DF45085557410AEAABDFEFAAFBC00BA007BC0000FFD542000557FE8A00",
INIT_2F => X"BAFFAEBDE10F7FBFDEBA007BFDE005D2AAABEFFB803DEAAAAD56ABEFAAD5575E",
INIT_30 => X"A105D554214551003FF45FF8400145FFD57FF55082E97555002E955550C55554",
INIT_31 => X"54AA5500021EF000028B55087BFDEBA042ABFE00F7AA821FF557FC0010F7D168",
INIT_32 => X"3FE10AEAAAAB4500557FF55082EA8AAA087FC20105504000AA597FC2010A2D15",
INIT_33 => X"E95410F7D57DE00FFFBC00AAFB8028A00007FE8A00A2803FF45F7AABDF55AA84",
INIT_34 => X"00000000000000000000000000000000000000000000055400BA5504155EFAAA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000007FFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(7),        -- Port A data input
DOA(0)   => data_read_a_lo(7),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(7),        -- Port B data input
DOB(0)   => data_read_b_lo(7),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_8_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00000648E2840112C00000418000002700500030B3132000400812082",
INIT_01 => X"A14008420008204D042100000212026840000000180800080200090048510204",
INIT_02 => X"080108000090000004655C040080000051000000000402400800000009000010",
INIT_03 => X"00000100803008D0842240024210810002800584488000103080894288800000",
INIT_04 => X"00009610A028B084000440C0040000040088323244280C950400808500321800",
INIT_05 => X"42800080400C8A09306420202804400402800035200A00020204283001114A00",
INIT_06 => X"2230400041404B141345A7C20426FFC01292214444081254002801A200821400",
INIT_07 => X"021810204214080069408200008C1010200018920E06C0000020DFFA453223D3",
INIT_08 => X"0084010110120008024000000000021F02040826400000008000440000240000",
INIT_09 => X"828D8880100040898128768820045142B0B902E815008080A0B13848A2200280",
INIT_0A => X"9148A4801C81C9C8100004590711800414002004402008013000403084090200",
INIT_0B => X"BC95C44522A002410040940084720450220089000100104DE924800030821452",
INIT_0C => X"0000400004000040000400004000220010200114AA4020004009092A0009E0A8",
INIT_0D => X"0BC4028430108150900408590109A00209642500120230200100220020400004",
INIT_0E => X"0010000600002210A320C89000005A142D0A16850B6294D10023420124240114",
INIT_0F => X"00000800008100020003C1FE00020080020003C1FE0002004401426008208041",
INIT_10 => X"E3F00000100080020003C1FE00020080020003C1FE000200080000081EA2F9EC",
INIT_11 => X"00081CB0FF3C000008000201000010001DA1F8FC0000080110080000010132C7",
INIT_12 => X"0B0BE6C00020040580040200000001004832CC19FCF81E000000010000200800",
INIT_13 => X"020000C31CF60001008000007F01FFE00004000200420000618E7B0000804000",
INIT_14 => X"000000F151F9EC0000040200401000200D547E3F00000800080001617AD80004",
INIT_15 => X"0100000822406E1B95A3F83000000008020040100000BAB87FB0000010080102",
INIT_16 => X"66D1A368C68D26000544D26A504AB12040022220640484000110184300002A02",
INIT_17 => X"6D1B46D1B46D1B46D1B46D1B46D0B42D0B42D0B42D0B42D0B42D1B46D1B46D1B",
INIT_18 => X"D1B42D0B42D0B42D0B42D1B46D1B46D1B46D1B42D0B42D0B42D0B42D0B42D0B4",
INIT_19 => X"442200000000000000000346D1B46D1B42D0B42D0B42D0B42D1B46D1B46D1B46",
INIT_1A => X"9E79E79E7B7F11E66C6FAD96D96520145052A1F5E2BD085122ED48F3AEB20840",
INIT_1B => X"C3E1F0F87C3E1F0F87C3E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7",
INIT_1C => X"FA2A6D4F87D3E1F4F87D3E1F4F87D3E1F4F87D3E1F4F87D3E1F4F87D3E1F4F87",
INIT_1D => X"FFFF84000AAFF80000000000000000000000000000000000000000000000401F",
INIT_1E => X"5455D557DFEF002AAAB55002E820AAAA840000000043DF55087BC01EF007FD75",
INIT_1F => X"AAAAFFAA95545552ABFE00087BC00AA082EBFE10A28028AAAAAFBC00AAF7D557",
INIT_20 => X"E8BFFA2FBFFFFFAAD5400AAFF843DFEFA2FBD54BA5555554BAAAFBC20BA5D7BE",
INIT_21 => X"AAAAAAF7D57FFEFF7D555555A2AEAAB55007FD74AAAAD57FF45002A975FF007B",
INIT_22 => X"556AABA5D2ABFFEFFFAA82000555555545AAFBE8A00082A97410F7D5555EFAAA",
INIT_23 => X"87BC2010AAD54014500516ABFFA2AABDF450055574AAA2802AA10FFFFFDE0008",
INIT_24 => X"000000000002ABDFEFFFAA801EFFFFBFDF550000175555504175450000155450",
INIT_25 => X"50075C71FF087BD75D7FF84050BAEB8000000000000000000000000000000000",
INIT_26 => X"BABEFFC70BAE3D155555415178FD7082EAAB550820870BAAA8407000140038F4",
INIT_27 => X"492B6F5C20825D7FE8A92FFA497545552AB8E10007FC50BA002ABFE00AA8A2AA",
INIT_28 => X"DF451C24955EF0875EFBD7B6F1FFFC7BEDB45082EB8E3DFFFAAFFD04AA415B52",
INIT_29 => X"92410EBD5505EFB6A0ADABAEBD578FFFEBD55557DBEA4AFB550871D7482AAD17",
INIT_2A => X"A2DA00FFFFFFE38085F6FA92552AB8FEFF7AA87000415B5057DAAFBE8A100820",
INIT_2B => X"0E17555000E17545007BC0000BED14217D005B6ABC7B6AABFFED0051574BAB68",
INIT_2C => X"000000000000000000000000000024BDFD7FFA4801D7F7F5FDF55000E1754541",
INIT_2D => X"A684174105D042AB550055555FF007BD7555F784174AAA280000000000000000",
INIT_2E => X"A082EBDE10AAAEA8ABAF7FFD54BAAAD15754508556AB45002AA8B450800174BA",
INIT_2F => X"EFAAFBC00BA007BC0000FFD542000557FE8A00F384175555D2EA8A00087BD74B",
INIT_30 => X"F45085557410AED17FF455D04155FF00557DF55FFD57DF55FFFBD5400A2AABDF",
INIT_31 => X"21EFA2FFEAA00000002010A2D5421FFFF803DEAAAAD56ABEFAAD5575EFF7803D",
INIT_32 => X"BDFEF0855554BAFFAEBDE10F7FBFDEBA007BFDE005D2AAABEFFBAE97410087BC",
INIT_33 => X"57FF55082E97555002E955550C2E95555087BC0010FFD1401EF087FE8B55FFAE",
INIT_34 => X"000000000000000000000000000000000000000000000003FF45FF8400145FFD",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000020000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(8),        -- Port A data input
DOA(0)   => data_read_a_lo(8),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(8),        -- Port B data input
DOB(0)   => data_read_b_lo(8),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_9_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00018248A2840112C00002C18000002300500030B3132000400812006",
INIT_01 => X"A1400802000020490000000000000240413C0A61590001D90213C90008510204",
INIT_02 => X"680108200010000054655C040080000041000000010402400800800009082011",
INIT_03 => X"00040100800020D0842240124210810042800504488000103081894288800000",
INIT_04 => X"00001410A00AA084000400C0060000040088323044201C850020820400101880",
INIT_05 => X"0200020040048A09202420000C00410402000025000800020804203000100800",
INIT_06 => X"22320400404048041144A7D2003A002012120004DC08125400A0008300821000",
INIT_07 => X"06181020421C08000940820000800010200018B20206C00000200002441223C1",
INIT_08 => X"0184010110120008004000000000061F02040826400008118000440000040000",
INIT_09 => X"8208888210004009010852882000510230A900A8040080800055086002200280",
INIT_0A => X"1402008004814948100004590111C004040120000020080121024012A4081200",
INIT_0B => X"2C91844522A0004100488000801200D00000880001000415E1248002103C2294",
INIT_0C => X"080040820408004082040800408202040020410402000000400809080508A080",
INIT_0D => X"0B4000803200C150108008490809A00219246101100220202102020820408204",
INIT_0E => X"00160006000120002120499020A04A14650A328519629651900142002404201E",
INIT_0F => X"0000080A20010002100000001402008002100000001402000001426008208041",
INIT_10 => X"0000000034008002800000001402008002800000001402008800000800000000",
INIT_11 => X"0008000000000000081500010000100800000000000008C10008000001200000",
INIT_12 => X"0088000000680005800002000000000000500000000000000004810010000800",
INIT_13 => X"02E8040200000003401F80004000000000040027000274000900000001A05D00",
INIT_14 => X"3B8000030000000000042B00009AB00008800000000008012BA010010000000D",
INIT_15 => X"0106520350000040100000000000010C0300009BA000200000000000105C0002",
INIT_16 => X"6651B328CA8D26540544924272EB91004002022024048400000098030A000A00",
INIT_17 => X"2509425094250942509425094250942509425094250942509425194651946519",
INIT_18 => X"5094250942509425094251946519465194651946519465194651946519465194",
INIT_19 => X"0480800000000000000001465194651946519465194651946509425094250942",
INIT_1A => X"34D34D34D1285B080201C92410480AB9A26667A46F345448020082E1C712A054",
INIT_1B => X"8341A0D068341A0D06834514514514514514514514514514514514514514D34D",
INIT_1C => X"F8B2B60D069349A0D068341A4D268341A4D268341A0D069349A0D069349A0D06",
INIT_1D => X"EFA2FFFFF555D000000000000000000000000000000000000000000000007FFF",
INIT_1E => X"F55087BC01EF007FD75FFFF84000AAFFD57DF45A280154BA5555401EFFFD5421",
INIT_1F => X"20AAAA843DFEF00517DEBA007BFDFEFFFD1575EF00557DF555D040000000043D",
INIT_20 => X"68AAAF7802AA00FFFBD7555087BC00AAF7D5575455D557DFEF002AAAB55002E8",
INIT_21 => X"A95545552ABFE00087BC00AA082EBFE10A28028AAAAAAABDF45F7803FFEF5555",
INIT_22 => X"FBC20BA5D7BEAAAAFFFBC00AA552E95545087BD54BA550417400085155555082",
INIT_23 => X"2FFFDF555D7BE8BFF5D51575EFA280175555D043DFEFA2FBD54BA5555554BAAA",
INIT_24 => X"00000000000557FF45002A975FF007BE8BFFA2FBFFFFFAAD5400AAFF8402000A",
INIT_25 => X"2415B471C7E3DF451EFBEFBFAF45490000000000000000000000000000000000",
INIT_26 => X"45490407000140038F450075C71FF087BD75D7FF84050BAEBDF78F45B6801048",
INIT_27 => X"FD7082EAAB550820870BAAA8438FFF00517DE82007FFAFEFE3DB505EF1C5B7AF",
INIT_28 => X"8F45F78A3DFD741516DAAAE38E2DA28EBFFD55451C7FC70BAE3D155555415178",
INIT_29 => X"1543808515756D1C2497545552AB8E10007FC50BA002ABFE00AA8A2AABABEAEB",
INIT_2A => X"FD04AA415B52492B6F5C20825D7FE8A92FFFFC20BA5D2E905550071D54825D0A",
INIT_2B => X"DB45082EB8002000AAFFFDF6D417FEABEF5D55505FFBE801256D490E3DFFFAAF",
INIT_2C => X"0000000000000000000000000000517DF451C24955EF0875EFBD7B6F1FFFC7BE",
INIT_2D => X"A2FBEAB45F78402010007BD5545AAFFD55EFF7FBE8B550000000000000000000",
INIT_2E => X"FAAFFC01FF557FE8B550004174105D042AB550055555FF007BD7555F784174AA",
INIT_2F => X"BAAAD15754508556AB45002AA8B450800174BAA68028BEF00517FE10007BE8BF",
INIT_30 => X"E10AAAEA8ABAF7AAAAB45F7AEBFF4508557FEAAAAAEBFEAAAAFFD5545557FD54",
INIT_31 => X"0145005557400552A954BA0051575EF5504175555D2EA8A00087BD74BA082EBD",
INIT_32 => X"021FF002ABDFEFAAFBC00BA007BC0000FFD542000557FE8A00F3FFC00BA552E8",
INIT_33 => X"57DF55FFD57DF55FFFBD5400A28400010A2FBFDFFF007FE8BFF5551401EFF784",
INIT_34 => X"000000000000000000000000000000000000000000000517FF455D04155FF005",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000040000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(9),        -- Port A data input
DOA(0)   => data_read_a_lo(9),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(9),        -- Port B data input
DOB(0)   => data_read_b_lo(9),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_10_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000B0001800002840002C0000281800020030000000033022000000180006",
INIT_01 => X"0000098218302849180060000C00424040000000080000080200090008510200",
INIT_02 => X"0801080200100000044008000080000041000000002002400800000009008010",
INIT_03 => X"0001000004000040000202000000000802006400088000003080040008C10000",
INIT_04 => X"0000100022008000000C08C00C00000400201830040000040000000400001820",
INIT_05 => X"0200000040000000248080210044000400000000000800000004004010000800",
INIT_06 => X"0030040000404004000006D00008002010100000880800001000000030829000",
INIT_07 => X"02100000021008000940800001800010200018920206C01020200002440003C0",
INIT_08 => X"0084010110120010004000000000021F00000024400000008000440080040000",
INIT_09 => X"8288880010100001200852882004404000000008800000100001004202000280",
INIT_0A => X"0000008000020008100004590111824004000100000008012000401084080200",
INIT_0B => X"AC04400022808001200014000040001082800000000010500000010400808000",
INIT_0C => X"002200002000020002200022000020000100011082442000480909220001E020",
INIT_0D => X"0080000010044000000080080001800200000400020011000000200002000220",
INIT_0E => X"001000020001000020010010248000200010000800040000008009040000002A",
INIT_0F => X"0000000A00010200800000001400008200800000001400000000024008208041",
INIT_10 => X"0000000024008200100000001400008200100000001400002800000000000000",
INIT_11 => X"0000000000000000001400012000200000000000000000C10008400080000000",
INIT_12 => X"8000000000480000040002040000001000000000000000000004800000002800",
INIT_13 => X"0000001000000002408000000000000000000025000200020000000001200000",
INIT_14 => X"0000040000000000000029000010000200000000000000012000001000000009",
INIT_15 => X"0100000000001000000000000000010401000010000000000000000000540002",
INIT_16 => X"00001400080002100544924002A000004000020000080000000010032A000000",
INIT_17 => X"4010040100401004010040100401004010040100401004010040000000000000",
INIT_18 => X"0000000000000000000001004010040100401004010040100401004010040100",
INIT_19 => X"1080800000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"8A28A28A28D532A0CCC2A28A28A7AA344854A07F069CB8930AFD6A1AAA902A14",
INIT_1B => X"4CA6532994CA6532994CA28A28A28A28A28A28A28A28A28A28A28A28A28A28A2",
INIT_1C => X"FB3CC772B94CA6532994CA6572B95CAE532994CA6532995CAE572B94CA653299",
INIT_1D => X"55A2AABFFEF0800000000000000000000000000000000000000000000000401F",
INIT_1E => X"4BA5555401EFFFD5421EFA2FFFFF555D003FE10AAFBE8AAAA2D540000F7D57DF",
INIT_1F => X"00AAFF8002155AAFFE8B45AAD540000087FFDF45FFFBC2010AAD57DF45A28015",
INIT_20 => X"D5400FFD568B555D00155EF08040000000043DF55087BC01EF007FD75FFFF840",
INIT_21 => X"43DFEF00517DEBA007BFDFEFFFD1575EF00557DF555D517FEBA082A801EFF7FB",
INIT_22 => X"2AAAB55002E820AAAA803FEBA082AAAAAAF7FBFDE00A2FBC0145005168A10AA8",
INIT_23 => X"FAEAAB55AAD568B455D00154BAFFFBD75EF5D7BC00AAF7D5575455D557DFEF00",
INIT_24 => X"000000000002ABDF45F7803FFEF555568AAAF7802AA00FFFBD7555082E82155F",
INIT_25 => X"AAAD547038EBD57DF7DA2AEB8FC7000000000000000000000000000000000000",
INIT_26 => X"38A2DF78F45B68010482415B471C7E3DF451EFBEFBFAF4549003DE10BEF5EDAA",
INIT_27 => X"1FF087BD75D7FF84050BAEB8002155BEF5EDB6DAADF470280075FFF45E3F1C70",
INIT_28 => X"DEAA0824851EFEBFBD2410EBD168B7D410A175C7000407000140038F450075C7",
INIT_29 => X"C2155005F68A10A28438FFF00517DE82007FFAFEFE3DB505EF1C5B7AF45495B7",
INIT_2A => X"155555415178FD7082EAAB550820870BAAA8038EAA0824A8AAAEBF5FAE28AAF1",
INIT_2B => X"FFD55451C2087155EBA4A8B7DAADF68B7D4104104AAF7F1D75EF557FC70BAE3D",
INIT_2C => X"00000000000000000000000000002EB8F45F78A3DFD741516DAAAE38E2DA28EB",
INIT_2D => X"00043FE00F7D17FEBAA2D5574BAAAD17DFEFA2AEAAB550000000000000000000",
INIT_2E => X"A00557FF45A2D5554AAA2FBEAB45F78402010007BD5545AAFFD55EFF7FBE8B55",
INIT_2F => X"105D042AB550055555FF007BD7555F784174AAA28002155FFD17FFFFA2FBD74B",
INIT_30 => X"1FF557FE8B55007FFDEAA0004175FFA2FBC2000AAD16ABFF002A975450004174",
INIT_31 => X"AABAAAD56AABAAAD140155087FEAA10A28028BEF00517FE10007BE8BFFAAFFC0",
INIT_32 => X"555EF557FD54BAAAD15754508556AB45002AA8B450800174BAA68428AAA08042",
INIT_33 => X"57FEAAAAAEBFEAAAAFFD5545550015555A2842ABEFAAFBE8BFF0004020AAFFD5",
INIT_34 => X"0000000000000000000000000000000000000000000002AAAB45F7AEBFF45085",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000047FFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(10),        -- Port A data input
DOA(0)   => data_read_a_lo(10),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(10),        -- Port B data input
DOB(0)   => data_read_b_lo(10),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_11_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10180B05A0010402840602C2D001019000000300000000330A20080EC180002",
INIT_01 => X"AB400984B830084C1820E0000C36424840000000080000088200000802112220",
INIT_02 => X"8801081438106400A4F55800008000004100000040CCE24208005000C9060032",
INIT_03 => X"000406A492E6E440842254D002108153432004800880000030C0315688C00006",
INIT_04 => X"00001201200090001205400000000094108C322644240C840008030440111800",
INIT_05 => X"222000444008010028404002A002009402400025080880000C04223000170900",
INIT_06 => X"0431018040014804920906C74B32002012121004540816544522008200821100",
INIT_07 => X"3A5B1220421408004A56E840008B90D0200018B60A0650D450FC800644A0438A",
INIT_08 => X"0485816170760268E04000000000323F42C50826490640D28088445B0E041900",
INIT_09 => X"820F8B2C100000808120308020024002B3B01AC9540080A623213008800A0280",
INIT_0A => X"10000080D80381881000045B0511D28D94012671272008013002000220001240",
INIT_0B => X"8811865D22BB384100E010908060349322008000A1001C49A9348498B0808010",
INIT_0C => X"50639504395063950639504395062CA821CA8210A0040000480808214001A020",
INIT_0D => X"088812203360410110A40008553980021040465602023269400A202863950439",
INIT_0E => X"01160006000101004A01811064B050204810240812241280D00200A08044290A",
INIT_0F => X"1B0482A01AAEC3602330CD2A02952DC3502330CB4A0318B41400024008208041",
INIT_10 => X"1630144C0155C3502330CD2A02952DC3602330CB4A0318B5600C587149B6D014",
INIT_11 => X"587083B6A51005956308D1E8202C436375908AA840AD4513437640F15245B455",
INIT_12 => X"67062F47B2872400044959BC42B1060F0D036B80B548523136C158878D8FE04E",
INIT_13 => X"7010A2699AAA3794392000D81852B0A050C224180062085134CD1719564E020C",
INIT_14 => X"400C50500D94C8121713C02B555101C90705D71009604140C0418CE0C378F0B2",
INIT_15 => X"27C828E024D8C50965A40821568A06113801505010334AA73AA0666DAC20AD57",
INIT_16 => X"048123408C0822040004C248604B2100400100084008001D0113920060CDC06A",
INIT_17 => X"4812048120481204812048120481204812048120481204812048120481204812",
INIT_18 => X"8020080200802008020081204812048120481204812048120481204812048120",
INIT_19 => X"1420000000000000000002008020080200802008020080200802008020080200",
INIT_1A => X"2082082082815220A4A380000002A8313044020C0605885026853A1082100A00",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000008208",
INIT_1C => X"F83F070000000000000100800000000000000000004020000000000000000000",
INIT_1D => X"EF0855400005500000000000000000000000000000000000000000000000401F",
INIT_1E => X"AAAA2D540000F7D57DF55A2AABFFEF0804155EFAA842ABEFA280155EFFFFBC01",
INIT_1F => X"FF555D51575FFA2FFD75FF550015400FFFBFFF4508514000000003FE10AAFBE8",
INIT_20 => X"155EF0051555FF0804155FFF7D57DF45A280154BA5555401EFFFD5421EFA2FFF",
INIT_21 => X"002155AAFFE8B45AAD540000087FFDF45FFFBC2010AAD568AAAAAD142145FF80",
INIT_22 => X"7FD75FFFF84000AAFF802ABFFA2AABFE1008001540008514215555003DFFFA28",
INIT_23 => X"85142010FFAE800AA5D7BFDF45F7FFEAA0000040000000043DF55087BC01EF00",
INIT_24 => X"00000000000517FEBA082A801EFF7FBD5400FFD568B555D00155EF085168B450",
INIT_25 => X"7BE8A155EFE3FBC71FF145B42038550000000000000000000000000000000000",
INIT_26 => X"381C003DE10BEF5EDAAAAAD547038EBD57DF7DA2AEB8FC70000175EFB6802DBC",
INIT_27 => X"1C7E3DF451EFBEFBFAF45495F575FFBEF5D05EF550E15400E3F1FFF7D085B420",
INIT_28 => X"8ABAB6D145145FF84155D7085B555C71404105C7F7DF78F45B68010482415B47",
INIT_29 => X"4515549003FFC7BE8002155BEF5EDB6DAADF470280075FFF45E3F1C7038A2DB6",
INIT_2A => X"038F450075C71FF087BD75D7FF84050BAEB8428BEFBEA4BDE28140A154380051",
INIT_2B => X"0A175C7005B6DB55145140000FFAE85082417FFFF7DE3F1EFA10140407000140",
INIT_2C => X"00000000000000000000000000005B7DEAA0824851EFEBFBD2410EBD168B7D41",
INIT_2D => X"0004175FFF7803DF45FFAE955EFAAFBD55EF557BC20AA5D00000000000000000",
INIT_2E => X"0AAD17DFEF007FC20AA5D043FE00F7D17FEBAA2D5574BAAAD17DFEFA2AEAAB55",
INIT_2F => X"45F78402010007BD5545AAFFD55EFF7FBE8B55007FD75FFF7D5401EF5D2E9741",
INIT_30 => X"F45A2D5554AAA2FBEAAAAFFD555545FF8015555007FD5545550400145FFFBEAB",
INIT_31 => X"DEAA5D2E974AA00515754500003FF55FF8002155FFD17FFFFA2FBD74BA00557F",
INIT_32 => X"7FE105D04174105D042AB550055555FF007BD7555F784174AAA2842ABEFFF803",
INIT_33 => X"BC2000AAD16ABFF002A97545007FFFF45555540000FFAE97410007BFFFFFA2D5",
INIT_34 => X"0000000000000000000000000000000000000000000007FFDEAA0004175FFA2F",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000040000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(11),        -- Port A data input
DOA(0)   => data_read_a_lo(11),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(11),        -- Port B data input
DOB(0)   => data_read_b_lo(11),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_12_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50080B01BC002006940202C0DE041196A83183000000023322287E0FC000006",
INIT_01 => X"0E000C048000C048400380000007026040000000080000088200002802153231",
INIT_02 => X"2809AD0E7D180040945008040090000061800000C0E2F66009DA3D11CB148015",
INIT_03 => X"210D050012F6F8D2108216E24842005B8A20640008800000B8E0141C28851006",
INIT_04 => X"0080100022408000060DE0000066630C70241827041000040800820480001AA4",
INIT_05 => X"0240000C400000003C808003E0C8001401000000040900020904004000070800",
INIT_06 => X"00300D800C1960C4400006E10B90002018184000100804005784000130821200",
INIT_07 => X"0652428112180C03E8E5A2C800A3F018200418927E06686450FF8006460003A0",
INIT_08 => X"09840903525281D4F460409000000E3F08D1202C5C26A0719CC96CC7BF462990",
INIT_09 => X"82488BAE10000040000410802008600843001E09F00000276F81020000230280",
INIT_0A => X"00000080000C000C100204593F11A489F480067D04D40C012400080000800240",
INIT_0B => X"0800021826933E03662802B300003C13E0000000460000000000010CE0000000",
INIT_0C => X"78419784197861978419784197860CBC30CBC20000000010400808056500A080",
INIT_0D => X"201E7F3F01F40401C17E800C7F33800200000357008C0249E2DE0D7841978619",
INIT_0E => X"0F500002200004005002001408400000000000000000000053A4096F80705FA0",
INIT_0F => X"1B17B2C53F2FC16691DB587201EDDF4162B1DB527201EDDC4607024100100020",
INIT_10 => X"F2A01D5CC9794162B1DB587201EDDF416691DB527201EDDD884272592D6246FC",
INIT_11 => X"7258E995D5A825DBA569F9FF02547068618CD3CC45B7863AE7EC00D4B122A67D",
INIT_12 => X"C6CCA5C33717461C045B5B182019473D19D7CCD856106F31A683621BDFC28800",
INIT_13 => X"FB10A652CC8E3538BBA01624E51AA6C0469AC5493F5688532966471A9C5F6208",
INIT_14 => X"40041E1F5759001B4AA1853E6D5144AA9C914C8608D2724A4C4118D992B866E2",
INIT_15 => X"AD9825682D4A36C0B0B4B85112B2C4A05D3E6D5051893335EB0072AA85A4F9B7",
INIT_16 => X"000008000000821000048260020000004001DC0800000010E7F70171401DE07E",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0100401004010040100400000000000000000000000000000000000000000000",
INIT_19 => X"1080800000000000000000040100401004010040100401004010040100401004",
INIT_1A => X"249249249120780800016A28A288028DCA30444409B054A88C5890486582A210",
INIT_1B => X"86432190C86432190C8641041041041041041041041041041041041041049249",
INIT_1C => X"FBC007592C964B2592C964B2592C964B2592C964B2592C964B2592C964B2592C",
INIT_1D => X"FF55002ABEF0800000000000000000000000000000000000000000000000401F",
INIT_1E => X"BEFA280155EFFFFBC01EF0855400005555421FF00042ABEFFF8400010082EAAB",
INIT_1F => X"FFEF08556AA10000028AAAFFD15541000002ABEFFFFBD54000004155EFAA842A",
INIT_20 => X"001FF00041554555557FE005D003FE10AAFBE8AAAA2D540000F7D57DF55A2AAB",
INIT_21 => X"1575FFA2FFD75FF550015400FFFBFFF45085140000005168AAA087BFFFFF5D04",
INIT_22 => X"D5421EFA2FFFFF555D0000145082E955FF0851555FF082AA8B55F7AEA8BEF555",
INIT_23 => X"000020BAAA801541055042ABEFFFFBD5410AAD57DF45A280154BA5555401EFFF",
INIT_24 => X"000000000005568AAAAAD142145FF80155EF0051555FF0804155FFF7842AA100",
INIT_25 => X"7EB80000280824ADBD7490E28BEF080000000000000000000000000000000000",
INIT_26 => X"101C00175EFB6802DBC7BE8A155EFE3FBC71FF145B42038555F401D71C0A2DBC",
INIT_27 => X"038EBD57DF7DA2AEB8FC7005F6AA381C0A2DA82FFDB5243800002FBD7EBFBD24",
INIT_28 => X"AA82147FF8FEF410E001FF000E17555555B7AE1041003DE10BEF5EDAAAAAD547",
INIT_29 => X"ADB45F7AEA8BEF555F575FFBEF5D05EF550E15400E3F1FFF7D085B420381C5B6",
INIT_2A => X"010482415B471C7E3DF451EFBEFBFAF4549000017D142E905EF1451525C7082A",
INIT_2B => X"04105C7F7842FA381C0A00082AA8A1041041002FBEFEBFBD2410AADF78F45B68",
INIT_2C => X"00000000000000000000000000005B68ABAB6D145145FF84155D7085B555C714",
INIT_2D => X"5D7BC01555D2EBFF55A284000AA08003FF55002AA8BEF0000000000000000000",
INIT_2E => X"A08003FF55A2FBC00105D04175FFF7803DF45FFAE955EFAAFBD55EF557BC20AA",
INIT_2F => X"00F7D17FEBAA2D5574BAAAD17DFEFA2AEAAB55007BE8AAA5D2EBDE00FFFFC00A",
INIT_30 => X"FEF007FC20AA5D7BE8A005D7FEABFF002E821FF082A97555557FE8A0000043FE",
INIT_31 => X"01EF5D5142145082EBFF55F7AAAABEF5D7FD75FFF7D5401EF5D2E97410AAD17D",
INIT_32 => X"C2010A2FBEAB45F78402010007BD5545AAFFD55EFF7FBE8B550004001FF5D2A8",
INIT_33 => X"015555007FD5545550400145FF843DEAA552A82010A2AA8000008043FFFFA2FB",
INIT_34 => X"0000000000000000000000000000000000000000000007BEAAAAFFD555545FF8",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000007FFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(12),        -- Port A data input
DOA(0)   => data_read_a_lo(12),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(12),        -- Port B data input
DOB(0)   => data_read_b_lo(12),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_13_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10110A0441812402840402822007818000E00700000000330A3000000008042",
INIT_01 => X"A1400984B830C848180260000C0042404001000008220008A200100802110200",
INIT_02 => X"88010C02801040002475580400800000410000000064024608134C0CC9018034",
INIT_03 => X"00010100926220D084234212421085084300648A0880000630C0654288C10000",
INIT_04 => X"0004122122029100100C00001200009C40A83A2044360C84190BAC04E0101820",
INIT_05 => X"027000004009050064C8C00104C10184034010250089C00EB004327064B60900",
INIT_06 => X"543000004080480492A946CE1032002012125804440812541027008230821380",
INIT_07 => X"0A581424525408000AE2AA8002BC00D020003896020658FC4030000246E543AE",
INIT_08 => X"04840101107200B80040210000002ABF02450A264002C8008000441680041900",
INIT_09 => X"825A98801000008001041080200B660E30B200C8840080808065102000280280",
INIT_0A => X"00000080C90391881000145B0111A30404016003A56008012C80080200801280",
INIT_0B => X"08088C5D2288004120E80290882400908000A000A1000809A93485D610000000",
INIT_0C => X"002000000000000002000000000000001000000000000000400808154100A080",
INIT_0D => X"08000000360401021280800E400B800610C84100014224200000000020000000",
INIT_0E => X"0086000600040D045E4195104D5854284A14250A12A512A8808289840084A020",
INIT_0F => X"0949E07A80948354B6E68982167061037496E683821670620681024000000000",
INIT_10 => X"8E510B456587037496E689821670610354B6E6838216706220431961CA985D48",
INIT_11 => X"196186A91674011CE61403562274AA49CD594CF00039C7C414B6509DA2265213",
INIT_12 => X"A983014780CC8604040424A5323845932E620295879818170304B2F5002C2043",
INIT_13 => X"451654B9104A328665603148895D44E0251142B42A3D8B2A5C8825194328A2E6",
INIT_14 => X"C06A6C6A465AA0091482382B17614F2202858EE300991415B45CD5306028F019",
INIT_15 => X"52E08DC8047F17D1C7C3C02128E587D6A02B17605A130A4E8BF002258850AC5D",
INIT_16 => X"84A123508508220808048240604B2100C00022084809000D000393722A140000",
INIT_17 => X"4A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A12",
INIT_18 => X"A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A128",
INIT_19 => X"154000000000000000000284A1284A1284A1284A1284A1284A1284A1284A1284",
INIT_1A => X"BAEBAEBAEBFF6FEFEFEEEAAAAAAFBF7DDF77F9FBEFBFF9F3F0FDFCFBEFBF1228",
INIT_1B => X"5FAFD7EBF5FAFD7EBF5FAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAE",
INIT_1C => X"F800077EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF",
INIT_1D => X"00FFD140155F780000000000000000000000000000000000000000000000401F",
INIT_1E => X"BEFFF8400010082EAABFF55002ABEF08556AAAA5D043FFFFAAAABDEAA557BFDE",
INIT_1F => X"000055043DEBAF7843FFFFF7AABDF55A2AA97400AAD540155A2D5421FF00042A",
INIT_20 => X"E8B45557FD7410552EAAABAAA84155EFAA842ABEFA280155EFFFFBC01EF08554",
INIT_21 => X"56AA10000028AAAFFD15541000002ABEFFFFBD5400005568A1055043DEBAAAFF",
INIT_22 => X"D57DF55A2AABFFEF085557545FFD17DEBAA2FFE8ABAAA8428A00087BD7555FFD",
INIT_23 => X"57BEAABA5D2ABDF450851420AA5D7FD5555A2803FE10AAFBE8AAAA2D540000F7",
INIT_24 => X"000000000005168AAA087BFFFFF5D04001FF00041554555557FE005D00001555",
INIT_25 => X"7AAA4B8E824971F8E38E3DF45155EB8000000000000000000000000000000000",
INIT_26 => X"55A2DF401D71C0A2DBC7EB80000280824ADBD7490E28BEF08516DA82410A3FFD",
INIT_27 => X"5EFE3FBC71FF145B42038550E38E92EB803FFD7EBA4BDF45AAAA90410BEDF451",
INIT_28 => X"FA38490A3FE92BEFFEAB45417FD24385D2AAFA82B680175EFB6802DBC7BE8A15",
INIT_29 => X"28A10007FD557DFFDF6AA381C0A2DA82FFDB5243800002FBD7EBFBD24101C556",
INIT_2A => X"5EDAAAAAD547038EBD57DF7DA2AEB8FC700515056DE3D17FE92BEF1EFA92AA84",
INIT_2B => X"5B7AE10410E00155497FEFABA4120B8F55085B400925D7FD557DA2803DE10BEF",
INIT_2C => X"00000000000000000000000000005B6AA82147FF8FEF410E001FF000E1755555",
INIT_2D => X"00517FE00082EBDF45AA8428A10085568ABAA2FBD7545AA80000000000000000",
INIT_2E => X"5AAAE82000F7FBD5545AAFBC01555D2EBFF55A284000AA08003FF55002AA8BEF",
INIT_2F => X"FFF7803DF45FFAE955EFAAFBD55EF557BC20AA5D2EA8A00A2803DF45AA843DF5",
INIT_30 => X"F55A2FBC00105D517FEAA082EBFE10F7FFE8B55087FC00BA552ABFE10F784175",
INIT_31 => X"FE10F7D57DE00AA842AA00007FD75FFF7FBE8AAA5D2EBDE00FFFFC00AA08003F",
INIT_32 => X"D55FFAA843FE00F7D17FEBAA2D5574BAAAD17DFEFA2AEAAB550051401FFA2D57",
INIT_33 => X"E821FF082A97555557FE8A00002E82155007BFDEAA08042AB45087FC0010557F",
INIT_34 => X"0000000000000000000000000000000000000000000007BE8A005D7FEABFF002",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000067FFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(13),        -- Port A data input
DOA(0)   => data_read_a_lo(13),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(13),        -- Port B data input
DOB(0)   => data_read_b_lo(13),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_14_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10020A000180000284008280000281800000030000000033022000000580002",
INIT_01 => X"A140098018300848184860000C20C24040000000084000084200000000110200",
INIT_02 => X"88010C5A8010A600A4F558040080000041000000022C024008003CCCC9028030",
INIT_03 => X"000103A7A00904D0842242024210810803006480088000003081054288C10000",
INIT_04 => X"0000120122009000100C00000000000400A83A2044200C840000800400101820",
INIT_05 => X"020000004008010024C0C0010040000402000025000800020004207000100800",
INIT_06 => X"0430000040004804920906C20022002012120004440812541020008230821000",
INIT_07 => X"2A5A14285A15080008768A80008000D0200018B202067AF100A0000244204382",
INIT_08 => X"04850101105205380040000000000A7F42840A264920406080004400A0040900",
INIT_09 => X"8208888010000080010010802000400230B000C8840080800021100000200280",
INIT_0A => X"00000080C8038188100004590111B68404012000016008012000000000000200",
INIT_0B => X"080084452280004120400000802000908000800001000009A924810410000000",
INIT_0C => X"000000000000200000000000000200000000000000000000400808000000A080",
INIT_0D => X"080000002204010010808008000B800210404100000220200000000020000200",
INIT_0E => X"0000000600000000020181100400502048102408122412808082098400042020",
INIT_0F => X"0480040A100A42008000161C140000420080001C1C1400003201024000000000",
INIT_10 => X"39600022260042001000161C140000420010001C1C140001604E8084341CBA34",
INIT_11 => X"8082580E2B8802201014800C220A21829A302F1C024010C001124020C8C1A8A0",
INIT_12 => X"CA60CA000048228404401004418012787124648157780120B8678C000801E04E",
INIT_13 => X"001072D04730000241000CB1325E78E0186030240000083B602398000120024A",
INIT_14 => X"001EF6F4163C480481506800004000CFD55196CB012481812049495C19400009",
INIT_15 => X"248800108B8FB61A0401200845594965000000400568D0CFB780055060500001",
INIT_16 => X"048123408408220000048240604B210040000008400800B0000090022A140068",
INIT_17 => X"4812048120481204812048120481204812048120481204812048120481204812",
INIT_18 => X"8120481204812048120481204812048120481204812048120481204812048120",
INIT_19 => X"1400000000000000000002048120481204812048120481204812048120481204",
INIT_1A => X"9E79E79E79FF3BEEEEEFE79E79EFAABCDA72E47F87BDF4EBAE7CFAFBEFB28200",
INIT_1B => X"CFE7F3F9FCFE7F3F9FCFE79E79E79E79E79E79E79E79E79E79E79E79E79E79E7",
INIT_1C => X"FBFFF83F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9F",
INIT_1D => X"555D5568A105D00000000000000000000000000000000000000000000000401F",
INIT_1E => X"FFFAAAABDEAA557BFDE00FFD140155F7D17DF45AAD157400007BEAAAAAAAE955",
INIT_1F => X"ABEF085155400FFD1420100055574AAA2AA800AAF784020AAF7D56AAAA5D043F",
INIT_20 => X"FFE105D7BD7545A284020BA0055421FF00042ABEFFF8400010082EAABFF55002",
INIT_21 => X"43DEBAF7843FFFFF7AABDF55A2AA97400AAD540155A28028B550051574005D7F",
INIT_22 => X"FBC01EF08554000055002AB455D51420100851421FF5D7FFDEBA085168B45FF8",
INIT_23 => X"AD140000002EBFFEFA2AAA8BEFF780021FF5504155EFAA842ABEFA280155EFFF",
INIT_24 => X"000000000005568A1055043DEBAAAFFE8B45557FD7410552EAAABAAA8017400A",
INIT_25 => X"01C71EDA82AAA0955455D556DA00490000000000000000000000000000000000",
INIT_26 => X"BAEBD16DA82410A3FFD7AAA4B8E824971F8E38E3DF45155EBD17FF6DAADB5040",
INIT_27 => X"0280824ADBD7490E28BEF085157428FFDB420101C55554AAAAA480082FF84000",
INIT_28 => X"AB7D0051504005D71F8E004975D556DB68405092085F401D71C0A2DBC7EB8000",
INIT_29 => X"FAEAA08516AB45E38E38E92EB803FFD7EBA4BDF45AAAA90410BEDF45155A28E2",
INIT_2A => X"02DBC7BE8A155EFE3FBC71FF145B42038550028B6D5D51420101C5B401EF417B",
INIT_2B => X"2AAFA82B68015400AADB40000082EBFFC7A2AEAFBC7EB80071FF5500175EFB68",
INIT_2C => X"0000000000000000000000000000556FA38490A3FE92BEFFEAB45417FD24385D",
INIT_2D => X"AAD17DFFFAAFFC200055557DE00A2801554555557FE100000000000000000000",
INIT_2E => X"AA28400000F784020BAAAD17FE00082EBDF45AA8428A10085568ABAA2FBD7545",
INIT_2F => X"555D2EBFF55A284000AA08003FF55002AA8BEF0051554AAFFFFC00105D55554B",
INIT_30 => X"000F7FBD5545AAAEAABFF0051400105D5568A000051575FFF78415410087BC01",
INIT_31 => X"2000557FC01EF007FEAABA00556AB55A2AEA8A00A2803DF45AA843DF55AAAE82",
INIT_32 => X"175FF5D04175FFF7803DF45FFAE955EFAAFBD55EF557BC20AA5D042ABFF55514",
INIT_33 => X"FE8B55087FC00BA552ABFE10F78415400A2FBC0010082EBDF55A2AABDF45A284",
INIT_34 => X"000000000000000000000000000000000000000000000517FEAA082EBFE10F7F",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000007FFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(14),        -- Port A data input
DOA(0)   => data_read_a_lo(14),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(14),        -- Port B data input
DOB(0)   => data_read_b_lo(14),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_15_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000A000000000284000280000001800020030000000033022000000180002",
INIT_01 => X"A140098018300848180060000C00424040000000080000080200000000110200",
INIT_02 => X"080108000010E60004E55800008000004100000000040240080000C009170016",
INIT_03 => X"0000000080000040842240000210810002000400888000003080014288C00000",
INIT_04 => X"0001100024A0800000440000000000040088322044200C840000011400151800",
INIT_05 => X"A200014C4000000020000000000B8094020000254C8800000514203000108800",
INIT_06 => X"0031042040804804100006EE4032002012120005540812540020008600831000",
INIT_07 => X"021912244A14080008408880008000D020001892020656300020000244000380",
INIT_08 => X"048501415032000800406180000002DF02440826400000008000440000043080",
INIT_09 => X"8208880110000000010010802000400230A000880400808000450200000B0280",
INIT_0A => X"00000080C003010810000459011182040400200003E0080120000000000002C0",
INIT_0B => X"080084452280004100400000800000100000800001000001A124800010000000",
INIT_0C => X"002000020000000000000000000200001000010000000000400808000020A000",
INIT_0D => X"08000000260001001280000C400B000200000000000220200000000020000200",
INIT_0E => X"008400060000000000010010040040000000000000201000000000000004A000",
INIT_0F => X"0000000000000202100000000000000202100000000000004600024000000000",
INIT_10 => X"0000000000000202800000000000000202800000000000002000000800000000",
INIT_11 => X"0008000000000000000000002000100800000000000000000000400001200000",
INIT_12 => X"00880000000006000400080C0000000000D08120280000000000000000002000",
INIT_13 => X"0010040200000000010000004020010000000000000008000900000000000200",
INIT_14 => X"0000000308801400000000000040000008822110000000000040100100000000",
INIT_15 => X"0080000000004840717050000000000000000040000020000000000000000001",
INIT_16 => X"000023000000220000048240404A010040000008000000000000000020C40000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"1400000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000200",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"F800000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"AA007BC2145F780000000000000000000000000000000000000000000000401F",
INIT_1E => X"400007BEAAAAAAAE955555D5568A105D7FC00000804154AA5D00001EFF78428A",
INIT_1F => X"0155F7FBD74AAAAD17DF45F7D1421EF0055400AA007FC2000F7D17DF45AAD157",
INIT_20 => X"BDFEF08517DF55A2FBEAB555D556AAAA5D043FFFFAAAABDEAA557BFDE00FFD14",
INIT_21 => X"155400FFD1420100055574AAA2AA800AAF784020AAF7FFFDF45FF84000BA552A",
INIT_22 => X"2EAABFF55002ABEF087BE8ABA555168B55AAFFEAB45F7843FF45082A801FF005",
INIT_23 => X"284000AA0055401550055574005D2E800AAA2D5421FF00042ABEFFF840001008",
INIT_24 => X"000000000000028B550051574005D7FFFE105D7BD7545A284020BA007FFFE10A",
INIT_25 => X"2550E021C7EB8028A821C7BC516DFF8000000000000000000000000000000000",
INIT_26 => X"28FFD17FF6DAADB504001C71EDA82AAA0955455D556DA004971C703814001248",
INIT_27 => X"E824971F8E38E3DF45155EBF1D5492BED17FF45E3DF471C70851400BA0071C50",
INIT_28 => X"FF7DEB8000092552ABFFEF08517DF6DB6FBE8B555D516DA82410A3FFD7AAA4B8",
INIT_29 => X"3DF551C20801C71C5157428FFDB420101C55554AAAAA480082FF84000BAEBF1F",
INIT_2A => X"A2DBC7EB80000280824ADBD7490E28BEF087FEFA8241516DB55A2FFEAB6DEB84",
INIT_2B => X"8405092087FF8E00BE8A02082005F47145085550428412A85082BEDF401D71C0",
INIT_2C => X"00000000000000000000000000000E2AB7D0051504005D71F8E004975D556DB6",
INIT_2D => X"0055554BA5504000105D2A80145AA842AA00557BD75EFF780000000000000000",
INIT_2E => X"50055420BA0055574BAF7D17DFFFAAFFC200055557DE00A2801554555557FE10",
INIT_2F => X"00082EBDF45AA8428A10085568ABAA2FBD7545AAD557410F7D57DF55AAFBD554",
INIT_30 => X"000F784020BAAAD57FFEFA28402010552ABDFFF08517FFFFF7FBEAB455D517FE",
INIT_31 => X"DF45AAFBE8BEFA2803FF455504001555551554AAFFFFC00105D55554BAA28400",
INIT_32 => X"95400F7FBC01555D2EBFF55A284000AA08003FF55002AA8BEF007FFDE1000557",
INIT_33 => X"568A000051575FFF78415410087FEAA10F7AE80000087BD55450855400BA002A",
INIT_34 => X"0000000000000000000000000000000000000000000002EAABFF0051400105D5",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000060000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(15),        -- Port A data input
DOA(0)   => data_read_a_lo(15),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(15),        -- Port B data input
DOB(0)   => data_read_b_lo(15),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_16_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"DA22C618B1000482B688B186588884862A400438255FC38381441205BA803003",
INIT_01 => X"8645A80028404C211203A952A90341080B173340412000E1005D628000820484",
INIT_02 => X"A101A9006DC1084833011850AAC55001349B10881802821808B4110007005E11",
INIT_03 => X"010108A802BB00080080006020020001A61036202800000D2410104200404550",
INIT_04 => X"8BFA58800005C40A46240252145148B38248030356415A4E62B6FC660F287240",
INIT_05 => X"0F05EA11E570000D610000000710296E542B6E3A825C15FB30A643695BFC2D56",
INIT_06 => X"00640044150C025A0000000901A054F2C0A8030140BCC0460050690A95C8383D",
INIT_07 => X"0288500102F85203E8010D0AA9BC4800015001219D0550077373CAA804000680",
INIT_08 => X"A2064193920A2004B51400001414091EAA14881C0002701881B120203B7A8012",
INIT_09 => X"C8204D02D965965200100104F2B0082251200000023153000C4400800000ACCA",
INIT_0A => X"000012C9000A0000D0A80000BF8028E87C1B9246002A8A562060410280081116",
INIT_0B => X"240014891801000495D40192D1000000000000A8A5AA80018120E00066000000",
INIT_0C => X"00088000880008800088000880008400044000400029011404008401CA809004",
INIT_0D => X"0140A80A5C8000102ED0044008004AD32400004001AB08C0031EDA7B08800088",
INIT_0E => X"04912AA28AA890BA00000024800480000000000000200802151025062C0BB400",
INIT_0F => X"1F554E11C596A64003195933741477264003195555B418687E35836020814004",
INIT_10 => X"0A499CF47DCB264003195933741597264003195555B4198843940076D296D003",
INIT_11 => X"00758486A556489347FE5F409CBC1362510695B6288743123C95251852041CD5",
INIT_12 => X"424EAE2992046EB70026486035600CEC45CBCA809654B48163CCC895E1E043D4",
INIT_13 => X"98E3A242DEA151848302BFD6D522B10C7EC71F6C1DB071D1216E078C4C1B1C74",
INIT_14 => X"037DAAABC982BE22267A2E2E4F44AA1DC5E37400C9EE1B7B638E8849D23C3832",
INIT_15 => X"2EE015998B28654565A003F0068E35352C1CAE48BFBF3A6C9B7B286B4DA8B93D",
INIT_16 => X"000009000040A8000452110A8442040D655602A102A0027E2C42320284086E6A",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"1451451451E96F2FC3C34F3CF3C2AC688AA263486D3260E34C0C3A7B451B0200",
INIT_1B => X"9F47A7D1E9F47A7D1E9F4D14D14D14D14D14D14D14D14D14D14D14D14D145145",
INIT_1C => X"F800007D3E9F4FA7D3E8F47A3D1E8F47A3D1E8F47A7D3E9F4FA7D3E9F4FA7D3E",
INIT_1D => X"FF00003FE005500000000000000000000000000000000000000000000000401F",
INIT_1E => X"4AA5D00001EFF78428AAA007BC2145F7843FFFFF7FBE8B45AAD568BFFFFAA975",
INIT_1F => X"8A105D2E974BAF7FBEAB45FFFFC00BAF780020005D2A95410FFFFC0000080415",
INIT_20 => X"821FFA2AAAAA00000417555FFD17DF45AAD157400007BEAAAAAAAE955555D556",
INIT_21 => X"BD74AAAAD17DF45F7D1421EF0055400AA007FC2000F78000010552E800AA002E",
INIT_22 => X"7BFDE00FFD140155F7AABDF55F7AE820AA08043FEBA5D55575FFF7AABFE00557",
INIT_23 => X"2FBE8B55FFFFD55FF557FC2000FF8015410FFD56AAAA5D043FFFFAAAABDEAA55",
INIT_24 => X"000000000007FFDF45FF84000BA552ABDFEF08517DF55A2FBEAB555D04154BAA",
INIT_25 => X"5B6DF6DBFFF7AA955C71C043FE10490000000000000000000000000000000000",
INIT_26 => X"38FFF1C7038140012482550E021C7EB8028A821C7BC516DFF8438FC7E3F1EAB5",
INIT_27 => X"A82AAA0955455D556DA00492490492F7FBE8B55FFF1C70BAF78A000005D20974",
INIT_28 => X"20285D2085092002A801FFB6AAA8A10080E1757DEBD17FF6DAADB504001C71ED",
INIT_29 => X"555FFE3AABFE005D71D5492BED17FF45E3DF471C70851400BA0071C5028FF840",
INIT_2A => X"A3FFD7AAA4B8E824971F8E38E3DF45155EBA4BAF6DE3AA8709208043FEBA555B",
INIT_2B => X"FBE8B555D04124BAB6FBE8B45E3FBD55D7557BC0028E38412428EBD16DA82410",
INIT_2C => X"000000000000000000000000000071FFF7DEB8000092552ABFFEF08517DF6DB6",
INIT_2D => X"F78428B55AAD168B55F7FFFDFEFFFAA9555555003DE000000000000000000000",
INIT_2E => X"AFFAE820105500154AAF7D5554BA5504000105D2A80145AA842AA00557BD75EF",
INIT_2F => X"FFAAFFC200055557DE00A2801554555557FE10000000010F7FBEAB45FFD1554A",
INIT_30 => X"0BA0055574BAF784000BA5D0017410082E801EFF7AEA8A10002E955FFA2D17DF",
INIT_31 => X"541000003DEBA557BD75EFA2AEBDE105D5557410F7D57DF55AAFBD5545005542",
INIT_32 => X"000AAAAD17FE00082EBDF45AA8428A10085568ABAA2FBD7545AA802ABEFA2AA9",
INIT_33 => X"ABDFFF08517FFFFF7FBEAB455D04020AAFFFBEAB45AAFFD55555D7FC20AAA280",
INIT_34 => X"000000000000000000000000000000000000000000000557FFEFA28402010552",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000020000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(16),        -- Port A data input
DOA(0)   => data_read_a_lo(16),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(16),        -- Port B data input
DOB(0)   => data_read_b_lo(16),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_17_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"5284CE4FB7BD2C8994A13392DBD02E14006B82AC7E800D44D3DD2FD5F9B961C0",
INIT_01 => X"F8ACD01F7E03FC6793F2199B39FC233C11D93AE6F3BB92B32091DBC339B24542",
INIT_02 => X"8F333007FD6808092A2AFA6667033DB50853379C10BFF70F1BD011110F205F18",
INIT_03 => X"294ADB4AFFCBF0DAD63ABF836B58EAFE060478202022234B2E0303FDC9E18339",
INIT_04 => X"DB7A40806FE4040840EBC563A0150A0926146FECB04196482236FC2005282AE1",
INIT_05 => X"0403DA0383200831C68206D7E6D0250834336D1E81500FDB306045255BFC2076",
INIT_06 => X"000A0E2D7D3EAFF15800100FBFB333C1CBC303163670497AFF00291B3C0E2015",
INIT_07 => X"451C581123AEE54DE8008B719E61C10BBA5DAAFA9DDA1194D51E067BB0000000",
INIT_08 => X"70320A9392083056C2270E004400091181168C4D14002A110C902481FC0B4212",
INIT_09 => X"0E28EFFC40C30E5F0182D0950190C0810BE00E9A76E4C7FD0E4700000B303806",
INIT_0A => X"C7DEF207000F00059D2ED56D7EED2ED3C9A86FB8013E7437823DF78CDB6CA60E",
INIT_0B => X"7C00319F8E853E64D73A08BFF0001D35682AC0CE8FCCC200A59BDD2FFE3F3EC7",
INIT_0C => X"7A7DE7A7DE7A7DE7A7DE7A7DE7A7DF3D3EF3D3C0030B889723782E816EC0A081",
INIT_0D => X"2D4CFEB69FF7A5F5AFFCCA787F7FE67C21800367451F8355EB9EDE7A7DE7A7DE",
INIT_0E => X"2C9F99FD0678B87A0003000D8D02E00000000000000040025D3C21463D6BFF25",
INIT_0F => X"232221ABD9CA854DFDD64A67D42C0F054DFDD64667D42C063E57A8F7B4594BB0",
INIT_10 => X"AEDAA504801F054DFDD64A67D42C0F054DFDD64667D42C07237DFE5865F6D2BF",
INIT_11 => X"FE58EAE7F5AB50D0806A9A2E0DFFF47DEDC496DA3181A0CC71440F9FBC3EFBB5",
INIT_12 => X"9C9C3FC95949AEFF556EF9C75E7DCF1EB1B6E6FCDC87CB35FC94B36AECF3A33D",
INIT_13 => X"382AF5B6AAAE594A4C0DBFDAD94AA669809809FEFAF4157ADB55572CA527056E",
INIT_14 => X"1AE33F32ADD543430808BABAF50E1A5EB4BAEA45A250202FE0ADD39387F92B29",
INIT_15 => X"669523E865D4B1293AB6B90BF2F0E30EDEFAFD0B3FBD72E9E90D20A003FBEBF4",
INIT_16 => X"00002F840000BCE0B6F67B3F845E017C833F6AAC02B002A2EFF22D4073DE83FB",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0600000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"9A69A69A6A4624C3434C0EBAEBA21B9001804F6E62029749701020B88A7CC0C0",
INIT_1B => X"41A0D46A341A0D46A341A69AEBA69A69AEBA69AEBA69A69AEBA69AEBA69A69A6",
INIT_1C => X"F8000046A351A8D46A351A8D46A351A8D46A351A8D068341A0D068341A0D0683",
INIT_1D => X"00F7D56ABFF55000000000000000000000000000000000000000000000007FFF",
INIT_1E => X"B45AAD568BFFFFAA975FF00003FE0055043FFFFFFFFFFFFFF7FBFDF55A284020",
INIT_1F => X"2145F7D568B45000002010552EBDF45A28028A00F7843FEBA55043FFFFF7FBE8",
INIT_20 => X"95410AAAEBFF55AAFFC00BAF7FFC00000804154AA5D00001EFF78428AAA007BC",
INIT_21 => X"E974BAF7FBEAB45FFFFC00BAF780020005D2A95410FFAE800105D2A95410002A",
INIT_22 => X"AE955555D5568A105D7FFFFEFA2D568BFFFFD57DE00F7AE800AAAAAABDFEF5D2",
INIT_23 => X"82A974105D003FF55F7802AAAAAAD168AAA5D517DF45AAD157400007BEAAAAAA",
INIT_24 => X"000000000000000010552E800AA002E821FFA2AAAAA00000417555FF8028B550",
INIT_25 => X"FE3F5FAF45AA8000038F7DB6FBD7490000000000000000000000000000000000",
INIT_26 => X"82490438FC7E3F1EAB55B6DF6DBFFF7AA955C71C043FE10490A3FFFFFFFFFDFE",
INIT_27 => X"1C7EB8028A821C7BC516DFFDF68B551C0E050384124BFF7DB68A28A38F7803DE",
INIT_28 => X"5000492495428082E95400AAA0BDF7DB6F5C70BAFFF1C7038140012482550E02",
INIT_29 => X"800BAB6AEBDFD75D2490492F7FBE8B55FFF1C70BAF78A000005D2097438FFAA8",
INIT_2A => X"B504001C71EDA82AAA0955455D556DA00497FFAFFFB6D56FBFFEBDB78E38F7AA",
INIT_2B => X"0E1757DEB8A2DB5514249243841003FF6DEB8028AAAB6D16FA8249517FF6DAAD",
INIT_2C => X"000000000000000000000000000004020285D2085092002A801FFB6AAA8A1008",
INIT_2D => X"002ABFFEFF7FBFDFFFAAD168B55AA80000BAF7FFFDF550000000000000000000",
INIT_2E => X"FFFAAA8AAAF7843FE10000428B55AAD168B55F7FFFDFEFFFAA9555555003DE00",
INIT_2F => X"BA5504000105D2A80145AA842AA00557BD75EFF7FBEAB45552E954BA08003DFF",
INIT_30 => X"0105500154AAF7AE974000800154AA002E95410AA843FFFFF7D5554BAF7D5554",
INIT_31 => X"FFEFAAFFE8ABAFFAA820BAF7AEBFF55550000010F7FBEAB45FFD1554AAFFAE82",
INIT_32 => X"7DE0000517DFFFAAFFC200055557DE00A2801554555557FE10007FEABEFFFD57",
INIT_33 => X"E801EFF7AEA8A10002E955FFA2AABFF455500020AA08003DFFFA28028AAAF7D1",
INIT_34 => X"00000000000000000000000000000000000000000000004000BA5D0017410082",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000067FFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(17),        -- Port A data input
DOA(0)   => data_read_a_lo(17),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(17),        -- Port B data input
DOB(0)   => data_read_b_lo(17),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_18_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"69844019080000A21A611406840014122A641074155FC28A2024001001801003",
INIT_01 => X"A643D920034004180005E9E3C90360C0041C0181002001602025800008440084",
INIT_02 => X"B7333980808408103F2000F81FC0FEDEAC2161B0B84D0002188011110C018041",
INIT_03 => X"0405D434003F2C020081587008020561E55116B0290000042B71240C800440F8",
INIT_04 => X"50805AC31007D6125724029216554A9847669903D640EC8E2001002604503004",
INIT_05 => X"07008000E0EA11803850C800010022660C1C0065003C0404002646DC20A02D40",
INIT_06 => X"8560000000022229A60B048048120FF040000000002C44D620F0228454C83810",
INIT_07 => X"058800A001D4033A004904087F9E3901218050018024110D6771C1F90C285682",
INIT_08 => X"F3020A82929A807B3731021400058C020000A9729400D10100420480202AC214",
INIT_09 => X"C820C802D86184A010180304307008025414204400220202F1A814A0080064C1",
INIT_0A => X"080003C32A10A19090C02010E10229440616900000022E0C6070000504102805",
INIT_0B => X"026226495446E2110AE44174112840880000060D7030C30B885200D274004008",
INIT_0C => X"840018400184001840018400184000C2000C200200301500C404C001B884B806",
INIT_0D => X"81010108003C000210020460801001FB3650D89888E06CAE1061018500184001",
INIT_0E => X"032007E281F840C00284A17210001060D8306C18360C1380A0260CB980840080",
INIT_0F => X"5D79BBEF8E50B041029075982BF3873041029079982BF39748AA0AC800014804",
INIT_10 => X"EA479BFD7F7F3041029075982BF3E73041029079982BF3F632C5F96D3C11555D",
INIT_11 => X"F96A595405FC7F1CFEBC7586C4100A53162B47FD7E39FFEECE1598702345156A",
INIT_12 => X"006FE037ACFB88083A99E06271BB0CA207DFDD5920057E0B001B0EBCC79932C5",
INIT_13 => X"5CA2A002DD51B6F7FC4A411D1E8D44517F14EAFE36E55150016EA8DB73E39464",
INIT_14 => X"953C30351452A13D55CFFA76E928E3891F148B30399F5FB7F28C800DFA06F5DF",
INIT_15 => X"5AC57DFEAEF1005475F1D1F608819CF0EE76E12C824ADD9089715F25FAF9DB84",
INIT_16 => X"0D834041A41A0000010180C02801680460FC900052FA10DC0006DA4881C11015",
INIT_17 => X"D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D836",
INIT_18 => X"8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360",
INIT_19 => X"00000000000000000000020D8360D8360D8360D8360D8360D8360D8360D8360D",
INIT_1A => X"8A28A28A2891182C8A82E0820825945DF675C0770B9E11807E54587BEF8B0000",
INIT_1B => X"44A2552A954AA5128944AAAA28A28A28AAAAAAA28A28A28AAAAAAA28A28A28A2",
INIT_1C => X"F80000128944A25128944A25128944A25128944A25128944A25128944A251289",
INIT_1D => X"BA5D04174AA0000000000000000000000000000000000000000000000000401F",
INIT_1E => X"FFFF7FBFDF55A28402000F7D56ABFF55043FFFFFFFFFFFFFFFFFFFFEFF7AE954",
INIT_1F => X"FE0055043FFFFFFFFFDFEFA2D56AB45AA8400145AA801741000043FFFFFFFFFF",
INIT_20 => X"FFFFFFF80021EF0855421EF00043FFFFF7FBE8B45AAD568BFFFFAA975FF00003",
INIT_21 => X"568B45000002010552EBDF45A28028A00F7843FEBA55557FFEFA2D168B55AAFB",
INIT_22 => X"8428AAA007BC2145F7D5400000004020AA5D2A82155F7AEBFEBAFFD56AA00A2D",
INIT_23 => X"82E954BA0004174AAAA8428B45082ABFEBAA2FFC00000804154AA5D00001EFF7",
INIT_24 => X"000000000002E800105D2A95410002A95410AAAEBFF55AAFFC00BAF7AE800100",
INIT_25 => X"FFFFBFDFEFFFAE954AA550415492140000000000000000000000000000000000",
INIT_26 => X"10140A3FFFFFFFFFDFEFE3F5FAF45AA8000038F7DB6FBD7490E3FFFFFFFFFFFF",
INIT_27 => X"BFFF7AA955C71C043FE1049043FFEFE3F1F8FD7AAD16FB6DBE8E00155BE80154",
INIT_28 => X"8FC7AAD56FB6DBEF1FAFD7E384001EF145B471C7140438FC7E3F1EAB55B6DF6D",
INIT_29 => X"BDE92FFD56FA28B6DF68B551C0E050384124BFF7DB68A28A38F7803DE82495B7",
INIT_2A => X"012482550E021C7EB8028A821C7BC516DFFD1420381C0A02082492A85155E3A4",
INIT_2B => X"F5C70BAFFAE870280024904BA1400174AABE8E28B7D1420BDEAAA2F1C7038140",
INIT_2C => X"00000000000000000000000000002A85000492495428082E95400AAA0BDF7DB6",
INIT_2D => X"002ABFFFFFFFFFFFEFF7FBFDFFFF7AA974BA5504154105500000000000000000",
INIT_2E => X"FF7AA82155F78015400552ABFFEFF7FBFDFFFAAD168B55AA80000BAF7FFFDF55",
INIT_2F => X"55AAD168B55F7FFFDFEFFFAA9555555003DE0000043DFEFA2D56AB45AAD57DFE",
INIT_30 => X"AAAF7843FE10007FEAB55A2D17FFEFFFD568B55A280021EF557FD7555550428B",
INIT_31 => X"2000002A95545A2843FE00F7D17FEAAF7FBEAB45552E954BA08003DFFFFFAAA8",
INIT_32 => X"3DEAAA2D5554BA5504000105D2A80145AA842AA00557BD75EFF7D1400AA5D2A8",
INIT_33 => X"E95410AA843FFFFF7D5554BAF7AE974BA0004020AA5D04154BAF7AEA8BEF5500",
INIT_34 => X"0000000000000000000000000000000000000000000002E974000800154AA002",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000020000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(18),        -- Port A data input
DOA(0)   => data_read_a_lo(18),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(18),        -- Port B data input
DOB(0)   => data_read_b_lo(18),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_19_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"042200000000000041088001001AA00000000000000000000000500802000003",
INIT_01 => X"200048000024000000000404000000000A22000800000800004A200000000001",
INIT_02 => X"032210008DEF00400060000001C008002489E0F0004037B00010101010000000",
INIT_03 => X"0000008128000000000000000000000024001620280000000000354200004008",
INIT_04 => X"000058800004C4024024001210001054B1C822009640000E2000002604003000",
INIT_05 => X"07008000E0200000000000000000200604000000001C04000026400000002C40",
INIT_06 => X"000000000000000100000000000001B040000000002C42010010200004C83810",
INIT_07 => X"0E0050A040041593104004500480090080A01120220140020420401800000000",
INIT_08 => X"130E409080188000021A0000100004082A140102B4020109801A4CE003710010",
INIT_09 => X"C80000005861840000000004301000B000000000001C1C0000000000000020C0",
INIT_0A => X"000002C30000000040500010301020400000000000022A040000000000000004",
INIT_0B => X"00000020001000022000000000000000000002F0001F00002024B20002000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"00108000EC000000000000000010004B20000000000000000000000000000000",
INIT_0E => X"0000006280180040000000000000000000000000000000000000000000000000",
INIT_0F => X"8084451B81A70AB3006BA0011400760AB3006BA0011400680F02096834820000",
INIT_10 => X"11204082248A0AB3006BA0011400160AB3006BA0011400084C780687DBA82800",
INIT_11 => X"068796E80A00802301BC0A7531EDD98E73B02800804620D030F873EB49F30B80",
INIT_12 => X"6B00000002044F091A860700FF9198AA115D5DA37F7A80C8A3604001C0664C78",
INIT_13 => X"98551AC9000000000314E01F9F30198600631448410A2A8D64800000081B0A93",
INIT_14 => X"2E00303842281C80A23004411AD661891F15148A4420804241526D6000000000",
INIT_15 => X"9D335F3D282000C6C5456C84850F61050C411AD6284FDA861682805A04A1046B",
INIT_16 => X"00000000000000000000000000000004600C0013800003088004202304366A4A",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"86186186186851046260A9A69A6039045DD1F863808633005010063A20C90000",
INIT_1B => X"D26930984C26130984C261861861869A61861861861869A61861861861861861",
INIT_1C => X"F800000984C26130984C26130984C26130984C26130984C26130984C26130984",
INIT_1D => X"BA5500020BA5D00000000000000000000000000000000000000000000000401F",
INIT_1E => X"FFFFFFFFFFEFF7AE954BA5D04174AA007BFFFFFFFFFFFFFFFFFFFFFFFFFAA954",
INIT_1F => X"ABFF557BFFFFFFFFFFFFFFFFFBFDFEFFFAA974BA5D517FFFF08043FFFFFFFFFF",
INIT_20 => X"6AB45AA8002000F7D5575455D043FFFFFFFFFFFFFF7FBFDF55A28402000F7D56",
INIT_21 => X"43FFFFFFFFFDFEFA2D56AB45AA8400145AA8017410007BFFFFFFFFFFFFEFF7D1",
INIT_22 => X"AA975FF00003FE00557BFFFFFFFFBFDF45AAD568B55F7AE955FFAA8402010080",
INIT_23 => X"7D168B55AAD17FFEFF7AE975FF00557FFFF5D043FFFFF7FBE8B45AAD568BFFFF",
INIT_24 => X"00000000000557FFEFA2D168B55AAFBFFFFFFF80021EF0855421EF002ABFFEFF",
INIT_25 => X"FFFFFFFFFFF7AA954BA550000082550000000000000000000000000000000000",
INIT_26 => X"C7080E3FFFFFFFFFFFFFFFFBFDFEFFFAE954AA5504154921471FFFFFFFFFFFFF",
INIT_27 => X"F45AA8000038F7DB6FBD74975FFFFFFFFFFFFEFF7FBFAFD7E3A4954BA555B7AF",
INIT_28 => X"FFFFF7FBF8FC7EBD568B55A28000000FFDF52545550A3FFFFFFFFFDFEFE3F5FA",
INIT_29 => X"955C7BE800000008043FFEFE3F1F8FD7AAD16FB6DBE8E00155BE8015410147FF",
INIT_2A => X"1EAB55B6DF6DBFFF7AA955C71C043FE10497BFDFC7E3F1FAF55A2DB6FB7DF7AE",
INIT_2B => X"5B471C71424B8FC7E3D56AB6DB6DF7AFC7EBA0955FF145B7AFC7410438FC7E3F",
INIT_2C => X"00000000000000000000000000005B78FC7AAD56FB6DBEF1FAFD7E384001EF14",
INIT_2D => X"55517FFFFFFFFFFFFFFFFFFFFEFF7AA974AA5500020005500000000000000000",
INIT_2E => X"5AA80154AA557BEAB45002ABFFFFFFFFFFFEFF7FBFDFFFF7AA974BA550415410",
INIT_2F => X"EFF7FBFDFFFAAD168B55AA80000BAF7FFFDF5500517FFFFFFFBFDFEFFFFFEAB4",
INIT_30 => X"155F78015400557BFDFEFF7FBEAB55A2D56AB55A28002000F7FFC2155552ABFF",
INIT_31 => X"8B45AAFBFFFFFFFAA95545F7840201000043DFEFA2D56AB45AAD57DFEFF7AA82",
INIT_32 => X"E8B55000428B55AAD168B55F7FFFDFEFFFAA9555555003DE00007FFDF45AAD56",
INIT_33 => X"568B55A280021EF557FD755555042AB55AAD16ABFFFFFBEAB45A280155EF557F",
INIT_34 => X"0000000000000000000000000000000000000000000007FEAB55A2D17FFEFFFD",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000040000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(19),        -- Port A data input
DOA(0)   => data_read_a_lo(19),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(19),        -- Port B data input
DOB(0)   => data_read_b_lo(19),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_20_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000003",
INIT_01 => X"A75FF80000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"14088080800008400F655001FFCFF80018FA8044000000000000011000000007",
INIT_03 => X"0000000000000000000000000000000024001660380000000000000000004FF8",
INIT_04 => X"000079800014CC02C034001600000000000000101EC0012EE0C0026E1E80F000",
INIT_05 => X"1F0FF433EFF0440C3902100002203F2EFC040388137C3E20C8EEC00284033CC0",
INIT_06 => X"00F00100002E22EB440012C809B2FFF7C8E8840155FDC0000010E40087D8787A",
INIT_07 => X"03B800000000000000008407FC800B0000000100600040000C205FF91C000F80",
INIT_08 => X"F28C0B0300020852000002101554021F00000000000000009049226020000200",
INIT_09 => X"D80000007BEFBC010002008FF7F00000000010018A81000041C401000004FFDF",
INIT_0A => X"00000ADF000000200000008000008028300100461003EAFE400000120000913F",
INIT_0B => X"0000000000000000000000000200200290000000000000000200000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000010001000000",
INIT_0D => X"00000100000010000002000080101FFB60000000000000000000000000000000",
INIT_0E => X"03007FE29FF800C00000001002040000000000000020480002E42429C0000080",
INIT_0F => X"0004D4E180010040000400000001E60040000400000001E6010003C000000000",
INIT_10 => X"000000094B1E0040000400000001E60040000400000001E60804000000400000",
INIT_11 => X"00002000000000033628000100100000004000000006170C0008001000004000",
INIT_12 => X"000000000295810000000A100020614148002000000000004307CC3CC0000804",
INIT_13 => X"5802000000000014AC000120200000000003F0D800020100000000000A4B0020",
INIT_14 => X"0020C0C00000000002E2D000001006204040000000005786C004000000000052",
INIT_15 => X"0100A0C0939BEE1810080200000E0CE0EC000010020000000000000AE8A00002",
INIT_16 => X"2008040400400C08080000000000049F6FFC0100000000000008008008000400",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0100000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0C30C30C320624C1090D0F3CF3CD038001801C10000804482A60D09008269020",
INIT_1B => X"90C86432190C86432190CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2C30C3",
INIT_1C => X"F80000432190C86432190C86432190C86432190C86432190C86432190C864321",
INIT_1D => X"AA5504020100800000000000000000000000000000000000000000000000401F",
INIT_1E => X"FFFFFFFFFFFFFFAA954BA5500020BA5D7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974",
INIT_1F => X"74AA00003FFFFFFFFFFFFFFFFFFFFFFF7AA974AA550002000007BFFFFFFFFFFF",
INIT_20 => X"FDFEFFFAE974AA5D003FE005D043FFFFFFFFFFFFFFFFFFFFEFF7AE954BA5D041",
INIT_21 => X"BFFFFFFFFFFFFFFFFFBFDFEFFFAA974BA5D517FFFF087FFFFFFFFFFFFFFFFFFF",
INIT_22 => X"8402000F7D56ABFF55003FFFFFFFFFFFFFF7FBFDFFFAA84000105D556AB55557",
INIT_23 => X"FFFFFFEFF7FBEAB55A28000010F7D16ABEF08043FFFFFFFFFFFFFF7FBFDF55A2",
INIT_24 => X"000000000007BFFFFFFFFFFFFEFF7D16AB45AA8002000F7D5575455D2EBFFFFF",
INIT_25 => X"FFFFFFFFFFFFAE974AA550400028000000000000000000000000000000000000",
INIT_26 => X"380071FFFFFFFFFFFFFFFFFFFFFFFF7AA954BA550000082557FFFFFFFFFFFFFF",
INIT_27 => X"FEFFFAE954AA55041549214043FFFFFFFFFFFFFFFFFFDFEFF7AE974BA5500050",
INIT_28 => X"FFFFFFFFFFFFFF7FBFDFFFFFAA974BA550038E285D0E3FFFFFFFFFFFFFFFFBFD",
INIT_29 => X"02028555F6FB7D5D75FFFFFFFFFFFFEFF7FBFAFD7E3A4954BA555B7AFC70871F",
INIT_2A => X"FFDFEFE3F5FAF45AA8000038F7DB6FBD7490E3FFFFFFFFFDFEFF7F1FAFC7A280",
INIT_2B => X"DF525455524BFFFFFFFBFDFC7E3F5E8B45A28402010FFDB6ABEF140A3FFFFFFF",
INIT_2C => X"00000000000000000000000000007FFFFFFF7FBF8FC7EBD568B55A28000000FF",
INIT_2D => X"557FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5504000BA0800000000000000000",
INIT_2E => X"FFFAE954BA5500174AA08517FFFFFFFFFFFFFFFFFFFFEFF7AA974AA550002000",
INIT_2F => X"FFFFFFFFFEFF7FBFDFFFF7AA974BA55041541055043FFFFFFFFFFFFFF7FBFDFE",
INIT_30 => X"4AA557BEAB4500557FFFFFFFFFDFEFF7FFFFFEFF7AE974AA550028AAA5D2ABFF",
INIT_31 => X"DFEFFFD568B55A284020BA557FFFFFF5D517FFFFFFFBFDFEFFFFFEAB45AA8015",
INIT_32 => X"EABEF5D2ABFFEFF7FBFDFFFAAD168B55AA80000BAF7FFFDF55002EBFFFFF7FBF",
INIT_33 => X"56AB55A28002000F7FFC215555043DFEFF7FBFFF55A2D16AB45AA8402000F7FB",
INIT_34 => X"0000000000000000000000000000000000000000000007BFDFEFF7FBEAB55A2D",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000007FFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(20),        -- Port A data input
DOA(0)   => data_read_a_lo(20),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(20),        -- Port B data input
DOB(0)   => data_read_b_lo(20),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_21_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"4A302428B824900A128C090A5C1800261500213C005FE812D10420054085A202",
INIT_01 => X"081FFE3440B609703B0427F801A40B8115BC4F655300340288A40D30040E4DD8",
INIT_02 => X"0109095C30C98809800000F9FFFFFFFF149FF1FCA4C0421B182E3490DF145FE4",
INIT_03 => X"084A76341244919000099486400026523C041660BA000100CC12701015007FF8",
INIT_04 => X"000079800014CC03C075161E001118653D2408041FC004AEF000816E1C11F541",
INIT_05 => X"3F0F807BFFE000240100004683103E7FFE02482553FC3C0204EFC25010143CC0",
INIT_06 => X"008808210996035A000006EC2E04FFFFC0A0000101FFE4036450E08247F87870",
INIT_07 => X"4003400812A156C002822987FC830F40134CC74D002016612DE87FFE00400804",
INIT_08 => X"F02348D2D00080C0C53400044114000000D022640B42406808790055043A8282",
INIT_09 => X"F84056387FEFBC110008420F7FF388B70A20389346FE9F26120200800008FDFF",
INIT_0A => X"4518DBFF00020004C0A6044901112A0908AA14601DE3EBFE0A812D8D5B742D3F",
INIT_0B => X"104032901CC63410ABD249C4B3007127080806FF917FC30010107688862A28C5",
INIT_0C => X"46C9146C9146C9146C9146C9146CC8A3648A3642003184822040D000D8C41807",
INIT_0D => X"201800500941044312000900D4621FFBE0008A94C822CA8919018206C9146C91",
INIT_0E => X"2029FFEADFF8050250010030165290008800440022201082401A002000C48000",
INIT_0F => X"18048A004A6C0D2820302C005A83480D1820302A009B02B101390C0CB2830816",
INIT_10 => X"1408904831400D1820302C005A83480D2820302A009B02B021A85C0941150013",
INIT_11 => X"5C08834600024D052C1051E0B92D400360520202682C19024B6164E300448510",
INIT_12 => X"6404093E22A2012418A9D1D44ADD9E0F174103820101C0B8160D5516259FA1A8",
INIT_13 => X"60D8AA288209E615100280DA0052000C5006402000206C55144104D510CC1B0D",
INIT_14 => X"0A0D50020C04023033C52009144231D902818100C90058010361AC808126C886",
INIT_15 => X"2202386454988140600C0181500A13E830011008B0374007000B4E0CD0002450",
INIT_16 => X"0080224004002000000703804008001F7FFF01B982B01258088C008CC41198A1",
INIT_17 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_18 => X"8020080200802008020080200802008020080200802008020080200802008020",
INIT_19 => X"0000000000000000000002008020080200802008020080200802008020080200",
INIT_1A => X"BEFBEFBEFBFF7FEFEFFFE79E79FFFF7CFF77FBFFEFBFF9F7E0FDF9EFEFBF0000",
INIT_1B => X"DFEFF7FBFDFEFF7FBFDFEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEF",
INIT_1C => X"F80000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"BA5D00020000800000000000000000000000000000000000000000000000401F",
INIT_1E => X"FFFFFFFFFFFFFFAE974AA550402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974",
INIT_1F => X"20BA5D7FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5D00020AA5D7FFFFFFFFFFFF",
INIT_20 => X"FFFFFF7AA974BA5D0402000557BFFFFFFFFFFFFFFFFFFFFFFFFFAA954BA55000",
INIT_21 => X"03FFFFFFFFFFFFFFFFFFFFFFF7AA974AA55000200000003FFFFFFFFFFFFFFFFF",
INIT_22 => X"AE954BA5D04174AA00003FFFFFFFFFFFFFFFFFFFFEFF7AE974BA5D00174BA000",
INIT_23 => X"FFFFFFFFFFFFFDFEFF7AE954AA5500174BA5D043FFFFFFFFFFFFFFFFFFFFEFF7",
INIT_24 => X"000000000007FFFFFFFFFFFFFFFFFFFFDFEFFFAE974AA5D003FE005D2EBFFFFF",
INIT_25 => X"FFFFFFFFFFFFAE974BA5D0000010000000000000000000000000000000000000",
INIT_26 => X"BA557FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550400028007FFFFFFFFFFFFFF",
INIT_27 => X"FFFF7AA954BA550000082557BFFFFFFFFFFFFFFFFFFFFFFFFFAA954BA5D00000",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFEFF7AA974AA5D04050005571FFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"954BA5D00154AA00043FFFFFFFFFFFFFFFFFFDFEFF7AE974BA55000503800003",
INIT_2A => X"FFFFFFFFFBFDFEFFFAE954AA550415492140E3FFFFFFFFFFFFFFFFFFDFEFF7AE",
INIT_2B => X"0038E285D2ABFFFFFFFFFFFFFFFFBFDFEFFFAA974BA5D00104925D0E3FFFFFFF",
INIT_2C => X"000000000000000000000000000071FFFFFFFFFFFFFFF7FBFDFFFFFAA974BA55",
INIT_2D => X"087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D00000100000000000000000000",
INIT_2E => X"FF7AA954BA5D00000BA5D7FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5504000BA",
INIT_2F => X"FFFFFFFFFFFFFFFFFFEFF7AA974AA550002000557BFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA5500174AA08043FFFFFFFFFFFFFFFFBFDFEFF7AE954AA5D041740055517FF",
INIT_31 => X"FFFFF7FBFDFFFFFAA974AA5D00174BA08043FFFFFFFFFFFFFF7FBFDFEFFFAE95",
INIT_32 => X"00010552ABFFFFFFFFFFFEFF7FBFDFFFF7AA974BA550415410552ABFFFFFFFFF",
INIT_33 => X"FFFFEFF7AE974AA550028AAA5D2EBFFFFFFFFFDFEFF7FBFFFFFF7AE954BA5D00",
INIT_34 => X"000000000000000000000000000000000000000000000557FFFFFFFFFDFEFF7F",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(21),        -- Port A data input
DOA(0)   => data_read_a_lo(21),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(21),        -- Port B data input
DOB(0)   => data_read_b_lo(21),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_22_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"5290F4CDE914905A14A43D33F488243E17122300F55FEB189B343A1140548380",
INIT_01 => X"A94007B259F6A975386262000C344BA9573C6FF57B18A5FB0ABFCD3C2C5F4F0C",
INIT_02 => X"877FE30EB378008D202551040030071869D0040180AC4B685F6E26FAA0810006",
INIT_03 => X"431965109E4481D6B5AAD6875AD6AB5A1815600802888808DEA83552954D3000",
INIT_04 => X"492C0020220001010E4916C884DCD607E5EC2A344103E48003D0800023D0072C",
INIT_05 => X"00107C441001100D620A06D683018001023D37E5088043620101179092540112",
INIT_06 => X"40111C2D50A46AE45281502E4A2200081ADA0E054402365774611E047020008E",
INIT_07 => X"680BD5AA4BF5C91F840C1710010344DB9A808FDFF3DE0313014A200754040180",
INIT_08 => X"0EA212D6D481ADF0CE47CA21544009007A64EBD64049D028B93D9561A48F6027",
INIT_09 => X"207246A80400015805060040080A2A0F4A82381B4000BFB65A0283800AA50020",
INIT_0A => X"4539C020E11810098D4067EFF9FF284D483E35602820110204804818CD280100",
INIT_0B => X"10081E9528963546278008AA800470370000A0004D0000002126F30C902A29C5",
INIT_0C => X"40E1540E1540E1540E1540E1540E4AA070AA07000A0000308000190168200281",
INIT_0D => X"6870A9CA0D458D131652A154D46B600085080B14009A2B2906504940E1540E15",
INIT_0E => X"448C00044000A1EC1C44140D101A54280A14050A028500A84F02842A24C594A0",
INIT_0F => X"38359E0C4E6C256690581800F1C3E82562B0581200F1C3F08145602280402080",
INIT_10 => X"100AB8581B602562B0581800F1C3E8256690581200F1C3F1238473F121000613",
INIT_11 => X"73F0E1050083750B3E4275F829547008600C030374361FA2CEE046D48122C438",
INIT_12 => X"C4CC012A66F61154C019511628756231018500C00203E1380615651607822384",
INIT_13 => X"608AA612C0096C37B00D1724801A0009C606D1221D104553096004B61BCC1128",
INIT_14 => X"12A41E0F0600035842E7601C2C4AC68A98810080AA825A890225189980254CDE",
INIT_15 => X"A89637E00D0A1080301401C390320188321C2C0B13890105800D520AF94870B0",
INIT_16 => X"88222F110111B281A54753AA004002601001918008C10912A4440B24E8B58234",
INIT_17 => X"8220882208822088220882208822088220882208822088220882208822088220",
INIT_18 => X"2008020080200802008020080200802008020080200802208822088220882208",
INIT_19 => X"1448000000001FFFFFFFFC802008020080200802008020080200802008020080",
INIT_1A => X"9E79E79E7BFF3FEFEBEEEFBEFBEFBEFDFEF7F47F8FBEF5EB7E6CFEFBEFBE8289",
INIT_1B => X"CFE7F3F9FCFE7F3F9FCFE79E79E79E79E79E79E79E79E79E79E79E79E79E79E7",
INIT_1C => X"F800003F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9F",
INIT_1D => X"BA5D04000000000000000000000000000000000000000000000000000000401F",
INIT_1E => X"FFFFFFFFFFFFFFAE974BA5D0002000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974",
INIT_1F => X"2010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA550000010007FFFFFFFFFFFF",
INIT_20 => X"FFFFFFFAE954AA5D00000AA007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA55040",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5D00020AA5D7FFFFFFFFFFFFFFFFFFF",
INIT_22 => X"AA954BA5500020BA5D7FFFFFFFFFFFFFFFFFFFFFFFFFFAA954BA5504000AA557",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFAA954BA5500000BA5D7BFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"00000000000003FFFFFFFFFFFFFFFFFFFFFFF7AA974BA5D040200055517FFFFF",
INIT_25 => X"FFFFFFFFFFFFAE974BA5D0402000080000000000000000000000000000000000",
INIT_26 => X"10087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0000010007FFFFFFFFFFFFFF",
INIT_27 => X"FFFFFAE974AA550400028007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA5500020",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFAE954AA5D00020BA087FFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"954BA5504020AA5D7BFFFFFFFFFFFFFFFFFFFFFFFFFAA954BA5D00000BA557FF",
INIT_2A => X"FFFFFFFFFFFFFFFF7AA954BA5500000825571FFFFFFFFFFFFFFFFFFFFFFFFFAA",
INIT_2B => X"040500055517FFFFFFFFFFFFFFFFFFFFFFF7AA974AA5D00070925D71FFFFFFFF",
INIT_2C => X"0000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFEFF7AA974AA5D",
INIT_2D => X"007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020000800000000000000000",
INIT_2E => X"FFFAE974AA550002000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0000010",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFAE954AA5504000BA087FFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA5D00000BA5D7BFFFFFFFFFFFFFFFFFFFFFFFFFAA954AA5D00020AA007FFFF",
INIT_31 => X"FFFFFFFFFFFEFF7AA974BA5504020BA557BFFFFFFFFFFFFFFFFFFFFFFFF7AA95",
INIT_32 => X"154105D517FFFFFFFFFFFFFFFFFFFFEFF7AA974AA55000200055517FFFFFFFFF",
INIT_33 => X"BFDFEFF7AE954AA5D041740055557FFFFFFFFFFFFFFFFFFDFEFF7AE974AA5D00",
INIT_34 => X"000000000000000000000000000000000000000000000043FFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000007FFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(22),        -- Port A data input
DOA(0)   => data_read_a_lo(22),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(22),        -- Port B data input
DOB(0)   => data_read_b_lo(22),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_23_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"EF20906D902424807BC8241BC81801B97D38AD3C0800103362A6741C80A12A02",
INIT_01 => X"001FFF8409F089003B4422000D80C80106804A7951C5B9D1C828043EA28838F9",
INIT_02 => X"073B8858218C2C50801000F9FFEFF8E72CA7F5FC2E048026496834D84721DFE0",
INIT_03 => X"2C4360101A4001001005080400401420350016E0BB222341C312000014006FF8",
INIT_04 => X"00017B810015DC03D034201E14000036486008101FC0002EE006297E1C05F561",
INIT_05 => X"BF0F817FFFE80100004044800080BEFFFC0248005FFC3C18A5FFC2444484BCC0",
INIT_06 => X"0400000409120338860900482404FFFFC000000001FFC0832050E00047F97870",
INIT_07 => X"200246801C41C3E81E872C8FFE900FC31348EFDF03BE15E22DA07FF92C204102",
INIT_08 => X"F6220280D2B025988311AB14155421006891A1089F6E200000022C140068EB90",
INIT_09 => X"F8001011FFEFBC80000000077FF184B03010004002FE000000201000000FFDFF",
INIT_0A => X"00001BFFA800808189A657EF81DD0C00079CD00837C3EBFD4201258112D4487F",
INIT_0B => X"24483890564084198AD249C433200180082A06FF907FC3081812048006000000",
INIT_0C => X"8608086080860808608086080860804304043042003184822150C000D8C41806",
INIT_0D => X"03000100200180480000095280001FFBF040C088CD20E0A21921828608086080",
INIT_0E => X"3821FFEAFFF805025E00853B92588000400020001000020A8018008002000014",
INIT_0F => X"486148484054395E27E428002A4200397E07E422002A420100382FCC30832A16",
INIT_10 => X"0C0788417000397E07E428002A4200395E27E422002A420110A51C01C0590401",
INIT_11 => X"1C01A2490040590C08120558C1759BE1C05A0400383808800DA1929F72864110",
INIT_12 => X"20000136006000215EA0A4833A32C8832050028603050014031B3950000C90A5",
INIT_13 => X"006658280009A2030108B14AC05C00112405222088B8332C140004D101800CE7",
INIT_14 => X"196B6808060201281004228996085F10020180C030880D11019CE4000026C00C",
INIT_15 => X"52A49DC7143F01C04240030720641E0A028996483A17204680410A04104A2659",
INIT_16 => X"0401000080080000000000002001201F7FFC0011C2F81A48080CA32800A01081",
INIT_17 => X"4010040100401004010040100401004010040100401004010040100401004010",
INIT_18 => X"0100401004010040100401004010040100401004010040100401004010040100",
INIT_19 => X"0000000000000000000000040100401004010040100401004010040100401004",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"F800000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"BA5D04020100000000000000000000000000000000000000000000000000401F",
INIT_1E => X"FFFFFFFFFFFFFFAE974BA5D0400000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974",
INIT_1F => X"2000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400010087FFFFFFFFFFFF",
INIT_20 => X"FFFFFFFAE974BA550002000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D000",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA550000010007FFFFFFFFFFFFFFFFFFF",
INIT_22 => X"AE974AA550402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550400000087",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFAE974AA550402000087FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5D00000AA007FFFFFFF",
INIT_25 => X"FFFFFFFFFFFFAE974BA5D0402010000000000000000000000000000000000000",
INIT_26 => X"10087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000087FFFFFFFFFFFFFF",
INIT_27 => X"FFFFFAE974BA5D0000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04000",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFAE974BA550002000007FFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974AA550400010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550002010087FF",
INIT_2A => X"FFFFFFFFFFFFFFFFFAE974AA550400028007FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_2B => X"00020BA087FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5D0402038007FFFFFFFFF",
INIT_2C => X"00000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5D",
INIT_2D => X"087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020100000000000000000000",
INIT_2E => X"FFFAE974BA5D0400000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D0000010007FFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4AA550002000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA550002010087FFFF",
INIT_31 => X"FFFFFFFFFFFFFFFAE954AA550400010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_32 => X"000AA087FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5504000BA087FFFFFFFFFFF",
INIT_33 => X"FFFFFFFFAA954AA5D00020AA007BFFFFFFFFFFFFFFFFFFFFFFFFFAA954AA5D04",
INIT_34 => X"0000000000000000000000000000000000000000000007BFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000007FFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(23),        -- Port A data input
DOA(0)   => data_read_a_lo(23),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(23),        -- Port B data input
DOB(0)   => data_read_b_lo(23),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_24_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100600007FFF000080108004000800020000840041000080808",
INIT_02 => X"172A00D000EF8210000000F9FFEFF8E7240FF1FC224087B1000639401D005FC0",
INIT_03 => X"00003A2E200811000000000400000000340016603A0000004860400014006FFF",
INIT_04 => X"000079800014CC03C034001E04010850300000101FC0002EE000006E1C00F500",
INIT_05 => X"1F0F8033FFE000000000000000003E2FFC024800137C3C0000EFC00000003CC0",
INIT_06 => X"0000000009120110020100002404FFFFC000000001FFC0000010E00007F87870",
INIT_07 => X"200102050840950002802C87FC800FCAA035400001B918600C207FF800000000",
INIT_08 => X"F6234AD280B02500063AC2840001610020408178B600C2400013649608730004",
INIT_09 => X"F80000007FEFBC00000000077FF000B00000000002FE0000000000000000FDFF",
INIT_0A => X"00001BFFA0000005501AA00000CE20000094000011C3EBFC020125811254083F",
INIT_0B => X"0040A040004000008012414433000100080806FD107FC3000000000006000000",
INIT_0C => X"0608006080060800608006080060800304003042003180822040C00090C41806",
INIT_0D => X"004800B0000000000000000000001FFBE0008080C820C0801801800608006080",
INIT_0E => X"2021FFEADFF80002080000000208800000000000000000020018000000000000",
INIT_0F => X"840009181008024A00043601100210024A00043C0110020901382CCCB28B0806",
INIT_10 => X"180040A03080024A00043601100210024A00043C01100209240C840C201D0210",
INIT_11 => X"840A604E0080820009908008341B000A8212070082002890010068320860C920",
INIT_12 => X"40600800082041205EC00044C1ACB66C37542082030281E0580001012811A40C",
INIT_13 => X"80B27A004300004103160DB3005E000618040C022000593D002180002090166B",
INIT_14 => X"2BBFF20406040084210C062000C2A2DDD00180C04504086002CD680C01000104",
INIT_15 => X"20804295C98F80400008040CC0582169022000C2876C40478002850016088001",
INIT_16 => X"0000000000000000000000000000001F7FFC001B823018F00880008805241060",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"9EF9EF9EFB263CC3090CABAEBAFF96857757B73E6089966B9EF9D5A220CC8000",
INIT_1B => X"C1E0F0783C1E0F0783C1EFBEFBEFBE79E79E79E79E79EFBEFBEFBEFBEFBEF9EF",
INIT_1C => X"F800000783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783",
INIT_1D => X"BA5D04020100800000000000000000000000000000000000000000000000401F",
INIT_1E => X"FFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974",
INIT_1F => X"0000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000087FFFFFFFFFFFF",
INIT_20 => X"FFFFFFFAE974BA5D0400000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400010087FFFFFFFFFFFFFFFFFFF",
INIT_22 => X"AE974BA5D0002000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0000010007",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFAE974BA5D0002000007FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA550002000007FFFFFFF",
INIT_25 => X"FFFFFFFFFFFFAE974BA5D0402010080000000000000000000000000000000000",
INIT_26 => X"00087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFF",
INIT_27 => X"FFFFFAE974BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000007FFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA5D0000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400010087FF",
INIT_2A => X"FFFFFFFFFFFFFFFFFAE974BA5D0000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_2B => X"0002000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA550002000087FFFFFFFFF",
INIT_2C => X"00000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA55",
INIT_2D => X"007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020100800000000000000000",
INIT_2E => X"FFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA5D0400000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000007FFFF",
INIT_31 => X"FFFFFFFFFFFFFFFAE974BA5D0000010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_32 => X"00010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0000010007FFFFFFFFFFF",
INIT_33 => X"FFFFFFFFAE974BA550002010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5500",
INIT_34 => X"0000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(24),        -- Port A data input
DOA(0)   => data_read_a_lo(24),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(24),        -- Port B data input
DOB(0)   => data_read_b_lo(24),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_25_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100200002000000080100004000000020000800041000080808",
INIT_02 => X"1000218000000800000000F9FFEFF8E738FFF1FC20400400000004455A375FE0",
INIT_03 => X"00002000000001000000000400000000340016623A0000004000000014006FFF",
INIT_04 => X"924279824C94CC1BE0B4001F20000000020380401FE0082EF000106E1C00F500",
INIT_05 => X"1F0F8033FFF048202582800100523E2FFE024820137C3C0040EFE02000003CE4",
INIT_06 => X"10DC00CC0992033A062116E82404FFFFC0E0801101FFC0000010E08A07FC7870",
INIT_07 => X"000000000000000002802C87FC800F8000000000019810600C207FFF3C410D84",
INIT_08 => X"FE8002000080281000008A0000014100200081000000000080480AE000000200",
INIT_09 => X"FC0020007FEFBE031018C31F7FFBAEBC0020008086FE0000100280800000FDFF",
INIT_0A => X"00001BFFE00301000000000000CC02000014000191C3EBFF4A7DF795965C6D3F",
INIT_0B => X"0040200000400000801243443B000100880806FD107FC3018000000006000000",
INIT_0C => X"0608006080060800608006080060800304003042003B99862444E61492C41806",
INIT_0D => X"00000000000000000000001280001FFBE0008080C820C4801801800608006080",
INIT_0E => X"3021FFEADFF805025C0304001E58906088304418222C108A009A090400000000",
INIT_0F => X"00000100100000480000200100000000480000200100000100380F0C30830A06",
INIT_10 => X"0000008000000048000020010000000048000020010000000004040000010000",
INIT_11 => X"0400004000000000008080000011000000020000000020000000001200000100",
INIT_12 => X"000000000800002018C010000020800000800122000000004004000008000004",
INIT_13 => X"0002080000000040000001020020000000000800200001040000000020000021",
INIT_14 => X"0021000008001000000800200000021000020100000000200004200000000100",
INIT_15 => X"0000008400000000605000000000200000200000020400000000000002008000",
INIT_16 => X"288226410410346010000000400A011F7FFE0031823010400800000800001840",
INIT_17 => X"8822088220882208822088220882208822088220882208822088220882208822",
INIT_18 => X"8220882208822088220882208822088220882208822088220882208822088220",
INIT_19 => X"00017FFFFFFFFFFFFFFFFE088220882208822088220882208822088220882208",
INIT_1A => X"2410492410A048029890AD34D35FDD144A50CB5462D14997BE09E760AED04040",
INIT_1B => X"8C46231188C46231188C49249249249249249249249241041041041041041049",
INIT_1C => X"F80000B158AC562B158AC562B158AC562B158AC562B158AC562B158AC562B158",
INIT_1D => X"BA5D040201000000000000000000000000000000000000000000000000007FFF",
INIT_1E => X"FFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974",
INIT_1F => X"2010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFF",
INIT_20 => X"FFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000087FFFFFFFFFFFFFFFFFFF",
INIT_22 => X"AE974BA5D0400000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000007",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFAE974BA5D0400000087FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000007FFFFFFF",
INIT_25 => X"FFFFFFFFFFFFAE974BA5D0402010000000000000000000000000000000000000",
INIT_26 => X"10087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFF",
INIT_27 => X"FFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA5D0402000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000087FF",
INIT_2A => X"FFFFFFFFFFFFFFFFFAE974BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_2B => X"0400000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000087FFFFFFFFF",
INIT_2C => X"00000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D",
INIT_2D => X"087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020100000000000000000000",
INIT_2E => X"FFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFF",
INIT_31 => X"FFFFFFFFFFFFFFFAE974BA5D0402000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_32 => X"02000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000087FFFFFFFFFFF",
INIT_33 => X"FFFFFFFFAE974BA5D0400000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_34 => X"0000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000007FFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(25),        -- Port A data input
DOA(0)   => data_read_a_lo(25),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(25),        -- Port B data input
DOB(0)   => data_read_b_lo(25),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_26_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"E9264EAB20190CA3BA4997AA9002AE9C001006B0778015CFA17E0811039879C7",
INIT_01 => X"F1FFF9BB1F773C7F9BB07DFFFDD863FC5FFF3FEFFBBF9FFB22FFFBC7B9F30686",
INIT_02 => X"1B33188302E708180F6FFBFFFFCFFFFF9C7FF7FC24350B99082400001D00DFD8",
INIT_03 => X"4A53D958C50000DCE7366303739CD98C27C57EF57980014F271807E3C9E9CFF8",
INIT_04 => X"DBFAFBD7FB1CDEBEF1BE17F7AC88042787FBFFF8FEE9FF7EE6F4C0EE1FFAF869",
INIT_05 => X"5F0FFEB3EFFEFFBDA7F7FED508707E2EFEBF6FFEB37C3FF302EEEDFF9B487CF6",
INIT_06 => X"AFBE564C71268F3BBF5FBFC2A427FFF7C3E3A74667FDDB7FB870FF30FFDEF87F",
INIT_07 => X"03BC18306396FBEC14489737FDC00B13BB79DFDB83BF4112AF205FFBDD3AFB93",
INIT_08 => X"F21E4391909B381B0B1F8E041051831FA3068D77E000030021324620C0B9C206",
INIT_09 => X"DE89ECC0FBEFBEBF30B8D79FF7F451F33CFD60FE8FFFDF58003B1D4223B4FFDF",
INIT_0A => X"8ED6BFDF3EB3EBF9DDBCE7FDC1DF8A760F3EB980580BFAFFF37DF7B9DF7DCB3F",
INIT_0B => X"6EE6F5E7FAC4C03DB856CD4CF73AC1FC98884FFF19FFC71FEFED7B251E35768E",
INIT_0C => X"06BC606BC606BC606BC606BC606BD3035E3035C62B7BB987666DEF8A90CCFA8F",
INIT_0D => X"CF6100C0E60FB9FC3A80EF69A04DFFFF7FF5F9A0DC33E9B41D01D207BC606BC6",
INIT_0E => X"7027FFFF9FF8FAFAA3ADEBFB9726BAF5FD7AFEBD7F7EFFD7ACDB7F947F0EA035",
INIT_0F => X"E020080A40403E8BD8002000FC02003E8BD8002000FC02010979AFFE36C36B86",
INIT_10 => X"000EE00034003E8BD8002000FC02003E8BD8002000FC020037B0040A00010003",
INIT_11 => X"040C00400003D80008160400FD81341C00020003B80008C00801EF0285380100",
INIT_12 => X"90981038406809677FA080468C46A81080581002000780C8001C8100201037B0",
INIT_13 => X"00F90D162001C803411FC0024080001F80040026C0807C868B1000E401A01F11",
INIT_14 => X"3F810503A00003E020042AC080CEB01228A80000F600080123E232130407080D",
INIT_15 => X"0087520750001064180807868000110C02C080CFA0042400000F8800105B0201",
INIT_16 => X"7FDFF7EFEEFF3EEC3FF7FBFFBCB7FFFFEFFE00BFF7FEBF420800EC0CBEE61F81",
INIT_17 => X"FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F",
INIT_18 => X"D7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5",
INIT_19 => X"43237FFFFFFFFFFFFFFFFF5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5F",
INIT_1A => X"A69A61861BAF15EAA6AFC38E38EA3AD8ADE7A48F0B366429F434AA9FC376DAE4",
INIT_1B => X"C26130984C26130984C261861861861861861861861861861861861861861869",
INIT_1C => X"F800000984C26130984C26130984C26130984C26130984C26130984C26130984",
INIT_1D => X"BA5D04020100000000000000000000000000000000000000000000000000401F",
INIT_1E => X"FFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974",
INIT_1F => X"2010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFF",
INIT_20 => X"FFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFF",
INIT_22 => X"AE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFF",
INIT_25 => X"FFFFFFFFFFFFAE974BA5D0402010000000000000000000000000000000000000",
INIT_26 => X"10007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFF",
INIT_27 => X"FFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FF",
INIT_2A => X"FFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_2B => X"0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFF",
INIT_2C => X"00000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D",
INIT_2D => X"007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020100000000000000000000",
INIT_2E => X"FFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFF",
INIT_31 => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_32 => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_33 => X"FFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_34 => X"0000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(26),        -- Port A data input
DOA(0)   => data_read_a_lo(26),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(26),        -- Port B data input
DOB(0)   => data_read_b_lo(26),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_27_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"00080A40000A41248002029000050A088000008242A0004404480002000A1155",
INIT_01 => X"F1FFF1C11F781C129C107DFFFE0860941E81258CA2B71C2220EC1B86E1A00002",
INIT_02 => X"4000002100000014400FF6FFFF0FFFFF8007F1FC211100014200800000887FC0",
INIT_03 => X"0842D85841000098C63061026318C18404C459757000015F00088BE3C0618FF8",
INIT_04 => X"DBEAE5D6D91C2EBCE1B21EA72C00000007FBE7C8F8E9EF79E6D440E91FDAE061",
INIT_05 => X"5C8FFCB38FF6B68984B5BCE408347E28FEBF6FEEB3723F7102E8EDBF8A4872F6",
INIT_06 => X"AB98420C71408D113956AFD0842FFFC7C3032646EFF1DB7FA868FE30EF1CE47E",
INIT_07 => X"10041830600640C415004637FC4003021259CFDB01BF80028E001FF8251AB9D1",
INIT_08 => X"F200822020842203000082050000110023068D03000002820000000840000005",
INIT_09 => X"1C852440E3DF7E2FB0B8E717C7F411F3BC6D60B60FFDDE480018AC4AA3B0FD1F",
INIT_0A => X"18109E1F16B16B71092CE7ED81CF403601229880400BE0FC137FF7A0FF75813F",
INIT_0B => X"86F7D5E382A440349816DD4C755AC16C1A884FFE18FFD757E7ED7A211E81C098",
INIT_0C => X"061A2061A2061A2061A2061A2061E1030D1030D6A37FB9872E65E6AA90CD5AAF",
INIT_0D => X"8FC10080A20ED1D41880CC61A044DFFC6EB5BCA0DE31F8B41C01E0071A2061A2",
INIT_0E => X"2023FFE91FF98AEAA1AC6AC9A3A4AAD5B56ADAB56D5AFD572C597B147506203E",
INIT_0F => X"E020000260403C8948002000EC0000BC8948002000EC00010878AC3CB8AB8857",
INIT_10 => X"000EE0000400BC8948002000EC0000BC8948002000EC000097B0040200010003",
INIT_11 => X"040400400003D80000070400DD81041400020003B80000410801AF0204180100",
INIT_12 => X"101010384008086378A080428C46A80080081002000780C800188000301017B0",
INIT_13 => X"02E909042001C800409FC0020080001F80000007C0807484821000E400205D11",
INIT_14 => X"3F810100A00003E020000BC0808EB01020280000F60000002BA2220204070801",
INIT_15 => X"0007520750000024080807868000100403C0808FA0040400000F8800001F0200",
INIT_16 => X"5B5EF3AF6AF6389C2FE128971AB2DDDF8FFE0031B776BF4208006C0C92621F81",
INIT_17 => X"B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D",
INIT_18 => X"56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5",
INIT_19 => X"43A3FFFFFFFFFFFFFFFFFD5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B",
INIT_1A => X"0000000001E0080397908000000A48710B4080240E543021B438A010825238B4",
INIT_1B => X"0804020100804020100800000000000000000000000000000000000000008200",
INIT_1C => X"F80000A05028140A05028140A05028140A05028140A05028140A05028140A050",
INIT_1D => X"BA5D04020100000000000000000000000000000000000000000000000000401F",
INIT_1E => X"FFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974",
INIT_1F => X"2010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFF",
INIT_20 => X"FFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFF",
INIT_22 => X"AE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFF",
INIT_25 => X"FFFFFFFFFFFFAE974BA5D0402010000000000000000000000000000000000000",
INIT_26 => X"10007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFF",
INIT_27 => X"FFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FF",
INIT_2A => X"FFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_2B => X"0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFF",
INIT_2C => X"00000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D",
INIT_2D => X"007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020100000000000000000000",
INIT_2E => X"FFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_31 => X"FFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_32 => X"02010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFF",
INIT_33 => X"FFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_34 => X"0000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000007FFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(27),        -- Port A data input
DOA(0)   => data_read_a_lo(27),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(27),        -- Port B data input
DOB(0)   => data_read_b_lo(27),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_28_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"02200AA400180030808802A900002A08001280A08A801044104A1000001818C3",
INIT_01 => X"50A00011460214428114180000882214413D0A71592A01D92213D28005210202",
INIT_02 => X"1444428102100884000AA30200000000C1000401041108404400022220800000",
INIT_03 => X"461080404900000C6314A900318C52A40051081000888806108802A141288001",
INIT_04 => X"00800040110102000902002000888400081045A8A00003C00000500000080008",
INIT_05 => X"0000000000024CA0A0101800032000400000000B800000014000000B08180000",
INIT_06 => X"814016012000C405280200008001000011110012220009A88800009A88000000",
INIT_07 => X"0004891224228810080010200040001020800000004000008200000240081400",
INIT_08 => X"00A010040401080308400821155540001122448142491008A004912040840221",
INIT_09 => X"0020405000000124058200408000880004440004080160C8100A858009940000",
INIT_0A => X"4D29400002002038104000000020003204000880082800010000000C0000E400",
INIT_0B => X"12220122A000416811040000400800081022C0000080000206CB0821082B694D",
INIT_0C => X"80B0280B0280B0280B0280B0280B01405814058009000421833010800A000200",
INIT_0D => X"C4210040860B188C0A8065302005A004039010280001001600200081B0280B02",
INIT_0E => X"500600010000280000802050010660001000080004004900204020105302A000",
INIT_0F => X"0000000A00000081480000001400000081480000001400000800C01082082210",
INIT_10 => X"0000000024000081480000001400000081480000001400000010000200000000",
INIT_11 => X"0004000000000000001400000080041400000000000000C00000010004180000",
INIT_12 => X"1010100000480802A40000000400000080081000000000000004800000000010",
INIT_13 => X"0001010420000002400040000080000000000024400000808210000001200010",
INIT_14 => X"04000100A0000000000028400004000020280000000000012002020204000009",
INIT_15 => X"0001000000000024080000000000010400400004000004000000000000510000",
INIT_16 => X"0108408420430E699AA42A1508104EA08000000810020000000044001AC20500",
INIT_17 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_18 => X"0040100401004010040100401004010040100401004010040100401004010040",
INIT_19 => X"1708000000000000000000010040100401004010040100401004010040100401",
INIT_1A => X"20820820800D41A8283AC618618EF1088160885001234B96061CCDEC4D205061",
INIT_1B => X"0C06030180C06030180C08208208208208208208208208208208208208208208",
INIT_1C => X"F80000B0582C160B0582C160B0582C160B0582C160B0582C160B0582C160B058",
INIT_1D => X"BA5D04020100000000000000000000000000000000000000000000000000401F",
INIT_1E => X"FFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974",
INIT_1F => X"2010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFF",
INIT_20 => X"FFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFF",
INIT_22 => X"AE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFF",
INIT_25 => X"FFFFFFFFFFFFAE974BA5D0402010000000000000000000000000000000000000",
INIT_26 => X"10007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFF",
INIT_27 => X"FFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FF",
INIT_2A => X"FFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_2B => X"0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFF",
INIT_2C => X"00000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D",
INIT_2D => X"007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020100000000000000000000",
INIT_2E => X"FFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_31 => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_32 => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_33 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_34 => X"0000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000007FFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(28),        -- Port A data input
DOA(0)   => data_read_a_lo(28),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(28),        -- Port B data input
DOB(0)   => data_read_b_lo(28),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_29_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"79964E4BA01DACAB9E659792D00AAE160002829C7FDFEFCEE97C2815039D70C3",
INIT_01 => X"50BFF9AB0775343F9AB01DF80D5821FC0FFF3FEFD1AF9FF1207FFBC7B9720586",
INIT_02 => X"0B33180300E700080F6AAA7BFFC007189C7FF2FC003503980A0000001D00DFD8",
INIT_03 => X"0401D940CD0000C8421A2B03210868AC23403E903900010E271006A148A0C000",
INIT_04 => X"49B87A417315D20A313E17F1800000058013DDF8BE21F36E02F0D06E03E8F800",
INIT_05 => X"1F007E33E01A4D9C87525E5101603E6E023D27DA937C03E340EE25CB9B483C12",
INIT_06 => X"85AA06002026872BAE0B1282A005FFF001E1870223FC3BFC98101F109FC6780F",
INIT_07 => X"03BC081023B233E804488527FDC008019968D74982C94110AF204001BC285A82",
INIT_08 => X"001E4191901A101B031F84000000831FA1028575A000110800124600C039C002",
INIT_09 => X"C60888D0782082B50080508FF00048B124D4005C8AFF4158102914800110FFC0",
INIT_0A => X"8AD6ABC02A02A0B0CCB463B4C0748A720B1EA980100BFA02E204D2154D28AA3F",
INIT_0B => X"6A22B126DA40C03531440800C22800B8900042FF0180000ABFEF89250815568A",
INIT_0C => X"803468034680346803468034680353401A340180010A0801422829800A00A001",
INIT_0D => X"87410080C60AB0F42A804628200DBFFF13D05928040329160520528134680346",
INIT_0E => X"2006FFFF8000F8F80281A16A1504302058102C0816244B82A0CA25907D0AA015",
INIT_0F => X"0000080A40000283D80000001402000283D80000001402010901A7D694494192",
INIT_10 => X"0000000034000283D80000001402000283D80000001402002010000A00000000",
INIT_11 => X"000C000000000000081600002080341C00000000000008C00000410085380000",
INIT_12 => X"90981000006809076B2000040400001080581000000000000004810020002010",
INIT_13 => X"0011051620000003410040004080000000040026C00008828B10000001A00210",
INIT_14 => X"04000503A000000000042AC00044000228A8000000000801204212130400000D",
INIT_15 => X"0081000000001064180000000000010C02C000440000240000000000105B0001",
INIT_16 => X"258964C4A44A0C689FF3F9FFEC5D6DBFE0020096528A0B000000CC043EC60780",
INIT_17 => X"5816058160581605816058160581605816058160581605816058160581605816",
INIT_18 => X"8160581605816058160581605816058160581605816058160581605816058160",
INIT_19 => X"03017FFFFFFFFFFFFFFFFE058160581605816058160581605816058160581605",
INIT_1A => X"AEBAEBAEBFFF7FEFCFDF7FFFFFF5DE7CFCB773FFEFBFF3C7E1E779FFEFFF5060",
INIT_1B => X"FEFF7FBFDFEFF7FBFDFEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEEBAEB",
INIT_1C => X"F80000FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFD",
INIT_1D => X"BA5D04020100000000000000000000000000000000000000000000000000401F",
INIT_1E => X"FFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974",
INIT_1F => X"2010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFF",
INIT_20 => X"FFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFF",
INIT_22 => X"AE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFF",
INIT_25 => X"FFFFFFFFFFFFAE974BA5D0402010000000000000000000000000000000000000",
INIT_26 => X"10007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFF",
INIT_27 => X"FFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FF",
INIT_2A => X"FFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_2B => X"0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFF",
INIT_2C => X"00000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D",
INIT_2D => X"007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020100000000000000000000",
INIT_2E => X"FFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_31 => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_32 => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_33 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_34 => X"0000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(29),        -- Port A data input
DOA(0)   => data_read_a_lo(29),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(29),        -- Port B data input
DOB(0)   => data_read_b_lo(29),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_30_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"9E79E79E7BAF7DEBAFAFEFBEFBFFBFFDFFF7FCFF0FBFFDFF7EFDDFFFEFFE8000",
INIT_1B => X"CFE7F3F9FCFE7F3F9FCFE79E79E79E79E79E79E79E79E79E79E79E79E79E79E7",
INIT_1C => X"F800003F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9F",
INIT_1D => X"BA5D04020100000000000000000000000000000000000000000000000000401F",
INIT_1E => X"FFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974",
INIT_1F => X"2010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFF",
INIT_20 => X"FFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFF",
INIT_22 => X"AE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFF",
INIT_25 => X"FFFFFFFFFFFFAE974BA5D0402010000000000000000000000000000000000000",
INIT_26 => X"10007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFF",
INIT_27 => X"FFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FF",
INIT_2A => X"FFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_2B => X"0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFF",
INIT_2C => X"00000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D",
INIT_2D => X"007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020100000000000000000000",
INIT_2E => X"FFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_31 => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_32 => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_33 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_34 => X"0000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(30),        -- Port A data input
DOA(0)   => data_read_a_lo(30),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(30),        -- Port B data input
DOB(0)   => data_read_b_lo(30),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_31_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"129000008004A00804A40000400800020000000C005FEA005800200400050100",
INIT_01 => X"A15FF18019700810180065FFFC0040801E80258CA2951C2200EC0906A0804140",
INIT_02 => X"0000000000000011000550FDFF0FFFFF0007F1FC200000011000000000205FC0",
INIT_03 => X"08425818000000908428C0024210A30004045060302223490002014280410FF8",
INIT_04 => X"DB6A618248140C18E0B016872400000007EBA24058E1ECA8E2D400681FD0E061",
INIT_05 => X"1C0FFC338FF01009048084C400103E28FE3F6FE513703F7000E8E5B4825030F6",
INIT_06 => X"0098000C51000910100006C00426FFC7C202060445F1F2572060FE82671C607E",
INIT_07 => X"40001020400440C41C000617FC0003021259CFDB01BF00020C001FF804000980",
INIT_08 => X"F200020000802000000082044000010022048902000002000000000000000004",
INIT_09 => X"1C002400E3CF3E0B1118C31747F000B33820209206FC9E80000000000220FD1F",
INIT_0A => X"00001A1F00110101092CE7ED81CF0004012290000023E0FC027DF780DF74013F",
INIT_0B => X"044094C1028400548812494C31004124080886FE187FC301B124F20016000000",
INIT_0C => X"0608006080060800608006080060C00304003042023B99862444E60090C41887",
INIT_0D => X"0B400080200481501000884080405FF864008880CC30E8A01C01C00608006080",
INIT_0E => X"2021FFE81FF880EA000400098200C04080204010200810020C18090424040034",
INIT_0F => X"E020000040403C0800002000E800003C0800002000E8000100780C2C30830806",
INIT_10 => X"000EE00000003C0800002000E800003C0800002000E8000017A0040000010003",
INIT_11 => X"040000400003D80000020400DD01000000020003B80000000801AE0200000100",
INIT_12 => X"000000384000006118A080428846A80000000002000780C800180000201017A0",
INIT_13 => X"00E808000001C800001F80020000001F8000000280807404000000E400001D01",
INIT_14 => X"3B810000000003E020000280808AB01000000000F600000003A0200000070800",
INIT_15 => X"000652075000000000080786800010000280808BA0040000000F8800000A0200",
INIT_16 => X"080223010010308025410082404A015F0FFE003182701B420800280C80201A81",
INIT_17 => X"8020080200802008020080200802008020080200802008020080200802008020",
INIT_18 => X"0200802008020080200802008020080200802008020080200802008020080200",
INIT_19 => X"04017FFFFFFFFFFFFFFFFC080200802008020080200802008020080200802008",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000080",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"F800000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"BA5D04020100000000000000000000000000000000000000000000000000401F",
INIT_1E => X"FFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974",
INIT_1F => X"2010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFF",
INIT_20 => X"FFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFF",
INIT_22 => X"AE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFF",
INIT_25 => X"FFFFFFFFFFFFAE974BA5D0402010000000000000000000000000000000000000",
INIT_26 => X"10007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFF",
INIT_27 => X"FFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FF",
INIT_2A => X"FFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_2B => X"0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFF",
INIT_2C => X"00000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D",
INIT_2D => X"007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020100000000000000000000",
INIT_2E => X"FFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_31 => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_32 => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_33 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_34 => X"0000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(31),        -- Port A data input
DOA(0)   => data_read_a_lo(31),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(31),        -- Port B data input
DOB(0)   => data_read_b_lo(31),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_0_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"ED39BA795990D275FB4A6E96ACC4731DEA4598B0AFB54867F6EE4618C3749803",
INIT_01 => X"58A0047D8607944AC7DA180001ECA2544042106208408208C20022E9173734B3",
INIT_02 => X"9F775E7CB273E6CCA7DAAF00001000000478020113C9C38E09FB7CCCDD9F203E",
INIT_03 => X"441406267B4CB04443163C91110C58F24A31000B8028A810A3D0F8B169A01006",
INIT_04 => X"0005802424830120024121209088809DF81454ACA01E03501D0A3B91E00F0A00",
INIT_05 => X"E0F001CC00012034C20B0232838F80D001C0100AEC83C008EF101A034C8CC300",
INIT_06 => X"582541A028D584E40CB0583CCA0100000161F84322000DA8C40F003C80030780",
INIT_07 => X"2BF70E1C3BBBB1138AF7F888025340C0888430047040FEE182CA00044BC5827C",
INIT_08 => X"0CAFC1F1F07F0FE1C94F65B11555EAFFC1C306758B24197ABCDA467F2C9CF9B3",
INIT_09 => X"027BDA3B0000011420A61080800B6E4C464258094101606E5A47A2A2098B0200",
INIT_0A => X"40198000D1281220444210123820B43B40804CE9AFC800017D82082E2081B6C0",
INIT_0B => X"CA2E0B32B01A752B078412A24844B01302A26900C4801854069B0C888890A081",
INIT_0C => X"C0F33C0F73C0F33C0F73C0F33C0E39E0319E0710A9402011C22908B56A21A020",
INIT_0D => X"8429A95E954868AD0E52273F542580000808061C0389161F027039C1F33C0F73",
INIT_0E => X"5C94001120055704FC4A1624485E2489024481224091282C4300942A19439481",
INIT_0F => X"1C55D65C3E3F01F52FFC1E0013C1F801F52FFC1E0013C1F8090423D38A18E3B1",
INIT_10 => X"1C0118796BE001F567FC1E0013C1F801F567FC1E0013C1F9085DFBF7E15C0610",
INIT_11 => X"FBF7E30F00C0270F3751F1FD00FECBF7E25C0700463E17B2C7F811FD7ADECC38",
INIT_12 => X"6474190626D6491063597F9177B956EF378D33E4030061341F077C571F8F885D",
INIT_13 => X"E207F328E3082636B2807FFD80FE00007E03F7207D3E03F9167184131B5C40FE",
INIT_14 => X"047EFA0CAE06101C53E3647D3F144FCDD22B81C0098E57D9081FCE8C8520C4DA",
INIT_15 => X"FF31ADF08DBF81846A540049707E0FE3307D3F141FFB45478040570EED41F4FE",
INIT_16 => X"902C189601208A1502B4AA5584B4068000019A80098120BCA4C617635C938574",
INIT_17 => X"0240902409024090240902409024090240902409024090240902409024090240",
INIT_18 => X"2409024090240902409024090240902409024090240902409024090240902409",
INIT_19 => X"424A800000000000000000902409024090240902409024090240902409024090",
INIT_1A => X"08208208208831042720EE38E38AAF9C4C704DAB63A6D58B3C10BAE8E789AA09",
INIT_1B => X"0F87C3E1F0F87C3E1F0F82082082082082082082082082082082082082082082",
INIT_1C => X"F800003E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F",
INIT_1D => X"55557BD75EF5D00000000000000000000000000000000000000000000018401F",
INIT_1E => X"FEFA28428B455D0017410A28428AAAA2FBD54BAF7FFD55EF007FD75EFFFAE975",
INIT_1F => X"0145F7AEBFFFF08002AA10A2AABFEAAA2FFC0000AA843FE00AAFBE8B45AA803D",
INIT_20 => X"974AA5D7BFFE000804000BAAAAAAAB45557FFFEBAA2D5401450051401555D7FC",
INIT_21 => X"FD7410557FC21555D51574AAA2FFE8B455D7BD755555517FFEFA280021FF082E",
INIT_22 => X"AEBFE00A2803FEBA002A820AA0800174BA5D2EA8B45005168A10AA8028A10087",
INIT_23 => X"7FFE8B45FFFBC00005D003FF45557FC01FFFFAE95410AA80000005D003FEAAFF",
INIT_24 => X"00000000000557DF5500003DFEFFF84175EFA2AEA8A10000417410A2FFE8BEFF",
INIT_25 => X"F0075D75EFEBAE9554540754717F1F8000000000000000000000000000000000",
INIT_26 => X"47E00A2DB45AA8A3AFD7B68E2AB78550E12555F524AFE38B780154BAFFF1D54A",
INIT_27 => X"1D500002A150038038E285D7F78FD7000B6AB50B6AABDE12BEA0AF010B7D1F8F",
INIT_28 => X"D5C7AA854008700249243A412EBFF5542A43FE9257F1E816D557095EAAA2D140",
INIT_29 => X"EDBC0B680900AAF52B474385D75C502D157545A87AAD178A8002D1D21C5E8257",
INIT_2A => X"F6A150012A2F02AFFDF40E85F475451D502D152A82000E3A5D2150AB8F401471",
INIT_2B => X"51EAFEDB52E3F1EFFFF485A2DA3D5D24BD417FD7E9541242FE920AD082E10A28",
INIT_2C => X"00000000000000000000000000005AAF555080550E87B7A405B52AAD152BD001",
INIT_2D => X"FA69574BAF7D5555AF0D79D55FFA2AC97445057F405458500000000000000000",
INIT_2E => X"0FF16565B2FA9075F4F7B3EBDF50FEAEAAB55F7AEAABFF5D2A81151FB8635A02",
INIT_2F => X"4D5D51F5E08A394003A908B8410E707EF34A08D46F6ABE7082AAAAF2FAC77FE0",
INIT_30 => X"FAE8C798A11A0EAEF75F7AA84001A7052C95256803CE3AEB038662E5D8140601",
INIT_31 => X"A05051023F9A9D57B63BFBF906CB45FABC0954AF0151555AF58794040077D774",
INIT_32 => X"FEE5555BE48AB2A2AE0A0F20C43EAC562245B4E1870108B11020AD4AA05542A0",
INIT_33 => X"D407A97F6F35F498B96BEB12DAAB77558ABD5F5F0DA6BC9525688C1A2A0C06E9",
INIT_34 => X"8000000FF8000000FF8000000FF8000000FF8000000FF80F55E25C00A0BA7FBE",
INIT_35 => X"F8000000FF8000000FF8000000FF8000000FF8000000FF8000000FF8000000FF",
INIT_36 => X"000000000000000000000000000000000000000000000000000000000000000F",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000008000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(0),        -- Port A data input
DOA(0)   => data_read_a_hi(0),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(0),        -- Port B data input
DOB(0)   => data_read_b_hi(0),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_1_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"212C001411984004084D000508C53810A03D1450E839B003342114428A000807",
INIT_01 => X"08000010400A0008010600000084004000400002000000000000000000140000",
INIT_02 => X"484DEBA0111800C004400D000000000028800001CC404E6008B4933336880010",
INIT_03 => X"650C00000848A0423183089008C604224200000100A200002C280810098C0001",
INIT_04 => X"00000004208B00200E010800006667BE7000102C00080000040012010000080C",
INIT_05 => X"0080000000002020600100208D04414000800000000200004800080000800200",
INIT_06 => X"0820196100006044401008100208000008082010000000800488000000020400",
INIT_07 => X"1210C18306788C00894098000011000820001000104050004108000001008250",
INIT_08 => X"00A48903121780004C6000311555521F183060AC564BF818B5EDFDE004460030",
INIT_09 => X"02AD881200100140A0223480000458400000480840002002184581A020000200",
INIT_0A => X"140040001020020410000010082080010400002001041001B102002E20013600",
INIT_0B => X"0895400004201001010884000000901100800800000004140002008280A8A815",
INIT_0C => X"C8D00C8D00C8D40C8D40C8D00C8D20642A06468400000030480808020F08E008",
INIT_0D => X"20BC417C16004C0B83822109040180000801000910000003203220C8C40C8D40",
INIT_0E => X"5C96000000010200200802100022008100408020401020040100142200E0E08A",
INIT_0F => X"0000021E300B000000781E00140018000000781E00140018000002430E30E061",
INIT_10 => X"1C00000024E0000000781E00140018000000781E0014001908400005E11C0610",
INIT_11 => X"0003C30F00C000000155800D00000003E21C0700000000F00118000000468C38",
INIT_12 => X"60640900004A400081401A0000004041218503E4030060000004804318008840",
INIT_13 => X"A0001208C30800025200003D807E000000000725201600090461840001340002",
INIT_14 => X"0000F00C0E06100000012D2005100409520381C00000005920004C0C81200009",
INIT_15 => X"25000120850B8180625400400000010711200510004B41478040000005548016",
INIT_16 => X"10040002002080040000804000A0000000011A000100208C008611430A000040",
INIT_17 => X"0040100401004010040100401004010040100401004010040100401004010040",
INIT_18 => X"0401004010040100401004010040100401004010040100401004010040100401",
INIT_19 => X"5000800000000000000000100401004010040100401004010040100401004010",
INIT_1A => X"8A28A28A2AC8090C69606492492C09945235D5F7E2A5040B80E1C863A2958000",
INIT_1B => X"5BADD6EB75BADD6EB75BAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA28A2",
INIT_1C => X"FC00002E974BA5D2E974BA5D2E974BA5D2E974BA5D2E974BA5D2E974BA5D2E97",
INIT_1D => X"BA55556AAAAAA800000000000000000000000000000000000000000000607FFF",
INIT_1E => X"F45A2FBD75EFA2AE97555F7FBFFF45FFAE80010AAAABFFFFFF803FE10F7D17FE",
INIT_1F => X"8AAAF7FBD54AA002A955555D7FE8ABA082EBFEBAFFD555400557BD54BA5D7FFD",
INIT_20 => X"17555AA8028BEFAAAE97555082A80000AA802ABEFA2D568A005D5157400AA802",
INIT_21 => X"EBDFEF5D7FEAA00AAAABFEAA007BC0145FFFFFDF55AAFBC00105555400105504",
INIT_22 => X"D5575555D7FC2155F7AEA8BEFAAAA954BA557BD7410550428ABA5D5168ABA552",
INIT_23 => X"FD57DF45F7D568ABAF7AABFFFF082ABFFFFFFFFEAB55557FFFEBAAAD568B45A2",
INIT_24 => X"000000000002EBFFEFA280021FF082E974AA5D7BD74000804154BA082ABFF55F",
INIT_25 => X"7F78A3FE28E3D17DEAA485FE8E02B50000000000000000000000000000000000",
INIT_26 => X"6D5D75D54BA5D7BFFF7DA2FFD55EFAAA495545E175EFF57BF8FC2000BEA4BAE9",
INIT_27 => X"A28550E10405F7A4AFE38EAA0924921C2FD55455571E8A2A087BF8EAAEB8E001",
INIT_28 => X"7A28415A001684104155C5B6DF6DBEFBFAA07157428145A00AA8A2FBD7B6DF6A",
INIT_29 => X"AAABF1FFBC7010FF8A38FEF557FEAB78B6AAB8E971471C7010B7D168F47400A0",
INIT_2A => X"495EAAA2D16D1FDBED56A55557A43DE385FD4BFBD7B6A0BF492415FC20105D24",
INIT_2B => X"F5D717FE2AAAA56DEBD17FE3DF7FB7FEBFE38017EBA4A8EB8F6FFD5FE8B7D557",
INIT_2C => X"00000000000000000000000000002A3D5C7AA854008700249243A417FFF41542",
INIT_2D => X"AF2A00010F78028B15F7823FEAAA2D57DFBA007DFCA127B80000000000000000",
INIT_2E => X"A0869AAAB8A7C19C55550E8574BA557BFFFEFAAFBD55FFAA8416545A6FB60F47",
INIT_2F => X"10A2AEBFF55F7BAAA8565DBAC1112FFAC21A022A38C20B2552E975F758516AAA",
INIT_30 => X"01E7AD1FFF5575841DE08007FC2048002895755FFEFBCEE5FBAACB10085EE5DE",
INIT_31 => X"D4000D7FC00FC5D062BBA05ED5034472A02EABEA097BEAAFAF2863FA00DD5742",
INIT_32 => X"62B0A2F7AE8B5D5D51F5E18ABD5EAFFF2AF9554FF57EFBFA18D4FBFFF40FF809",
INIT_33 => X"C95256807DC31AA8114DE55F5BED201FFFED17DFBFF6963FCAAA2283CF140500",
INIT_34 => X"0000000000000000000000000000000000000000000002CB75F7AA84001A7052",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000008000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(1),        -- Port A data input
DOA(0)   => data_read_a_hi(1),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(1),        -- Port B data input
DOB(0)   => data_read_b_hi(1),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_2_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10E44660018259B2843913100062C98004802322D3E030235201006009B2816",
INIT_01 => X"8005A188084900481C8024A542400340404000720885800802000906E4910204",
INIT_02 => X"5C010802020408040C640850AA055254090541A111240A104A0000000908B510",
INIT_03 => X"0C1101108800004481060A001204102803156020218808002440850008C80550",
INIT_04 => X"8840C08122050400582812C21C0804040968987810688899444090C10A124A69",
INIT_05 => X"4885109105400129210040010340086856B141212252142242A068A080106372",
INIT_06 => X"047450004062400090000202000054C28012204400908281302852A6710AA420",
INIT_07 => X"121810000230089008408402A800011012D41D518044411005000AA8A5004390",
INIT_08 => X"A214110514163218085008010141421F02000124000010880000442080810201",
INIT_09 => X"0A09E89041451581B53A739C42A0C9223000004881708D80100331CA8A848E0A",
INIT_0A => X"1009020A30020008096A06B8C1208A000A9C20004820B0573165541CD5482216",
INIT_0B => X"ACC084404A8000490152D100344001108AA88B1D007291402802B1041632A011",
INIT_0C => X"8696086860869608686086920868004309043414A2191C24485C4D2A9A0DF823",
INIT_0D => X"484000804201C1102080215900038AD030014588D200F0221821808682086820",
INIT_0E => X"00002AA00AA80240A001010026824040C000201030000200C8980080260C201E",
INIT_0F => X"0000000A20001602900020001400002A029000200014000100280E6694490312",
INIT_10 => X"0000000024002A02900020001400001602900020001400002700000800010000",
INIT_11 => X"0008004000000000001500006C00300800020000000000C100014A0081200100",
INIT_12 => X"8088000000480005188000440840081000500002000000000004800010003420",
INIT_13 => X"0070041200000002411280004000000000000026000038020900000001201300",
INIT_14 => X"2A0004030000000000002A00004A100208800000000000012260101100000009",
INIT_15 => X"0084420300001040100000000000010402000049800020000000000000580001",
INIT_16 => X"040111000008001505448340606B21090556002E00000000000080002A040A00",
INIT_17 => X"401004010040300C0300C0300C0100401004010040300C0300C0300C01004010",
INIT_18 => X"0200400004000040000C0200C0200C0200400004000040300C0300C0300C0100",
INIT_19 => X"14A97C0FC0FC1F81F81F800C0200C0200C0200400004000040000C0200C0200C",
INIT_1A => X"0410410411823A4301040B2CB2CBACB002009C6B860185AA1491B0E2863EA015",
INIT_1B => X"8944A25128944A25128941041041041041041041041041041041041041041041",
INIT_1C => X"FC703F25128944A25128944A25128944A25128944A25128944A25128944A2512",
INIT_1D => X"AA0004001550000000000000000000000000000000000000000000000078401F",
INIT_1E => X"5FF5D003FE10F7D17FEBAF7D5420AA0855420AAAA843DFFFAAD1554005D7FD74",
INIT_1F => X"FF45AAFBC20AAF7D1575EF55517DF555D2EBFF45AAAAA8A10A2AE80010A2AA97",
INIT_20 => X"AABEFAAD1575EFAAAE974AA5D51554BA5D7FFFF45A2AA975EFA2FFD7555FFFBF",
INIT_21 => X"5554AA555555555557FE8ABA082EBFFFFAAAE95555552E974105D517DF55AAAA",
INIT_22 => X"D540000AA802AABAF7FFC2010AAAE821EF552E82010F7AABFE10FFD542145FFD",
INIT_23 => X"02E800AA08042AB45007FC00BAFFD168BEFF7FBC0010AA802ABEFAAD540000FF",
INIT_24 => X"000000000002E80010555540010550417555AA8028BEFAAAE821550851420AA0",
INIT_25 => X"7A2DF55400557FD54AA1D04001C5150000000000000000000000000000000000",
INIT_26 => X"D5F7A482000BEAE905C755003FE28E3D17DEAAE95F40002157F470AABE803AE9",
INIT_27 => X"5EFAAA495545E3F5EFF57F7FE80082FFDE105EF55517DFC5552ABDF45B6AEAFF",
INIT_28 => X"24105D5B7FF7DB6AAAABC7BEDB505EFBEA4070BA5FD0154BA5D7BFAF7DA2AE95",
INIT_29 => X"38E00B6DF68FEF4871D24BA495B5556D5571E8AAF082AB8EAAEB8E0016D5D2A9",
INIT_2A => X"E2FBD7B6DF47A00EBDB50000A380AAE28E80495038AAAEAF1D7410E80000FF84",
INIT_2B => X"FBC703AE2DF42AAA002A851C214003FF680071ED1EFEAF1EFFFDEAD1C5010AA8",
INIT_2C => X"00000000000000000000000000002087A28415A001684104155C5B68E2DBEFBF",
INIT_2D => X"51FBD74BAF7802AB05AAFBD5400557BD54AA5500021555100000000000000000",
INIT_2E => X"55D2ABDF55F782BEB47AFAD00010F7AA8215555003FEAAAAD57DEBAA2FDDC010",
INIT_2F => X"BA557BEABEFAAEBD55FFAA1456547A2D360F47AF7FC20B2F7FBC015D58517FF5",
INIT_30 => X"AB4A78016545540400010557BFDFFFF7822A955FFFFC20FFF3AE544108410174",
INIT_31 => X"D545002A800A8FF862BA00F2F9E8F0050D4420BA547FD75FF58516AAAA0828AA",
INIT_32 => X"35B57AB5155400A2AEBFF45FFFB404007FFBD550AAFACAAA122AA8954BAA2AE9",
INIT_33 => X"895755FFAEBCFE57BBA57002DF3C4AAAA002E954505C417FFFF08555555BAAD3",
INIT_34 => X"000000000000000000000000000000000000000000000061DE08007FC2048002",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000010000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(2),        -- Port A data input
DOA(0)   => data_read_a_hi(2),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(2),        -- Port B data input
DOB(0)   => data_read_b_hi(2),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_3_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"210C44A20020248B08431120001604B8156023104C40771B3430400A02380206",
INIT_01 => X"014C9A4250B0296D3C2422C992100B49404040028804A0080A000416A8D90A0C",
INIT_02 => X"4809A900031800444460589C66E331352180D468B8040E600C0081110B802CD0",
INIT_03 => X"6D0B6110880001D23583480648D60520330066810A80881068A808029CC56330",
INIT_04 => X"48221A066A09D03B348C1C1928DD5A4402A13868070940842640902107002D24",
INIT_05 => X"058318035328202004C1C4E50B44644B30A86D01014A0D224063090082100E34",
INIT_06 => X"08381A010040200AC2190ED2002ACD99881822104C5A40942048288234629414",
INIT_07 => X"0218408142740E2C0948C3066400071913209CC8004640100D003999552083D2",
INIT_08 => X"900409231292A8080C2000110001521F0810A92E7402F08AB0016CA000C60011",
INIT_09 => X"620C889014D30E4A210214D5099058808010605A81A41480102130C020A43A39",
INIT_0A => X"512850E61822020C899046740121820004102000402079CCA037A02C68552A35",
INIT_0B => X"8895000026A00141015290040460C0B4828289AC1011954C0026A20400882914",
INIT_0C => X"80CA080DA080DA080CA080CE080DB0402F040654A2442834C0092E228A0DF2AB",
INIT_0D => X"289080600E04C50206808059000999C98840C508D220108200202080DA080CA0",
INIT_0E => X"300E6660599802602209021204A050E1C850C428521C208480821D842085A03E",
INIT_0F => X"0000010000003202900000010000000A02900000010000008038666920920A24",
INIT_10 => X"0000008000002202900000010000001E02900000010000002380000800000000",
INIT_11 => X"0008000000000000008000002D00300800000000000020010001620081200000",
INIT_12 => X"8088000008001021C88000048800281000500000000000004000000000003600",
INIT_13 => X"00B8041200000040011980004000000000000803000068020900000020001B00",
INIT_14 => X"29800403000000000008030000C83002088000000000002002E0101100000100",
INIT_15 => X"00841003100010401000000000002000030000C38000200000000000020C0001",
INIT_16 => X"108722420420A0100006D34A404800185CCE0128410820000008008021C40A00",
INIT_17 => X"0872108721085218852188521885218852188521887210872108721087210872",
INIT_18 => X"8721086214872108621C852188421C852188421C852188721087210872108721",
INIT_19 => X"54A2EAA555AAB554AAB5561C852188421C852188421C85218842148721086214",
INIT_1A => X"0410410412881D0B0000092492480A981E063C638321450A08899A62C314A014",
INIT_1B => X"9D4EA753A9D4EA753A9D49249249249249249249249249249249249249241041",
INIT_1C => X"FAABC4351A8D46A351A8D46A351A8D46A351A8D46A351A8D46A351A8D46A351A",
INIT_1D => X"5500002AA100000000000000000000000000000000000000000000000000401F",
INIT_1E => X"FFFAAD1554005D7FD74AAA284001550055421EFAAFFD54AAF7D168B45AAAABDF",
INIT_1F => X"20AA080400155AAD5554AAF7802AB4500043DF45FFD168AAA0855420AAAA843D",
INIT_20 => X"021550855555FFAA84001FFAAAE80010A2AA955FF5D003FE10F7803FEBAFFD54",
INIT_21 => X"BC20AAA284175EF55517DF555D2EBFE00AA8028B45A2AE82155A2FBFFEBA0800",
INIT_22 => X"7BD7555FFFBFDF55AAFBD55EF5D2EBFE10085168ABAFFFBD54BAAAAE97400A2F",
INIT_23 => X"D0015410F7AAAAAAA55043DE00FFFFD5555AAAA954AA5D7FFFF45AAAA975EF00",
INIT_24 => X"0000000000004174105D517DF55AAAAAABEFAAD1575EFAAAE974AA5D00175555",
INIT_25 => X"2EBD56DB7DBEAEBFF551C042AA101D0000000000000000000000000000000000",
INIT_26 => X"D75D5B470AABE8A3AFD7A2DF55400557FD54AABC04001C51551471D7AAF1D05D",
INIT_27 => X"E28E3D17DEAAEBDF40002550F47155AADB50492EB842FB5508043FF55EBD56AB",
INIT_28 => X"017DAAFFFAE821C0A0717D1C5B575FFB68E82557FD2082000BEAE905C755003F",
INIT_29 => X"D74BAE3AE85480FFFFC00AABE8E105C755517DF40552ABDF45B6AEAFFD5F7A48",
INIT_2A => X"FFAF7DA2AE905EF0075D5545E3F5EFF57F7D5C55D7492E90E3808756DA92EBFF",
INIT_2B => X"F5C7092FF801756D490A10438EBA4B8E9241043AE10EAF5C5547FF80954AA5D7",
INIT_2C => X"00000000000000000000000000000E124105D5B7FF7DB6AAAABC7BEDB505EFBE",
INIT_2D => X"515157555AAD142040A2D57FFFFFFAEBFF555D0028A005100000000000000000",
INIT_2E => X"500003FF55AAFD6AB455157D74BAF7AAA8B45AAFBD54005D7BD54AAF78002155",
INIT_2F => X"10F7AA8215555003FEAAAAC53DEB8A2FDDC01051AE955F7AAFBC0000AF843FF5",
INIT_30 => X"F51F782BCB47ABAE801FFAAFBEAA105D2E955FF557BD74EFFBACD41577B84000",
INIT_31 => X"0AAA00557FEA8A2FDD64BAAF8282012AFFEC20BAF7AA8015558517FF555D2ABD",
INIT_32 => X"48547AE04174BA557BEABEFA2AA951FF88554214FA2D3EAF57AFFDD7555082AA",
INIT_33 => X"22A955FFFFC21FFF3BE40412DE02955FF082A820AAAB842AA00000028AB0AAFF",
INIT_34 => X"0000000000000000000000000000000000000000000002A80010557BFDFFFF78",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000008000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(3),        -- Port A data input
DOA(0)   => data_read_a_hi(3),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(3),        -- Port B data input
DOB(0)   => data_read_b_hi(3),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_4_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10804002061080A284201081034809800A00230340007833522C82D04A16006",
INIT_01 => X"804399801838084C0420450E1E104348403008418984014902030006A0910204",
INIT_02 => X"480108A200000000446418E01E80F00A4104311868240200080000000988A390",
INIT_03 => X"065140108800004080064A0002001128270072E03000000030808D00888100F0",
INIT_04 => X"9100EB836A155C1AF0B81CD60433B944022AB8385AC0D4B8E02010E81C32E821",
INIT_05 => X"5C0F20B36F08000024C084C501441C4CF01C489533483C8042EAC190001074C4",
INIT_06 => X"0034420151620118120106902406C3C7800201448DD9D2871020F2AA375A6071",
INIT_07 => X"12181000023480040840C001E080030032009700024641000C00187A442007C2",
INIT_08 => X"8084830110160218004000001101121F220000260000108AA000440880000000",
INIT_09 => X"5A8C881063DF3E839008F29F407448F200B020DA841CA2001001008882046647",
INIT_0A => X"C61504C1380101801900439001FD8804041400001002003C230B6715A4786E0F",
INIT_0B => X"ACD1240522E000098100D104B26041348A088078116C105DA006D10416BE3002",
INIT_0C => X"8608086180860808608086180860A0434C0430D4A25F3182CC4D5D221A09E821",
INIT_0D => X"0BC28081080549504400A8080009B878184044881222D1821821A08628086180",
INIT_0E => X"20481E0E18790012820001100200D02048300418022C1282809A09040415002A",
INIT_0F => X"0000010020005E0090000001000000C6009000000100000000380E6C30830806",
INIT_10 => X"000000800000D20090000001000000EE0090000001000000A6A2000000000000",
INIT_11 => X"0000000000000000008100003B00200800000000000020010002EA0080200000",
INIT_12 => X"80800000080000211D80000C0044281000400000000000004000000010003282",
INIT_13 => X"03B00410000000400121800000000000000008020000B8020800000020006F00",
INIT_14 => X"59000402000000000008020000C9000200800000000000200FC0101000000100",
INIT_15 => X"008A500100001040000000000000200002000042E00000000000000002080001",
INIT_16 => X"08820440040802500104C34820E3031B63C20530C01800410009009821040A00",
INIT_17 => X"C832008020C812008220C81200802048320880204832008020C8320082204812",
INIT_18 => X"8120481208822008020C812048320880208802048320C8120882204812088020",
INIT_19 => X"10A3A5930C9A6CB261934E048320C81200822008220C81204832008020882204",
INIT_1A => X"8A28A28A2BD30264686668A28A2605145031C03F028000A1C2ED7831A2822250",
INIT_1B => X"51A8D46A351A8D46A351AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA28A2",
INIT_1C => X"F94304068341A0D068341A0D068341A0D068341A0D068341A0D068341A0D0683",
INIT_1D => X"BAAA84154005500000000000000000000000000000000000000000000000401F",
INIT_1E => X"4AAF7D168B45AAAABDF55A2802AA1000002ABFF087FFDF5508003FEBA087FD54",
INIT_1F => X"015500002AABA082E954005500021FF5D2EBFF5500003DF455555421EFAAFFD5",
INIT_20 => X"174BAA2AABDE0055517FF555555420AAAA843DFFFAAD1554005D7FD74AAAA840",
INIT_21 => X"400155AAD1554AAF7802AB4500043DF45FFD168BEF080028BFF0855555455500",
INIT_22 => X"803FEBAFFD5420BA085168A00007BFDE10085168ABA0055574BA5555554BA5D0",
INIT_23 => X"02A97545F7D1555EF55043DF5555517DEAA5D0400010A2AA955FF55003FE10F7",
INIT_24 => X"000000000002A82155A2FBFFEBA0800021550855555FFAA84001FFAAFBEAB450",
INIT_25 => X"5080A3AEAA007BD2482BE84124285C0000000000000000000000000000000000",
INIT_26 => X"381451471D7AAFBD0492EBD56DB7DBEAEBFF55BC042AA101D0A28BC7007FFDF4",
INIT_27 => X"400557FD54AABE84001C5550A28ABA1424974004100021FF492AB8F7D1C0438E",
INIT_28 => X"8BEF005557545490012482B6A0BAE2849557AFED1C5F470AABE8A3AFD7A2DF55",
INIT_29 => X"504924955524AA140E0717DAADB50492EB842FB5508043FF55EBD56ABD75D042",
INIT_2A => X"A905C755003FE28E3803DEAAEBDF40002557F6DA101475FDE10145F68A921C55",
INIT_2B => X"DF425575D7BEFB55002097555FFD5401EF5D043AF6D405F78E3A1C2002000BEA",
INIT_2C => X"0000000000000000000000000000208017DAAFFFAE821C0A0717D1C5B575FFB6",
INIT_2D => X"512EAAB45007FFFF55082EA8AAA087FC2010F784000AA5900000000000000000",
INIT_2E => X"F002EA8BEF5D0428ABA595557555AAFBC2000A2D57FFFFF7AEBFF55FF8028A00",
INIT_2F => X"BAF7AAA8B45AAFBD54005D7BD54AAF78002155512AAAA085D04174100800021F",
INIT_30 => X"F55AAFD6AB4551002ABEF005555555000402000FF802ABAA04552ABFF597FD74",
INIT_31 => X"DE005D7BE8AA85555400100879560AA592F955FFAAFBC0000AF843FF5500003F",
INIT_32 => X"FCABA598400010F7AA8215555003FEAAAA843DEB0A2FD5600051537DE005D557",
INIT_33 => X"E955FF557BD75EFFBBCD415521FBFDF45000417545FFD5421FF5D0428BEF0079",
INIT_34 => X"00000000000000000000000000000000000000000000004001FFAAFBEAA105D2",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000010000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(4),        -- Port A data input
DOA(0)   => data_read_a_hi(4),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(4),        -- Port B data input
DOB(0)   => data_read_b_hi(4),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_5_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50DB4A0791B1B4B694369283C81F9996A091832112004AB37B20E07C0C1E006",
INIT_01 => X"085FBC448000804C446A00000034826841280A00084000C8C212802EE2953235",
INIT_02 => X"C809AD5CB118E640A4D018FC011FF0002080000082C8C66609DB7DDDCB1F2036",
INIT_03 => X"250907263E4C90D210835C82484205720B20640A88800000B8E0F810A8C4500E",
INIT_04 => X"4005102126898100064D20001044429C7824382C0416C087198AB916E0551A24",
INIT_05 => X"A370C14CA0E101094008002389CFE2F20D7D7A114CB5C20AE514178054948912",
INIT_06 => X"547319A1499121D4C0A046FC4E06C030581859058C2404844437118630839B88",
INIT_07 => X"2A53468D1A758C038AFFEA9FE39348C9204C389672407EF120EA5806E6C543AC",
INIT_08 => X"8C05896372728FE0C420619000003AFF48D1222E5D26F06ABCC96CD72C463990",
INIT_09 => X"82DE9AB9182080C801041080300F6F0E42821809C2FEA0B65A212282002B029F",
INIT_0A => X"1688E480D10A90049026145B3830B64944904569E7E00A002C836D35B68D26C0",
INIT_0B => X"88990E14269AB54B078092E6BD4431138A00AEFDD567DA480816848C94180846",
INIT_0C => X"C0591C0791C0491C0791C0591C06A8E0248E03D68860A0106119883D6AE1A0A4",
INIT_0D => X"23D829FA654184533252095E542387F81008071C1BAAD68B027029C0491C0691",
INIT_0E => X"0CA7FE0227FC25847C4395166C5844480204011210A11028C380802A24C89494",
INIT_0F => X"1C55D65E3E3C017C37FC3E0017C1F8017C37FC3E0017C1F90005024108308061",
INIT_10 => X"1C0118796FE0017CA7FC3E0017C1F8017CA7FC3E0017C1F9100DFFF5E15D0610",
INIT_11 => X"FFF3E34F00C0270F3755F1F8007FCBEBE25E0700463E17F2C7E014FF7AE6CD38",
INIT_12 => X"64E4090626DE40100459759173BBD6EF37C523E6030061341F07FC571F8F800D",
INIT_13 => X"E0A6FE28C3082636F201BFFF807E00007E03F7243D38337D1C6184131B7C1DEF",
INIT_14 => X"397FFA0E0E06101C53E36C3D3E884FDDD28381C0098E57D923BDFC8C8120C4DB",
INIT_15 => X"FA36FDF58DBF81C062540049707E0FE7303D3E03BFFF41478040570EED50F4F8",
INIT_16 => X"88212B100901A2349004C26A624A21040FC190050A2110B8ACC40B204A119074",
INIT_17 => X"C20080230802108C2008C22080210882108C220842208821088210842208C200",
INIT_18 => X"20084220842208C2008823080230802108823084220842008821080230842008",
INIT_19 => X"54C1892596D34924B2DA6884220842008C20084220802108821080230802308C",
INIT_1A => X"BEFBEFBEFB7F7FE7EFEEE79E79EFAF2DDA73FBDCEDBFF9D3F0FDE0DB6DBF6218",
INIT_1B => X"DEEF77BBDDEEF77BBDDEEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEF",
INIT_1C => X"FAF3167BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBD",
INIT_1D => X"BA5D2ABFFEFFF80000000000000000000000000000000000000000000000401F",
INIT_1E => X"F5508003FEBA087FD54BA0804154005555574AAA2802AA10FFFFFDE0008556AA",
INIT_1F => X"AA1000003FEBA00002AABA5D2EBFEBAAAD16AABAF7AAA8BFFAA802ABFF087FFD",
INIT_20 => X"E8B45FF80001555D2E955FFFFD5421EFAAFFD54AAF7D168B45AAAABDF55AA802",
INIT_21 => X"02AABA082E954005500021FF5D2EBFF5500003DE005555575EFA2D142145A2FF",
INIT_22 => X"7FD74AAAA840014500517FFEF007BEABFF5D7FC00BA5D5568AAAF7AAAAAAAAA8",
INIT_23 => X"2FBEAA105D2E97410FFD16AAAA5D2ABDEBAFFD5420AAAA843DFFFAAD1554005D",
INIT_24 => X"000000000000028BFF0855555455500174BAA2AABDE0055517FF555504154BAA",
INIT_25 => X"0FFFFFFE38085F6FA92552AB8FEFF78000000000000000000000000000000000",
INIT_26 => X"C7B68A28BC70075FDF45080A3AEAA007BD24821E84124285C51574BAB68A2DA0",
INIT_27 => X"B7DBEAEBFF55BE842AA105D0A38EBA1C0428A925D2AB8EBABEDB6AA92F7AAA8B",
INIT_28 => X"75EFA2DB45145B6F5EFB6DF78E05145552A925FFFFD1471D7AAFBD0492EBD56D",
INIT_29 => X"68AAAF7AAAAA82BE8A28A921424974004100021FF492AB8F7D1C0438E38145B5",
INIT_2A => X"A3AFD7A2DF55400557FD54AABE84001C555517DFC70875EABC7557FC20AA415F",
INIT_2B => X"043AFED1C0E10492B6FFEFA105D2A95410FFDB6FABA542ABAE2AF7DF470AABE8",
INIT_2C => X"00000000000000000000000000000428BEF005557545490012482B6A0BAE2849",
INIT_2D => X"5955554BAFFAEBDE10F7FBFDEBA007BFDE005D2AAABEFFB80000000000000000",
INIT_2E => X"AF7FBE8A00FFAEAAB45F3AAAAB4500557FF55082EA8AAA087FC20105504000AA",
INIT_2F => X"55AAFBC2000A2D57FFFFF7AEBFF55FF8028A00512AA8AAA5D0028A005D2AA8AB",
INIT_30 => X"BEF5D0428ABA597FD55FFA2FFD5555FFD57FFEFFFAA97545552A821EFFBD5575",
INIT_31 => X"8B55557FC0012087FEAABAF7AAAAA10F3AAAAA005D04174100800021FF002EA8",
INIT_32 => X"A8ABAFBFFD74BAF7AAA8B45AAFBD54005D7BD54AAF7800015551517DF4500516",
INIT_33 => X"402000FF802AAAA04452ABFF592E80010FFFFFFE005D2A95410F7FFFFEBA5D2E",
INIT_34 => X"000000000000000000000000000000000000000000000002ABEF005555555000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000060000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(5),        -- Port A data input
DOA(0)   => data_read_a_hi(5),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(5),        -- Port B data input
DOB(0)   => data_read_b_hi(5),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_6_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10804B0061A010A2840012C030028180004003220200403302301C0381A0086",
INIT_01 => X"A70041CA3839684D18A160000C52424841000000090800090210080008110204",
INIT_02 => X"080108200C1000004465480400C0080100000000010432400800800009882050",
INIT_03 => X"040001008C2340D0842208624210802182800584488000103080014E08C10000",
INIT_04 => X"00101611A029B08410044800000000040088122A44281C040400900500001800",
INIT_05 => X"02800000400C820934E4A0002900404402820024000A00824004283011200A00",
INIT_06 => X"2632000004084804134DA7C011A83FC012122100C80812D00308010000829400",
INIT_07 => X"02181020423088002940C2401D0480112000100004404014602447F805326393",
INIT_08 => X"7004812130160008304000000000021F020408244000108A0000440003040000",
INIT_09 => X"020C889010104088A000348037F05840303902E814000010341108802020FF40",
INIT_0A => X"86C8B5DF1C83C9C8900000100220C244840021100017E2FD200000A40001223F",
INIT_0B => X"88D1804122A088018152D144317205502A880C00107FD75DE922005026A62A15",
INIT_0C => X"B6284B6284B6184B6184B6384B62825B0425B0568075A0826849C8229AC5F8AE",
INIT_0D => X"03C440C054048850A300A8480009A0020865A588DA20F1A2D92D82B6084B6084",
INIT_0E => X"031001E0800122100321C89214A01A742D3A168D1B4686D100234B442428C034",
INIT_0F => X"000008AB80030202800000001402068202800000001402067400026000000000",
INIT_10 => X"00000000341E8202100000001402068202100000001402062840000800000000",
INIT_11 => X"0008000000000000083C00052000300000000000000008CD0018400081000000",
INIT_12 => X"800800000069A48584000A0400000010001000000000000000048128C0002840",
INIT_13 => X"1A480012000000034C1E000040000000000400FE000644020100000001A34000",
INIT_14 => X"02800401000000000004BA000112B0020800000000000807E80000110000000D",
INIT_15 => X"0500020250001000100000000000010CCE000198000020000000000010F80006",
INIT_16 => X"62D18468CE8402440404D24A3081B020603E0A20640C8400010298432A002A00",
INIT_17 => X"ED3B4ED0B42D1B4ED3B42D0B42D1B4ED2B42D0B46D3B4ED2B42D1B46D3B4AD2B",
INIT_18 => X"D0B46D3B4AD0B46D1B4AD3B4ED0B42D1B4ED2B4ED1B42D0B4AD3B4ED0B42D0B4",
INIT_19 => X"002331C618E38E38C31C7346D3B4AD2B46D1B42D2B4ED2B42D1B46D2B4AD1B42",
INIT_1A => X"8E38E38E39DB3B676F66EFBEFBEFAFBC5E73FC7F87A7D4ABFE7CFAFBE7BF8040",
INIT_1B => X"CFE7F3F9FCFE7F3F9FCFE38E38E38E38E38E38E38E38E38E38E38E38E38E38E3",
INIT_1C => X"FF75A43F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9F",
INIT_1D => X"BA5D7BEAAAAFF80000000000000000000000000000000000000000000060401F",
INIT_1E => X"A10FFFFFDE0008556AABA5D2ABFFEFFF843DFEFA2FBD54BA5555554BAAAFBC20",
INIT_1F => X"5400550428AAAAA84021FF007BD54BAAAD17DEBA0855421455555574AAA2802A",
INIT_20 => X"17400AAFBE8ABAF7FFD54AAAA802ABFF087FFDF5508003FEBA087FD54BA00041",
INIT_21 => X"03FEBA00002AABA5D2EBFEBAAAD16AABAF7AAA8BFFAAD1554BA002A95555A284",
INIT_22 => X"AABDF55AA802AA100000001EF087FEAA00FFFBD5545080417555A2D17FE10000",
INIT_23 => X"2803DFEF0855401FF082EA8B555D7FC21FFFFD5421EFAAFFD54AAF7D168B45AA",
INIT_24 => X"0000000000055575EFA2D142145A2FFE8B45FF80001555D2E955FFFF843DEAAA",
INIT_25 => X"A415B52492B6F5C20825D7FE8A92FF8000000000000000000000000000000000",
INIT_26 => X"555551574BAB68A2DA00FFFFFFE38085F6FA92552AB8FEFF78E3DFFFAAFFD04A",
INIT_27 => X"EAA007BD24821C04124281C0E2DA82BE8E001EF147BD2482BED57AE921451421",
INIT_28 => X"24AA14209557DA28E15400BEF1EFA92FFFFD24BAB68A28BC70075FDF45080A3A",
INIT_29 => X"17545B6D178E281C0A38EBA1C0428A925D2AB8EBABEDB6AA92F7AAA8BC7B6D55",
INIT_2A => X"BD0492EBD56DB7DBEAEBFF55BE842AA105D0E071FF0071EDA38F7F1D55550004",
INIT_2B => X"2A925FFFF8E3DE82BE8E38FFF0851401C70824A8B555C7FC2147F7D1471D7AAF",
INIT_2C => X"00000000000000000000000000005B575EFA2DB45145B6F5EFB6DF78E0514555",
INIT_2D => X"FBAABDFEFAAFBC00BA007BC0000FFD542000557FE8A00F380000000000000000",
INIT_2E => X"0F7D168A105D55421455155554BAFFAEBDE10F7FBFDEBA007BFDE005D2AAABEF",
INIT_2F => X"4500557FF55082EA8AAA087FC20105504000AA592ABFE00F7AA821FF557FC001",
INIT_30 => X"A00FFAEAAB45F3D5400BA5504155EFAAAE95410F7D57DE00FFFBC00AAFBAAAAB",
INIT_31 => X"FEAAF7D157545080417545F7D56AAAA592AA8AAA5D0028A005D2AA8ABAF7FBE8",
INIT_32 => X"C2145F3D557555AAFBC2000A2D57FFFFF7AEBFF55FF8028A00512E975FF08557",
INIT_33 => X"57FFEFFFAA97545552A821EFFBAABDE00F7AAAABEF005542155000028B555D7F",
INIT_34 => X"0000000000000000000000000000000000000000000007FD55FFA2FFD5555FFD",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000048000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(6),        -- Port A data input
DOA(0)   => data_read_a_hi(6),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(6),        -- Port B data input
DOB(0)   => data_read_b_hi(6),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_7_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10840B0048225802842102C02450418800002300500030B313300C418992002",
INIT_01 => X"A34009C23838684D1C20E0000E11426840000000080000080200090000510200",
INIT_02 => X"4801082048100000446558040080000041000000000622400800000009000010",
INIT_03 => X"040001818CA144D0842248424210812102000400088000003080014688800000",
INIT_04 => X"000010002041800000048000000000040088322944200C850001940400301800",
INIT_05 => X"0200000040004100280040204104004402000025000800065004203030320800",
INIT_06 => X"0430060044084804900806D1112A002012120004440812D40120008200829001",
INIT_07 => X"02181020423408002940C24001A4A010200018920646C10C7035000244004380",
INIT_08 => X"008481213016020C204000000000121F020408264000100AA000440012040000",
INIT_09 => X"820C899410000000A100348020005902B1A0048825008091350100CAA0200280",
INIT_0A => X"50140A0010058188100004590331C9C4A400231200340C012100002400012200",
INIT_0B => X"1811C44D22A1884141600411800008104080890023000009A926801050001C00",
INIT_0C => X"9002C9002C9022C9022C9022C903064809648080204020004009080A0A00E088",
INIT_0D => X"0880144434A0010012280008031980036000014A0046206241A4069002C9002C",
INIT_0E => X"0216000200010000000081102080400040002000002010000004008080048A00",
INIT_0F => X"038A2881210382000000001E003E0582000000001E003E042283424000000000",
INIT_10 => X"60700706901982000000001E003E0582000000001E003E046840000000009864",
INIT_11 => X"00000000330C00F0C8210807200000000000581C01C1C809201C400000000001",
INIT_12 => X"0000C2419121028C00020A2400000000000080082C180603A0E003A090406840",
INIT_13 => X"14E8000004321189085F8000000061E001FC00C00207740000021908C4829D00",
INIT_14 => X"BB800000009864038C14800201BAB000000026130071A80613A0000018483224",
INIT_15 => X"0546520350000600812058100F81C018880201BBA0000008239020F110800806",
INIT_16 => X"24003300080022140444D268624B210040004A08000000044222900320C84008",
INIT_17 => X"4010040100402000000000000003004010040100000000000000100401004010",
INIT_18 => X"0000C01004010000000001004010040000000004010040300400000000000200",
INIT_19 => X"54A2C208200010410400000800000000040100C01000000000100C0100400000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000002A10",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FAF8800000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"55002E820AAAA80000000000000000000000000000000000000000000000401F",
INIT_1E => X"4BA5555554BAAAFBC20BA5D7BEAAAAFFFBC00AAF7D5575455D557DFEF002AAAB",
INIT_1F => X"FFEFFFAAAAAAAF7D57FFEFF7D555555A2AEAAB55007FD74AAAA843DFEFA2FBD5",
INIT_20 => X"FDF550000175555504175450055574AAA2802AA10FFFFFDE0008556AABA5D2AB",
INIT_21 => X"428AAAAA84021FF007BD54BAAAD17DEBA085542145552ABDFEFFFAA801EFFFFB",
INIT_22 => X"7FD54BA000415400557BD74BAFFD140000082A975EF00003DF55555168A00000",
INIT_23 => X"5557FEAAA2843FF55A2AEA8B55AAAABDEAAFF802ABFF087FFDF5508003FEBA08",
INIT_24 => X"0000000000051554BA002A95555A28417400AAFBE8ABAF7FFD54AAAAAEA8ABA5",
INIT_25 => X"5415178FD7082EAAB550820870BAAA8000000000000000000000000000000000",
INIT_26 => X"82AA8E3DFFFAAFFD04AA415B52492B6F5C20825D7FE8A92FFFFC70BAE3D15555",
INIT_27 => X"E38085F6FA92552AB8FEFF7A0ADABAEBD578FFFEBD55557DBEA4AFB550871D74",
INIT_28 => X"DFD7FFA4801D7F7F5FDF55000E17545410E175550051574BAB68A2DA00FFFFFF",
INIT_29 => X"3AF55415F6DA38080E2DA82BE8E001EF147BD2482BED57AE921451421555524B",
INIT_2A => X"5FDF45080A3AEAA007BD24821C04124281C7BD2482E3D1450381C20905EF0800",
INIT_2B => X"FFD24BAB6A4A8A82495F78E92AA843DF45BEAAAFB55ABA0BDE02EB8A28BC7007",
INIT_2C => X"000000000000000000000000000055524AA14209557DA28E15400BEF1EFA92FF",
INIT_2D => X"F3FFD54BAAAD15754508556AB45002AA8B450800174BAA680000000000000000",
INIT_2E => X"FF7803DF45085557410AEAABDFEFAAFBC00BA007BC0000FFD542000557FE8A00",
INIT_2F => X"BAFFAEBDE10F7FBFDEBA007BFDE005D2AAABEFFB803DEAAAAD56ABEFAAD5575E",
INIT_30 => X"A105D554214551003FF45FF8400145FFD57FF55082E97555002E955550C55554",
INIT_31 => X"54AA5500021EF000028B55087BFDEBA042ABFE00F7AA821FF557FC0010F7D168",
INIT_32 => X"3FE10AEAAAAB4500557FF55082EA8AAA087FC20105504000AA597FC2010A2D15",
INIT_33 => X"E95410F7D57DE00FFFBC00AAFB8028A00007FE8A00A2803FF45F7AABDF55AA84",
INIT_34 => X"00000000000000000000000000000000000000000000055400BA5504155EFAAA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000007FFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(7),        -- Port A data input
DOA(0)   => data_read_a_hi(7),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(7),        -- Port B data input
DOB(0)   => data_read_b_hi(7),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_8_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00000648E2840112C00000418000002700500030B3132000400812082",
INIT_01 => X"A14008420008204D042100000212026840000000180800080200090048510204",
INIT_02 => X"080108000090000004655C040080000051000000000402400800000009000010",
INIT_03 => X"00000100803008D0842240024210810002800584488000103080894288800000",
INIT_04 => X"00009610A028B084000440C0040000040088323244280C950400808500321800",
INIT_05 => X"42800080400C8A09306420202804400402800035200A00020204283001114A00",
INIT_06 => X"2230400041404B141345A7C20426FFC01292214444081254002801A200821400",
INIT_07 => X"021810204214080069408200008C1010200018920E06C0000020DFFA453223D3",
INIT_08 => X"0084010110120008024000000000021F02040826400000008000440000240000",
INIT_09 => X"828D8880100040898128768820045142B0B902E815008080A0B13848A2200280",
INIT_0A => X"9148A4801C81C9C8100004590711800414002004402008013000403084090200",
INIT_0B => X"BC95C44522A002410040940084720450220089000100104DE924800030821452",
INIT_0C => X"0000400004000040000400004000220010200114AA4020004009092A0009E0A8",
INIT_0D => X"0BC4028430108150900408590109A00209642500120230200100220020400004",
INIT_0E => X"0010000600002210A320C89000005A142D0A16850B6294D10023420124240114",
INIT_0F => X"00000800008100020003C1FE00020080020003C1FE0002004401426008208041",
INIT_10 => X"E3F00000100080020003C1FE00020080020003C1FE000200080000081EA2F9EC",
INIT_11 => X"00081CB0FF3C000008000201000010001DA1F8FC0000080110080000010132C7",
INIT_12 => X"0B0BE6C00020040580040200000001004832CC19FCF81E000000010000200800",
INIT_13 => X"020000C31CF60001008000007F01FFE00004000200420000618E7B0000804000",
INIT_14 => X"000000F151F9EC0000040200401000200D547E3F00000800080001617AD80004",
INIT_15 => X"0100000822406E1B95A3F83000000008020040100000BAB87FB0000010080102",
INIT_16 => X"66D1A368C68D26000544D26A504AB12040022220640484000110184300002A02",
INIT_17 => X"6D1B46D1B46D1B46D1B46D1B46D0B42D0B42D0B42D0B42D0B42D1B46D1B46D1B",
INIT_18 => X"D1B42D0B42D0B42D0B42D1B46D1B46D1B46D1B42D0B42D0B42D0B42D0B42D0B4",
INIT_19 => X"442200000000000000000346D1B46D1B42D0B42D0B42D0B42D1B46D1B46D1B46",
INIT_1A => X"9E79E79E7B7F11E66C6FAD96D96520145052A1F5E2BD085122ED48F3AEB20840",
INIT_1B => X"C3E1F0F87C3E1F0F87C3E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7",
INIT_1C => X"FA2A6D4F87D3E1F4F87D3E1F4F87D3E1F4F87D3E1F4F87D3E1F4F87D3E1F4F87",
INIT_1D => X"FFFF84000AAFF80000000000000000000000000000000000000000000000401F",
INIT_1E => X"5455D557DFEF002AAAB55002E820AAAA840000000043DF55087BC01EF007FD75",
INIT_1F => X"AAAAFFAA95545552ABFE00087BC00AA082EBFE10A28028AAAAAFBC00AAF7D557",
INIT_20 => X"E8BFFA2FBFFFFFAAD5400AAFF843DFEFA2FBD54BA5555554BAAAFBC20BA5D7BE",
INIT_21 => X"AAAAAAF7D57FFEFF7D555555A2AEAAB55007FD74AAAAD57FF45002A975FF007B",
INIT_22 => X"556AABA5D2ABFFEFFFAA82000555555545AAFBE8A00082A97410F7D5555EFAAA",
INIT_23 => X"87BC2010AAD54014500516ABFFA2AABDF450055574AAA2802AA10FFFFFDE0008",
INIT_24 => X"000000000002ABDFEFFFAA801EFFFFBFDF550000175555504175450000155450",
INIT_25 => X"50075C71FF087BD75D7FF84050BAEB8000000000000000000000000000000000",
INIT_26 => X"BABEFFC70BAE3D155555415178FD7082EAAB550820870BAAA8407000140038F4",
INIT_27 => X"492B6F5C20825D7FE8A92FFA497545552AB8E10007FC50BA002ABFE00AA8A2AA",
INIT_28 => X"DF451C24955EF0875EFBD7B6F1FFFC7BEDB45082EB8E3DFFFAAFFD04AA415B52",
INIT_29 => X"92410EBD5505EFB6A0ADABAEBD578FFFEBD55557DBEA4AFB550871D7482AAD17",
INIT_2A => X"A2DA00FFFFFFE38085F6FA92552AB8FEFF7AA87000415B5057DAAFBE8A100820",
INIT_2B => X"0E17555000E17545007BC0000BED14217D005B6ABC7B6AABFFED0051574BAB68",
INIT_2C => X"000000000000000000000000000024BDFD7FFA4801D7F7F5FDF55000E1754541",
INIT_2D => X"A684174105D042AB550055555FF007BD7555F784174AAA280000000000000000",
INIT_2E => X"A082EBDE10AAAEA8ABAF7FFD54BAAAD15754508556AB45002AA8B450800174BA",
INIT_2F => X"EFAAFBC00BA007BC0000FFD542000557FE8A00F384175555D2EA8A00087BD74B",
INIT_30 => X"F45085557410AED17FF455D04155FF00557DF55FFD57DF55FFFBD5400A2AABDF",
INIT_31 => X"21EFA2FFEAA00000002010A2D5421FFFF803DEAAAAD56ABEFAAD5575EFF7803D",
INIT_32 => X"BDFEF0855554BAFFAEBDE10F7FBFDEBA007BFDE005D2AAABEFFBAE97410087BC",
INIT_33 => X"57FF55082E97555002E955550C2E95555087BC0010FFD1401EF087FE8B55FFAE",
INIT_34 => X"000000000000000000000000000000000000000000000003FF45FF8400145FFD",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000020000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(8),        -- Port A data input
DOA(0)   => data_read_a_hi(8),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(8),        -- Port B data input
DOB(0)   => data_read_b_hi(8),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_9_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00018248A2840112C00002C18000002300500030B3132000400812006",
INIT_01 => X"A1400802000020490000000000000240413C0A61590001D90213C90008510204",
INIT_02 => X"680108200010000054655C040080000041000000010402400800800009082011",
INIT_03 => X"00040100800020D0842240124210810042800504488000103081894288800000",
INIT_04 => X"00001410A00AA084000400C0060000040088323044201C850020820400101880",
INIT_05 => X"0200020040048A09202420000C00410402000025000800020804203000100800",
INIT_06 => X"22320400404048041144A7D2003A002012120004DC08125400A0008300821000",
INIT_07 => X"06181020421C08000940820000800010200018B20206C00000200002441223C1",
INIT_08 => X"0184010110120008004000000000061F02040826400008118000440000040000",
INIT_09 => X"8208888210004009010852882000510230A900A8040080800055086002200280",
INIT_0A => X"1402008004814948100004590111C004040120000020080121024012A4081200",
INIT_0B => X"2C91844522A0004100488000801200D00000880001000415E1248002103C2294",
INIT_0C => X"080040820408004082040800408202040020410402000000400809080508A080",
INIT_0D => X"0B4000803200C150108008490809A00219246101100220202102020820408204",
INIT_0E => X"00160006000120002120499020A04A14650A328519629651900142002404201E",
INIT_0F => X"0000080A20010002100000001402008002100000001402000001426008208041",
INIT_10 => X"0000000034008002800000001402008002800000001402008800000800000000",
INIT_11 => X"0008000000000000081500010000100800000000000008C10008000001200000",
INIT_12 => X"0088000000680005800002000000000000500000000000000004810010000800",
INIT_13 => X"02E8040200000003401F80004000000000040027000274000900000001A05D00",
INIT_14 => X"3B8000030000000000042B00009AB00008800000000008012BA010010000000D",
INIT_15 => X"0106520350000040100000000000010C0300009BA000200000000000105C0002",
INIT_16 => X"6651B328CA8D26540544924272EB91004002022024048400000098030A000A00",
INIT_17 => X"2509425094250942509425094250942509425094250942509425194651946519",
INIT_18 => X"5094250942509425094251946519465194651946519465194651946519465194",
INIT_19 => X"0480800000000000000001465194651946519465194651946509425094250942",
INIT_1A => X"34D34D34D1285B080201C92410480AB9A26667A46F345448020082E1C712A054",
INIT_1B => X"8341A0D068341A0D06834514514514514514514514514514514514514514D34D",
INIT_1C => X"F8B2B60D069349A0D068341A4D268341A4D268341A0D069349A0D069349A0D06",
INIT_1D => X"EFA2FFFFF555D000000000000000000000000000000000000000000000007FFF",
INIT_1E => X"F55087BC01EF007FD75FFFF84000AAFFD57DF45A280154BA5555401EFFFD5421",
INIT_1F => X"20AAAA843DFEF00517DEBA007BFDFEFFFD1575EF00557DF555D040000000043D",
INIT_20 => X"68AAAF7802AA00FFFBD7555087BC00AAF7D5575455D557DFEF002AAAB55002E8",
INIT_21 => X"A95545552ABFE00087BC00AA082EBFE10A28028AAAAAAABDF45F7803FFEF5555",
INIT_22 => X"FBC20BA5D7BEAAAAFFFBC00AA552E95545087BD54BA550417400085155555082",
INIT_23 => X"2FFFDF555D7BE8BFF5D51575EFA280175555D043DFEFA2FBD54BA5555554BAAA",
INIT_24 => X"00000000000557FF45002A975FF007BE8BFFA2FBFFFFFAAD5400AAFF8402000A",
INIT_25 => X"2415B471C7E3DF451EFBEFBFAF45490000000000000000000000000000000000",
INIT_26 => X"45490407000140038F450075C71FF087BD75D7FF84050BAEBDF78F45B6801048",
INIT_27 => X"FD7082EAAB550820870BAAA8438FFF00517DE82007FFAFEFE3DB505EF1C5B7AF",
INIT_28 => X"8F45F78A3DFD741516DAAAE38E2DA28EBFFD55451C7FC70BAE3D155555415178",
INIT_29 => X"1543808515756D1C2497545552AB8E10007FC50BA002ABFE00AA8A2AABABEAEB",
INIT_2A => X"FD04AA415B52492B6F5C20825D7FE8A92FFFFC20BA5D2E905550071D54825D0A",
INIT_2B => X"DB45082EB8002000AAFFFDF6D417FEABEF5D55505FFBE801256D490E3DFFFAAF",
INIT_2C => X"0000000000000000000000000000517DF451C24955EF0875EFBD7B6F1FFFC7BE",
INIT_2D => X"A2FBEAB45F78402010007BD5545AAFFD55EFF7FBE8B550000000000000000000",
INIT_2E => X"FAAFFC01FF557FE8B550004174105D042AB550055555FF007BD7555F784174AA",
INIT_2F => X"BAAAD15754508556AB45002AA8B450800174BAA68028BEF00517FE10007BE8BF",
INIT_30 => X"E10AAAEA8ABAF7AAAAB45F7AEBFF4508557FEAAAAAEBFEAAAAFFD5545557FD54",
INIT_31 => X"0145005557400552A954BA0051575EF5504175555D2EA8A00087BD74BA082EBD",
INIT_32 => X"021FF002ABDFEFAAFBC00BA007BC0000FFD542000557FE8A00F3FFC00BA552E8",
INIT_33 => X"57DF55FFD57DF55FFFBD5400A28400010A2FBFDFFF007FE8BFF5551401EFF784",
INIT_34 => X"000000000000000000000000000000000000000000000517FF455D04155FF005",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000040000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(9),        -- Port A data input
DOA(0)   => data_read_a_hi(9),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(9),        -- Port B data input
DOB(0)   => data_read_b_hi(9),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_10_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000B0001800002840002C0000281800020030000000033022000000180006",
INIT_01 => X"0000098218302849180060000C00424040000000080000080200090008510200",
INIT_02 => X"0801080200100000044008000080000041000000002002400800000009008010",
INIT_03 => X"0001000004000040000202000000000802006400088000003080040008C10000",
INIT_04 => X"0000100022008000000C08C00C00000400201830040000040000000400001820",
INIT_05 => X"0200000040000000248080210044000400000000000800000004004010000800",
INIT_06 => X"0030040000404004000006D00008002010100000880800001000000030829000",
INIT_07 => X"02100000021008000940800001800010200018920206C01020200002440003C0",
INIT_08 => X"0084010110120010004000000000021F00000024400000008000440080040000",
INIT_09 => X"8288880010100001200852882004404000000008800000100001004202000280",
INIT_0A => X"0000008000020008100004590111824004000100000008012000401084080200",
INIT_0B => X"AC04400022808001200014000040001082800000000010500000010400808000",
INIT_0C => X"002200002000020002200022000020000100011082442000480909220001E020",
INIT_0D => X"0080000010044000000080080001800200000400020011000000200002000220",
INIT_0E => X"001000020001000020010010248000200010000800040000008009040000002A",
INIT_0F => X"0000000A00010200800000001400008200800000001400000000024008208041",
INIT_10 => X"0000000024008200100000001400008200100000001400002800000000000000",
INIT_11 => X"0000000000000000001400012000200000000000000000C10008400080000000",
INIT_12 => X"8000000000480000040002040000001000000000000000000004800000002800",
INIT_13 => X"0000001000000002408000000000000000000025000200020000000001200000",
INIT_14 => X"0000040000000000000029000010000200000000000000012000001000000009",
INIT_15 => X"0100000000001000000000000000010401000010000000000000000000540002",
INIT_16 => X"00001400080002100544924002A000004000020000080000000010032A000000",
INIT_17 => X"4010040100401004010040100401004010040100401004010040000000000000",
INIT_18 => X"0000000000000000000001004010040100401004010040100401004010040100",
INIT_19 => X"1080800000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"8A28A28A28D532A0CCC2A28A28A7AA344854A07F069CB8930AFD6A1AAA902A14",
INIT_1B => X"4CA6532994CA6532994CA28A28A28A28A28A28A28A28A28A28A28A28A28A28A2",
INIT_1C => X"FB3CC772B94CA6532994CA6572B95CAE532994CA6532995CAE572B94CA653299",
INIT_1D => X"55A2AABFFEF0800000000000000000000000000000000000000000000000401F",
INIT_1E => X"4BA5555401EFFFD5421EFA2FFFFF555D003FE10AAFBE8AAAA2D540000F7D57DF",
INIT_1F => X"00AAFF8002155AAFFE8B45AAD540000087FFDF45FFFBC2010AAD57DF45A28015",
INIT_20 => X"D5400FFD568B555D00155EF08040000000043DF55087BC01EF007FD75FFFF840",
INIT_21 => X"43DFEF00517DEBA007BFDFEFFFD1575EF00557DF555D517FEBA082A801EFF7FB",
INIT_22 => X"2AAAB55002E820AAAA803FEBA082AAAAAAF7FBFDE00A2FBC0145005168A10AA8",
INIT_23 => X"FAEAAB55AAD568B455D00154BAFFFBD75EF5D7BC00AAF7D5575455D557DFEF00",
INIT_24 => X"000000000002ABDF45F7803FFEF555568AAAF7802AA00FFFBD7555082E82155F",
INIT_25 => X"AAAD547038EBD57DF7DA2AEB8FC7000000000000000000000000000000000000",
INIT_26 => X"38A2DF78F45B68010482415B471C7E3DF451EFBEFBFAF4549003DE10BEF5EDAA",
INIT_27 => X"1FF087BD75D7FF84050BAEB8002155BEF5EDB6DAADF470280075FFF45E3F1C70",
INIT_28 => X"DEAA0824851EFEBFBD2410EBD168B7D410A175C7000407000140038F450075C7",
INIT_29 => X"C2155005F68A10A28438FFF00517DE82007FFAFEFE3DB505EF1C5B7AF45495B7",
INIT_2A => X"155555415178FD7082EAAB550820870BAAA8038EAA0824A8AAAEBF5FAE28AAF1",
INIT_2B => X"FFD55451C2087155EBA4A8B7DAADF68B7D4104104AAF7F1D75EF557FC70BAE3D",
INIT_2C => X"00000000000000000000000000002EB8F45F78A3DFD741516DAAAE38E2DA28EB",
INIT_2D => X"00043FE00F7D17FEBAA2D5574BAAAD17DFEFA2AEAAB550000000000000000000",
INIT_2E => X"A00557FF45A2D5554AAA2FBEAB45F78402010007BD5545AAFFD55EFF7FBE8B55",
INIT_2F => X"105D042AB550055555FF007BD7555F784174AAA28002155FFD17FFFFA2FBD74B",
INIT_30 => X"1FF557FE8B55007FFDEAA0004175FFA2FBC2000AAD16ABFF002A975450004174",
INIT_31 => X"AABAAAD56AABAAAD140155087FEAA10A28028BEF00517FE10007BE8BFFAAFFC0",
INIT_32 => X"555EF557FD54BAAAD15754508556AB45002AA8B450800174BAA68428AAA08042",
INIT_33 => X"57FEAAAAAEBFEAAAAFFD5545550015555A2842ABEFAAFBE8BFF0004020AAFFD5",
INIT_34 => X"0000000000000000000000000000000000000000000002AAAB45F7AEBFF45085",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000047FFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(10),        -- Port A data input
DOA(0)   => data_read_a_hi(10),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(10),        -- Port B data input
DOB(0)   => data_read_b_hi(10),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_11_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10180B05A0010402840602C2D001019000000300000000330A20080EC180002",
INIT_01 => X"AB400984B830084C1820E0000C36424840000000080000088200000802112220",
INIT_02 => X"8801081438106400A4F55800008000004100000040CCE24208005000C9060032",
INIT_03 => X"000406A492E6E440842254D002108153432004800880000030C0315688C00006",
INIT_04 => X"00001201200090001205400000000094108C322644240C840008030440111800",
INIT_05 => X"222000444008010028404002A002009402400025080880000C04223000170900",
INIT_06 => X"0431018040014804920906C74B32002012121004540816544522008200821100",
INIT_07 => X"3A5B1220421408004A56E840008B90D0200018B60A0650D450FC800644A0438A",
INIT_08 => X"0485816170760268E04000000000323F42C50826490640D28088445B0E041900",
INIT_09 => X"820F8B2C100000808120308020024002B3B01AC9540080A623213008800A0280",
INIT_0A => X"10000080D80381881000045B0511D28D94012671272008013002000220001240",
INIT_0B => X"8811865D22BB384100E010908060349322008000A1001C49A9348498B0808010",
INIT_0C => X"50639504395063950639504395062CA821CA8210A0040000480808214001A020",
INIT_0D => X"088812203360410110A40008553980021040465602023269400A202863950439",
INIT_0E => X"01160006000101004A01811064B050204810240812241280D00200A08044290A",
INIT_0F => X"1B0482A01AAEC3602330CD2A02952DC3502330CB4A0318B41400024008208041",
INIT_10 => X"1630144C0155C3502330CD2A02952DC3602330CB4A0318B5600C587149B6D014",
INIT_11 => X"587083B6A51005956308D1E8202C436375908AA840AD4513437640F15245B455",
INIT_12 => X"67062F47B2872400044959BC42B1060F0D036B80B548523136C158878D8FE04E",
INIT_13 => X"7010A2699AAA3794392000D81852B0A050C224180062085134CD1719564E020C",
INIT_14 => X"400C50500D94C8121713C02B555101C90705D71009604140C0418CE0C378F0B2",
INIT_15 => X"27C828E024D8C50965A40821568A06113801505010334AA73AA0666DAC20AD57",
INIT_16 => X"048123408C0822040004C248604B2100400100084008001D0113920060CDC06A",
INIT_17 => X"4812048120481204812048120481204812048120481204812048120481204812",
INIT_18 => X"8020080200802008020081204812048120481204812048120481204812048120",
INIT_19 => X"1420000000000000000002008020080200802008020080200802008020080200",
INIT_1A => X"2082082082815220A4A380000002A8313044020C0605885026853A1082100A00",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000008208",
INIT_1C => X"F83F070000000000000100800000000000000000004020000000000000000000",
INIT_1D => X"EF0855400005500000000000000000000000000000000000000000000000401F",
INIT_1E => X"AAAA2D540000F7D57DF55A2AABFFEF0804155EFAA842ABEFA280155EFFFFBC01",
INIT_1F => X"FF555D51575FFA2FFD75FF550015400FFFBFFF4508514000000003FE10AAFBE8",
INIT_20 => X"155EF0051555FF0804155FFF7D57DF45A280154BA5555401EFFFD5421EFA2FFF",
INIT_21 => X"002155AAFFE8B45AAD540000087FFDF45FFFBC2010AAD568AAAAAD142145FF80",
INIT_22 => X"7FD75FFFF84000AAFF802ABFFA2AABFE1008001540008514215555003DFFFA28",
INIT_23 => X"85142010FFAE800AA5D7BFDF45F7FFEAA0000040000000043DF55087BC01EF00",
INIT_24 => X"00000000000517FEBA082A801EFF7FBD5400FFD568B555D00155EF085168B450",
INIT_25 => X"7BE8A155EFE3FBC71FF145B42038550000000000000000000000000000000000",
INIT_26 => X"381C003DE10BEF5EDAAAAAD547038EBD57DF7DA2AEB8FC70000175EFB6802DBC",
INIT_27 => X"1C7E3DF451EFBEFBFAF45495F575FFBEF5D05EF550E15400E3F1FFF7D085B420",
INIT_28 => X"8ABAB6D145145FF84155D7085B555C71404105C7F7DF78F45B68010482415B47",
INIT_29 => X"4515549003FFC7BE8002155BEF5EDB6DAADF470280075FFF45E3F1C7038A2DB6",
INIT_2A => X"038F450075C71FF087BD75D7FF84050BAEB8428BEFBEA4BDE28140A154380051",
INIT_2B => X"0A175C7005B6DB55145140000FFAE85082417FFFF7DE3F1EFA10140407000140",
INIT_2C => X"00000000000000000000000000005B7DEAA0824851EFEBFBD2410EBD168B7D41",
INIT_2D => X"0004175FFF7803DF45FFAE955EFAAFBD55EF557BC20AA5D00000000000000000",
INIT_2E => X"0AAD17DFEF007FC20AA5D043FE00F7D17FEBAA2D5574BAAAD17DFEFA2AEAAB55",
INIT_2F => X"45F78402010007BD5545AAFFD55EFF7FBE8B55007FD75FFF7D5401EF5D2E9741",
INIT_30 => X"F45A2D5554AAA2FBEAAAAFFD555545FF8015555007FD5545550400145FFFBEAB",
INIT_31 => X"DEAA5D2E974AA00515754500003FF55FF8002155FFD17FFFFA2FBD74BA00557F",
INIT_32 => X"7FE105D04174105D042AB550055555FF007BD7555F784174AAA2842ABEFFF803",
INIT_33 => X"BC2000AAD16ABFF002A97545007FFFF45555540000FFAE97410007BFFFFFA2D5",
INIT_34 => X"0000000000000000000000000000000000000000000007FFDEAA0004175FFA2F",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000040000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(11),        -- Port A data input
DOA(0)   => data_read_a_hi(11),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(11),        -- Port B data input
DOB(0)   => data_read_b_hi(11),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_12_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50080B01BC002006940202C0DE041196A83183000000023322287E0FC000006",
INIT_01 => X"0E000C048000C048400380000007026040000000080000088200002802153231",
INIT_02 => X"2809AD0E7D180040945008040090000061800000C0E2F66009DA3D11CB148015",
INIT_03 => X"210D050012F6F8D2108216E24842005B8A20640008800000B8E0141C28851006",
INIT_04 => X"0080100022408000060DE0000066630C70241827041000040800820480001AA4",
INIT_05 => X"0240000C400000003C808003E0C8001401000000040900020904004000070800",
INIT_06 => X"00300D800C1960C4400006E10B90002018184000100804005784000130821200",
INIT_07 => X"0652428112180C03E8E5A2C800A3F018200418927E06686450FF8006460003A0",
INIT_08 => X"09840903525281D4F460409000000E3F08D1202C5C26A0719CC96CC7BF462990",
INIT_09 => X"82488BAE10000040000410802008600843001E09F00000276F81020000230280",
INIT_0A => X"00000080000C000C100204593F11A489F480067D04D40C012400080000800240",
INIT_0B => X"0800021826933E03662802B300003C13E0000000460000000000010CE0000000",
INIT_0C => X"78419784197861978419784197860CBC30CBC20000000010400808056500A080",
INIT_0D => X"201E7F3F01F40401C17E800C7F33800200000357008C0249E2DE0D7841978619",
INIT_0E => X"0F500002200004005002001408400000000000000000000053A4096F80705FA0",
INIT_0F => X"1B17B2C53F2FC16691DB587201EDDF4162B1DB527201EDDC4607024100100020",
INIT_10 => X"F2A01D5CC9794162B1DB587201EDDF416691DB527201EDDD884272592D6246FC",
INIT_11 => X"7258E995D5A825DBA569F9FF02547068618CD3CC45B7863AE7EC00D4B122A67D",
INIT_12 => X"C6CCA5C33717461C045B5B182019473D19D7CCD856106F31A683621BDFC28800",
INIT_13 => X"FB10A652CC8E3538BBA01624E51AA6C0469AC5493F5688532966471A9C5F6208",
INIT_14 => X"40041E1F5759001B4AA1853E6D5144AA9C914C8608D2724A4C4118D992B866E2",
INIT_15 => X"AD9825682D4A36C0B0B4B85112B2C4A05D3E6D5051893335EB0072AA85A4F9B7",
INIT_16 => X"000008000000821000048260020000004001DC0800000010E7F70171401DE07E",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0100401004010040100400000000000000000000000000000000000000000000",
INIT_19 => X"1080800000000000000000040100401004010040100401004010040100401004",
INIT_1A => X"249249249120780800016A28A288028DCA30444409B054A88C5890486582A210",
INIT_1B => X"86432190C86432190C8641041041041041041041041041041041041041049249",
INIT_1C => X"FBC007592C964B2592C964B2592C964B2592C964B2592C964B2592C964B2592C",
INIT_1D => X"FF55002ABEF0800000000000000000000000000000000000000000000000401F",
INIT_1E => X"BEFA280155EFFFFBC01EF0855400005555421FF00042ABEFFF8400010082EAAB",
INIT_1F => X"FFEF08556AA10000028AAAFFD15541000002ABEFFFFBD54000004155EFAA842A",
INIT_20 => X"001FF00041554555557FE005D003FE10AAFBE8AAAA2D540000F7D57DF55A2AAB",
INIT_21 => X"1575FFA2FFD75FF550015400FFFBFFF45085140000005168AAA087BFFFFF5D04",
INIT_22 => X"D5421EFA2FFFFF555D0000145082E955FF0851555FF082AA8B55F7AEA8BEF555",
INIT_23 => X"000020BAAA801541055042ABEFFFFBD5410AAD57DF45A280154BA5555401EFFF",
INIT_24 => X"000000000005568AAAAAD142145FF80155EF0051555FF0804155FFF7842AA100",
INIT_25 => X"7EB80000280824ADBD7490E28BEF080000000000000000000000000000000000",
INIT_26 => X"101C00175EFB6802DBC7BE8A155EFE3FBC71FF145B42038555F401D71C0A2DBC",
INIT_27 => X"038EBD57DF7DA2AEB8FC7005F6AA381C0A2DA82FFDB5243800002FBD7EBFBD24",
INIT_28 => X"AA82147FF8FEF410E001FF000E17555555B7AE1041003DE10BEF5EDAAAAAD547",
INIT_29 => X"ADB45F7AEA8BEF555F575FFBEF5D05EF550E15400E3F1FFF7D085B420381C5B6",
INIT_2A => X"010482415B471C7E3DF451EFBEFBFAF4549000017D142E905EF1451525C7082A",
INIT_2B => X"04105C7F7842FA381C0A00082AA8A1041041002FBEFEBFBD2410AADF78F45B68",
INIT_2C => X"00000000000000000000000000005B68ABAB6D145145FF84155D7085B555C714",
INIT_2D => X"5D7BC01555D2EBFF55A284000AA08003FF55002AA8BEF0000000000000000000",
INIT_2E => X"A08003FF55A2FBC00105D04175FFF7803DF45FFAE955EFAAFBD55EF557BC20AA",
INIT_2F => X"00F7D17FEBAA2D5574BAAAD17DFEFA2AEAAB55007BE8AAA5D2EBDE00FFFFC00A",
INIT_30 => X"FEF007FC20AA5D7BE8A005D7FEABFF002E821FF082A97555557FE8A0000043FE",
INIT_31 => X"01EF5D5142145082EBFF55F7AAAABEF5D7FD75FFF7D5401EF5D2E97410AAD17D",
INIT_32 => X"C2010A2FBEAB45F78402010007BD5545AAFFD55EFF7FBE8B550004001FF5D2A8",
INIT_33 => X"015555007FD5545550400145FF843DEAA552A82010A2AA8000008043FFFFA2FB",
INIT_34 => X"0000000000000000000000000000000000000000000007BEAAAAFFD555545FF8",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000007FFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(12),        -- Port A data input
DOA(0)   => data_read_a_hi(12),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(12),        -- Port B data input
DOB(0)   => data_read_b_hi(12),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_13_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10110A0441812402840402822007818000E00700000000330A3000000008042",
INIT_01 => X"A1400984B830C848180260000C0042404001000008220008A200100802110200",
INIT_02 => X"88010C02801040002475580400800000410000000064024608134C0CC9018034",
INIT_03 => X"00010100926220D084234212421085084300648A0880000630C0654288C10000",
INIT_04 => X"0004122122029100100C00001200009C40A83A2044360C84190BAC04E0101820",
INIT_05 => X"027000004009050064C8C00104C10184034010250089C00EB004327064B60900",
INIT_06 => X"543000004080480492A946CE1032002012125804440812541027008230821380",
INIT_07 => X"0A581424525408000AE2AA8002BC00D020003896020658FC4030000246E543AE",
INIT_08 => X"04840101107200B80040210000002ABF02450A264002C8008000441680041900",
INIT_09 => X"825A98801000008001041080200B660E30B200C8840080808065102000280280",
INIT_0A => X"00000080C90391881000145B0111A30404016003A56008012C80080200801280",
INIT_0B => X"08088C5D2288004120E80290882400908000A000A1000809A93485D610000000",
INIT_0C => X"002000000000000002000000000000001000000000000000400808154100A080",
INIT_0D => X"08000000360401021280800E400B800610C84100014224200000000020000000",
INIT_0E => X"0086000600040D045E4195104D5854284A14250A12A512A8808289840084A020",
INIT_0F => X"0949E07A80948354B6E68982167061037496E683821670620681024000000000",
INIT_10 => X"8E510B456587037496E689821670610354B6E6838216706220431961CA985D48",
INIT_11 => X"196186A91674011CE61403562274AA49CD594CF00039C7C414B6509DA2265213",
INIT_12 => X"A983014780CC8604040424A5323845932E620295879818170304B2F5002C2043",
INIT_13 => X"451654B9104A328665603148895D44E0251142B42A3D8B2A5C8825194328A2E6",
INIT_14 => X"C06A6C6A465AA0091482382B17614F2202858EE300991415B45CD5306028F019",
INIT_15 => X"52E08DC8047F17D1C7C3C02128E587D6A02B17605A130A4E8BF002258850AC5D",
INIT_16 => X"84A123508508220808048240604B2100C00022084809000D000393722A140000",
INIT_17 => X"4A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A12",
INIT_18 => X"A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A128",
INIT_19 => X"154000000000000000000284A1284A1284A1284A1284A1284A1284A1284A1284",
INIT_1A => X"BAEBAEBAEBFF6FEFEFEEEAAAAAAFBF7DDF77F9FBEFBFF9F3F0FDFCFBEFBF1228",
INIT_1B => X"5FAFD7EBF5FAFD7EBF5FAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAE",
INIT_1C => X"F800077EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF",
INIT_1D => X"00FFD140155F780000000000000000000000000000000000000000000000401F",
INIT_1E => X"BEFFF8400010082EAABFF55002ABEF08556AAAA5D043FFFFAAAABDEAA557BFDE",
INIT_1F => X"000055043DEBAF7843FFFFF7AABDF55A2AA97400AAD540155A2D5421FF00042A",
INIT_20 => X"E8B45557FD7410552EAAABAAA84155EFAA842ABEFA280155EFFFFBC01EF08554",
INIT_21 => X"56AA10000028AAAFFD15541000002ABEFFFFBD5400005568A1055043DEBAAAFF",
INIT_22 => X"D57DF55A2AABFFEF085557545FFD17DEBAA2FFE8ABAAA8428A00087BD7555FFD",
INIT_23 => X"57BEAABA5D2ABDF450851420AA5D7FD5555A2803FE10AAFBE8AAAA2D540000F7",
INIT_24 => X"000000000005168AAA087BFFFFF5D04001FF00041554555557FE005D00001555",
INIT_25 => X"7AAA4B8E824971F8E38E3DF45155EB8000000000000000000000000000000000",
INIT_26 => X"55A2DF401D71C0A2DBC7EB80000280824ADBD7490E28BEF08516DA82410A3FFD",
INIT_27 => X"5EFE3FBC71FF145B42038550E38E92EB803FFD7EBA4BDF45AAAA90410BEDF451",
INIT_28 => X"FA38490A3FE92BEFFEAB45417FD24385D2AAFA82B680175EFB6802DBC7BE8A15",
INIT_29 => X"28A10007FD557DFFDF6AA381C0A2DA82FFDB5243800002FBD7EBFBD24101C556",
INIT_2A => X"5EDAAAAAD547038EBD57DF7DA2AEB8FC700515056DE3D17FE92BEF1EFA92AA84",
INIT_2B => X"5B7AE10410E00155497FEFABA4120B8F55085B400925D7FD557DA2803DE10BEF",
INIT_2C => X"00000000000000000000000000005B6AA82147FF8FEF410E001FF000E1755555",
INIT_2D => X"00517FE00082EBDF45AA8428A10085568ABAA2FBD7545AA80000000000000000",
INIT_2E => X"5AAAE82000F7FBD5545AAFBC01555D2EBFF55A284000AA08003FF55002AA8BEF",
INIT_2F => X"FFF7803DF45FFAE955EFAAFBD55EF557BC20AA5D2EA8A00A2803DF45AA843DF5",
INIT_30 => X"F55A2FBC00105D517FEAA082EBFE10F7FFE8B55087FC00BA552ABFE10F784175",
INIT_31 => X"FE10F7D57DE00AA842AA00007FD75FFF7FBE8AAA5D2EBDE00FFFFC00AA08003F",
INIT_32 => X"D55FFAA843FE00F7D17FEBAA2D5574BAAAD17DFEFA2AEAAB550051401FFA2D57",
INIT_33 => X"E821FF082A97555557FE8A00002E82155007BFDEAA08042AB45087FC0010557F",
INIT_34 => X"0000000000000000000000000000000000000000000007BE8A005D7FEABFF002",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000067FFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(13),        -- Port A data input
DOA(0)   => data_read_a_hi(13),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(13),        -- Port B data input
DOB(0)   => data_read_b_hi(13),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_14_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10020A000180000284008280000281800000030000000033022000000580002",
INIT_01 => X"A140098018300848184860000C20C24040000000084000084200000000110200",
INIT_02 => X"88010C5A8010A600A4F558040080000041000000022C024008003CCCC9028030",
INIT_03 => X"000103A7A00904D0842242024210810803006480088000003081054288C10000",
INIT_04 => X"0000120122009000100C00000000000400A83A2044200C840000800400101820",
INIT_05 => X"020000004008010024C0C0010040000402000025000800020004207000100800",
INIT_06 => X"0430000040004804920906C20022002012120004440812541020008230821000",
INIT_07 => X"2A5A14285A15080008768A80008000D0200018B202067AF100A0000244204382",
INIT_08 => X"04850101105205380040000000000A7F42840A264920406080004400A0040900",
INIT_09 => X"8208888010000080010010802000400230B000C8840080800021100000200280",
INIT_0A => X"00000080C8038188100004590111B68404012000016008012000000000000200",
INIT_0B => X"080084452280004120400000802000908000800001000009A924810410000000",
INIT_0C => X"000000000000200000000000000200000000000000000000400808000000A080",
INIT_0D => X"080000002204010010808008000B800210404100000220200000000020000200",
INIT_0E => X"0000000600000000020181100400502048102408122412808082098400042020",
INIT_0F => X"0480040A100A42008000161C140000420080001C1C1400003201024000000000",
INIT_10 => X"39600022260042001000161C140000420010001C1C140001604E8084341CBA34",
INIT_11 => X"8082580E2B8802201014800C220A21829A302F1C024010C001124020C8C1A8A0",
INIT_12 => X"CA60CA000048228404401004418012787124648157780120B8678C000801E04E",
INIT_13 => X"001072D04730000241000CB1325E78E0186030240000083B602398000120024A",
INIT_14 => X"001EF6F4163C480481506800004000CFD55196CB012481812049495C19400009",
INIT_15 => X"248800108B8FB61A0401200845594965000000400568D0CFB780055060500001",
INIT_16 => X"048123408408220000048240604B210040000008400800B0000090022A140068",
INIT_17 => X"4812048120481204812048120481204812048120481204812048120481204812",
INIT_18 => X"8120481204812048120481204812048120481204812048120481204812048120",
INIT_19 => X"1400000000000000000002048120481204812048120481204812048120481204",
INIT_1A => X"9E79E79E79FF3BEEEEEFE79E79EFAABCDA72E47F87BDF4EBAE7CFAFBEFB28200",
INIT_1B => X"CFE7F3F9FCFE7F3F9FCFE79E79E79E79E79E79E79E79E79E79E79E79E79E79E7",
INIT_1C => X"FBFFF83F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9F",
INIT_1D => X"555D5568A105D00000000000000000000000000000000000000000000000401F",
INIT_1E => X"FFFAAAABDEAA557BFDE00FFD140155F7D17DF45AAD157400007BEAAAAAAAE955",
INIT_1F => X"ABEF085155400FFD1420100055574AAA2AA800AAF784020AAF7D56AAAA5D043F",
INIT_20 => X"FFE105D7BD7545A284020BA0055421FF00042ABEFFF8400010082EAABFF55002",
INIT_21 => X"43DEBAF7843FFFFF7AABDF55A2AA97400AAD540155A28028B550051574005D7F",
INIT_22 => X"FBC01EF08554000055002AB455D51420100851421FF5D7FFDEBA085168B45FF8",
INIT_23 => X"AD140000002EBFFEFA2AAA8BEFF780021FF5504155EFAA842ABEFA280155EFFF",
INIT_24 => X"000000000005568A1055043DEBAAAFFE8B45557FD7410552EAAABAAA8017400A",
INIT_25 => X"01C71EDA82AAA0955455D556DA00490000000000000000000000000000000000",
INIT_26 => X"BAEBD16DA82410A3FFD7AAA4B8E824971F8E38E3DF45155EBD17FF6DAADB5040",
INIT_27 => X"0280824ADBD7490E28BEF085157428FFDB420101C55554AAAAA480082FF84000",
INIT_28 => X"AB7D0051504005D71F8E004975D556DB68405092085F401D71C0A2DBC7EB8000",
INIT_29 => X"FAEAA08516AB45E38E38E92EB803FFD7EBA4BDF45AAAA90410BEDF45155A28E2",
INIT_2A => X"02DBC7BE8A155EFE3FBC71FF145B42038550028B6D5D51420101C5B401EF417B",
INIT_2B => X"2AAFA82B68015400AADB40000082EBFFC7A2AEAFBC7EB80071FF5500175EFB68",
INIT_2C => X"0000000000000000000000000000556FA38490A3FE92BEFFEAB45417FD24385D",
INIT_2D => X"AAD17DFFFAAFFC200055557DE00A2801554555557FE100000000000000000000",
INIT_2E => X"AA28400000F784020BAAAD17FE00082EBDF45AA8428A10085568ABAA2FBD7545",
INIT_2F => X"555D2EBFF55A284000AA08003FF55002AA8BEF0051554AAFFFFC00105D55554B",
INIT_30 => X"000F7FBD5545AAAEAABFF0051400105D5568A000051575FFF78415410087BC01",
INIT_31 => X"2000557FC01EF007FEAABA00556AB55A2AEA8A00A2803DF45AA843DF55AAAE82",
INIT_32 => X"175FF5D04175FFF7803DF45FFAE955EFAAFBD55EF557BC20AA5D042ABFF55514",
INIT_33 => X"FE8B55087FC00BA552ABFE10F78415400A2FBC0010082EBDF55A2AABDF45A284",
INIT_34 => X"000000000000000000000000000000000000000000000517FEAA082EBFE10F7F",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000007FFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(14),        -- Port A data input
DOA(0)   => data_read_a_hi(14),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(14),        -- Port B data input
DOB(0)   => data_read_b_hi(14),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_15_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000A000000000284000280000001800020030000000033022000000180002",
INIT_01 => X"A140098018300848180060000C00424040000000080000080200000000110200",
INIT_02 => X"080108000010E60004E55800008000004100000000040240080000C009170016",
INIT_03 => X"0000000080000040842240000210810002000400888000003080014288C00000",
INIT_04 => X"0001100024A0800000440000000000040088322044200C840000011400151800",
INIT_05 => X"A200014C4000000020000000000B8094020000254C8800000514203000108800",
INIT_06 => X"0031042040804804100006EE4032002012120005540812540020008600831000",
INIT_07 => X"021912244A14080008408880008000D020001892020656300020000244000380",
INIT_08 => X"048501415032000800406180000002DF02440826400000008000440000043080",
INIT_09 => X"8208880110000000010010802000400230A000880400808000450200000B0280",
INIT_0A => X"00000080C003010810000459011182040400200003E0080120000000000002C0",
INIT_0B => X"080084452280004100400000800000100000800001000001A124800010000000",
INIT_0C => X"002000020000000000000000000200001000010000000000400808000020A000",
INIT_0D => X"08000000260001001280000C400B000200000000000220200000000020000200",
INIT_0E => X"008400060000000000010010040040000000000000201000000000000004A000",
INIT_0F => X"0000000000000202100000000000000202100000000000004600024000000000",
INIT_10 => X"0000000000000202800000000000000202800000000000002000000800000000",
INIT_11 => X"0008000000000000000000002000100800000000000000000000400001200000",
INIT_12 => X"00880000000006000400080C0000000000D08120280000000000000000002000",
INIT_13 => X"0010040200000000010000004020010000000000000008000900000000000200",
INIT_14 => X"0000000308801400000000000040000008822110000000000040100100000000",
INIT_15 => X"0080000000004840717050000000000000000040000020000000000000000001",
INIT_16 => X"000023000000220000048240404A010040000008000000000000000020C40000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"1400000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000200",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"F800000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"AA007BC2145F780000000000000000000000000000000000000000000000401F",
INIT_1E => X"400007BEAAAAAAAE955555D5568A105D7FC00000804154AA5D00001EFF78428A",
INIT_1F => X"0155F7FBD74AAAAD17DF45F7D1421EF0055400AA007FC2000F7D17DF45AAD157",
INIT_20 => X"BDFEF08517DF55A2FBEAB555D556AAAA5D043FFFFAAAABDEAA557BFDE00FFD14",
INIT_21 => X"155400FFD1420100055574AAA2AA800AAF784020AAF7FFFDF45FF84000BA552A",
INIT_22 => X"2EAABFF55002ABEF087BE8ABA555168B55AAFFEAB45F7843FF45082A801FF005",
INIT_23 => X"284000AA0055401550055574005D2E800AAA2D5421FF00042ABEFFF840001008",
INIT_24 => X"000000000000028B550051574005D7FFFE105D7BD7545A284020BA007FFFE10A",
INIT_25 => X"2550E021C7EB8028A821C7BC516DFF8000000000000000000000000000000000",
INIT_26 => X"28FFD17FF6DAADB504001C71EDA82AAA0955455D556DA004971C703814001248",
INIT_27 => X"E824971F8E38E3DF45155EBF1D5492BED17FF45E3DF471C70851400BA0071C50",
INIT_28 => X"FF7DEB8000092552ABFFEF08517DF6DB6FBE8B555D516DA82410A3FFD7AAA4B8",
INIT_29 => X"3DF551C20801C71C5157428FFDB420101C55554AAAAA480082FF84000BAEBF1F",
INIT_2A => X"A2DBC7EB80000280824ADBD7490E28BEF087FEFA8241516DB55A2FFEAB6DEB84",
INIT_2B => X"8405092087FF8E00BE8A02082005F47145085550428412A85082BEDF401D71C0",
INIT_2C => X"00000000000000000000000000000E2AB7D0051504005D71F8E004975D556DB6",
INIT_2D => X"0055554BA5504000105D2A80145AA842AA00557BD75EFF780000000000000000",
INIT_2E => X"50055420BA0055574BAF7D17DFFFAAFFC200055557DE00A2801554555557FE10",
INIT_2F => X"00082EBDF45AA8428A10085568ABAA2FBD7545AAD557410F7D57DF55AAFBD554",
INIT_30 => X"000F784020BAAAD57FFEFA28402010552ABDFFF08517FFFFF7FBEAB455D517FE",
INIT_31 => X"DF45AAFBE8BEFA2803FF455504001555551554AAFFFFC00105D55554BAA28400",
INIT_32 => X"95400F7FBC01555D2EBFF55A284000AA08003FF55002AA8BEF007FFDE1000557",
INIT_33 => X"568A000051575FFF78415410087FEAA10F7AE80000087BD55450855400BA002A",
INIT_34 => X"0000000000000000000000000000000000000000000002EAABFF0051400105D5",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000060000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(15),        -- Port A data input
DOA(0)   => data_read_a_hi(15),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(15),        -- Port B data input
DOB(0)   => data_read_b_hi(15),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_16_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"DA22C618B1000482B688B186588884862A400438255FC38381441205BA803003",
INIT_01 => X"8645A80028404C211203A952A90341080B173340412000E1005D628000820484",
INIT_02 => X"A101A9006DC1084833011850AAC55001349B10881802821808B4110007005E11",
INIT_03 => X"010108A802BB00080080006020020001A61036202800000D2410104200404550",
INIT_04 => X"8BFA58800005C40A46240252145148B38248030356415A4E62B6FC660F287240",
INIT_05 => X"0F05EA11E570000D610000000710296E542B6E3A825C15FB30A643695BFC2D56",
INIT_06 => X"00640044150C025A0000000901A054F2C0A8030140BCC0460050690A95C8383D",
INIT_07 => X"0288500102F85203E8010D0AA9BC4800015001219D0550077373CAA804000680",
INIT_08 => X"A2064193920A2004B51400001414091EAA14881C0002701881B120203B7A8012",
INIT_09 => X"C8204D02D965965200100104F2B0082251200000023153000C4400800000ACCA",
INIT_0A => X"000012C9000A0000D0A80000BF8028E87C1B9246002A8A562060410280081116",
INIT_0B => X"240014891801000495D40192D1000000000000A8A5AA80018120E00066000000",
INIT_0C => X"00088000880008800088000880008400044000400029011404008401CA809004",
INIT_0D => X"0140A80A5C8000102ED0044008004AD32400004001AB08C0031EDA7B08800088",
INIT_0E => X"04912AA28AA890BA00000024800480000000000000200802151025062C0BB400",
INIT_0F => X"1F554E11C596A64003195933741477264003195555B418687E35836020814004",
INIT_10 => X"0A499CF47DCB264003195933741597264003195555B4198843940076D296D003",
INIT_11 => X"00758486A556489347FE5F409CBC1362510695B6288743123C95251852041CD5",
INIT_12 => X"424EAE2992046EB70026486035600CEC45CBCA809654B48163CCC895E1E043D4",
INIT_13 => X"98E3A242DEA151848302BFD6D522B10C7EC71F6C1DB071D1216E078C4C1B1C74",
INIT_14 => X"037DAAABC982BE22267A2E2E4F44AA1DC5E37400C9EE1B7B638E8849D23C3832",
INIT_15 => X"2EE015998B28654565A003F0068E35352C1CAE48BFBF3A6C9B7B286B4DA8B93D",
INIT_16 => X"000009000040A8000452110A8442040D655602A102A0027E2C42320284086E6A",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"1451451451E96F2FC3C34F3CF3C2AC688AA263486D3260E34C0C3A7B451B0200",
INIT_1B => X"9F47A7D1E9F47A7D1E9F4D14D14D14D14D14D14D14D14D14D14D14D14D145145",
INIT_1C => X"F800007D3E9F4FA7D3E8F47A3D1E8F47A3D1E8F47A7D3E9F4FA7D3E9F4FA7D3E",
INIT_1D => X"FF00003FE005500000000000000000000000000000000000000000000000401F",
INIT_1E => X"4AA5D00001EFF78428AAA007BC2145F7843FFFFF7FBE8B45AAD568BFFFFAA975",
INIT_1F => X"8A105D2E974BAF7FBEAB45FFFFC00BAF780020005D2A95410FFFFC0000080415",
INIT_20 => X"821FFA2AAAAA00000417555FFD17DF45AAD157400007BEAAAAAAAE955555D556",
INIT_21 => X"BD74AAAAD17DF45F7D1421EF0055400AA007FC2000F78000010552E800AA002E",
INIT_22 => X"7BFDE00FFD140155F7AABDF55F7AE820AA08043FEBA5D55575FFF7AABFE00557",
INIT_23 => X"2FBE8B55FFFFD55FF557FC2000FF8015410FFD56AAAA5D043FFFFAAAABDEAA55",
INIT_24 => X"000000000007FFDF45FF84000BA552ABDFEF08517DF55A2FBEAB555D04154BAA",
INIT_25 => X"5B6DF6DBFFF7AA955C71C043FE10490000000000000000000000000000000000",
INIT_26 => X"38FFF1C7038140012482550E021C7EB8028A821C7BC516DFF8438FC7E3F1EAB5",
INIT_27 => X"A82AAA0955455D556DA00492490492F7FBE8B55FFF1C70BAF78A000005D20974",
INIT_28 => X"20285D2085092002A801FFB6AAA8A10080E1757DEBD17FF6DAADB504001C71ED",
INIT_29 => X"555FFE3AABFE005D71D5492BED17FF45E3DF471C70851400BA0071C5028FF840",
INIT_2A => X"A3FFD7AAA4B8E824971F8E38E3DF45155EBA4BAF6DE3AA8709208043FEBA555B",
INIT_2B => X"FBE8B555D04124BAB6FBE8B45E3FBD55D7557BC0028E38412428EBD16DA82410",
INIT_2C => X"000000000000000000000000000071FFF7DEB8000092552ABFFEF08517DF6DB6",
INIT_2D => X"F78428B55AAD168B55F7FFFDFEFFFAA9555555003DE000000000000000000000",
INIT_2E => X"AFFAE820105500154AAF7D5554BA5504000105D2A80145AA842AA00557BD75EF",
INIT_2F => X"FFAAFFC200055557DE00A2801554555557FE10000000010F7FBEAB45FFD1554A",
INIT_30 => X"0BA0055574BAF784000BA5D0017410082E801EFF7AEA8A10002E955FFA2D17DF",
INIT_31 => X"541000003DEBA557BD75EFA2AEBDE105D5557410F7D57DF55AAFBD5545005542",
INIT_32 => X"000AAAAD17FE00082EBDF45AA8428A10085568ABAA2FBD7545AA802ABEFA2AA9",
INIT_33 => X"ABDFFF08517FFFFF7FBEAB455D04020AAFFFBEAB45AAFFD55555D7FC20AAA280",
INIT_34 => X"000000000000000000000000000000000000000000000557FFEFA28402010552",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000020000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(16),        -- Port A data input
DOA(0)   => data_read_a_hi(16),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(16),        -- Port B data input
DOB(0)   => data_read_b_hi(16),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_17_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"5284CE4FB7BD2C8994A13392DBD02E14006B82AC7E800D44D3DD2FD5F9B961C0",
INIT_01 => X"F8ACD01F7E03FC6793F2199B39FC233C11D93AE6F3BB92B32091DBC339B24542",
INIT_02 => X"8F333007FD6808092A2AFA6667033DB50853379C10BFF70F1BD011110F205F18",
INIT_03 => X"294ADB4AFFCBF0DAD63ABF836B58EAFE060478202022234B2E0303FDC9E18339",
INIT_04 => X"DB7A40806FE4040840EBC563A0150A0926146FECB04196482236FC2005282AE1",
INIT_05 => X"0403DA0383200831C68206D7E6D0250834336D1E81500FDB306045255BFC2076",
INIT_06 => X"000A0E2D7D3EAFF15800100FBFB333C1CBC303163670497AFF00291B3C0E2015",
INIT_07 => X"451C581123AEE54DE8008B719E61C10BBA5DAAFA9DDA1194D51E067BB0000000",
INIT_08 => X"70320A9392083056C2270E004400091181168C4D14002A110C902481FC0B4212",
INIT_09 => X"0E28EFFC40C30E5F0182D0950190C0810BE00E9A76E4C7FD0E4700000B303806",
INIT_0A => X"C7DEF207000F00059D2ED56D7EED2ED3C9A86FB8013E7437823DF78CDB6CA60E",
INIT_0B => X"7C00319F8E853E64D73A08BFF0001D35682AC0CE8FCCC200A59BDD2FFE3F3EC7",
INIT_0C => X"7A7DE7A7DE7A7DE7A7DE7A7DE7A7DF3D3EF3D3C0030B889723782E816EC0A081",
INIT_0D => X"2D4CFEB69FF7A5F5AFFCCA787F7FE67C21800367451F8355EB9EDE7A7DE7A7DE",
INIT_0E => X"2C9F99FD0678B87A0003000D8D02E00000000000000040025D3C21463D6BFF25",
INIT_0F => X"232221ABD9CA854DFDD64A67D42C0F054DFDD64667D42C063E57A8F7B4594BB0",
INIT_10 => X"AEDAA504801F054DFDD64A67D42C0F054DFDD64667D42C07237DFE5865F6D2BF",
INIT_11 => X"FE58EAE7F5AB50D0806A9A2E0DFFF47DEDC496DA3181A0CC71440F9FBC3EFBB5",
INIT_12 => X"9C9C3FC95949AEFF556EF9C75E7DCF1EB1B6E6FCDC87CB35FC94B36AECF3A33D",
INIT_13 => X"382AF5B6AAAE594A4C0DBFDAD94AA669809809FEFAF4157ADB55572CA527056E",
INIT_14 => X"1AE33F32ADD543430808BABAF50E1A5EB4BAEA45A250202FE0ADD39387F92B29",
INIT_15 => X"669523E865D4B1293AB6B90BF2F0E30EDEFAFD0B3FBD72E9E90D20A003FBEBF4",
INIT_16 => X"00002F840000BCE0B6F67B3F845E017C833F6AAC02B002A2EFF22D4073DE83FB",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0600000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"9A69A69A6A4624C3434C0EBAEBA21B9001804F6E62029749701020B88A7CC0C0",
INIT_1B => X"41A0D46A341A0D46A341A69AEBA69A69AEBA69AEBA69A69AEBA69AEBA69A69A6",
INIT_1C => X"F8000046A351A8D46A351A8D46A351A8D46A351A8D068341A0D068341A0D0683",
INIT_1D => X"00F7D56ABFF55000000000000000000000000000000000000000000000007FFF",
INIT_1E => X"B45AAD568BFFFFAA975FF00003FE0055043FFFFFFFFFFFFFF7FBFDF55A284020",
INIT_1F => X"2145F7D568B45000002010552EBDF45A28028A00F7843FEBA55043FFFFF7FBE8",
INIT_20 => X"95410AAAEBFF55AAFFC00BAF7FFC00000804154AA5D00001EFF78428AAA007BC",
INIT_21 => X"E974BAF7FBEAB45FFFFC00BAF780020005D2A95410FFAE800105D2A95410002A",
INIT_22 => X"AE955555D5568A105D7FFFFEFA2D568BFFFFD57DE00F7AE800AAAAAABDFEF5D2",
INIT_23 => X"82A974105D003FF55F7802AAAAAAD168AAA5D517DF45AAD157400007BEAAAAAA",
INIT_24 => X"000000000000000010552E800AA002E821FFA2AAAAA00000417555FF8028B550",
INIT_25 => X"FE3F5FAF45AA8000038F7DB6FBD7490000000000000000000000000000000000",
INIT_26 => X"82490438FC7E3F1EAB55B6DF6DBFFF7AA955C71C043FE10490A3FFFFFFFFFDFE",
INIT_27 => X"1C7EB8028A821C7BC516DFFDF68B551C0E050384124BFF7DB68A28A38F7803DE",
INIT_28 => X"5000492495428082E95400AAA0BDF7DB6F5C70BAFFF1C7038140012482550E02",
INIT_29 => X"800BAB6AEBDFD75D2490492F7FBE8B55FFF1C70BAF78A000005D2097438FFAA8",
INIT_2A => X"B504001C71EDA82AAA0955455D556DA00497FFAFFFB6D56FBFFEBDB78E38F7AA",
INIT_2B => X"0E1757DEB8A2DB5514249243841003FF6DEB8028AAAB6D16FA8249517FF6DAAD",
INIT_2C => X"000000000000000000000000000004020285D2085092002A801FFB6AAA8A1008",
INIT_2D => X"002ABFFEFF7FBFDFFFAAD168B55AA80000BAF7FFFDF550000000000000000000",
INIT_2E => X"FFFAAA8AAAF7843FE10000428B55AAD168B55F7FFFDFEFFFAA9555555003DE00",
INIT_2F => X"BA5504000105D2A80145AA842AA00557BD75EFF7FBEAB45552E954BA08003DFF",
INIT_30 => X"0105500154AAF7AE974000800154AA002E95410AA843FFFFF7D5554BAF7D5554",
INIT_31 => X"FFEFAAFFE8ABAFFAA820BAF7AEBFF55550000010F7FBEAB45FFD1554AAFFAE82",
INIT_32 => X"7DE0000517DFFFAAFFC200055557DE00A2801554555557FE10007FEABEFFFD57",
INIT_33 => X"E801EFF7AEA8A10002E955FFA2AABFF455500020AA08003DFFFA28028AAAF7D1",
INIT_34 => X"00000000000000000000000000000000000000000000004000BA5D0017410082",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000067FFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(17),        -- Port A data input
DOA(0)   => data_read_a_hi(17),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(17),        -- Port B data input
DOB(0)   => data_read_b_hi(17),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_18_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"69844019080000A21A611406840014122A641074155FC28A2024001001801003",
INIT_01 => X"A643D920034004180005E9E3C90360C0041C0181002001602025800008440084",
INIT_02 => X"B7333980808408103F2000F81FC0FEDEAC2161B0B84D0002188011110C018041",
INIT_03 => X"0405D434003F2C020081587008020561E55116B0290000042B71240C800440F8",
INIT_04 => X"50805AC31007D6125724029216554A9847669903D640EC8E2001002604503004",
INIT_05 => X"07008000E0EA11803850C800010022660C1C0065003C0404002646DC20A02D40",
INIT_06 => X"8560000000022229A60B048048120FF040000000002C44D620F0228454C83810",
INIT_07 => X"058800A001D4033A004904087F9E3901218050018024110D6771C1F90C285682",
INIT_08 => X"F3020A82929A807B3731021400058C020000A9729400D10100420480202AC214",
INIT_09 => X"C820C802D86184A010180304307008025414204400220202F1A814A0080064C1",
INIT_0A => X"080003C32A10A19090C02010E10229440616900000022E0C6070000504102805",
INIT_0B => X"026226495446E2110AE44174112840880000060D7030C30B885200D274004008",
INIT_0C => X"840018400184001840018400184000C2000C200200301500C404C001B884B806",
INIT_0D => X"81010108003C000210020460801001FB3650D89888E06CAE1061018500184001",
INIT_0E => X"032007E281F840C00284A17210001060D8306C18360C1380A0260CB980840080",
INIT_0F => X"5D79BBEF8E50B041029075982BF3873041029079982BF39748AA0AC800014804",
INIT_10 => X"EA479BFD7F7F3041029075982BF3E73041029079982BF3F632C5F96D3C11555D",
INIT_11 => X"F96A595405FC7F1CFEBC7586C4100A53162B47FD7E39FFEECE1598702345156A",
INIT_12 => X"006FE037ACFB88083A99E06271BB0CA207DFDD5920057E0B001B0EBCC79932C5",
INIT_13 => X"5CA2A002DD51B6F7FC4A411D1E8D44517F14EAFE36E55150016EA8DB73E39464",
INIT_14 => X"953C30351452A13D55CFFA76E928E3891F148B30399F5FB7F28C800DFA06F5DF",
INIT_15 => X"5AC57DFEAEF1005475F1D1F608819CF0EE76E12C824ADD9089715F25FAF9DB84",
INIT_16 => X"0D834041A41A0000010180C02801680460FC900052FA10DC0006DA4881C11015",
INIT_17 => X"D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D836",
INIT_18 => X"8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360",
INIT_19 => X"00000000000000000000020D8360D8360D8360D8360D8360D8360D8360D8360D",
INIT_1A => X"8A28A28A2891182C8A82E0820825945DF675C0770B9E11807E54587BEF8B0000",
INIT_1B => X"44A2552A954AA5128944AAAA28A28A28AAAAAAA28A28A28AAAAAAA28A28A28A2",
INIT_1C => X"F80000128944A25128944A25128944A25128944A25128944A25128944A251289",
INIT_1D => X"BA5D04174AA0000000000000000000000000000000000000000000000000401F",
INIT_1E => X"FFFF7FBFDF55A28402000F7D56ABFF55043FFFFFFFFFFFFFFFFFFFFEFF7AE954",
INIT_1F => X"FE0055043FFFFFFFFFDFEFA2D56AB45AA8400145AA801741000043FFFFFFFFFF",
INIT_20 => X"FFFFFFF80021EF0855421EF00043FFFFF7FBE8B45AAD568BFFFFAA975FF00003",
INIT_21 => X"568B45000002010552EBDF45A28028A00F7843FEBA55557FFEFA2D168B55AAFB",
INIT_22 => X"8428AAA007BC2145F7D5400000004020AA5D2A82155F7AEBFEBAFFD56AA00A2D",
INIT_23 => X"82E954BA0004174AAAA8428B45082ABFEBAA2FFC00000804154AA5D00001EFF7",
INIT_24 => X"000000000002E800105D2A95410002A95410AAAEBFF55AAFFC00BAF7AE800100",
INIT_25 => X"FFFFBFDFEFFFAE954AA550415492140000000000000000000000000000000000",
INIT_26 => X"10140A3FFFFFFFFFDFEFE3F5FAF45AA8000038F7DB6FBD7490E3FFFFFFFFFFFF",
INIT_27 => X"BFFF7AA955C71C043FE1049043FFEFE3F1F8FD7AAD16FB6DBE8E00155BE80154",
INIT_28 => X"8FC7AAD56FB6DBEF1FAFD7E384001EF145B471C7140438FC7E3F1EAB55B6DF6D",
INIT_29 => X"BDE92FFD56FA28B6DF68B551C0E050384124BFF7DB68A28A38F7803DE82495B7",
INIT_2A => X"012482550E021C7EB8028A821C7BC516DFFD1420381C0A02082492A85155E3A4",
INIT_2B => X"F5C70BAFFAE870280024904BA1400174AABE8E28B7D1420BDEAAA2F1C7038140",
INIT_2C => X"00000000000000000000000000002A85000492495428082E95400AAA0BDF7DB6",
INIT_2D => X"002ABFFFFFFFFFFFEFF7FBFDFFFF7AA974BA5504154105500000000000000000",
INIT_2E => X"FF7AA82155F78015400552ABFFEFF7FBFDFFFAAD168B55AA80000BAF7FFFDF55",
INIT_2F => X"55AAD168B55F7FFFDFEFFFAA9555555003DE0000043DFEFA2D56AB45AAD57DFE",
INIT_30 => X"AAAF7843FE10007FEAB55A2D17FFEFFFD568B55A280021EF557FD7555550428B",
INIT_31 => X"2000002A95545A2843FE00F7D17FEAAF7FBEAB45552E954BA08003DFFFFFAAA8",
INIT_32 => X"3DEAAA2D5554BA5504000105D2A80145AA842AA00557BD75EFF7D1400AA5D2A8",
INIT_33 => X"E95410AA843FFFFF7D5554BAF7AE974BA0004020AA5D04154BAF7AEA8BEF5500",
INIT_34 => X"0000000000000000000000000000000000000000000002E974000800154AA002",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000020000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(18),        -- Port A data input
DOA(0)   => data_read_a_hi(18),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(18),        -- Port B data input
DOB(0)   => data_read_b_hi(18),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_19_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"042200000000000041088001001AA00000000000000000000000500802000003",
INIT_01 => X"200048000024000000000404000000000A22000800000800004A200000000001",
INIT_02 => X"032210008DEF00400060000001C008002489E0F0004037B00010101010000000",
INIT_03 => X"0000008128000000000000000000000024001620280000000000354200004008",
INIT_04 => X"000058800004C4024024001210001054B1C822009640000E2000002604003000",
INIT_05 => X"07008000E0200000000000000000200604000000001C04000026400000002C40",
INIT_06 => X"000000000000000100000000000001B040000000002C42010010200004C83810",
INIT_07 => X"0E0050A040041593104004500480090080A01120220140020420401800000000",
INIT_08 => X"130E409080188000021A0000100004082A140102B4020109801A4CE003710010",
INIT_09 => X"C80000005861840000000004301000B000000000001C1C0000000000000020C0",
INIT_0A => X"000002C30000000040500010301020400000000000022A040000000000000004",
INIT_0B => X"00000020001000022000000000000000000002F0001F00002024B20002000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"00108000EC000000000000000010004B20000000000000000000000000000000",
INIT_0E => X"0000006280180040000000000000000000000000000000000000000000000000",
INIT_0F => X"8084451B81A70AB3006BA0011400760AB3006BA0011400680F02096834820000",
INIT_10 => X"11204082248A0AB3006BA0011400160AB3006BA0011400084C780687DBA82800",
INIT_11 => X"068796E80A00802301BC0A7531EDD98E73B02800804620D030F873EB49F30B80",
INIT_12 => X"6B00000002044F091A860700FF9198AA115D5DA37F7A80C8A3604001C0664C78",
INIT_13 => X"98551AC9000000000314E01F9F30198600631448410A2A8D64800000081B0A93",
INIT_14 => X"2E00303842281C80A23004411AD661891F15148A4420804241526D6000000000",
INIT_15 => X"9D335F3D282000C6C5456C84850F61050C411AD6284FDA861682805A04A1046B",
INIT_16 => X"00000000000000000000000000000004600C0013800003088004202304366A4A",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"86186186186851046260A9A69A6039045DD1F863808633005010063A20C90000",
INIT_1B => X"D26930984C26130984C261861861869A61861861861869A61861861861861861",
INIT_1C => X"F800000984C26130984C26130984C26130984C26130984C26130984C26130984",
INIT_1D => X"BA5500020BA5D00000000000000000000000000000000000000000000000401F",
INIT_1E => X"FFFFFFFFFFEFF7AE954BA5D04174AA007BFFFFFFFFFFFFFFFFFFFFFFFFFAA954",
INIT_1F => X"ABFF557BFFFFFFFFFFFFFFFFFBFDFEFFFAA974BA5D517FFFF08043FFFFFFFFFF",
INIT_20 => X"6AB45AA8002000F7D5575455D043FFFFFFFFFFFFFF7FBFDF55A28402000F7D56",
INIT_21 => X"43FFFFFFFFFDFEFA2D56AB45AA8400145AA8017410007BFFFFFFFFFFFFEFF7D1",
INIT_22 => X"AA975FF00003FE00557BFFFFFFFFBFDF45AAD568B55F7AE955FFAA8402010080",
INIT_23 => X"7D168B55AAD17FFEFF7AE975FF00557FFFF5D043FFFFF7FBE8B45AAD568BFFFF",
INIT_24 => X"00000000000557FFEFA2D168B55AAFBFFFFFFF80021EF0855421EF002ABFFEFF",
INIT_25 => X"FFFFFFFFFFF7AA954BA550000082550000000000000000000000000000000000",
INIT_26 => X"C7080E3FFFFFFFFFFFFFFFFBFDFEFFFAE954AA5504154921471FFFFFFFFFFFFF",
INIT_27 => X"F45AA8000038F7DB6FBD74975FFFFFFFFFFFFEFF7FBFAFD7E3A4954BA555B7AF",
INIT_28 => X"FFFFF7FBF8FC7EBD568B55A28000000FFDF52545550A3FFFFFFFFFDFEFE3F5FA",
INIT_29 => X"955C7BE800000008043FFEFE3F1F8FD7AAD16FB6DBE8E00155BE8015410147FF",
INIT_2A => X"1EAB55B6DF6DBFFF7AA955C71C043FE10497BFDFC7E3F1FAF55A2DB6FB7DF7AE",
INIT_2B => X"5B471C71424B8FC7E3D56AB6DB6DF7AFC7EBA0955FF145B7AFC7410438FC7E3F",
INIT_2C => X"00000000000000000000000000005B78FC7AAD56FB6DBEF1FAFD7E384001EF14",
INIT_2D => X"55517FFFFFFFFFFFFFFFFFFFFEFF7AA974AA5500020005500000000000000000",
INIT_2E => X"5AA80154AA557BEAB45002ABFFFFFFFFFFFEFF7FBFDFFFF7AA974BA550415410",
INIT_2F => X"EFF7FBFDFFFAAD168B55AA80000BAF7FFFDF5500517FFFFFFFBFDFEFFFFFEAB4",
INIT_30 => X"155F78015400557BFDFEFF7FBEAB55A2D56AB55A28002000F7FFC2155552ABFF",
INIT_31 => X"8B45AAFBFFFFFFFAA95545F7840201000043DFEFA2D56AB45AAD57DFEFF7AA82",
INIT_32 => X"E8B55000428B55AAD168B55F7FFFDFEFFFAA9555555003DE00007FFDF45AAD56",
INIT_33 => X"568B55A280021EF557FD755555042AB55AAD16ABFFFFFBEAB45A280155EF557F",
INIT_34 => X"0000000000000000000000000000000000000000000007FEAB55A2D17FFEFFFD",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000040000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(19),        -- Port A data input
DOA(0)   => data_read_a_hi(19),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(19),        -- Port B data input
DOB(0)   => data_read_b_hi(19),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_20_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000003",
INIT_01 => X"A75FF80000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"14088080800008400F655001FFCFF80018FA8044000000000000011000000007",
INIT_03 => X"0000000000000000000000000000000024001660380000000000000000004FF8",
INIT_04 => X"000079800014CC02C034001600000000000000101EC0012EE0C0026E1E80F000",
INIT_05 => X"1F0FF433EFF0440C3902100002203F2EFC040388137C3E20C8EEC00284033CC0",
INIT_06 => X"00F00100002E22EB440012C809B2FFF7C8E8840155FDC0000010E40087D8787A",
INIT_07 => X"03B800000000000000008407FC800B0000000100600040000C205FF91C000F80",
INIT_08 => X"F28C0B0300020852000002101554021F00000000000000009049226020000200",
INIT_09 => X"D80000007BEFBC010002008FF7F00000000010018A81000041C401000004FFDF",
INIT_0A => X"00000ADF000000200000008000008028300100461003EAFE400000120000913F",
INIT_0B => X"0000000000000000000000000200200290000000000000000200000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000010001000000",
INIT_0D => X"00000100000010000002000080101FFB60000000000000000000000000000000",
INIT_0E => X"03007FE29FF800C00000001002040000000000000020480002E42429C0000080",
INIT_0F => X"0004D4E180010040000400000001E60040000400000001E6010003C000000000",
INIT_10 => X"000000094B1E0040000400000001E60040000400000001E60804000000400000",
INIT_11 => X"00002000000000033628000100100000004000000006170C0008001000004000",
INIT_12 => X"000000000295810000000A100020614148002000000000004307CC3CC0000804",
INIT_13 => X"5802000000000014AC000120200000000003F0D800020100000000000A4B0020",
INIT_14 => X"0020C0C00000000002E2D000001006204040000000005786C004000000000052",
INIT_15 => X"0100A0C0939BEE1810080200000E0CE0EC000010020000000000000AE8A00002",
INIT_16 => X"2008040400400C08080000000000049F6FFC0100000000000008008008000400",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0100000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0C30C30C320624C1090D0F3CF3CD038001801C10000804482A60D09008269020",
INIT_1B => X"90C86432190C86432190CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2C30C3",
INIT_1C => X"F80000432190C86432190C86432190C86432190C86432190C86432190C864321",
INIT_1D => X"AA5504020100800000000000000000000000000000000000000000000000401F",
INIT_1E => X"FFFFFFFFFFFFFFAA954BA5500020BA5D7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974",
INIT_1F => X"74AA00003FFFFFFFFFFFFFFFFFFFFFFF7AA974AA550002000007BFFFFFFFFFFF",
INIT_20 => X"FDFEFFFAE974AA5D003FE005D043FFFFFFFFFFFFFFFFFFFFEFF7AE954BA5D041",
INIT_21 => X"BFFFFFFFFFFFFFFFFFBFDFEFFFAA974BA5D517FFFF087FFFFFFFFFFFFFFFFFFF",
INIT_22 => X"8402000F7D56ABFF55003FFFFFFFFFFFFFF7FBFDFFFAA84000105D556AB55557",
INIT_23 => X"FFFFFFEFF7FBEAB55A28000010F7D16ABEF08043FFFFFFFFFFFFFF7FBFDF55A2",
INIT_24 => X"000000000007BFFFFFFFFFFFFEFF7D16AB45AA8002000F7D5575455D2EBFFFFF",
INIT_25 => X"FFFFFFFFFFFFAE974AA550400028000000000000000000000000000000000000",
INIT_26 => X"380071FFFFFFFFFFFFFFFFFFFFFFFF7AA954BA550000082557FFFFFFFFFFFFFF",
INIT_27 => X"FEFFFAE954AA55041549214043FFFFFFFFFFFFFFFFFFDFEFF7AE974BA5500050",
INIT_28 => X"FFFFFFFFFFFFFF7FBFDFFFFFAA974BA550038E285D0E3FFFFFFFFFFFFFFFFBFD",
INIT_29 => X"02028555F6FB7D5D75FFFFFFFFFFFFEFF7FBFAFD7E3A4954BA555B7AFC70871F",
INIT_2A => X"FFDFEFE3F5FAF45AA8000038F7DB6FBD7490E3FFFFFFFFFDFEFF7F1FAFC7A280",
INIT_2B => X"DF525455524BFFFFFFFBFDFC7E3F5E8B45A28402010FFDB6ABEF140A3FFFFFFF",
INIT_2C => X"00000000000000000000000000007FFFFFFF7FBF8FC7EBD568B55A28000000FF",
INIT_2D => X"557FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5504000BA0800000000000000000",
INIT_2E => X"FFFAE954BA5500174AA08517FFFFFFFFFFFFFFFFFFFFEFF7AA974AA550002000",
INIT_2F => X"FFFFFFFFFEFF7FBFDFFFF7AA974BA55041541055043FFFFFFFFFFFFFF7FBFDFE",
INIT_30 => X"4AA557BEAB4500557FFFFFFFFFDFEFF7FFFFFEFF7AE974AA550028AAA5D2ABFF",
INIT_31 => X"DFEFFFD568B55A284020BA557FFFFFF5D517FFFFFFFBFDFEFFFFFEAB45AA8015",
INIT_32 => X"EABEF5D2ABFFEFF7FBFDFFFAAD168B55AA80000BAF7FFFDF55002EBFFFFF7FBF",
INIT_33 => X"56AB55A28002000F7FFC215555043DFEFF7FBFFF55A2D16AB45AA8402000F7FB",
INIT_34 => X"0000000000000000000000000000000000000000000007BFDFEFF7FBEAB55A2D",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000007FFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(20),        -- Port A data input
DOA(0)   => data_read_a_hi(20),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(20),        -- Port B data input
DOB(0)   => data_read_b_hi(20),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_21_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"4A302428B824900A128C090A5C1800261500213C005FE812D10420054085A202",
INIT_01 => X"081FFE3440B609703B0427F801A40B8115BC4F655300340288A40D30040E4DD8",
INIT_02 => X"0109095C30C98809800000F9FFFFFFFF149FF1FCA4C0421B182E3490DF145FE4",
INIT_03 => X"084A76341244919000099486400026523C041660BA000100CC12701015007FF8",
INIT_04 => X"000079800014CC03C075161E001118653D2408041FC004AEF000816E1C11F541",
INIT_05 => X"3F0F807BFFE000240100004683103E7FFE02482553FC3C0204EFC25010143CC0",
INIT_06 => X"008808210996035A000006EC2E04FFFFC0A0000101FFE4036450E08247F87870",
INIT_07 => X"4003400812A156C002822987FC830F40134CC74D002016612DE87FFE00400804",
INIT_08 => X"F02348D2D00080C0C53400044114000000D022640B42406808790055043A8282",
INIT_09 => X"F84056387FEFBC110008420F7FF388B70A20389346FE9F26120200800008FDFF",
INIT_0A => X"4518DBFF00020004C0A6044901112A0908AA14601DE3EBFE0A812D8D5B742D3F",
INIT_0B => X"104032901CC63410ABD249C4B3007127080806FF917FC30010107688862A28C5",
INIT_0C => X"46C9146C9146C9146C9146C9146CC8A3648A3642003184822040D000D8C41807",
INIT_0D => X"201800500941044312000900D4621FFBE0008A94C822CA8919018206C9146C91",
INIT_0E => X"2029FFEADFF8050250010030165290008800440022201082401A002000C48000",
INIT_0F => X"18048A004A6C0D2820302C005A83480D1820302A009B02B101390C0CB2830816",
INIT_10 => X"1408904831400D1820302C005A83480D2820302A009B02B021A85C0941150013",
INIT_11 => X"5C08834600024D052C1051E0B92D400360520202682C19024B6164E300448510",
INIT_12 => X"6404093E22A2012418A9D1D44ADD9E0F174103820101C0B8160D5516259FA1A8",
INIT_13 => X"60D8AA288209E615100280DA0052000C5006402000206C55144104D510CC1B0D",
INIT_14 => X"0A0D50020C04023033C52009144231D902818100C90058010361AC808126C886",
INIT_15 => X"2202386454988140600C0181500A13E830011008B0374007000B4E0CD0002450",
INIT_16 => X"0080224004002000000703804008001F7FFF01B982B01258088C008CC41198A1",
INIT_17 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_18 => X"8020080200802008020080200802008020080200802008020080200802008020",
INIT_19 => X"0000000000000000000002008020080200802008020080200802008020080200",
INIT_1A => X"BEFBEFBEFBFF7FEFEFFFE79E79FFFF7CFF77FBFFEFBFF9F7E0FDF9EFEFBF0000",
INIT_1B => X"DFEFF7FBFDFEFF7FBFDFEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEF",
INIT_1C => X"F80000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"BA5D00020000800000000000000000000000000000000000000000000000401F",
INIT_1E => X"FFFFFFFFFFFFFFAE974AA550402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974",
INIT_1F => X"20BA5D7FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5D00020AA5D7FFFFFFFFFFFF",
INIT_20 => X"FFFFFF7AA974BA5D0402000557BFFFFFFFFFFFFFFFFFFFFFFFFFAA954BA55000",
INIT_21 => X"03FFFFFFFFFFFFFFFFFFFFFFF7AA974AA55000200000003FFFFFFFFFFFFFFFFF",
INIT_22 => X"AE954BA5D04174AA00003FFFFFFFFFFFFFFFFFFFFEFF7AE974BA5D00174BA000",
INIT_23 => X"FFFFFFFFFFFFFDFEFF7AE954AA5500174BA5D043FFFFFFFFFFFFFFFFFFFFEFF7",
INIT_24 => X"000000000007FFFFFFFFFFFFFFFFFFFFDFEFFFAE974AA5D003FE005D2EBFFFFF",
INIT_25 => X"FFFFFFFFFFFFAE974BA5D0000010000000000000000000000000000000000000",
INIT_26 => X"BA557FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550400028007FFFFFFFFFFFFFF",
INIT_27 => X"FFFF7AA954BA550000082557BFFFFFFFFFFFFFFFFFFFFFFFFFAA954BA5D00000",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFEFF7AA974AA5D04050005571FFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"954BA5D00154AA00043FFFFFFFFFFFFFFFFFFDFEFF7AE974BA55000503800003",
INIT_2A => X"FFFFFFFFFBFDFEFFFAE954AA550415492140E3FFFFFFFFFFFFFFFFFFDFEFF7AE",
INIT_2B => X"0038E285D2ABFFFFFFFFFFFFFFFFBFDFEFFFAA974BA5D00104925D0E3FFFFFFF",
INIT_2C => X"000000000000000000000000000071FFFFFFFFFFFFFFF7FBFDFFFFFAA974BA55",
INIT_2D => X"087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D00000100000000000000000000",
INIT_2E => X"FF7AA954BA5D00000BA5D7FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5504000BA",
INIT_2F => X"FFFFFFFFFFFFFFFFFFEFF7AA974AA550002000557BFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA5500174AA08043FFFFFFFFFFFFFFFFBFDFEFF7AE954AA5D041740055517FF",
INIT_31 => X"FFFFF7FBFDFFFFFAA974AA5D00174BA08043FFFFFFFFFFFFFF7FBFDFEFFFAE95",
INIT_32 => X"00010552ABFFFFFFFFFFFEFF7FBFDFFFF7AA974BA550415410552ABFFFFFFFFF",
INIT_33 => X"FFFFEFF7AE974AA550028AAA5D2EBFFFFFFFFFDFEFF7FBFFFFFF7AE954BA5D00",
INIT_34 => X"000000000000000000000000000000000000000000000557FFFFFFFFFDFEFF7F",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(21),        -- Port A data input
DOA(0)   => data_read_a_hi(21),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(21),        -- Port B data input
DOB(0)   => data_read_b_hi(21),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_22_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"5290F4CDE914905A14A43D33F488243E17122300F55FEB189B343A1140548380",
INIT_01 => X"A94007B259F6A975386262000C344BA9573C6FF57B18A5FB0ABFCD3C2C5F4F0C",
INIT_02 => X"877FE30EB378008D202551040030071869D0040180AC4B685F6E26FAA0810006",
INIT_03 => X"431965109E4481D6B5AAD6875AD6AB5A1815600802888808DEA83552954D3000",
INIT_04 => X"492C0020220001010E4916C884DCD607E5EC2A344103E48003D0800023D0072C",
INIT_05 => X"00107C441001100D620A06D683018001023D37E5088043620101179092540112",
INIT_06 => X"40111C2D50A46AE45281502E4A2200081ADA0E054402365774611E047020008E",
INIT_07 => X"680BD5AA4BF5C91F840C1710010344DB9A808FDFF3DE0313014A200754040180",
INIT_08 => X"0EA212D6D481ADF0CE47CA21544009007A64EBD64049D028B93D9561A48F6027",
INIT_09 => X"207246A80400015805060040080A2A0F4A82381B4000BFB65A0283800AA50020",
INIT_0A => X"4539C020E11810098D4067EFF9FF284D483E35602820110204804818CD280100",
INIT_0B => X"10081E9528963546278008AA800470370000A0004D0000002126F30C902A29C5",
INIT_0C => X"40E1540E1540E1540E1540E1540E4AA070AA07000A0000308000190168200281",
INIT_0D => X"6870A9CA0D458D131652A154D46B600085080B14009A2B2906504940E1540E15",
INIT_0E => X"448C00044000A1EC1C44140D101A54280A14050A028500A84F02842A24C594A0",
INIT_0F => X"38359E0C4E6C256690581800F1C3E82562B0581200F1C3F08145602280402080",
INIT_10 => X"100AB8581B602562B0581800F1C3E8256690581200F1C3F1238473F121000613",
INIT_11 => X"73F0E1050083750B3E4275F829547008600C030374361FA2CEE046D48122C438",
INIT_12 => X"C4CC012A66F61154C019511628756231018500C00203E1380615651607822384",
INIT_13 => X"608AA612C0096C37B00D1724801A0009C606D1221D104553096004B61BCC1128",
INIT_14 => X"12A41E0F0600035842E7601C2C4AC68A98810080AA825A890225189980254CDE",
INIT_15 => X"A89637E00D0A1080301401C390320188321C2C0B13890105800D520AF94870B0",
INIT_16 => X"88222F110111B281A54753AA004002601001918008C10912A4440B24E8B58234",
INIT_17 => X"8220882208822088220882208822088220882208822088220882208822088220",
INIT_18 => X"2008020080200802008020080200802008020080200802208822088220882208",
INIT_19 => X"1448000000001FFFFFFFFC802008020080200802008020080200802008020080",
INIT_1A => X"9E79E79E7BFF3FEFEBEEEFBEFBEFBEFDFEF7F47F8FBEF5EB7E6CFEFBEFBE8289",
INIT_1B => X"CFE7F3F9FCFE7F3F9FCFE79E79E79E79E79E79E79E79E79E79E79E79E79E79E7",
INIT_1C => X"F800003F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9F",
INIT_1D => X"BA5D04000000000000000000000000000000000000000000000000000000401F",
INIT_1E => X"FFFFFFFFFFFFFFAE974BA5D0002000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974",
INIT_1F => X"2010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA550000010007FFFFFFFFFFFF",
INIT_20 => X"FFFFFFFAE954AA5D00000AA007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA55040",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5D00020AA5D7FFFFFFFFFFFFFFFFFFF",
INIT_22 => X"AA954BA5500020BA5D7FFFFFFFFFFFFFFFFFFFFFFFFFFAA954BA5504000AA557",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFAA954BA5500000BA5D7BFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"00000000000003FFFFFFFFFFFFFFFFFFFFFFF7AA974BA5D040200055517FFFFF",
INIT_25 => X"FFFFFFFFFFFFAE974BA5D0402000080000000000000000000000000000000000",
INIT_26 => X"10087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0000010007FFFFFFFFFFFFFF",
INIT_27 => X"FFFFFAE974AA550400028007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA5500020",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFAE954AA5D00020BA087FFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"954BA5504020AA5D7BFFFFFFFFFFFFFFFFFFFFFFFFFAA954BA5D00000BA557FF",
INIT_2A => X"FFFFFFFFFFFFFFFF7AA954BA5500000825571FFFFFFFFFFFFFFFFFFFFFFFFFAA",
INIT_2B => X"040500055517FFFFFFFFFFFFFFFFFFFFFFF7AA974AA5D00070925D71FFFFFFFF",
INIT_2C => X"0000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFEFF7AA974AA5D",
INIT_2D => X"007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020000800000000000000000",
INIT_2E => X"FFFAE974AA550002000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0000010",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFAE954AA5504000BA087FFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA5D00000BA5D7BFFFFFFFFFFFFFFFFFFFFFFFFFAA954AA5D00020AA007FFFF",
INIT_31 => X"FFFFFFFFFFFEFF7AA974BA5504020BA557BFFFFFFFFFFFFFFFFFFFFFFFF7AA95",
INIT_32 => X"154105D517FFFFFFFFFFFFFFFFFFFFEFF7AA974AA55000200055517FFFFFFFFF",
INIT_33 => X"BFDFEFF7AE954AA5D041740055557FFFFFFFFFFFFFFFFFFDFEFF7AE974AA5D00",
INIT_34 => X"000000000000000000000000000000000000000000000043FFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000007FFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(22),        -- Port A data input
DOA(0)   => data_read_a_hi(22),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(22),        -- Port B data input
DOB(0)   => data_read_b_hi(22),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_23_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"EF20906D902424807BC8241BC81801B97D38AD3C0800103362A6741C80A12A02",
INIT_01 => X"001FFF8409F089003B4422000D80C80106804A7951C5B9D1C828043EA28838F9",
INIT_02 => X"073B8858218C2C50801000F9FFEFF8E72CA7F5FC2E048026496834D84721DFE0",
INIT_03 => X"2C4360101A4001001005080400401420350016E0BB222341C312000014006FF8",
INIT_04 => X"00017B810015DC03D034201E14000036486008101FC0002EE006297E1C05F561",
INIT_05 => X"BF0F817FFFE80100004044800080BEFFFC0248005FFC3C18A5FFC2444484BCC0",
INIT_06 => X"0400000409120338860900482404FFFFC000000001FFC0832050E00047F97870",
INIT_07 => X"200246801C41C3E81E872C8FFE900FC31348EFDF03BE15E22DA07FF92C204102",
INIT_08 => X"F6220280D2B025988311AB14155421006891A1089F6E200000022C140068EB90",
INIT_09 => X"F8001011FFEFBC80000000077FF184B03010004002FE000000201000000FFDFF",
INIT_0A => X"00001BFFA800808189A657EF81DD0C00079CD00837C3EBFD4201258112D4487F",
INIT_0B => X"24483890564084198AD249C433200180082A06FF907FC3081812048006000000",
INIT_0C => X"8608086080860808608086080860804304043042003184822150C000D8C41806",
INIT_0D => X"03000100200180480000095280001FFBF040C088CD20E0A21921828608086080",
INIT_0E => X"3821FFEAFFF805025E00853B92588000400020001000020A8018008002000014",
INIT_0F => X"486148484054395E27E428002A4200397E07E422002A420100382FCC30832A16",
INIT_10 => X"0C0788417000397E07E428002A4200395E27E422002A420110A51C01C0590401",
INIT_11 => X"1C01A2490040590C08120558C1759BE1C05A0400383808800DA1929F72864110",
INIT_12 => X"20000136006000215EA0A4833A32C8832050028603050014031B3950000C90A5",
INIT_13 => X"006658280009A2030108B14AC05C00112405222088B8332C140004D101800CE7",
INIT_14 => X"196B6808060201281004228996085F10020180C030880D11019CE4000026C00C",
INIT_15 => X"52A49DC7143F01C04240030720641E0A028996483A17204680410A04104A2659",
INIT_16 => X"0401000080080000000000002001201F7FFC0011C2F81A48080CA32800A01081",
INIT_17 => X"4010040100401004010040100401004010040100401004010040100401004010",
INIT_18 => X"0100401004010040100401004010040100401004010040100401004010040100",
INIT_19 => X"0000000000000000000000040100401004010040100401004010040100401004",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"F800000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"BA5D04020100000000000000000000000000000000000000000000000000401F",
INIT_1E => X"FFFFFFFFFFFFFFAE974BA5D0400000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974",
INIT_1F => X"2000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400010087FFFFFFFFFFFF",
INIT_20 => X"FFFFFFFAE974BA550002000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D000",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA550000010007FFFFFFFFFFFFFFFFFFF",
INIT_22 => X"AE974AA550402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550400000087",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFAE974AA550402000087FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5D00000AA007FFFFFFF",
INIT_25 => X"FFFFFFFFFFFFAE974BA5D0402010000000000000000000000000000000000000",
INIT_26 => X"10087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000087FFFFFFFFFFFFFF",
INIT_27 => X"FFFFFAE974BA5D0000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04000",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFAE974BA550002000007FFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974AA550400010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550002010087FF",
INIT_2A => X"FFFFFFFFFFFFFFFFFAE974AA550400028007FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_2B => X"00020BA087FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5D0402038007FFFFFFFFF",
INIT_2C => X"00000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5D",
INIT_2D => X"087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020100000000000000000000",
INIT_2E => X"FFFAE974BA5D0400000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D0000010007FFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4AA550002000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA550002010087FFFF",
INIT_31 => X"FFFFFFFFFFFFFFFAE954AA550400010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_32 => X"000AA087FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5504000BA087FFFFFFFFFFF",
INIT_33 => X"FFFFFFFFAA954AA5D00020AA007BFFFFFFFFFFFFFFFFFFFFFFFFFAA954AA5D04",
INIT_34 => X"0000000000000000000000000000000000000000000007BFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000007FFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(23),        -- Port A data input
DOA(0)   => data_read_a_hi(23),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(23),        -- Port B data input
DOB(0)   => data_read_b_hi(23),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_24_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100600007FFF000080108004000800020000840041000080808",
INIT_02 => X"172A00D000EF8210000000F9FFEFF8E7240FF1FC224087B1000639401D005FC0",
INIT_03 => X"00003A2E200811000000000400000000340016603A0000004860400014006FFF",
INIT_04 => X"000079800014CC03C034001E04010850300000101FC0002EE000006E1C00F500",
INIT_05 => X"1F0F8033FFE000000000000000003E2FFC024800137C3C0000EFC00000003CC0",
INIT_06 => X"0000000009120110020100002404FFFFC000000001FFC0000010E00007F87870",
INIT_07 => X"200102050840950002802C87FC800FCAA035400001B918600C207FF800000000",
INIT_08 => X"F6234AD280B02500063AC2840001610020408178B600C2400013649608730004",
INIT_09 => X"F80000007FEFBC00000000077FF000B00000000002FE0000000000000000FDFF",
INIT_0A => X"00001BFFA0000005501AA00000CE20000094000011C3EBFC020125811254083F",
INIT_0B => X"0040A040004000008012414433000100080806FD107FC3000000000006000000",
INIT_0C => X"0608006080060800608006080060800304003042003180822040C00090C41806",
INIT_0D => X"004800B0000000000000000000001FFBE0008080C820C0801801800608006080",
INIT_0E => X"2021FFEADFF80002080000000208800000000000000000020018000000000000",
INIT_0F => X"840009181008024A00043601100210024A00043C0110020901382CCCB28B0806",
INIT_10 => X"180040A03080024A00043601100210024A00043C01100209240C840C201D0210",
INIT_11 => X"840A604E0080820009908008341B000A8212070082002890010068320860C920",
INIT_12 => X"40600800082041205EC00044C1ACB66C37542082030281E0580001012811A40C",
INIT_13 => X"80B27A004300004103160DB3005E000618040C022000593D002180002090166B",
INIT_14 => X"2BBFF20406040084210C062000C2A2DDD00180C04504086002CD680C01000104",
INIT_15 => X"20804295C98F80400008040CC0582169022000C2876C40478002850016088001",
INIT_16 => X"0000000000000000000000000000001F7FFC001B823018F00880008805241060",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"9EF9EF9EFB263CC3090CABAEBAFF96857757B73E6089966B9EF9D5A220CC8000",
INIT_1B => X"C1E0F0783C1E0F0783C1EFBEFBEFBE79E79E79E79E79EFBEFBEFBEFBEFBEF9EF",
INIT_1C => X"F800000783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783",
INIT_1D => X"BA5D04020100800000000000000000000000000000000000000000000000401F",
INIT_1E => X"FFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974",
INIT_1F => X"0000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000087FFFFFFFFFFFF",
INIT_20 => X"FFFFFFFAE974BA5D0400000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400010087FFFFFFFFFFFFFFFFFFF",
INIT_22 => X"AE974BA5D0002000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0000010007",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFAE974BA5D0002000007FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA550002000007FFFFFFF",
INIT_25 => X"FFFFFFFFFFFFAE974BA5D0402010080000000000000000000000000000000000",
INIT_26 => X"00087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFF",
INIT_27 => X"FFFFFAE974BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000007FFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA5D0000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400010087FF",
INIT_2A => X"FFFFFFFFFFFFFFFFFAE974BA5D0000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_2B => X"0002000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA550002000087FFFFFFFFF",
INIT_2C => X"00000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA55",
INIT_2D => X"007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020100800000000000000000",
INIT_2E => X"FFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA5D0400000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000007FFFF",
INIT_31 => X"FFFFFFFFFFFFFFFAE974BA5D0000010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_32 => X"00010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0000010007FFFFFFFFFFF",
INIT_33 => X"FFFFFFFFAE974BA550002010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5500",
INIT_34 => X"0000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(24),        -- Port A data input
DOA(0)   => data_read_a_hi(24),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(24),        -- Port B data input
DOB(0)   => data_read_b_hi(24),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_25_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100200002000000080100004000000020000800041000080808",
INIT_02 => X"1000218000000800000000F9FFEFF8E738FFF1FC20400400000004455A375FE0",
INIT_03 => X"00002000000001000000000400000000340016623A0000004000000014006FFF",
INIT_04 => X"924279824C94CC1BE0B4001F20000000020380401FE0082EF000106E1C00F500",
INIT_05 => X"1F0F8033FFF048202582800100523E2FFE024820137C3C0040EFE02000003CE4",
INIT_06 => X"10DC00CC0992033A062116E82404FFFFC0E0801101FFC0000010E08A07FC7870",
INIT_07 => X"000000000000000002802C87FC800F8000000000019810600C207FFF3C410D84",
INIT_08 => X"FE8002000080281000008A0000014100200081000000000080480AE000000200",
INIT_09 => X"FC0020007FEFBE031018C31F7FFBAEBC0020008086FE0000100280800000FDFF",
INIT_0A => X"00001BFFE00301000000000000CC02000014000191C3EBFF4A7DF795965C6D3F",
INIT_0B => X"0040200000400000801243443B000100880806FD107FC3018000000006000000",
INIT_0C => X"0608006080060800608006080060800304003042003B99862444E61492C41806",
INIT_0D => X"00000000000000000000001280001FFBE0008080C820C4801801800608006080",
INIT_0E => X"3021FFEADFF805025C0304001E58906088304418222C108A009A090400000000",
INIT_0F => X"00000100100000480000200100000000480000200100000100380F0C30830A06",
INIT_10 => X"0000008000000048000020010000000048000020010000000004040000010000",
INIT_11 => X"0400004000000000008080000011000000020000000020000000001200000100",
INIT_12 => X"000000000800002018C010000020800000800122000000004004000008000004",
INIT_13 => X"0002080000000040000001020020000000000800200001040000000020000021",
INIT_14 => X"0021000008001000000800200000021000020100000000200004200000000100",
INIT_15 => X"0000008400000000605000000000200000200000020400000000000002008000",
INIT_16 => X"288226410410346010000000400A011F7FFE0031823010400800000800001840",
INIT_17 => X"8822088220882208822088220882208822088220882208822088220882208822",
INIT_18 => X"8220882208822088220882208822088220882208822088220882208822088220",
INIT_19 => X"00017FFFFFFFFFFFFFFFFE088220882208822088220882208822088220882208",
INIT_1A => X"2410492410A048029890AD34D35FDD144A50CB5462D14997BE09E760AED04040",
INIT_1B => X"8C46231188C46231188C49249249249249249249249241041041041041041049",
INIT_1C => X"F80000B158AC562B158AC562B158AC562B158AC562B158AC562B158AC562B158",
INIT_1D => X"BA5D040201000000000000000000000000000000000000000000000000007FFF",
INIT_1E => X"FFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974",
INIT_1F => X"2010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFF",
INIT_20 => X"FFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000087FFFFFFFFFFFFFFFFFFF",
INIT_22 => X"AE974BA5D0400000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000007",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFAE974BA5D0400000087FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000007FFFFFFF",
INIT_25 => X"FFFFFFFFFFFFAE974BA5D0402010000000000000000000000000000000000000",
INIT_26 => X"10087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFF",
INIT_27 => X"FFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA5D0402000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000087FF",
INIT_2A => X"FFFFFFFFFFFFFFFFFAE974BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_2B => X"0400000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000087FFFFFFFFF",
INIT_2C => X"00000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D",
INIT_2D => X"087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020100000000000000000000",
INIT_2E => X"FFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFF",
INIT_31 => X"FFFFFFFFFFFFFFFAE974BA5D0402000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_32 => X"02000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000087FFFFFFFFFFF",
INIT_33 => X"FFFFFFFFAE974BA5D0400000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_34 => X"0000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000007FFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(25),        -- Port A data input
DOA(0)   => data_read_a_hi(25),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(25),        -- Port B data input
DOB(0)   => data_read_b_hi(25),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_26_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"E9264EAB20190CA3BA4997AA9002AE9C001006B0778015CFA17E0811039879C7",
INIT_01 => X"F1FFF9BB1F773C7F9BB07DFFFDD863FC5FFF3FEFFBBF9FFB22FFFBC7B9F30686",
INIT_02 => X"1B33188302E708180F6FFBFFFFCFFFFF9C7FF7FC24350B99082400001D00DFD8",
INIT_03 => X"4A53D958C50000DCE7366303739CD98C27C57EF57980014F271807E3C9E9CFF8",
INIT_04 => X"DBFAFBD7FB1CDEBEF1BE17F7AC88042787FBFFF8FEE9FF7EE6F4C0EE1FFAF869",
INIT_05 => X"5F0FFEB3EFFEFFBDA7F7FED508707E2EFEBF6FFEB37C3FF302EEEDFF9B487CF6",
INIT_06 => X"AFBE564C71268F3BBF5FBFC2A427FFF7C3E3A74667FDDB7FB870FF30FFDEF87F",
INIT_07 => X"03BC18306396FBEC14489737FDC00B13BB79DFDB83BF4112AF205FFBDD3AFB93",
INIT_08 => X"F21E4391909B381B0B1F8E041051831FA3068D77E000030021324620C0B9C206",
INIT_09 => X"DE89ECC0FBEFBEBF30B8D79FF7F451F33CFD60FE8FFFDF58003B1D4223B4FFDF",
INIT_0A => X"8ED6BFDF3EB3EBF9DDBCE7FDC1DF8A760F3EB980580BFAFFF37DF7B9DF7DCB3F",
INIT_0B => X"6EE6F5E7FAC4C03DB856CD4CF73AC1FC98884FFF19FFC71FEFED7B251E35768E",
INIT_0C => X"06BC606BC606BC606BC606BC606BD3035E3035C62B7BB987666DEF8A90CCFA8F",
INIT_0D => X"CF6100C0E60FB9FC3A80EF69A04DFFFF7FF5F9A0DC33E9B41D01D207BC606BC6",
INIT_0E => X"7027FFFF9FF8FAFAA3ADEBFB9726BAF5FD7AFEBD7F7EFFD7ACDB7F947F0EA035",
INIT_0F => X"E020080A40403E8BD8002000FC02003E8BD8002000FC02010979AFFE36C36B86",
INIT_10 => X"000EE00034003E8BD8002000FC02003E8BD8002000FC020037B0040A00010003",
INIT_11 => X"040C00400003D80008160400FD81341C00020003B80008C00801EF0285380100",
INIT_12 => X"90981038406809677FA080468C46A81080581002000780C8001C8100201037B0",
INIT_13 => X"00F90D162001C803411FC0024080001F80040026C0807C868B1000E401A01F11",
INIT_14 => X"3F810503A00003E020042AC080CEB01228A80000F600080123E232130407080D",
INIT_15 => X"0087520750001064180807868000110C02C080CFA0042400000F8800105B0201",
INIT_16 => X"7FDFF7EFEEFF3EEC3FF7FBFFBCB7FFFFEFFE00BFF7FEBF420800EC0CBEE61F81",
INIT_17 => X"FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F",
INIT_18 => X"D7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5",
INIT_19 => X"43237FFFFFFFFFFFFFFFFF5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5F",
INIT_1A => X"A69A61861BAF15EAA6AFC38E38EA3AD8ADE7A48F0B366429F434AA9FC376DAE4",
INIT_1B => X"C26130984C26130984C261861861861861861861861861861861861861861869",
INIT_1C => X"F800000984C26130984C26130984C26130984C26130984C26130984C26130984",
INIT_1D => X"BA5D04020100000000000000000000000000000000000000000000000000401F",
INIT_1E => X"FFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974",
INIT_1F => X"2010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFF",
INIT_20 => X"FFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFF",
INIT_22 => X"AE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFF",
INIT_25 => X"FFFFFFFFFFFFAE974BA5D0402010000000000000000000000000000000000000",
INIT_26 => X"10007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFF",
INIT_27 => X"FFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FF",
INIT_2A => X"FFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_2B => X"0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFF",
INIT_2C => X"00000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D",
INIT_2D => X"007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020100000000000000000000",
INIT_2E => X"FFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFF",
INIT_31 => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_32 => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_33 => X"FFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_34 => X"0000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(26),        -- Port A data input
DOA(0)   => data_read_a_hi(26),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(26),        -- Port B data input
DOB(0)   => data_read_b_hi(26),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_27_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"00080A40000A41248002029000050A088000008242A0004404480002000A1155",
INIT_01 => X"F1FFF1C11F781C129C107DFFFE0860941E81258CA2B71C2220EC1B86E1A00002",
INIT_02 => X"4000002100000014400FF6FFFF0FFFFF8007F1FC211100014200800000887FC0",
INIT_03 => X"0842D85841000098C63061026318C18404C459757000015F00088BE3C0618FF8",
INIT_04 => X"DBEAE5D6D91C2EBCE1B21EA72C00000007FBE7C8F8E9EF79E6D440E91FDAE061",
INIT_05 => X"5C8FFCB38FF6B68984B5BCE408347E28FEBF6FEEB3723F7102E8EDBF8A4872F6",
INIT_06 => X"AB98420C71408D113956AFD0842FFFC7C3032646EFF1DB7FA868FE30EF1CE47E",
INIT_07 => X"10041830600640C415004637FC4003021259CFDB01BF80028E001FF8251AB9D1",
INIT_08 => X"F200822020842203000082050000110023068D03000002820000000840000005",
INIT_09 => X"1C852440E3DF7E2FB0B8E717C7F411F3BC6D60B60FFDDE480018AC4AA3B0FD1F",
INIT_0A => X"18109E1F16B16B71092CE7ED81CF403601229880400BE0FC137FF7A0FF75813F",
INIT_0B => X"86F7D5E382A440349816DD4C755AC16C1A884FFE18FFD757E7ED7A211E81C098",
INIT_0C => X"061A2061A2061A2061A2061A2061E1030D1030D6A37FB9872E65E6AA90CD5AAF",
INIT_0D => X"8FC10080A20ED1D41880CC61A044DFFC6EB5BCA0DE31F8B41C01E0071A2061A2",
INIT_0E => X"2023FFE91FF98AEAA1AC6AC9A3A4AAD5B56ADAB56D5AFD572C597B147506203E",
INIT_0F => X"E020000260403C8948002000EC0000BC8948002000EC00010878AC3CB8AB8857",
INIT_10 => X"000EE0000400BC8948002000EC0000BC8948002000EC000097B0040200010003",
INIT_11 => X"040400400003D80000070400DD81041400020003B80000410801AF0204180100",
INIT_12 => X"101010384008086378A080428C46A80080081002000780C800188000301017B0",
INIT_13 => X"02E909042001C800409FC0020080001F80000007C0807484821000E400205D11",
INIT_14 => X"3F810100A00003E020000BC0808EB01020280000F60000002BA2220204070801",
INIT_15 => X"0007520750000024080807868000100403C0808FA0040400000F8800001F0200",
INIT_16 => X"5B5EF3AF6AF6389C2FE128971AB2DDDF8FFE0031B776BF4208006C0C92621F81",
INIT_17 => X"B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D",
INIT_18 => X"56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5",
INIT_19 => X"43A3FFFFFFFFFFFFFFFFFD5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B",
INIT_1A => X"0000000001E0080397908000000A48710B4080240E543021B438A010825238B4",
INIT_1B => X"0804020100804020100800000000000000000000000000000000000000008200",
INIT_1C => X"F80000A05028140A05028140A05028140A05028140A05028140A05028140A050",
INIT_1D => X"BA5D04020100000000000000000000000000000000000000000000000000401F",
INIT_1E => X"FFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974",
INIT_1F => X"2010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFF",
INIT_20 => X"FFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFF",
INIT_22 => X"AE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFF",
INIT_25 => X"FFFFFFFFFFFFAE974BA5D0402010000000000000000000000000000000000000",
INIT_26 => X"10007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFF",
INIT_27 => X"FFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FF",
INIT_2A => X"FFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_2B => X"0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFF",
INIT_2C => X"00000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D",
INIT_2D => X"007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020100000000000000000000",
INIT_2E => X"FFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_31 => X"FFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_32 => X"02010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFF",
INIT_33 => X"FFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_34 => X"0000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000007FFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(27),        -- Port A data input
DOA(0)   => data_read_a_hi(27),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(27),        -- Port B data input
DOB(0)   => data_read_b_hi(27),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_28_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"02200AA400180030808802A900002A08001280A08A801044104A1000001818C3",
INIT_01 => X"50A00011460214428114180000882214413D0A71592A01D92213D28005210202",
INIT_02 => X"1444428102100884000AA30200000000C1000401041108404400022220800000",
INIT_03 => X"461080404900000C6314A900318C52A40051081000888806108802A141288001",
INIT_04 => X"00800040110102000902002000888400081045A8A00003C00000500000080008",
INIT_05 => X"0000000000024CA0A0101800032000400000000B800000014000000B08180000",
INIT_06 => X"814016012000C405280200008001000011110012220009A88800009A88000000",
INIT_07 => X"0004891224228810080010200040001020800000004000008200000240081400",
INIT_08 => X"00A010040401080308400821155540001122448142491008A004912040840221",
INIT_09 => X"0020405000000124058200408000880004440004080160C8100A858009940000",
INIT_0A => X"4D29400002002038104000000020003204000880082800010000000C0000E400",
INIT_0B => X"12220122A000416811040000400800081022C0000080000206CB0821082B694D",
INIT_0C => X"80B0280B0280B0280B0280B0280B01405814058009000421833010800A000200",
INIT_0D => X"C4210040860B188C0A8065302005A004039010280001001600200081B0280B02",
INIT_0E => X"500600010000280000802050010660001000080004004900204020105302A000",
INIT_0F => X"0000000A00000081480000001400000081480000001400000800C01082082210",
INIT_10 => X"0000000024000081480000001400000081480000001400000010000200000000",
INIT_11 => X"0004000000000000001400000080041400000000000000C00000010004180000",
INIT_12 => X"1010100000480802A40000000400000080081000000000000004800000000010",
INIT_13 => X"0001010420000002400040000080000000000024400000808210000001200010",
INIT_14 => X"04000100A0000000000028400004000020280000000000012002020204000009",
INIT_15 => X"0001000000000024080000000000010400400004000004000000000000510000",
INIT_16 => X"0108408420430E699AA42A1508104EA08000000810020000000044001AC20500",
INIT_17 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_18 => X"0040100401004010040100401004010040100401004010040100401004010040",
INIT_19 => X"1708000000000000000000010040100401004010040100401004010040100401",
INIT_1A => X"20820820800D41A8283AC618618EF1088160885001234B96061CCDEC4D205061",
INIT_1B => X"0C06030180C06030180C08208208208208208208208208208208208208208208",
INIT_1C => X"F80000B0582C160B0582C160B0582C160B0582C160B0582C160B0582C160B058",
INIT_1D => X"BA5D04020100000000000000000000000000000000000000000000000000401F",
INIT_1E => X"FFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974",
INIT_1F => X"2010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFF",
INIT_20 => X"FFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFF",
INIT_22 => X"AE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFF",
INIT_25 => X"FFFFFFFFFFFFAE974BA5D0402010000000000000000000000000000000000000",
INIT_26 => X"10007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFF",
INIT_27 => X"FFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FF",
INIT_2A => X"FFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_2B => X"0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFF",
INIT_2C => X"00000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D",
INIT_2D => X"007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020100000000000000000000",
INIT_2E => X"FFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_31 => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_32 => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_33 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_34 => X"0000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000007FFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(28),        -- Port A data input
DOA(0)   => data_read_a_hi(28),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(28),        -- Port B data input
DOB(0)   => data_read_b_hi(28),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_29_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"79964E4BA01DACAB9E659792D00AAE160002829C7FDFEFCEE97C2815039D70C3",
INIT_01 => X"50BFF9AB0775343F9AB01DF80D5821FC0FFF3FEFD1AF9FF1207FFBC7B9720586",
INIT_02 => X"0B33180300E700080F6AAA7BFFC007189C7FF2FC003503980A0000001D00DFD8",
INIT_03 => X"0401D940CD0000C8421A2B03210868AC23403E903900010E271006A148A0C000",
INIT_04 => X"49B87A417315D20A313E17F1800000058013DDF8BE21F36E02F0D06E03E8F800",
INIT_05 => X"1F007E33E01A4D9C87525E5101603E6E023D27DA937C03E340EE25CB9B483C12",
INIT_06 => X"85AA06002026872BAE0B1282A005FFF001E1870223FC3BFC98101F109FC6780F",
INIT_07 => X"03BC081023B233E804488527FDC008019968D74982C94110AF204001BC285A82",
INIT_08 => X"001E4191901A101B031F84000000831FA1028575A000110800124600C039C002",
INIT_09 => X"C60888D0782082B50080508FF00048B124D4005C8AFF4158102914800110FFC0",
INIT_0A => X"8AD6ABC02A02A0B0CCB463B4C0748A720B1EA980100BFA02E204D2154D28AA3F",
INIT_0B => X"6A22B126DA40C03531440800C22800B8900042FF0180000ABFEF89250815568A",
INIT_0C => X"803468034680346803468034680353401A340180010A0801422829800A00A001",
INIT_0D => X"87410080C60AB0F42A804628200DBFFF13D05928040329160520528134680346",
INIT_0E => X"2006FFFF8000F8F80281A16A1504302058102C0816244B82A0CA25907D0AA015",
INIT_0F => X"0000080A40000283D80000001402000283D80000001402010901A7D694494192",
INIT_10 => X"0000000034000283D80000001402000283D80000001402002010000A00000000",
INIT_11 => X"000C000000000000081600002080341C00000000000008C00000410085380000",
INIT_12 => X"90981000006809076B2000040400001080581000000000000004810020002010",
INIT_13 => X"0011051620000003410040004080000000040026C00008828B10000001A00210",
INIT_14 => X"04000503A000000000042AC00044000228A8000000000801204212130400000D",
INIT_15 => X"0081000000001064180000000000010C02C000440000240000000000105B0001",
INIT_16 => X"258964C4A44A0C689FF3F9FFEC5D6DBFE0020096528A0B000000CC043EC60780",
INIT_17 => X"5816058160581605816058160581605816058160581605816058160581605816",
INIT_18 => X"8160581605816058160581605816058160581605816058160581605816058160",
INIT_19 => X"03017FFFFFFFFFFFFFFFFE058160581605816058160581605816058160581605",
INIT_1A => X"AEBAEBAEBFFF7FEFCFDF7FFFFFF5DE7CFCB773FFEFBFF3C7E1E779FFEFFF5060",
INIT_1B => X"FEFF7FBFDFEFF7FBFDFEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEEBAEB",
INIT_1C => X"F80000FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFD",
INIT_1D => X"BA5D04020100000000000000000000000000000000000000000000000000401F",
INIT_1E => X"FFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974",
INIT_1F => X"2010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFF",
INIT_20 => X"FFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFF",
INIT_22 => X"AE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFF",
INIT_25 => X"FFFFFFFFFFFFAE974BA5D0402010000000000000000000000000000000000000",
INIT_26 => X"10007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFF",
INIT_27 => X"FFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FF",
INIT_2A => X"FFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_2B => X"0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFF",
INIT_2C => X"00000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D",
INIT_2D => X"007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020100000000000000000000",
INIT_2E => X"FFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_31 => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_32 => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_33 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_34 => X"0000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(29),        -- Port A data input
DOA(0)   => data_read_a_hi(29),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(29),        -- Port B data input
DOB(0)   => data_read_b_hi(29),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_30_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"9E79E79E7BAF7DEBAFAFEFBEFBFFBFFDFFF7FCFF0FBFFDFF7EFDDFFFEFFE8000",
INIT_1B => X"CFE7F3F9FCFE7F3F9FCFE79E79E79E79E79E79E79E79E79E79E79E79E79E79E7",
INIT_1C => X"F800003F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9F",
INIT_1D => X"BA5D04020100000000000000000000000000000000000000000000000000401F",
INIT_1E => X"FFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974",
INIT_1F => X"2010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFF",
INIT_20 => X"FFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFF",
INIT_22 => X"AE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFF",
INIT_25 => X"FFFFFFFFFFFFAE974BA5D0402010000000000000000000000000000000000000",
INIT_26 => X"10007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFF",
INIT_27 => X"FFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FF",
INIT_2A => X"FFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_2B => X"0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFF",
INIT_2C => X"00000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D",
INIT_2D => X"007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020100000000000000000000",
INIT_2E => X"FFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_31 => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_32 => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_33 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_34 => X"0000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(30),        -- Port A data input
DOA(0)   => data_read_a_hi(30),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(30),        -- Port B data input
DOB(0)   => data_read_b_hi(30),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_31_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"129000008004A00804A40000400800020000000C005FEA005800200400050100",
INIT_01 => X"A15FF18019700810180065FFFC0040801E80258CA2951C2200EC0906A0804140",
INIT_02 => X"0000000000000011000550FDFF0FFFFF0007F1FC200000011000000000205FC0",
INIT_03 => X"08425818000000908428C0024210A30004045060302223490002014280410FF8",
INIT_04 => X"DB6A618248140C18E0B016872400000007EBA24058E1ECA8E2D400681FD0E061",
INIT_05 => X"1C0FFC338FF01009048084C400103E28FE3F6FE513703F7000E8E5B4825030F6",
INIT_06 => X"0098000C51000910100006C00426FFC7C202060445F1F2572060FE82671C607E",
INIT_07 => X"40001020400440C41C000617FC0003021259CFDB01BF00020C001FF804000980",
INIT_08 => X"F200020000802000000082044000010022048902000002000000000000000004",
INIT_09 => X"1C002400E3CF3E0B1118C31747F000B33820209206FC9E80000000000220FD1F",
INIT_0A => X"00001A1F00110101092CE7ED81CF0004012290000023E0FC027DF780DF74013F",
INIT_0B => X"044094C1028400548812494C31004124080886FE187FC301B124F20016000000",
INIT_0C => X"0608006080060800608006080060C00304003042023B99862444E60090C41887",
INIT_0D => X"0B400080200481501000884080405FF864008880CC30E8A01C01C00608006080",
INIT_0E => X"2021FFE81FF880EA000400098200C04080204010200810020C18090424040034",
INIT_0F => X"E020000040403C0800002000E800003C0800002000E8000100780C2C30830806",
INIT_10 => X"000EE00000003C0800002000E800003C0800002000E8000017A0040000010003",
INIT_11 => X"040000400003D80000020400DD01000000020003B80000000801AE0200000100",
INIT_12 => X"000000384000006118A080428846A80000000002000780C800180000201017A0",
INIT_13 => X"00E808000001C800001F80020000001F8000000280807404000000E400001D01",
INIT_14 => X"3B810000000003E020000280808AB01000000000F600000003A0200000070800",
INIT_15 => X"000652075000000000080786800010000280808BA0040000000F8800000A0200",
INIT_16 => X"080223010010308025410082404A015F0FFE003182701B420800280C80201A81",
INIT_17 => X"8020080200802008020080200802008020080200802008020080200802008020",
INIT_18 => X"0200802008020080200802008020080200802008020080200802008020080200",
INIT_19 => X"04017FFFFFFFFFFFFFFFFC080200802008020080200802008020080200802008",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000080",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"F800000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"BA5D04020100000000000000000000000000000000000000000000000000401F",
INIT_1E => X"FFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974",
INIT_1F => X"2010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFF",
INIT_20 => X"FFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFF",
INIT_22 => X"AE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFF",
INIT_25 => X"FFFFFFFFFFFFAE974BA5D0402010000000000000000000000000000000000000",
INIT_26 => X"10007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFF",
INIT_27 => X"FFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FF",
INIT_2A => X"FFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_2B => X"0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFF",
INIT_2C => X"00000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D",
INIT_2D => X"007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020100000000000000000000",
INIT_2E => X"FFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_31 => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_32 => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_33 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_34 => X"0000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(31),        -- Port A data input
DOA(0)   => data_read_a_hi(31),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(31),        -- Port B data input
DOB(0)   => data_read_b_hi(31),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_0_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"ED39BA795990D275FB4A6E96ACC4731DEA4598B0AFB54867F6EE4618C3749803",
INIT_01 => X"58A0047D8607944AC7DA180001ECA2544042106208408208C20022E9173734B3",
INIT_02 => X"9F775E7CB273E6CCA7DAAF00001000000478020113C9C38E09FB7CCCDD9F203E",
INIT_03 => X"441406267B4CB04443163C91110C58F24A31000B8028A810A3D0F8B169A01006",
INIT_04 => X"0005802424830120024121209088809DF81454ACA01E03501D0A3B91E00F0A00",
INIT_05 => X"E0F001CC00012034C20B0232838F80D001C0100AEC83C008EF101A034C8CC300",
INIT_06 => X"582541A028D584E40CB0583CCA0100000161F84322000DA8C40F003C80030780",
INIT_07 => X"2BF70E1C3BBBB1138AF7F888025340C0888430047040FEE182CA00044BC5827C",
INIT_08 => X"0CAFC1F1F07F0FE1C94F65B11555EAFFC1C306758B24197ABCDA467F2C9CF9B3",
INIT_09 => X"027BDA3B0000011420A61080800B6E4C464258094101606E5A47A2A2098B0200",
INIT_0A => X"40198000D1281220444210123820B43B40804CE9AFC800017D82082E2081B6C0",
INIT_0B => X"CA2E0B32B01A752B078412A24844B01302A26900C4801854069B0C888890A081",
INIT_0C => X"C0F33C0F73C0F33C0F73C0F33C0E39E0319E0710A9402011C22908B56A21A020",
INIT_0D => X"8429A95E954868AD0E52273F542580000808061C0389161F027039C1F33C0F73",
INIT_0E => X"5C94001120055704FC4A1624485E2489024481224091282C4300942A19439481",
INIT_0F => X"1C55D65C3E3F01F52FFC1E0013C1F801F52FFC1E0013C1F8090423D38A18E3B1",
INIT_10 => X"1C0118796BE001F567FC1E0013C1F801F567FC1E0013C1F9085DFBF7E15C0610",
INIT_11 => X"FBF7E30F00C0270F3751F1FD00FECBF7E25C0700463E17B2C7F811FD7ADECC38",
INIT_12 => X"6474190626D6491063597F9177B956EF378D33E4030061341F077C571F8F885D",
INIT_13 => X"E207F328E3082636B2807FFD80FE00007E03F7207D3E03F9167184131B5C40FE",
INIT_14 => X"047EFA0CAE06101C53E3647D3F144FCDD22B81C0098E57D9081FCE8C8520C4DA",
INIT_15 => X"FF31ADF08DBF81846A540049707E0FE3307D3F141FFB45478040570EED41F4FE",
INIT_16 => X"902C189601208A1502B4AA5584B4068000019A80098120BCA4C617635C938574",
INIT_17 => X"0240902409024090240902409024090240902409024090240902409024090240",
INIT_18 => X"2409024090240902409024090240902409024090240902409024090240902409",
INIT_19 => X"424A800000000000000000902409024090240902409024090240902409024090",
INIT_1A => X"08208208208831042720EE38E38AAF9C4C704DAB63A6D58B3C10BAE8E789AA09",
INIT_1B => X"0F87C3E1F0F87C3E1F0F82082082082082082082082082082082082082082082",
INIT_1C => X"F800003E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F",
INIT_1D => X"55557BD75EF5D00000000000000000000000000000000000000000000018401F",
INIT_1E => X"FEFA28428B455D0017410A28428AAAA2FBD54BAF7FFD55EF007FD75EFFFAE975",
INIT_1F => X"0145F7AEBFFFF08002AA10A2AABFEAAA2FFC0000AA843FE00AAFBE8B45AA803D",
INIT_20 => X"974AA5D7BFFE000804000BAAAAAAAB45557FFFEBAA2D5401450051401555D7FC",
INIT_21 => X"FD7410557FC21555D51574AAA2FFE8B455D7BD755555517FFEFA280021FF082E",
INIT_22 => X"AEBFE00A2803FEBA002A820AA0800174BA5D2EA8B45005168A10AA8028A10087",
INIT_23 => X"7FFE8B45FFFBC00005D003FF45557FC01FFFFAE95410AA80000005D003FEAAFF",
INIT_24 => X"00000000000557DF5500003DFEFFF84175EFA2AEA8A10000417410A2FFE8BEFF",
INIT_25 => X"F0075D75EFEBAE9554540754717F1F8000000000000000000000000000000000",
INIT_26 => X"47E00A2DB45AA8A3AFD7B68E2AB78550E12555F524AFE38B780154BAFFF1D54A",
INIT_27 => X"1D500002A150038038E285D7F78FD7000B6AB50B6AABDE12BEA0AF010B7D1F8F",
INIT_28 => X"D5C7AA854008700249243A412EBFF5542A43FE9257F1E816D557095EAAA2D140",
INIT_29 => X"EDBC0B680900AAF52B474385D75C502D157545A87AAD178A8002D1D21C5E8257",
INIT_2A => X"F6A150012A2F02AFFDF40E85F475451D502D152A82000E3A5D2150AB8F401471",
INIT_2B => X"51EAFEDB52E3F1EFFFF485A2DA3D5D24BD417FD7E9541242FE920AD082E10A28",
INIT_2C => X"00000000000000000000000000005AAF555080550E87B7A405B52AAD152BD001",
INIT_2D => X"FA69574BAF7D5555AF0D79D55FFA2AC97445057F405458500000000000000000",
INIT_2E => X"0FF16565B2FA9075F4F7B3EBDF50FEAEAAB55F7AEAABFF5D2A81151FB8635A02",
INIT_2F => X"4D5D51F5E08A394003A908B8410E707EF34A08D46F6ABE7082AAAAF2FAC77FE0",
INIT_30 => X"FAE8C798A11A0EAEF75F7AA84001A7052C95256803CE3AEB038662E5D8140601",
INIT_31 => X"A05051023F9A9D57B63BFBF906CB45FABC0954AF0151555AF58794040077D774",
INIT_32 => X"FEE5555BE48AB2A2AE0A0F20C43EAC562245B4E1870108B11020AD4AA05542A0",
INIT_33 => X"D407A97F6F35F498B96BEB12DAAB77558ABD5F5F0DA6BC9525688C1A2A0C06E9",
INIT_34 => X"8000000FF8000000FF8000000FF8000000FF8000000FF80F55E25C00A0BA7FBE",
INIT_35 => X"F8000000FF8000000FF8000000FF8000000FF8000000FF8000000FF8000000FF",
INIT_36 => X"000000000000000000000000000000000000000000000000000000000000000F",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000008000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(0),        -- Port A data input
DOA(0)   => data_read_a_lo_256(0),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(0),        -- Port B data input
DOB(0)   => data_read_b_lo_256(0),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_1_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"212C001411984004084D000508C53810A03D1450E839B003342114428A000807",
INIT_01 => X"08000010400A0008010600000084004000400002000000000000000000140000",
INIT_02 => X"484DEBA0111800C004400D000000000028800001CC404E6008B4933336880010",
INIT_03 => X"650C00000848A0423183089008C604224200000100A200002C280810098C0001",
INIT_04 => X"00000004208B00200E010800006667BE7000102C00080000040012010000080C",
INIT_05 => X"0080000000002020600100208D04414000800000000200004800080000800200",
INIT_06 => X"0820196100006044401008100208000008082010000000800488000000020400",
INIT_07 => X"1210C18306788C00894098000011000820001000104050004108000001008250",
INIT_08 => X"00A48903121780004C6000311555521F183060AC564BF818B5EDFDE004460030",
INIT_09 => X"02AD881200100140A0223480000458400000480840002002184581A020000200",
INIT_0A => X"140040001020020410000010082080010400002001041001B102002E20013600",
INIT_0B => X"0895400004201001010884000000901100800800000004140002008280A8A815",
INIT_0C => X"C8D00C8D00C8D40C8D40C8D00C8D20642A06468400000030480808020F08E008",
INIT_0D => X"20BC417C16004C0B83822109040180000801000910000003203220C8C40C8D40",
INIT_0E => X"5C96000000010200200802100022008100408020401020040100142200E0E08A",
INIT_0F => X"0000021E300B000000781E00140018000000781E00140018000002430E30E061",
INIT_10 => X"1C00000024E0000000781E00140018000000781E0014001908400005E11C0610",
INIT_11 => X"0003C30F00C000000155800D00000003E21C0700000000F00118000000468C38",
INIT_12 => X"60640900004A400081401A0000004041218503E4030060000004804318008840",
INIT_13 => X"A0001208C30800025200003D807E000000000725201600090461840001340002",
INIT_14 => X"0000F00C0E06100000012D2005100409520381C00000005920004C0C81200009",
INIT_15 => X"25000120850B8180625400400000010711200510004B41478040000005548016",
INIT_16 => X"10040002002080040000804000A0000000011A000100208C008611430A000040",
INIT_17 => X"0040100401004010040100401004010040100401004010040100401004010040",
INIT_18 => X"0401004010040100401004010040100401004010040100401004010040100401",
INIT_19 => X"5000800000000000000000100401004010040100401004010040100401004010",
INIT_1A => X"8A28A28A2AC8090C69606492492C09945235D5F7E2A5040B80E1C863A2958000",
INIT_1B => X"5BADD6EB75BADD6EB75BAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA28A2",
INIT_1C => X"FC00002E974BA5D2E974BA5D2E974BA5D2E974BA5D2E974BA5D2E974BA5D2E97",
INIT_1D => X"BA55556AAAAAA800000000000000000000000000000000000000000000607FFF",
INIT_1E => X"F45A2FBD75EFA2AE97555F7FBFFF45FFAE80010AAAABFFFFFF803FE10F7D17FE",
INIT_1F => X"8AAAF7FBD54AA002A955555D7FE8ABA082EBFEBAFFD555400557BD54BA5D7FFD",
INIT_20 => X"17555AA8028BEFAAAE97555082A80000AA802ABEFA2D568A005D5157400AA802",
INIT_21 => X"EBDFEF5D7FEAA00AAAABFEAA007BC0145FFFFFDF55AAFBC00105555400105504",
INIT_22 => X"D5575555D7FC2155F7AEA8BEFAAAA954BA557BD7410550428ABA5D5168ABA552",
INIT_23 => X"FD57DF45F7D568ABAF7AABFFFF082ABFFFFFFFFEAB55557FFFEBAAAD568B45A2",
INIT_24 => X"000000000002EBFFEFA280021FF082E974AA5D7BD74000804154BA082ABFF55F",
INIT_25 => X"7F78A3FE28E3D17DEAA485FE8E02B50000000000000000000000000000000000",
INIT_26 => X"6D5D75D54BA5D7BFFF7DA2FFD55EFAAA495545E175EFF57BF8FC2000BEA4BAE9",
INIT_27 => X"A28550E10405F7A4AFE38EAA0924921C2FD55455571E8A2A087BF8EAAEB8E001",
INIT_28 => X"7A28415A001684104155C5B6DF6DBEFBFAA07157428145A00AA8A2FBD7B6DF6A",
INIT_29 => X"AAABF1FFBC7010FF8A38FEF557FEAB78B6AAB8E971471C7010B7D168F47400A0",
INIT_2A => X"495EAAA2D16D1FDBED56A55557A43DE385FD4BFBD7B6A0BF492415FC20105D24",
INIT_2B => X"F5D717FE2AAAA56DEBD17FE3DF7FB7FEBFE38017EBA4A8EB8F6FFD5FE8B7D557",
INIT_2C => X"00000000000000000000000000002A3D5C7AA854008700249243A417FFF41542",
INIT_2D => X"AF2A00010F78028B15F7823FEAAA2D57DFBA007DFCA127B80000000000000000",
INIT_2E => X"A0869AAAB8A7C19C55550E8574BA557BFFFEFAAFBD55FFAA8416545A6FB60F47",
INIT_2F => X"10A2AEBFF55F7BAAA8565DBAC1112FFAC21A022A38C20B2552E975F758516AAA",
INIT_30 => X"01E7AD1FFF5575841DE08007FC2048002895755FFEFBCEE5FBAACB10085EE5DE",
INIT_31 => X"D4000D7FC00FC5D062BBA05ED5034472A02EABEA097BEAAFAF2863FA00DD5742",
INIT_32 => X"62B0A2F7AE8B5D5D51F5E18ABD5EAFFF2AF9554FF57EFBFA18D4FBFFF40FF809",
INIT_33 => X"C95256807DC31AA8114DE55F5BED201FFFED17DFBFF6963FCAAA2283CF140500",
INIT_34 => X"0000000000000000000000000000000000000000000002CB75F7AA84001A7052",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000008000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(1),        -- Port A data input
DOA(0)   => data_read_a_lo_256(1),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(1),        -- Port B data input
DOB(0)   => data_read_b_lo_256(1),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_2_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10E44660018259B2843913100062C98004802322D3E030235201006009B2816",
INIT_01 => X"8005A188084900481C8024A542400340404000720885800802000906E4910204",
INIT_02 => X"5C010802020408040C640850AA055254090541A111240A104A0000000908B510",
INIT_03 => X"0C1101108800004481060A001204102803156020218808002440850008C80550",
INIT_04 => X"8840C08122050400582812C21C0804040968987810688899444090C10A124A69",
INIT_05 => X"4885109105400129210040010340086856B141212252142242A068A080106372",
INIT_06 => X"047450004062400090000202000054C28012204400908281302852A6710AA420",
INIT_07 => X"121810000230089008408402A800011012D41D518044411005000AA8A5004390",
INIT_08 => X"A214110514163218085008010141421F02000124000010880000442080810201",
INIT_09 => X"0A09E89041451581B53A739C42A0C9223000004881708D80100331CA8A848E0A",
INIT_0A => X"1009020A30020008096A06B8C1208A000A9C20004820B0573165541CD5482216",
INIT_0B => X"ACC084404A8000490152D100344001108AA88B1D007291402802B1041632A011",
INIT_0C => X"8696086860869608686086920868004309043414A2191C24485C4D2A9A0DF823",
INIT_0D => X"484000804201C1102080215900038AD030014588D200F0221821808682086820",
INIT_0E => X"00002AA00AA80240A001010026824040C000201030000200C8980080260C201E",
INIT_0F => X"0000000A20001602900020001400002A029000200014000100280E6694490312",
INIT_10 => X"0000000024002A02900020001400001602900020001400002700000800010000",
INIT_11 => X"0008004000000000001500006C00300800020000000000C100014A0081200100",
INIT_12 => X"8088000000480005188000440840081000500002000000000004800010003420",
INIT_13 => X"0070041200000002411280004000000000000026000038020900000001201300",
INIT_14 => X"2A0004030000000000002A00004A100208800000000000012260101100000009",
INIT_15 => X"0084420300001040100000000000010402000049800020000000000000580001",
INIT_16 => X"040111000008001505448340606B21090556002E00000000000080002A040A00",
INIT_17 => X"401004010040300C0300C0300C0100401004010040300C0300C0300C01004010",
INIT_18 => X"0200400004000040000C0200C0200C0200400004000040300C0300C0300C0100",
INIT_19 => X"14A97C0FC0FC1F81F81F800C0200C0200C0200400004000040000C0200C0200C",
INIT_1A => X"0410410411823A4301040B2CB2CBACB002009C6B860185AA1491B0E2863EA015",
INIT_1B => X"8944A25128944A25128941041041041041041041041041041041041041041041",
INIT_1C => X"FC703F25128944A25128944A25128944A25128944A25128944A25128944A2512",
INIT_1D => X"AA0004001550000000000000000000000000000000000000000000000078401F",
INIT_1E => X"5FF5D003FE10F7D17FEBAF7D5420AA0855420AAAA843DFFFAAD1554005D7FD74",
INIT_1F => X"FF45AAFBC20AAF7D1575EF55517DF555D2EBFF45AAAAA8A10A2AE80010A2AA97",
INIT_20 => X"AABEFAAD1575EFAAAE974AA5D51554BA5D7FFFF45A2AA975EFA2FFD7555FFFBF",
INIT_21 => X"5554AA555555555557FE8ABA082EBFFFFAAAE95555552E974105D517DF55AAAA",
INIT_22 => X"D540000AA802AABAF7FFC2010AAAE821EF552E82010F7AABFE10FFD542145FFD",
INIT_23 => X"02E800AA08042AB45007FC00BAFFD168BEFF7FBC0010AA802ABEFAAD540000FF",
INIT_24 => X"000000000002E80010555540010550417555AA8028BEFAAAE821550851420AA0",
INIT_25 => X"7A2DF55400557FD54AA1D04001C5150000000000000000000000000000000000",
INIT_26 => X"D5F7A482000BEAE905C755003FE28E3D17DEAAE95F40002157F470AABE803AE9",
INIT_27 => X"5EFAAA495545E3F5EFF57F7FE80082FFDE105EF55517DFC5552ABDF45B6AEAFF",
INIT_28 => X"24105D5B7FF7DB6AAAABC7BEDB505EFBEA4070BA5FD0154BA5D7BFAF7DA2AE95",
INIT_29 => X"38E00B6DF68FEF4871D24BA495B5556D5571E8AAF082AB8EAAEB8E0016D5D2A9",
INIT_2A => X"E2FBD7B6DF47A00EBDB50000A380AAE28E80495038AAAEAF1D7410E80000FF84",
INIT_2B => X"FBC703AE2DF42AAA002A851C214003FF680071ED1EFEAF1EFFFDEAD1C5010AA8",
INIT_2C => X"00000000000000000000000000002087A28415A001684104155C5B68E2DBEFBF",
INIT_2D => X"51FBD74BAF7802AB05AAFBD5400557BD54AA5500021555100000000000000000",
INIT_2E => X"55D2ABDF55F782BEB47AFAD00010F7AA8215555003FEAAAAD57DEBAA2FDDC010",
INIT_2F => X"BA557BEABEFAAEBD55FFAA1456547A2D360F47AF7FC20B2F7FBC015D58517FF5",
INIT_30 => X"AB4A78016545540400010557BFDFFFF7822A955FFFFC20FFF3AE544108410174",
INIT_31 => X"D545002A800A8FF862BA00F2F9E8F0050D4420BA547FD75FF58516AAAA0828AA",
INIT_32 => X"35B57AB5155400A2AEBFF45FFFB404007FFBD550AAFACAAA122AA8954BAA2AE9",
INIT_33 => X"895755FFAEBCFE57BBA57002DF3C4AAAA002E954505C417FFFF08555555BAAD3",
INIT_34 => X"000000000000000000000000000000000000000000000061DE08007FC2048002",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000010000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(2),        -- Port A data input
DOA(0)   => data_read_a_lo_256(2),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(2),        -- Port B data input
DOB(0)   => data_read_b_lo_256(2),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_3_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"210C44A20020248B08431120001604B8156023104C40771B3430400A02380206",
INIT_01 => X"014C9A4250B0296D3C2422C992100B49404040028804A0080A000416A8D90A0C",
INIT_02 => X"4809A900031800444460589C66E331352180D468B8040E600C0081110B802CD0",
INIT_03 => X"6D0B6110880001D23583480648D60520330066810A80881068A808029CC56330",
INIT_04 => X"48221A066A09D03B348C1C1928DD5A4402A13868070940842640902107002D24",
INIT_05 => X"058318035328202004C1C4E50B44644B30A86D01014A0D224063090082100E34",
INIT_06 => X"08381A010040200AC2190ED2002ACD99881822104C5A40942048288234629414",
INIT_07 => X"0218408142740E2C0948C3066400071913209CC8004640100D003999552083D2",
INIT_08 => X"900409231292A8080C2000110001521F0810A92E7402F08AB0016CA000C60011",
INIT_09 => X"620C889014D30E4A210214D5099058808010605A81A41480102130C020A43A39",
INIT_0A => X"512850E61822020C899046740121820004102000402079CCA037A02C68552A35",
INIT_0B => X"8895000026A00141015290040460C0B4828289AC1011954C0026A20400882914",
INIT_0C => X"80CA080DA080DA080CA080CE080DB0402F040654A2442834C0092E228A0DF2AB",
INIT_0D => X"289080600E04C50206808059000999C98840C508D220108200202080DA080CA0",
INIT_0E => X"300E6660599802602209021204A050E1C850C428521C208480821D842085A03E",
INIT_0F => X"0000010000003202900000010000000A02900000010000008038666920920A24",
INIT_10 => X"0000008000002202900000010000001E02900000010000002380000800000000",
INIT_11 => X"0008000000000000008000002D00300800000000000020010001620081200000",
INIT_12 => X"8088000008001021C88000048800281000500000000000004000000000003600",
INIT_13 => X"00B8041200000040011980004000000000000803000068020900000020001B00",
INIT_14 => X"29800403000000000008030000C83002088000000000002002E0101100000100",
INIT_15 => X"00841003100010401000000000002000030000C38000200000000000020C0001",
INIT_16 => X"108722420420A0100006D34A404800185CCE0128410820000008008021C40A00",
INIT_17 => X"0872108721085218852188521885218852188521887210872108721087210872",
INIT_18 => X"8721086214872108621C852188421C852188421C852188721087210872108721",
INIT_19 => X"54A2EAA555AAB554AAB5561C852188421C852188421C85218842148721086214",
INIT_1A => X"0410410412881D0B0000092492480A981E063C638321450A08899A62C314A014",
INIT_1B => X"9D4EA753A9D4EA753A9D49249249249249249249249249249249249249241041",
INIT_1C => X"FAABC4351A8D46A351A8D46A351A8D46A351A8D46A351A8D46A351A8D46A351A",
INIT_1D => X"5500002AA100000000000000000000000000000000000000000000000000401F",
INIT_1E => X"FFFAAD1554005D7FD74AAA284001550055421EFAAFFD54AAF7D168B45AAAABDF",
INIT_1F => X"20AA080400155AAD5554AAF7802AB4500043DF45FFD168AAA0855420AAAA843D",
INIT_20 => X"021550855555FFAA84001FFAAAE80010A2AA955FF5D003FE10F7803FEBAFFD54",
INIT_21 => X"BC20AAA284175EF55517DF555D2EBFE00AA8028B45A2AE82155A2FBFFEBA0800",
INIT_22 => X"7BD7555FFFBFDF55AAFBD55EF5D2EBFE10085168ABAFFFBD54BAAAAE97400A2F",
INIT_23 => X"D0015410F7AAAAAAA55043DE00FFFFD5555AAAA954AA5D7FFFF45AAAA975EF00",
INIT_24 => X"0000000000004174105D517DF55AAAAAABEFAAD1575EFAAAE974AA5D00175555",
INIT_25 => X"2EBD56DB7DBEAEBFF551C042AA101D0000000000000000000000000000000000",
INIT_26 => X"D75D5B470AABE8A3AFD7A2DF55400557FD54AABC04001C51551471D7AAF1D05D",
INIT_27 => X"E28E3D17DEAAEBDF40002550F47155AADB50492EB842FB5508043FF55EBD56AB",
INIT_28 => X"017DAAFFFAE821C0A0717D1C5B575FFB68E82557FD2082000BEAE905C755003F",
INIT_29 => X"D74BAE3AE85480FFFFC00AABE8E105C755517DF40552ABDF45B6AEAFFD5F7A48",
INIT_2A => X"FFAF7DA2AE905EF0075D5545E3F5EFF57F7D5C55D7492E90E3808756DA92EBFF",
INIT_2B => X"F5C7092FF801756D490A10438EBA4B8E9241043AE10EAF5C5547FF80954AA5D7",
INIT_2C => X"00000000000000000000000000000E124105D5B7FF7DB6AAAABC7BEDB505EFBE",
INIT_2D => X"515157555AAD142040A2D57FFFFFFAEBFF555D0028A005100000000000000000",
INIT_2E => X"500003FF55AAFD6AB455157D74BAF7AAA8B45AAFBD54005D7BD54AAF78002155",
INIT_2F => X"10F7AA8215555003FEAAAAC53DEB8A2FDDC01051AE955F7AAFBC0000AF843FF5",
INIT_30 => X"F51F782BCB47ABAE801FFAAFBEAA105D2E955FF557BD74EFFBACD41577B84000",
INIT_31 => X"0AAA00557FEA8A2FDD64BAAF8282012AFFEC20BAF7AA8015558517FF555D2ABD",
INIT_32 => X"48547AE04174BA557BEABEFA2AA951FF88554214FA2D3EAF57AFFDD7555082AA",
INIT_33 => X"22A955FFFFC21FFF3BE40412DE02955FF082A820AAAB842AA00000028AB0AAFF",
INIT_34 => X"0000000000000000000000000000000000000000000002A80010557BFDFFFF78",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000008000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(3),        -- Port A data input
DOA(0)   => data_read_a_lo_256(3),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(3),        -- Port B data input
DOB(0)   => data_read_b_lo_256(3),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_4_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10804002061080A284201081034809800A00230340007833522C82D04A16006",
INIT_01 => X"804399801838084C0420450E1E104348403008418984014902030006A0910204",
INIT_02 => X"480108A200000000446418E01E80F00A4104311868240200080000000988A390",
INIT_03 => X"065140108800004080064A0002001128270072E03000000030808D00888100F0",
INIT_04 => X"9100EB836A155C1AF0B81CD60433B944022AB8385AC0D4B8E02010E81C32E821",
INIT_05 => X"5C0F20B36F08000024C084C501441C4CF01C489533483C8042EAC190001074C4",
INIT_06 => X"0034420151620118120106902406C3C7800201448DD9D2871020F2AA375A6071",
INIT_07 => X"12181000023480040840C001E080030032009700024641000C00187A442007C2",
INIT_08 => X"8084830110160218004000001101121F220000260000108AA000440880000000",
INIT_09 => X"5A8C881063DF3E839008F29F407448F200B020DA841CA2001001008882046647",
INIT_0A => X"C61504C1380101801900439001FD8804041400001002003C230B6715A4786E0F",
INIT_0B => X"ACD1240522E000098100D104B26041348A088078116C105DA006D10416BE3002",
INIT_0C => X"8608086180860808608086180860A0434C0430D4A25F3182CC4D5D221A09E821",
INIT_0D => X"0BC28081080549504400A8080009B878184044881222D1821821A08628086180",
INIT_0E => X"20481E0E18790012820001100200D02048300418022C1282809A09040415002A",
INIT_0F => X"0000010020005E0090000001000000C6009000000100000000380E6C30830806",
INIT_10 => X"000000800000D20090000001000000EE0090000001000000A6A2000000000000",
INIT_11 => X"0000000000000000008100003B00200800000000000020010002EA0080200000",
INIT_12 => X"80800000080000211D80000C0044281000400000000000004000000010003282",
INIT_13 => X"03B00410000000400121800000000000000008020000B8020800000020006F00",
INIT_14 => X"59000402000000000008020000C9000200800000000000200FC0101000000100",
INIT_15 => X"008A500100001040000000000000200002000042E00000000000000002080001",
INIT_16 => X"08820440040802500104C34820E3031B63C20530C01800410009009821040A00",
INIT_17 => X"C832008020C812008220C81200802048320880204832008020C8320082204812",
INIT_18 => X"8120481208822008020C812048320880208802048320C8120882204812088020",
INIT_19 => X"10A3A5930C9A6CB261934E048320C81200822008220C81204832008020882204",
INIT_1A => X"8A28A28A2BD30264686668A28A2605145031C03F028000A1C2ED7831A2822250",
INIT_1B => X"51A8D46A351A8D46A351AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA28A2",
INIT_1C => X"F94304068341A0D068341A0D068341A0D068341A0D068341A0D068341A0D0683",
INIT_1D => X"BAAA84154005500000000000000000000000000000000000000000000000401F",
INIT_1E => X"4AAF7D168B45AAAABDF55A2802AA1000002ABFF087FFDF5508003FEBA087FD54",
INIT_1F => X"015500002AABA082E954005500021FF5D2EBFF5500003DF455555421EFAAFFD5",
INIT_20 => X"174BAA2AABDE0055517FF555555420AAAA843DFFFAAD1554005D7FD74AAAA840",
INIT_21 => X"400155AAD1554AAF7802AB4500043DF45FFD168BEF080028BFF0855555455500",
INIT_22 => X"803FEBAFFD5420BA085168A00007BFDE10085168ABA0055574BA5555554BA5D0",
INIT_23 => X"02A97545F7D1555EF55043DF5555517DEAA5D0400010A2AA955FF55003FE10F7",
INIT_24 => X"000000000002A82155A2FBFFEBA0800021550855555FFAA84001FFAAFBEAB450",
INIT_25 => X"5080A3AEAA007BD2482BE84124285C0000000000000000000000000000000000",
INIT_26 => X"381451471D7AAFBD0492EBD56DB7DBEAEBFF55BC042AA101D0A28BC7007FFDF4",
INIT_27 => X"400557FD54AABE84001C5550A28ABA1424974004100021FF492AB8F7D1C0438E",
INIT_28 => X"8BEF005557545490012482B6A0BAE2849557AFED1C5F470AABE8A3AFD7A2DF55",
INIT_29 => X"504924955524AA140E0717DAADB50492EB842FB5508043FF55EBD56ABD75D042",
INIT_2A => X"A905C755003FE28E3803DEAAEBDF40002557F6DA101475FDE10145F68A921C55",
INIT_2B => X"DF425575D7BEFB55002097555FFD5401EF5D043AF6D405F78E3A1C2002000BEA",
INIT_2C => X"0000000000000000000000000000208017DAAFFFAE821C0A0717D1C5B575FFB6",
INIT_2D => X"512EAAB45007FFFF55082EA8AAA087FC2010F784000AA5900000000000000000",
INIT_2E => X"F002EA8BEF5D0428ABA595557555AAFBC2000A2D57FFFFF7AEBFF55FF8028A00",
INIT_2F => X"BAF7AAA8B45AAFBD54005D7BD54AAF78002155512AAAA085D04174100800021F",
INIT_30 => X"F55AAFD6AB4551002ABEF005555555000402000FF802ABAA04552ABFF597FD74",
INIT_31 => X"DE005D7BE8AA85555400100879560AA592F955FFAAFBC0000AF843FF5500003F",
INIT_32 => X"FCABA598400010F7AA8215555003FEAAAA843DEB0A2FD5600051537DE005D557",
INIT_33 => X"E955FF557BD75EFFBBCD415521FBFDF45000417545FFD5421FF5D0428BEF0079",
INIT_34 => X"00000000000000000000000000000000000000000000004001FFAAFBEAA105D2",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000010000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(4),        -- Port A data input
DOA(0)   => data_read_a_lo_256(4),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(4),        -- Port B data input
DOB(0)   => data_read_b_lo_256(4),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_5_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50DB4A0791B1B4B694369283C81F9996A091832112004AB37B20E07C0C1E006",
INIT_01 => X"085FBC448000804C446A00000034826841280A00084000C8C212802EE2953235",
INIT_02 => X"C809AD5CB118E640A4D018FC011FF0002080000082C8C66609DB7DDDCB1F2036",
INIT_03 => X"250907263E4C90D210835C82484205720B20640A88800000B8E0F810A8C4500E",
INIT_04 => X"4005102126898100064D20001044429C7824382C0416C087198AB916E0551A24",
INIT_05 => X"A370C14CA0E101094008002389CFE2F20D7D7A114CB5C20AE514178054948912",
INIT_06 => X"547319A1499121D4C0A046FC4E06C030581859058C2404844437118630839B88",
INIT_07 => X"2A53468D1A758C038AFFEA9FE39348C9204C389672407EF120EA5806E6C543AC",
INIT_08 => X"8C05896372728FE0C420619000003AFF48D1222E5D26F06ABCC96CD72C463990",
INIT_09 => X"82DE9AB9182080C801041080300F6F0E42821809C2FEA0B65A212282002B029F",
INIT_0A => X"1688E480D10A90049026145B3830B64944904569E7E00A002C836D35B68D26C0",
INIT_0B => X"88990E14269AB54B078092E6BD4431138A00AEFDD567DA480816848C94180846",
INIT_0C => X"C0591C0791C0491C0791C0591C06A8E0248E03D68860A0106119883D6AE1A0A4",
INIT_0D => X"23D829FA654184533252095E542387F81008071C1BAAD68B027029C0491C0691",
INIT_0E => X"0CA7FE0227FC25847C4395166C5844480204011210A11028C380802A24C89494",
INIT_0F => X"1C55D65E3E3C017C37FC3E0017C1F8017C37FC3E0017C1F90005024108308061",
INIT_10 => X"1C0118796FE0017CA7FC3E0017C1F8017CA7FC3E0017C1F9100DFFF5E15D0610",
INIT_11 => X"FFF3E34F00C0270F3755F1F8007FCBEBE25E0700463E17F2C7E014FF7AE6CD38",
INIT_12 => X"64E4090626DE40100459759173BBD6EF37C523E6030061341F07FC571F8F800D",
INIT_13 => X"E0A6FE28C3082636F201BFFF807E00007E03F7243D38337D1C6184131B7C1DEF",
INIT_14 => X"397FFA0E0E06101C53E36C3D3E884FDDD28381C0098E57D923BDFC8C8120C4DB",
INIT_15 => X"FA36FDF58DBF81C062540049707E0FE7303D3E03BFFF41478040570EED50F4F8",
INIT_16 => X"88212B100901A2349004C26A624A21040FC190050A2110B8ACC40B204A119074",
INIT_17 => X"C20080230802108C2008C22080210882108C220842208821088210842208C200",
INIT_18 => X"20084220842208C2008823080230802108823084220842008821080230842008",
INIT_19 => X"54C1892596D34924B2DA6884220842008C20084220802108821080230802308C",
INIT_1A => X"BEFBEFBEFB7F7FE7EFEEE79E79EFAF2DDA73FBDCEDBFF9D3F0FDE0DB6DBF6218",
INIT_1B => X"DEEF77BBDDEEF77BBDDEEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEF",
INIT_1C => X"FAF3167BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBD",
INIT_1D => X"BA5D2ABFFEFFF80000000000000000000000000000000000000000000000401F",
INIT_1E => X"F5508003FEBA087FD54BA0804154005555574AAA2802AA10FFFFFDE0008556AA",
INIT_1F => X"AA1000003FEBA00002AABA5D2EBFEBAAAD16AABAF7AAA8BFFAA802ABFF087FFD",
INIT_20 => X"E8B45FF80001555D2E955FFFFD5421EFAAFFD54AAF7D168B45AAAABDF55AA802",
INIT_21 => X"02AABA082E954005500021FF5D2EBFF5500003DE005555575EFA2D142145A2FF",
INIT_22 => X"7FD74AAAA840014500517FFEF007BEABFF5D7FC00BA5D5568AAAF7AAAAAAAAA8",
INIT_23 => X"2FBEAA105D2E97410FFD16AAAA5D2ABDEBAFFD5420AAAA843DFFFAAD1554005D",
INIT_24 => X"000000000000028BFF0855555455500174BAA2AABDE0055517FF555504154BAA",
INIT_25 => X"0FFFFFFE38085F6FA92552AB8FEFF78000000000000000000000000000000000",
INIT_26 => X"C7B68A28BC70075FDF45080A3AEAA007BD24821E84124285C51574BAB68A2DA0",
INIT_27 => X"B7DBEAEBFF55BE842AA105D0A38EBA1C0428A925D2AB8EBABEDB6AA92F7AAA8B",
INIT_28 => X"75EFA2DB45145B6F5EFB6DF78E05145552A925FFFFD1471D7AAFBD0492EBD56D",
INIT_29 => X"68AAAF7AAAAA82BE8A28A921424974004100021FF492AB8F7D1C0438E38145B5",
INIT_2A => X"A3AFD7A2DF55400557FD54AABE84001C555517DFC70875EABC7557FC20AA415F",
INIT_2B => X"043AFED1C0E10492B6FFEFA105D2A95410FFDB6FABA542ABAE2AF7DF470AABE8",
INIT_2C => X"00000000000000000000000000000428BEF005557545490012482B6A0BAE2849",
INIT_2D => X"5955554BAFFAEBDE10F7FBFDEBA007BFDE005D2AAABEFFB80000000000000000",
INIT_2E => X"AF7FBE8A00FFAEAAB45F3AAAAB4500557FF55082EA8AAA087FC20105504000AA",
INIT_2F => X"55AAFBC2000A2D57FFFFF7AEBFF55FF8028A00512AA8AAA5D0028A005D2AA8AB",
INIT_30 => X"BEF5D0428ABA597FD55FFA2FFD5555FFD57FFEFFFAA97545552A821EFFBD5575",
INIT_31 => X"8B55557FC0012087FEAABAF7AAAAA10F3AAAAA005D04174100800021FF002EA8",
INIT_32 => X"A8ABAFBFFD74BAF7AAA8B45AAFBD54005D7BD54AAF7800015551517DF4500516",
INIT_33 => X"402000FF802AAAA04452ABFF592E80010FFFFFFE005D2A95410F7FFFFEBA5D2E",
INIT_34 => X"000000000000000000000000000000000000000000000002ABEF005555555000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000060000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(5),        -- Port A data input
DOA(0)   => data_read_a_lo_256(5),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(5),        -- Port B data input
DOB(0)   => data_read_b_lo_256(5),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_6_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10804B0061A010A2840012C030028180004003220200403302301C0381A0086",
INIT_01 => X"A70041CA3839684D18A160000C52424841000000090800090210080008110204",
INIT_02 => X"080108200C1000004465480400C0080100000000010432400800800009882050",
INIT_03 => X"040001008C2340D0842208624210802182800584488000103080014E08C10000",
INIT_04 => X"00101611A029B08410044800000000040088122A44281C040400900500001800",
INIT_05 => X"02800000400C820934E4A0002900404402820024000A00824004283011200A00",
INIT_06 => X"2632000004084804134DA7C011A83FC012122100C80812D00308010000829400",
INIT_07 => X"02181020423088002940C2401D0480112000100004404014602447F805326393",
INIT_08 => X"7004812130160008304000000000021F020408244000108A0000440003040000",
INIT_09 => X"020C889010104088A000348037F05840303902E814000010341108802020FF40",
INIT_0A => X"86C8B5DF1C83C9C8900000100220C244840021100017E2FD200000A40001223F",
INIT_0B => X"88D1804122A088018152D144317205502A880C00107FD75DE922005026A62A15",
INIT_0C => X"B6284B6284B6184B6184B6384B62825B0425B0568075A0826849C8229AC5F8AE",
INIT_0D => X"03C440C054048850A300A8480009A0020865A588DA20F1A2D92D82B6084B6084",
INIT_0E => X"031001E0800122100321C89214A01A742D3A168D1B4686D100234B442428C034",
INIT_0F => X"000008AB80030202800000001402068202800000001402067400026000000000",
INIT_10 => X"00000000341E8202100000001402068202100000001402062840000800000000",
INIT_11 => X"0008000000000000083C00052000300000000000000008CD0018400081000000",
INIT_12 => X"800800000069A48584000A0400000010001000000000000000048128C0002840",
INIT_13 => X"1A480012000000034C1E000040000000000400FE000644020100000001A34000",
INIT_14 => X"02800401000000000004BA000112B0020800000000000807E80000110000000D",
INIT_15 => X"0500020250001000100000000000010CCE000198000020000000000010F80006",
INIT_16 => X"62D18468CE8402440404D24A3081B020603E0A20640C8400010298432A002A00",
INIT_17 => X"ED3B4ED0B42D1B4ED3B42D0B42D1B4ED2B42D0B46D3B4ED2B42D1B46D3B4AD2B",
INIT_18 => X"D0B46D3B4AD0B46D1B4AD3B4ED0B42D1B4ED2B4ED1B42D0B4AD3B4ED0B42D0B4",
INIT_19 => X"002331C618E38E38C31C7346D3B4AD2B46D1B42D2B4ED2B42D1B46D2B4AD1B42",
INIT_1A => X"8E38E38E39DB3B676F66EFBEFBEFAFBC5E73FC7F87A7D4ABFE7CFAFBE7BF8040",
INIT_1B => X"CFE7F3F9FCFE7F3F9FCFE38E38E38E38E38E38E38E38E38E38E38E38E38E38E3",
INIT_1C => X"FF75A43F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9F",
INIT_1D => X"BA5D7BEAAAAFF80000000000000000000000000000000000000000000060401F",
INIT_1E => X"A10FFFFFDE0008556AABA5D2ABFFEFFF843DFEFA2FBD54BA5555554BAAAFBC20",
INIT_1F => X"5400550428AAAAA84021FF007BD54BAAAD17DEBA0855421455555574AAA2802A",
INIT_20 => X"17400AAFBE8ABAF7FFD54AAAA802ABFF087FFDF5508003FEBA087FD54BA00041",
INIT_21 => X"03FEBA00002AABA5D2EBFEBAAAD16AABAF7AAA8BFFAAD1554BA002A95555A284",
INIT_22 => X"AABDF55AA802AA100000001EF087FEAA00FFFBD5545080417555A2D17FE10000",
INIT_23 => X"2803DFEF0855401FF082EA8B555D7FC21FFFFD5421EFAAFFD54AAF7D168B45AA",
INIT_24 => X"0000000000055575EFA2D142145A2FFE8B45FF80001555D2E955FFFF843DEAAA",
INIT_25 => X"A415B52492B6F5C20825D7FE8A92FF8000000000000000000000000000000000",
INIT_26 => X"555551574BAB68A2DA00FFFFFFE38085F6FA92552AB8FEFF78E3DFFFAAFFD04A",
INIT_27 => X"EAA007BD24821C04124281C0E2DA82BE8E001EF147BD2482BED57AE921451421",
INIT_28 => X"24AA14209557DA28E15400BEF1EFA92FFFFD24BAB68A28BC70075FDF45080A3A",
INIT_29 => X"17545B6D178E281C0A38EBA1C0428A925D2AB8EBABEDB6AA92F7AAA8BC7B6D55",
INIT_2A => X"BD0492EBD56DB7DBEAEBFF55BE842AA105D0E071FF0071EDA38F7F1D55550004",
INIT_2B => X"2A925FFFF8E3DE82BE8E38FFF0851401C70824A8B555C7FC2147F7D1471D7AAF",
INIT_2C => X"00000000000000000000000000005B575EFA2DB45145B6F5EFB6DF78E0514555",
INIT_2D => X"FBAABDFEFAAFBC00BA007BC0000FFD542000557FE8A00F380000000000000000",
INIT_2E => X"0F7D168A105D55421455155554BAFFAEBDE10F7FBFDEBA007BFDE005D2AAABEF",
INIT_2F => X"4500557FF55082EA8AAA087FC20105504000AA592ABFE00F7AA821FF557FC001",
INIT_30 => X"A00FFAEAAB45F3D5400BA5504155EFAAAE95410F7D57DE00FFFBC00AAFBAAAAB",
INIT_31 => X"FEAAF7D157545080417545F7D56AAAA592AA8AAA5D0028A005D2AA8ABAF7FBE8",
INIT_32 => X"C2145F3D557555AAFBC2000A2D57FFFFF7AEBFF55FF8028A00512E975FF08557",
INIT_33 => X"57FFEFFFAA97545552A821EFFBAABDE00F7AAAABEF005542155000028B555D7F",
INIT_34 => X"0000000000000000000000000000000000000000000007FD55FFA2FFD5555FFD",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000048000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(6),        -- Port A data input
DOA(0)   => data_read_a_lo_256(6),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(6),        -- Port B data input
DOB(0)   => data_read_b_lo_256(6),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_7_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10840B0048225802842102C02450418800002300500030B313300C418992002",
INIT_01 => X"A34009C23838684D1C20E0000E11426840000000080000080200090000510200",
INIT_02 => X"4801082048100000446558040080000041000000000622400800000009000010",
INIT_03 => X"040001818CA144D0842248424210812102000400088000003080014688800000",
INIT_04 => X"000010002041800000048000000000040088322944200C850001940400301800",
INIT_05 => X"0200000040004100280040204104004402000025000800065004203030320800",
INIT_06 => X"0430060044084804900806D1112A002012120004440812D40120008200829001",
INIT_07 => X"02181020423408002940C24001A4A010200018920646C10C7035000244004380",
INIT_08 => X"008481213016020C204000000000121F020408264000100AA000440012040000",
INIT_09 => X"820C899410000000A100348020005902B1A0048825008091350100CAA0200280",
INIT_0A => X"50140A0010058188100004590331C9C4A400231200340C012100002400012200",
INIT_0B => X"1811C44D22A1884141600411800008104080890023000009A926801050001C00",
INIT_0C => X"9002C9002C9022C9022C9022C903064809648080204020004009080A0A00E088",
INIT_0D => X"0880144434A0010012280008031980036000014A0046206241A4069002C9002C",
INIT_0E => X"0216000200010000000081102080400040002000002010000004008080048A00",
INIT_0F => X"038A2881210382000000001E003E0582000000001E003E042283424000000000",
INIT_10 => X"60700706901982000000001E003E0582000000001E003E046840000000009864",
INIT_11 => X"00000000330C00F0C8210807200000000000581C01C1C809201C400000000001",
INIT_12 => X"0000C2419121028C00020A2400000000000080082C180603A0E003A090406840",
INIT_13 => X"14E8000004321189085F8000000061E001FC00C00207740000021908C4829D00",
INIT_14 => X"BB800000009864038C14800201BAB000000026130071A80613A0000018483224",
INIT_15 => X"0546520350000600812058100F81C018880201BBA0000008239020F110800806",
INIT_16 => X"24003300080022140444D268624B210040004A08000000044222900320C84008",
INIT_17 => X"4010040100402000000000000003004010040100000000000000100401004010",
INIT_18 => X"0000C01004010000000001004010040000000004010040300400000000000200",
INIT_19 => X"54A2C208200010410400000800000000040100C01000000000100C0100400000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000002A10",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FAF8800000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"55002E820AAAA80000000000000000000000000000000000000000000000401F",
INIT_1E => X"4BA5555554BAAAFBC20BA5D7BEAAAAFFFBC00AAF7D5575455D557DFEF002AAAB",
INIT_1F => X"FFEFFFAAAAAAAF7D57FFEFF7D555555A2AEAAB55007FD74AAAA843DFEFA2FBD5",
INIT_20 => X"FDF550000175555504175450055574AAA2802AA10FFFFFDE0008556AABA5D2AB",
INIT_21 => X"428AAAAA84021FF007BD54BAAAD17DEBA085542145552ABDFEFFFAA801EFFFFB",
INIT_22 => X"7FD54BA000415400557BD74BAFFD140000082A975EF00003DF55555168A00000",
INIT_23 => X"5557FEAAA2843FF55A2AEA8B55AAAABDEAAFF802ABFF087FFDF5508003FEBA08",
INIT_24 => X"0000000000051554BA002A95555A28417400AAFBE8ABAF7FFD54AAAAAEA8ABA5",
INIT_25 => X"5415178FD7082EAAB550820870BAAA8000000000000000000000000000000000",
INIT_26 => X"82AA8E3DFFFAAFFD04AA415B52492B6F5C20825D7FE8A92FFFFC70BAE3D15555",
INIT_27 => X"E38085F6FA92552AB8FEFF7A0ADABAEBD578FFFEBD55557DBEA4AFB550871D74",
INIT_28 => X"DFD7FFA4801D7F7F5FDF55000E17545410E175550051574BAB68A2DA00FFFFFF",
INIT_29 => X"3AF55415F6DA38080E2DA82BE8E001EF147BD2482BED57AE921451421555524B",
INIT_2A => X"5FDF45080A3AEAA007BD24821C04124281C7BD2482E3D1450381C20905EF0800",
INIT_2B => X"FFD24BAB6A4A8A82495F78E92AA843DF45BEAAAFB55ABA0BDE02EB8A28BC7007",
INIT_2C => X"000000000000000000000000000055524AA14209557DA28E15400BEF1EFA92FF",
INIT_2D => X"F3FFD54BAAAD15754508556AB45002AA8B450800174BAA680000000000000000",
INIT_2E => X"FF7803DF45085557410AEAABDFEFAAFBC00BA007BC0000FFD542000557FE8A00",
INIT_2F => X"BAFFAEBDE10F7FBFDEBA007BFDE005D2AAABEFFB803DEAAAAD56ABEFAAD5575E",
INIT_30 => X"A105D554214551003FF45FF8400145FFD57FF55082E97555002E955550C55554",
INIT_31 => X"54AA5500021EF000028B55087BFDEBA042ABFE00F7AA821FF557FC0010F7D168",
INIT_32 => X"3FE10AEAAAAB4500557FF55082EA8AAA087FC20105504000AA597FC2010A2D15",
INIT_33 => X"E95410F7D57DE00FFFBC00AAFB8028A00007FE8A00A2803FF45F7AABDF55AA84",
INIT_34 => X"00000000000000000000000000000000000000000000055400BA5504155EFAAA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000007FFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(7),        -- Port A data input
DOA(0)   => data_read_a_lo_256(7),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(7),        -- Port B data input
DOB(0)   => data_read_b_lo_256(7),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_8_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00000648E2840112C00000418000002700500030B3132000400812082",
INIT_01 => X"A14008420008204D042100000212026840000000180800080200090048510204",
INIT_02 => X"080108000090000004655C040080000051000000000402400800000009000010",
INIT_03 => X"00000100803008D0842240024210810002800584488000103080894288800000",
INIT_04 => X"00009610A028B084000440C0040000040088323244280C950400808500321800",
INIT_05 => X"42800080400C8A09306420202804400402800035200A00020204283001114A00",
INIT_06 => X"2230400041404B141345A7C20426FFC01292214444081254002801A200821400",
INIT_07 => X"021810204214080069408200008C1010200018920E06C0000020DFFA453223D3",
INIT_08 => X"0084010110120008024000000000021F02040826400000008000440000240000",
INIT_09 => X"828D8880100040898128768820045142B0B902E815008080A0B13848A2200280",
INIT_0A => X"9148A4801C81C9C8100004590711800414002004402008013000403084090200",
INIT_0B => X"BC95C44522A002410040940084720450220089000100104DE924800030821452",
INIT_0C => X"0000400004000040000400004000220010200114AA4020004009092A0009E0A8",
INIT_0D => X"0BC4028430108150900408590109A00209642500120230200100220020400004",
INIT_0E => X"0010000600002210A320C89000005A142D0A16850B6294D10023420124240114",
INIT_0F => X"00000800008100020003C1FE00020080020003C1FE0002004401426008208041",
INIT_10 => X"E3F00000100080020003C1FE00020080020003C1FE000200080000081EA2F9EC",
INIT_11 => X"00081CB0FF3C000008000201000010001DA1F8FC0000080110080000010132C7",
INIT_12 => X"0B0BE6C00020040580040200000001004832CC19FCF81E000000010000200800",
INIT_13 => X"020000C31CF60001008000007F01FFE00004000200420000618E7B0000804000",
INIT_14 => X"000000F151F9EC0000040200401000200D547E3F00000800080001617AD80004",
INIT_15 => X"0100000822406E1B95A3F83000000008020040100000BAB87FB0000010080102",
INIT_16 => X"66D1A368C68D26000544D26A504AB12040022220640484000110184300002A02",
INIT_17 => X"6D1B46D1B46D1B46D1B46D1B46D0B42D0B42D0B42D0B42D0B42D1B46D1B46D1B",
INIT_18 => X"D1B42D0B42D0B42D0B42D1B46D1B46D1B46D1B42D0B42D0B42D0B42D0B42D0B4",
INIT_19 => X"442200000000000000000346D1B46D1B42D0B42D0B42D0B42D1B46D1B46D1B46",
INIT_1A => X"9E79E79E7B7F11E66C6FAD96D96520145052A1F5E2BD085122ED48F3AEB20840",
INIT_1B => X"C3E1F0F87C3E1F0F87C3E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7",
INIT_1C => X"FA2A6D4F87D3E1F4F87D3E1F4F87D3E1F4F87D3E1F4F87D3E1F4F87D3E1F4F87",
INIT_1D => X"FFFF84000AAFF80000000000000000000000000000000000000000000000401F",
INIT_1E => X"5455D557DFEF002AAAB55002E820AAAA840000000043DF55087BC01EF007FD75",
INIT_1F => X"AAAAFFAA95545552ABFE00087BC00AA082EBFE10A28028AAAAAFBC00AAF7D557",
INIT_20 => X"E8BFFA2FBFFFFFAAD5400AAFF843DFEFA2FBD54BA5555554BAAAFBC20BA5D7BE",
INIT_21 => X"AAAAAAF7D57FFEFF7D555555A2AEAAB55007FD74AAAAD57FF45002A975FF007B",
INIT_22 => X"556AABA5D2ABFFEFFFAA82000555555545AAFBE8A00082A97410F7D5555EFAAA",
INIT_23 => X"87BC2010AAD54014500516ABFFA2AABDF450055574AAA2802AA10FFFFFDE0008",
INIT_24 => X"000000000002ABDFEFFFAA801EFFFFBFDF550000175555504175450000155450",
INIT_25 => X"50075C71FF087BD75D7FF84050BAEB8000000000000000000000000000000000",
INIT_26 => X"BABEFFC70BAE3D155555415178FD7082EAAB550820870BAAA8407000140038F4",
INIT_27 => X"492B6F5C20825D7FE8A92FFA497545552AB8E10007FC50BA002ABFE00AA8A2AA",
INIT_28 => X"DF451C24955EF0875EFBD7B6F1FFFC7BEDB45082EB8E3DFFFAAFFD04AA415B52",
INIT_29 => X"92410EBD5505EFB6A0ADABAEBD578FFFEBD55557DBEA4AFB550871D7482AAD17",
INIT_2A => X"A2DA00FFFFFFE38085F6FA92552AB8FEFF7AA87000415B5057DAAFBE8A100820",
INIT_2B => X"0E17555000E17545007BC0000BED14217D005B6ABC7B6AABFFED0051574BAB68",
INIT_2C => X"000000000000000000000000000024BDFD7FFA4801D7F7F5FDF55000E1754541",
INIT_2D => X"A684174105D042AB550055555FF007BD7555F784174AAA280000000000000000",
INIT_2E => X"A082EBDE10AAAEA8ABAF7FFD54BAAAD15754508556AB45002AA8B450800174BA",
INIT_2F => X"EFAAFBC00BA007BC0000FFD542000557FE8A00F384175555D2EA8A00087BD74B",
INIT_30 => X"F45085557410AED17FF455D04155FF00557DF55FFD57DF55FFFBD5400A2AABDF",
INIT_31 => X"21EFA2FFEAA00000002010A2D5421FFFF803DEAAAAD56ABEFAAD5575EFF7803D",
INIT_32 => X"BDFEF0855554BAFFAEBDE10F7FBFDEBA007BFDE005D2AAABEFFBAE97410087BC",
INIT_33 => X"57FF55082E97555002E955550C2E95555087BC0010FFD1401EF087FE8B55FFAE",
INIT_34 => X"000000000000000000000000000000000000000000000003FF45FF8400145FFD",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000020000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(8),        -- Port A data input
DOA(0)   => data_read_a_lo_256(8),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(8),        -- Port B data input
DOB(0)   => data_read_b_lo_256(8),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_9_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00018248A2840112C00002C18000002300500030B3132000400812006",
INIT_01 => X"A1400802000020490000000000000240413C0A61590001D90213C90008510204",
INIT_02 => X"680108200010000054655C040080000041000000010402400800800009082011",
INIT_03 => X"00040100800020D0842240124210810042800504488000103081894288800000",
INIT_04 => X"00001410A00AA084000400C0060000040088323044201C850020820400101880",
INIT_05 => X"0200020040048A09202420000C00410402000025000800020804203000100800",
INIT_06 => X"22320400404048041144A7D2003A002012120004DC08125400A0008300821000",
INIT_07 => X"06181020421C08000940820000800010200018B20206C00000200002441223C1",
INIT_08 => X"0184010110120008004000000000061F02040826400008118000440000040000",
INIT_09 => X"8208888210004009010852882000510230A900A8040080800055086002200280",
INIT_0A => X"1402008004814948100004590111C004040120000020080121024012A4081200",
INIT_0B => X"2C91844522A0004100488000801200D00000880001000415E1248002103C2294",
INIT_0C => X"080040820408004082040800408202040020410402000000400809080508A080",
INIT_0D => X"0B4000803200C150108008490809A00219246101100220202102020820408204",
INIT_0E => X"00160006000120002120499020A04A14650A328519629651900142002404201E",
INIT_0F => X"0000080A20010002100000001402008002100000001402000001426008208041",
INIT_10 => X"0000000034008002800000001402008002800000001402008800000800000000",
INIT_11 => X"0008000000000000081500010000100800000000000008C10008000001200000",
INIT_12 => X"0088000000680005800002000000000000500000000000000004810010000800",
INIT_13 => X"02E8040200000003401F80004000000000040027000274000900000001A05D00",
INIT_14 => X"3B8000030000000000042B00009AB00008800000000008012BA010010000000D",
INIT_15 => X"0106520350000040100000000000010C0300009BA000200000000000105C0002",
INIT_16 => X"6651B328CA8D26540544924272EB91004002022024048400000098030A000A00",
INIT_17 => X"2509425094250942509425094250942509425094250942509425194651946519",
INIT_18 => X"5094250942509425094251946519465194651946519465194651946519465194",
INIT_19 => X"0480800000000000000001465194651946519465194651946509425094250942",
INIT_1A => X"34D34D34D1285B080201C92410480AB9A26667A46F345448020082E1C712A054",
INIT_1B => X"8341A0D068341A0D06834514514514514514514514514514514514514514D34D",
INIT_1C => X"F8B2B60D069349A0D068341A4D268341A4D268341A0D069349A0D069349A0D06",
INIT_1D => X"EFA2FFFFF555D000000000000000000000000000000000000000000000007FFF",
INIT_1E => X"F55087BC01EF007FD75FFFF84000AAFFD57DF45A280154BA5555401EFFFD5421",
INIT_1F => X"20AAAA843DFEF00517DEBA007BFDFEFFFD1575EF00557DF555D040000000043D",
INIT_20 => X"68AAAF7802AA00FFFBD7555087BC00AAF7D5575455D557DFEF002AAAB55002E8",
INIT_21 => X"A95545552ABFE00087BC00AA082EBFE10A28028AAAAAAABDF45F7803FFEF5555",
INIT_22 => X"FBC20BA5D7BEAAAAFFFBC00AA552E95545087BD54BA550417400085155555082",
INIT_23 => X"2FFFDF555D7BE8BFF5D51575EFA280175555D043DFEFA2FBD54BA5555554BAAA",
INIT_24 => X"00000000000557FF45002A975FF007BE8BFFA2FBFFFFFAAD5400AAFF8402000A",
INIT_25 => X"2415B471C7E3DF451EFBEFBFAF45490000000000000000000000000000000000",
INIT_26 => X"45490407000140038F450075C71FF087BD75D7FF84050BAEBDF78F45B6801048",
INIT_27 => X"FD7082EAAB550820870BAAA8438FFF00517DE82007FFAFEFE3DB505EF1C5B7AF",
INIT_28 => X"8F45F78A3DFD741516DAAAE38E2DA28EBFFD55451C7FC70BAE3D155555415178",
INIT_29 => X"1543808515756D1C2497545552AB8E10007FC50BA002ABFE00AA8A2AABABEAEB",
INIT_2A => X"FD04AA415B52492B6F5C20825D7FE8A92FFFFC20BA5D2E905550071D54825D0A",
INIT_2B => X"DB45082EB8002000AAFFFDF6D417FEABEF5D55505FFBE801256D490E3DFFFAAF",
INIT_2C => X"0000000000000000000000000000517DF451C24955EF0875EFBD7B6F1FFFC7BE",
INIT_2D => X"A2FBEAB45F78402010007BD5545AAFFD55EFF7FBE8B550000000000000000000",
INIT_2E => X"FAAFFC01FF557FE8B550004174105D042AB550055555FF007BD7555F784174AA",
INIT_2F => X"BAAAD15754508556AB45002AA8B450800174BAA68028BEF00517FE10007BE8BF",
INIT_30 => X"E10AAAEA8ABAF7AAAAB45F7AEBFF4508557FEAAAAAEBFEAAAAFFD5545557FD54",
INIT_31 => X"0145005557400552A954BA0051575EF5504175555D2EA8A00087BD74BA082EBD",
INIT_32 => X"021FF002ABDFEFAAFBC00BA007BC0000FFD542000557FE8A00F3FFC00BA552E8",
INIT_33 => X"57DF55FFD57DF55FFFBD5400A28400010A2FBFDFFF007FE8BFF5551401EFF784",
INIT_34 => X"000000000000000000000000000000000000000000000517FF455D04155FF005",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000040000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(9),        -- Port A data input
DOA(0)   => data_read_a_lo_256(9),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(9),        -- Port B data input
DOB(0)   => data_read_b_lo_256(9),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_10_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000B0001800002840002C0000281800020030000000033022000000180006",
INIT_01 => X"0000098218302849180060000C00424040000000080000080200090008510200",
INIT_02 => X"0801080200100000044008000080000041000000002002400800000009008010",
INIT_03 => X"0001000004000040000202000000000802006400088000003080040008C10000",
INIT_04 => X"0000100022008000000C08C00C00000400201830040000040000000400001820",
INIT_05 => X"0200000040000000248080210044000400000000000800000004004010000800",
INIT_06 => X"0030040000404004000006D00008002010100000880800001000000030829000",
INIT_07 => X"02100000021008000940800001800010200018920206C01020200002440003C0",
INIT_08 => X"0084010110120010004000000000021F00000024400000008000440080040000",
INIT_09 => X"8288880010100001200852882004404000000008800000100001004202000280",
INIT_0A => X"0000008000020008100004590111824004000100000008012000401084080200",
INIT_0B => X"AC04400022808001200014000040001082800000000010500000010400808000",
INIT_0C => X"002200002000020002200022000020000100011082442000480909220001E020",
INIT_0D => X"0080000010044000000080080001800200000400020011000000200002000220",
INIT_0E => X"001000020001000020010010248000200010000800040000008009040000002A",
INIT_0F => X"0000000A00010200800000001400008200800000001400000000024008208041",
INIT_10 => X"0000000024008200100000001400008200100000001400002800000000000000",
INIT_11 => X"0000000000000000001400012000200000000000000000C10008400080000000",
INIT_12 => X"8000000000480000040002040000001000000000000000000004800000002800",
INIT_13 => X"0000001000000002408000000000000000000025000200020000000001200000",
INIT_14 => X"0000040000000000000029000010000200000000000000012000001000000009",
INIT_15 => X"0100000000001000000000000000010401000010000000000000000000540002",
INIT_16 => X"00001400080002100544924002A000004000020000080000000010032A000000",
INIT_17 => X"4010040100401004010040100401004010040100401004010040000000000000",
INIT_18 => X"0000000000000000000001004010040100401004010040100401004010040100",
INIT_19 => X"1080800000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"8A28A28A28D532A0CCC2A28A28A7AA344854A07F069CB8930AFD6A1AAA902A14",
INIT_1B => X"4CA6532994CA6532994CA28A28A28A28A28A28A28A28A28A28A28A28A28A28A2",
INIT_1C => X"FB3CC772B94CA6532994CA6572B95CAE532994CA6532995CAE572B94CA653299",
INIT_1D => X"55A2AABFFEF0800000000000000000000000000000000000000000000000401F",
INIT_1E => X"4BA5555401EFFFD5421EFA2FFFFF555D003FE10AAFBE8AAAA2D540000F7D57DF",
INIT_1F => X"00AAFF8002155AAFFE8B45AAD540000087FFDF45FFFBC2010AAD57DF45A28015",
INIT_20 => X"D5400FFD568B555D00155EF08040000000043DF55087BC01EF007FD75FFFF840",
INIT_21 => X"43DFEF00517DEBA007BFDFEFFFD1575EF00557DF555D517FEBA082A801EFF7FB",
INIT_22 => X"2AAAB55002E820AAAA803FEBA082AAAAAAF7FBFDE00A2FBC0145005168A10AA8",
INIT_23 => X"FAEAAB55AAD568B455D00154BAFFFBD75EF5D7BC00AAF7D5575455D557DFEF00",
INIT_24 => X"000000000002ABDF45F7803FFEF555568AAAF7802AA00FFFBD7555082E82155F",
INIT_25 => X"AAAD547038EBD57DF7DA2AEB8FC7000000000000000000000000000000000000",
INIT_26 => X"38A2DF78F45B68010482415B471C7E3DF451EFBEFBFAF4549003DE10BEF5EDAA",
INIT_27 => X"1FF087BD75D7FF84050BAEB8002155BEF5EDB6DAADF470280075FFF45E3F1C70",
INIT_28 => X"DEAA0824851EFEBFBD2410EBD168B7D410A175C7000407000140038F450075C7",
INIT_29 => X"C2155005F68A10A28438FFF00517DE82007FFAFEFE3DB505EF1C5B7AF45495B7",
INIT_2A => X"155555415178FD7082EAAB550820870BAAA8038EAA0824A8AAAEBF5FAE28AAF1",
INIT_2B => X"FFD55451C2087155EBA4A8B7DAADF68B7D4104104AAF7F1D75EF557FC70BAE3D",
INIT_2C => X"00000000000000000000000000002EB8F45F78A3DFD741516DAAAE38E2DA28EB",
INIT_2D => X"00043FE00F7D17FEBAA2D5574BAAAD17DFEFA2AEAAB550000000000000000000",
INIT_2E => X"A00557FF45A2D5554AAA2FBEAB45F78402010007BD5545AAFFD55EFF7FBE8B55",
INIT_2F => X"105D042AB550055555FF007BD7555F784174AAA28002155FFD17FFFFA2FBD74B",
INIT_30 => X"1FF557FE8B55007FFDEAA0004175FFA2FBC2000AAD16ABFF002A975450004174",
INIT_31 => X"AABAAAD56AABAAAD140155087FEAA10A28028BEF00517FE10007BE8BFFAAFFC0",
INIT_32 => X"555EF557FD54BAAAD15754508556AB45002AA8B450800174BAA68428AAA08042",
INIT_33 => X"57FEAAAAAEBFEAAAAFFD5545550015555A2842ABEFAAFBE8BFF0004020AAFFD5",
INIT_34 => X"0000000000000000000000000000000000000000000002AAAB45F7AEBFF45085",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000047FFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(10),        -- Port A data input
DOA(0)   => data_read_a_lo_256(10),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(10),        -- Port B data input
DOB(0)   => data_read_b_lo_256(10),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_11_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10180B05A0010402840602C2D001019000000300000000330A20080EC180002",
INIT_01 => X"AB400984B830084C1820E0000C36424840000000080000088200000802112220",
INIT_02 => X"8801081438106400A4F55800008000004100000040CCE24208005000C9060032",
INIT_03 => X"000406A492E6E440842254D002108153432004800880000030C0315688C00006",
INIT_04 => X"00001201200090001205400000000094108C322644240C840008030440111800",
INIT_05 => X"222000444008010028404002A002009402400025080880000C04223000170900",
INIT_06 => X"0431018040014804920906C74B32002012121004540816544522008200821100",
INIT_07 => X"3A5B1220421408004A56E840008B90D0200018B60A0650D450FC800644A0438A",
INIT_08 => X"0485816170760268E04000000000323F42C50826490640D28088445B0E041900",
INIT_09 => X"820F8B2C100000808120308020024002B3B01AC9540080A623213008800A0280",
INIT_0A => X"10000080D80381881000045B0511D28D94012671272008013002000220001240",
INIT_0B => X"8811865D22BB384100E010908060349322008000A1001C49A9348498B0808010",
INIT_0C => X"50639504395063950639504395062CA821CA8210A0040000480808214001A020",
INIT_0D => X"088812203360410110A40008553980021040465602023269400A202863950439",
INIT_0E => X"01160006000101004A01811064B050204810240812241280D00200A08044290A",
INIT_0F => X"1B0482A01AAEC3602330CD2A02952DC3502330CB4A0318B41400024008208041",
INIT_10 => X"1630144C0155C3502330CD2A02952DC3602330CB4A0318B5600C587149B6D014",
INIT_11 => X"587083B6A51005956308D1E8202C436375908AA840AD4513437640F15245B455",
INIT_12 => X"67062F47B2872400044959BC42B1060F0D036B80B548523136C158878D8FE04E",
INIT_13 => X"7010A2699AAA3794392000D81852B0A050C224180062085134CD1719564E020C",
INIT_14 => X"400C50500D94C8121713C02B555101C90705D71009604140C0418CE0C378F0B2",
INIT_15 => X"27C828E024D8C50965A40821568A06113801505010334AA73AA0666DAC20AD57",
INIT_16 => X"048123408C0822040004C248604B2100400100084008001D0113920060CDC06A",
INIT_17 => X"4812048120481204812048120481204812048120481204812048120481204812",
INIT_18 => X"8020080200802008020081204812048120481204812048120481204812048120",
INIT_19 => X"1420000000000000000002008020080200802008020080200802008020080200",
INIT_1A => X"2082082082815220A4A380000002A8313044020C0605885026853A1082100A00",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000008208",
INIT_1C => X"F83F070000000000000100800000000000000000004020000000000000000000",
INIT_1D => X"EF0855400005500000000000000000000000000000000000000000000000401F",
INIT_1E => X"AAAA2D540000F7D57DF55A2AABFFEF0804155EFAA842ABEFA280155EFFFFBC01",
INIT_1F => X"FF555D51575FFA2FFD75FF550015400FFFBFFF4508514000000003FE10AAFBE8",
INIT_20 => X"155EF0051555FF0804155FFF7D57DF45A280154BA5555401EFFFD5421EFA2FFF",
INIT_21 => X"002155AAFFE8B45AAD540000087FFDF45FFFBC2010AAD568AAAAAD142145FF80",
INIT_22 => X"7FD75FFFF84000AAFF802ABFFA2AABFE1008001540008514215555003DFFFA28",
INIT_23 => X"85142010FFAE800AA5D7BFDF45F7FFEAA0000040000000043DF55087BC01EF00",
INIT_24 => X"00000000000517FEBA082A801EFF7FBD5400FFD568B555D00155EF085168B450",
INIT_25 => X"7BE8A155EFE3FBC71FF145B42038550000000000000000000000000000000000",
INIT_26 => X"381C003DE10BEF5EDAAAAAD547038EBD57DF7DA2AEB8FC70000175EFB6802DBC",
INIT_27 => X"1C7E3DF451EFBEFBFAF45495F575FFBEF5D05EF550E15400E3F1FFF7D085B420",
INIT_28 => X"8ABAB6D145145FF84155D7085B555C71404105C7F7DF78F45B68010482415B47",
INIT_29 => X"4515549003FFC7BE8002155BEF5EDB6DAADF470280075FFF45E3F1C7038A2DB6",
INIT_2A => X"038F450075C71FF087BD75D7FF84050BAEB8428BEFBEA4BDE28140A154380051",
INIT_2B => X"0A175C7005B6DB55145140000FFAE85082417FFFF7DE3F1EFA10140407000140",
INIT_2C => X"00000000000000000000000000005B7DEAA0824851EFEBFBD2410EBD168B7D41",
INIT_2D => X"0004175FFF7803DF45FFAE955EFAAFBD55EF557BC20AA5D00000000000000000",
INIT_2E => X"0AAD17DFEF007FC20AA5D043FE00F7D17FEBAA2D5574BAAAD17DFEFA2AEAAB55",
INIT_2F => X"45F78402010007BD5545AAFFD55EFF7FBE8B55007FD75FFF7D5401EF5D2E9741",
INIT_30 => X"F45A2D5554AAA2FBEAAAAFFD555545FF8015555007FD5545550400145FFFBEAB",
INIT_31 => X"DEAA5D2E974AA00515754500003FF55FF8002155FFD17FFFFA2FBD74BA00557F",
INIT_32 => X"7FE105D04174105D042AB550055555FF007BD7555F784174AAA2842ABEFFF803",
INIT_33 => X"BC2000AAD16ABFF002A97545007FFFF45555540000FFAE97410007BFFFFFA2D5",
INIT_34 => X"0000000000000000000000000000000000000000000007FFDEAA0004175FFA2F",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000040000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(11),        -- Port A data input
DOA(0)   => data_read_a_lo_256(11),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(11),        -- Port B data input
DOB(0)   => data_read_b_lo_256(11),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_12_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50080B01BC002006940202C0DE041196A83183000000023322287E0FC000006",
INIT_01 => X"0E000C048000C048400380000007026040000000080000088200002802153231",
INIT_02 => X"2809AD0E7D180040945008040090000061800000C0E2F66009DA3D11CB148015",
INIT_03 => X"210D050012F6F8D2108216E24842005B8A20640008800000B8E0141C28851006",
INIT_04 => X"0080100022408000060DE0000066630C70241827041000040800820480001AA4",
INIT_05 => X"0240000C400000003C808003E0C8001401000000040900020904004000070800",
INIT_06 => X"00300D800C1960C4400006E10B90002018184000100804005784000130821200",
INIT_07 => X"0652428112180C03E8E5A2C800A3F018200418927E06686450FF8006460003A0",
INIT_08 => X"09840903525281D4F460409000000E3F08D1202C5C26A0719CC96CC7BF462990",
INIT_09 => X"82488BAE10000040000410802008600843001E09F00000276F81020000230280",
INIT_0A => X"00000080000C000C100204593F11A489F480067D04D40C012400080000800240",
INIT_0B => X"0800021826933E03662802B300003C13E0000000460000000000010CE0000000",
INIT_0C => X"78419784197861978419784197860CBC30CBC20000000010400808056500A080",
INIT_0D => X"201E7F3F01F40401C17E800C7F33800200000357008C0249E2DE0D7841978619",
INIT_0E => X"0F500002200004005002001408400000000000000000000053A4096F80705FA0",
INIT_0F => X"1B17B2C53F2FC16691DB587201EDDF4162B1DB527201EDDC4607024100100020",
INIT_10 => X"F2A01D5CC9794162B1DB587201EDDF416691DB527201EDDD884272592D6246FC",
INIT_11 => X"7258E995D5A825DBA569F9FF02547068618CD3CC45B7863AE7EC00D4B122A67D",
INIT_12 => X"C6CCA5C33717461C045B5B182019473D19D7CCD856106F31A683621BDFC28800",
INIT_13 => X"FB10A652CC8E3538BBA01624E51AA6C0469AC5493F5688532966471A9C5F6208",
INIT_14 => X"40041E1F5759001B4AA1853E6D5144AA9C914C8608D2724A4C4118D992B866E2",
INIT_15 => X"AD9825682D4A36C0B0B4B85112B2C4A05D3E6D5051893335EB0072AA85A4F9B7",
INIT_16 => X"000008000000821000048260020000004001DC0800000010E7F70171401DE07E",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0100401004010040100400000000000000000000000000000000000000000000",
INIT_19 => X"1080800000000000000000040100401004010040100401004010040100401004",
INIT_1A => X"249249249120780800016A28A288028DCA30444409B054A88C5890486582A210",
INIT_1B => X"86432190C86432190C8641041041041041041041041041041041041041049249",
INIT_1C => X"FBC007592C964B2592C964B2592C964B2592C964B2592C964B2592C964B2592C",
INIT_1D => X"FF55002ABEF0800000000000000000000000000000000000000000000000401F",
INIT_1E => X"BEFA280155EFFFFBC01EF0855400005555421FF00042ABEFFF8400010082EAAB",
INIT_1F => X"FFEF08556AA10000028AAAFFD15541000002ABEFFFFBD54000004155EFAA842A",
INIT_20 => X"001FF00041554555557FE005D003FE10AAFBE8AAAA2D540000F7D57DF55A2AAB",
INIT_21 => X"1575FFA2FFD75FF550015400FFFBFFF45085140000005168AAA087BFFFFF5D04",
INIT_22 => X"D5421EFA2FFFFF555D0000145082E955FF0851555FF082AA8B55F7AEA8BEF555",
INIT_23 => X"000020BAAA801541055042ABEFFFFBD5410AAD57DF45A280154BA5555401EFFF",
INIT_24 => X"000000000005568AAAAAD142145FF80155EF0051555FF0804155FFF7842AA100",
INIT_25 => X"7EB80000280824ADBD7490E28BEF080000000000000000000000000000000000",
INIT_26 => X"101C00175EFB6802DBC7BE8A155EFE3FBC71FF145B42038555F401D71C0A2DBC",
INIT_27 => X"038EBD57DF7DA2AEB8FC7005F6AA381C0A2DA82FFDB5243800002FBD7EBFBD24",
INIT_28 => X"AA82147FF8FEF410E001FF000E17555555B7AE1041003DE10BEF5EDAAAAAD547",
INIT_29 => X"ADB45F7AEA8BEF555F575FFBEF5D05EF550E15400E3F1FFF7D085B420381C5B6",
INIT_2A => X"010482415B471C7E3DF451EFBEFBFAF4549000017D142E905EF1451525C7082A",
INIT_2B => X"04105C7F7842FA381C0A00082AA8A1041041002FBEFEBFBD2410AADF78F45B68",
INIT_2C => X"00000000000000000000000000005B68ABAB6D145145FF84155D7085B555C714",
INIT_2D => X"5D7BC01555D2EBFF55A284000AA08003FF55002AA8BEF0000000000000000000",
INIT_2E => X"A08003FF55A2FBC00105D04175FFF7803DF45FFAE955EFAAFBD55EF557BC20AA",
INIT_2F => X"00F7D17FEBAA2D5574BAAAD17DFEFA2AEAAB55007BE8AAA5D2EBDE00FFFFC00A",
INIT_30 => X"FEF007FC20AA5D7BE8A005D7FEABFF002E821FF082A97555557FE8A0000043FE",
INIT_31 => X"01EF5D5142145082EBFF55F7AAAABEF5D7FD75FFF7D5401EF5D2E97410AAD17D",
INIT_32 => X"C2010A2FBEAB45F78402010007BD5545AAFFD55EFF7FBE8B550004001FF5D2A8",
INIT_33 => X"015555007FD5545550400145FF843DEAA552A82010A2AA8000008043FFFFA2FB",
INIT_34 => X"0000000000000000000000000000000000000000000007BEAAAAFFD555545FF8",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000007FFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(12),        -- Port A data input
DOA(0)   => data_read_a_lo_256(12),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(12),        -- Port B data input
DOB(0)   => data_read_b_lo_256(12),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_13_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10110A0441812402840402822007818000E00700000000330A3000000008042",
INIT_01 => X"A1400984B830C848180260000C0042404001000008220008A200100802110200",
INIT_02 => X"88010C02801040002475580400800000410000000064024608134C0CC9018034",
INIT_03 => X"00010100926220D084234212421085084300648A0880000630C0654288C10000",
INIT_04 => X"0004122122029100100C00001200009C40A83A2044360C84190BAC04E0101820",
INIT_05 => X"027000004009050064C8C00104C10184034010250089C00EB004327064B60900",
INIT_06 => X"543000004080480492A946CE1032002012125804440812541027008230821380",
INIT_07 => X"0A581424525408000AE2AA8002BC00D020003896020658FC4030000246E543AE",
INIT_08 => X"04840101107200B80040210000002ABF02450A264002C8008000441680041900",
INIT_09 => X"825A98801000008001041080200B660E30B200C8840080808065102000280280",
INIT_0A => X"00000080C90391881000145B0111A30404016003A56008012C80080200801280",
INIT_0B => X"08088C5D2288004120E80290882400908000A000A1000809A93485D610000000",
INIT_0C => X"002000000000000002000000000000001000000000000000400808154100A080",
INIT_0D => X"08000000360401021280800E400B800610C84100014224200000000020000000",
INIT_0E => X"0086000600040D045E4195104D5854284A14250A12A512A8808289840084A020",
INIT_0F => X"0949E07A80948354B6E68982167061037496E683821670620681024000000000",
INIT_10 => X"8E510B456587037496E689821670610354B6E6838216706220431961CA985D48",
INIT_11 => X"196186A91674011CE61403562274AA49CD594CF00039C7C414B6509DA2265213",
INIT_12 => X"A983014780CC8604040424A5323845932E620295879818170304B2F5002C2043",
INIT_13 => X"451654B9104A328665603148895D44E0251142B42A3D8B2A5C8825194328A2E6",
INIT_14 => X"C06A6C6A465AA0091482382B17614F2202858EE300991415B45CD5306028F019",
INIT_15 => X"52E08DC8047F17D1C7C3C02128E587D6A02B17605A130A4E8BF002258850AC5D",
INIT_16 => X"84A123508508220808048240604B2100C00022084809000D000393722A140000",
INIT_17 => X"4A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A12",
INIT_18 => X"A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A128",
INIT_19 => X"154000000000000000000284A1284A1284A1284A1284A1284A1284A1284A1284",
INIT_1A => X"BAEBAEBAEBFF6FEFEFEEEAAAAAAFBF7DDF77F9FBEFBFF9F3F0FDFCFBEFBF1228",
INIT_1B => X"5FAFD7EBF5FAFD7EBF5FAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAE",
INIT_1C => X"F800077EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF",
INIT_1D => X"00FFD140155F780000000000000000000000000000000000000000000000401F",
INIT_1E => X"BEFFF8400010082EAABFF55002ABEF08556AAAA5D043FFFFAAAABDEAA557BFDE",
INIT_1F => X"000055043DEBAF7843FFFFF7AABDF55A2AA97400AAD540155A2D5421FF00042A",
INIT_20 => X"E8B45557FD7410552EAAABAAA84155EFAA842ABEFA280155EFFFFBC01EF08554",
INIT_21 => X"56AA10000028AAAFFD15541000002ABEFFFFBD5400005568A1055043DEBAAAFF",
INIT_22 => X"D57DF55A2AABFFEF085557545FFD17DEBAA2FFE8ABAAA8428A00087BD7555FFD",
INIT_23 => X"57BEAABA5D2ABDF450851420AA5D7FD5555A2803FE10AAFBE8AAAA2D540000F7",
INIT_24 => X"000000000005168AAA087BFFFFF5D04001FF00041554555557FE005D00001555",
INIT_25 => X"7AAA4B8E824971F8E38E3DF45155EB8000000000000000000000000000000000",
INIT_26 => X"55A2DF401D71C0A2DBC7EB80000280824ADBD7490E28BEF08516DA82410A3FFD",
INIT_27 => X"5EFE3FBC71FF145B42038550E38E92EB803FFD7EBA4BDF45AAAA90410BEDF451",
INIT_28 => X"FA38490A3FE92BEFFEAB45417FD24385D2AAFA82B680175EFB6802DBC7BE8A15",
INIT_29 => X"28A10007FD557DFFDF6AA381C0A2DA82FFDB5243800002FBD7EBFBD24101C556",
INIT_2A => X"5EDAAAAAD547038EBD57DF7DA2AEB8FC700515056DE3D17FE92BEF1EFA92AA84",
INIT_2B => X"5B7AE10410E00155497FEFABA4120B8F55085B400925D7FD557DA2803DE10BEF",
INIT_2C => X"00000000000000000000000000005B6AA82147FF8FEF410E001FF000E1755555",
INIT_2D => X"00517FE00082EBDF45AA8428A10085568ABAA2FBD7545AA80000000000000000",
INIT_2E => X"5AAAE82000F7FBD5545AAFBC01555D2EBFF55A284000AA08003FF55002AA8BEF",
INIT_2F => X"FFF7803DF45FFAE955EFAAFBD55EF557BC20AA5D2EA8A00A2803DF45AA843DF5",
INIT_30 => X"F55A2FBC00105D517FEAA082EBFE10F7FFE8B55087FC00BA552ABFE10F784175",
INIT_31 => X"FE10F7D57DE00AA842AA00007FD75FFF7FBE8AAA5D2EBDE00FFFFC00AA08003F",
INIT_32 => X"D55FFAA843FE00F7D17FEBAA2D5574BAAAD17DFEFA2AEAAB550051401FFA2D57",
INIT_33 => X"E821FF082A97555557FE8A00002E82155007BFDEAA08042AB45087FC0010557F",
INIT_34 => X"0000000000000000000000000000000000000000000007BE8A005D7FEABFF002",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000067FFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(13),        -- Port A data input
DOA(0)   => data_read_a_lo_256(13),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(13),        -- Port B data input
DOB(0)   => data_read_b_lo_256(13),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_14_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10020A000180000284008280000281800000030000000033022000000580002",
INIT_01 => X"A140098018300848184860000C20C24040000000084000084200000000110200",
INIT_02 => X"88010C5A8010A600A4F558040080000041000000022C024008003CCCC9028030",
INIT_03 => X"000103A7A00904D0842242024210810803006480088000003081054288C10000",
INIT_04 => X"0000120122009000100C00000000000400A83A2044200C840000800400101820",
INIT_05 => X"020000004008010024C0C0010040000402000025000800020004207000100800",
INIT_06 => X"0430000040004804920906C20022002012120004440812541020008230821000",
INIT_07 => X"2A5A14285A15080008768A80008000D0200018B202067AF100A0000244204382",
INIT_08 => X"04850101105205380040000000000A7F42840A264920406080004400A0040900",
INIT_09 => X"8208888010000080010010802000400230B000C8840080800021100000200280",
INIT_0A => X"00000080C8038188100004590111B68404012000016008012000000000000200",
INIT_0B => X"080084452280004120400000802000908000800001000009A924810410000000",
INIT_0C => X"000000000000200000000000000200000000000000000000400808000000A080",
INIT_0D => X"080000002204010010808008000B800210404100000220200000000020000200",
INIT_0E => X"0000000600000000020181100400502048102408122412808082098400042020",
INIT_0F => X"0480040A100A42008000161C140000420080001C1C1400003201024000000000",
INIT_10 => X"39600022260042001000161C140000420010001C1C140001604E8084341CBA34",
INIT_11 => X"8082580E2B8802201014800C220A21829A302F1C024010C001124020C8C1A8A0",
INIT_12 => X"CA60CA000048228404401004418012787124648157780120B8678C000801E04E",
INIT_13 => X"001072D04730000241000CB1325E78E0186030240000083B602398000120024A",
INIT_14 => X"001EF6F4163C480481506800004000CFD55196CB012481812049495C19400009",
INIT_15 => X"248800108B8FB61A0401200845594965000000400568D0CFB780055060500001",
INIT_16 => X"048123408408220000048240604B210040000008400800B0000090022A140068",
INIT_17 => X"4812048120481204812048120481204812048120481204812048120481204812",
INIT_18 => X"8120481204812048120481204812048120481204812048120481204812048120",
INIT_19 => X"1400000000000000000002048120481204812048120481204812048120481204",
INIT_1A => X"9E79E79E79FF3BEEEEEFE79E79EFAABCDA72E47F87BDF4EBAE7CFAFBEFB28200",
INIT_1B => X"CFE7F3F9FCFE7F3F9FCFE79E79E79E79E79E79E79E79E79E79E79E79E79E79E7",
INIT_1C => X"FBFFF83F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9F",
INIT_1D => X"555D5568A105D00000000000000000000000000000000000000000000000401F",
INIT_1E => X"FFFAAAABDEAA557BFDE00FFD140155F7D17DF45AAD157400007BEAAAAAAAE955",
INIT_1F => X"ABEF085155400FFD1420100055574AAA2AA800AAF784020AAF7D56AAAA5D043F",
INIT_20 => X"FFE105D7BD7545A284020BA0055421FF00042ABEFFF8400010082EAABFF55002",
INIT_21 => X"43DEBAF7843FFFFF7AABDF55A2AA97400AAD540155A28028B550051574005D7F",
INIT_22 => X"FBC01EF08554000055002AB455D51420100851421FF5D7FFDEBA085168B45FF8",
INIT_23 => X"AD140000002EBFFEFA2AAA8BEFF780021FF5504155EFAA842ABEFA280155EFFF",
INIT_24 => X"000000000005568A1055043DEBAAAFFE8B45557FD7410552EAAABAAA8017400A",
INIT_25 => X"01C71EDA82AAA0955455D556DA00490000000000000000000000000000000000",
INIT_26 => X"BAEBD16DA82410A3FFD7AAA4B8E824971F8E38E3DF45155EBD17FF6DAADB5040",
INIT_27 => X"0280824ADBD7490E28BEF085157428FFDB420101C55554AAAAA480082FF84000",
INIT_28 => X"AB7D0051504005D71F8E004975D556DB68405092085F401D71C0A2DBC7EB8000",
INIT_29 => X"FAEAA08516AB45E38E38E92EB803FFD7EBA4BDF45AAAA90410BEDF45155A28E2",
INIT_2A => X"02DBC7BE8A155EFE3FBC71FF145B42038550028B6D5D51420101C5B401EF417B",
INIT_2B => X"2AAFA82B68015400AADB40000082EBFFC7A2AEAFBC7EB80071FF5500175EFB68",
INIT_2C => X"0000000000000000000000000000556FA38490A3FE92BEFFEAB45417FD24385D",
INIT_2D => X"AAD17DFFFAAFFC200055557DE00A2801554555557FE100000000000000000000",
INIT_2E => X"AA28400000F784020BAAAD17FE00082EBDF45AA8428A10085568ABAA2FBD7545",
INIT_2F => X"555D2EBFF55A284000AA08003FF55002AA8BEF0051554AAFFFFC00105D55554B",
INIT_30 => X"000F7FBD5545AAAEAABFF0051400105D5568A000051575FFF78415410087BC01",
INIT_31 => X"2000557FC01EF007FEAABA00556AB55A2AEA8A00A2803DF45AA843DF55AAAE82",
INIT_32 => X"175FF5D04175FFF7803DF45FFAE955EFAAFBD55EF557BC20AA5D042ABFF55514",
INIT_33 => X"FE8B55087FC00BA552ABFE10F78415400A2FBC0010082EBDF55A2AABDF45A284",
INIT_34 => X"000000000000000000000000000000000000000000000517FEAA082EBFE10F7F",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000007FFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(14),        -- Port A data input
DOA(0)   => data_read_a_lo_256(14),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(14),        -- Port B data input
DOB(0)   => data_read_b_lo_256(14),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_15_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000A000000000284000280000001800020030000000033022000000180002",
INIT_01 => X"A140098018300848180060000C00424040000000080000080200000000110200",
INIT_02 => X"080108000010E60004E55800008000004100000000040240080000C009170016",
INIT_03 => X"0000000080000040842240000210810002000400888000003080014288C00000",
INIT_04 => X"0001100024A0800000440000000000040088322044200C840000011400151800",
INIT_05 => X"A200014C4000000020000000000B8094020000254C8800000514203000108800",
INIT_06 => X"0031042040804804100006EE4032002012120005540812540020008600831000",
INIT_07 => X"021912244A14080008408880008000D020001892020656300020000244000380",
INIT_08 => X"048501415032000800406180000002DF02440826400000008000440000043080",
INIT_09 => X"8208880110000000010010802000400230A000880400808000450200000B0280",
INIT_0A => X"00000080C003010810000459011182040400200003E0080120000000000002C0",
INIT_0B => X"080084452280004100400000800000100000800001000001A124800010000000",
INIT_0C => X"002000020000000000000000000200001000010000000000400808000020A000",
INIT_0D => X"08000000260001001280000C400B000200000000000220200000000020000200",
INIT_0E => X"008400060000000000010010040040000000000000201000000000000004A000",
INIT_0F => X"0000000000000202100000000000000202100000000000004600024000000000",
INIT_10 => X"0000000000000202800000000000000202800000000000002000000800000000",
INIT_11 => X"0008000000000000000000002000100800000000000000000000400001200000",
INIT_12 => X"00880000000006000400080C0000000000D08120280000000000000000002000",
INIT_13 => X"0010040200000000010000004020010000000000000008000900000000000200",
INIT_14 => X"0000000308801400000000000040000008822110000000000040100100000000",
INIT_15 => X"0080000000004840717050000000000000000040000020000000000000000001",
INIT_16 => X"000023000000220000048240404A010040000008000000000000000020C40000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"1400000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000200",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"F800000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"AA007BC2145F780000000000000000000000000000000000000000000000401F",
INIT_1E => X"400007BEAAAAAAAE955555D5568A105D7FC00000804154AA5D00001EFF78428A",
INIT_1F => X"0155F7FBD74AAAAD17DF45F7D1421EF0055400AA007FC2000F7D17DF45AAD157",
INIT_20 => X"BDFEF08517DF55A2FBEAB555D556AAAA5D043FFFFAAAABDEAA557BFDE00FFD14",
INIT_21 => X"155400FFD1420100055574AAA2AA800AAF784020AAF7FFFDF45FF84000BA552A",
INIT_22 => X"2EAABFF55002ABEF087BE8ABA555168B55AAFFEAB45F7843FF45082A801FF005",
INIT_23 => X"284000AA0055401550055574005D2E800AAA2D5421FF00042ABEFFF840001008",
INIT_24 => X"000000000000028B550051574005D7FFFE105D7BD7545A284020BA007FFFE10A",
INIT_25 => X"2550E021C7EB8028A821C7BC516DFF8000000000000000000000000000000000",
INIT_26 => X"28FFD17FF6DAADB504001C71EDA82AAA0955455D556DA004971C703814001248",
INIT_27 => X"E824971F8E38E3DF45155EBF1D5492BED17FF45E3DF471C70851400BA0071C50",
INIT_28 => X"FF7DEB8000092552ABFFEF08517DF6DB6FBE8B555D516DA82410A3FFD7AAA4B8",
INIT_29 => X"3DF551C20801C71C5157428FFDB420101C55554AAAAA480082FF84000BAEBF1F",
INIT_2A => X"A2DBC7EB80000280824ADBD7490E28BEF087FEFA8241516DB55A2FFEAB6DEB84",
INIT_2B => X"8405092087FF8E00BE8A02082005F47145085550428412A85082BEDF401D71C0",
INIT_2C => X"00000000000000000000000000000E2AB7D0051504005D71F8E004975D556DB6",
INIT_2D => X"0055554BA5504000105D2A80145AA842AA00557BD75EFF780000000000000000",
INIT_2E => X"50055420BA0055574BAF7D17DFFFAAFFC200055557DE00A2801554555557FE10",
INIT_2F => X"00082EBDF45AA8428A10085568ABAA2FBD7545AAD557410F7D57DF55AAFBD554",
INIT_30 => X"000F784020BAAAD57FFEFA28402010552ABDFFF08517FFFFF7FBEAB455D517FE",
INIT_31 => X"DF45AAFBE8BEFA2803FF455504001555551554AAFFFFC00105D55554BAA28400",
INIT_32 => X"95400F7FBC01555D2EBFF55A284000AA08003FF55002AA8BEF007FFDE1000557",
INIT_33 => X"568A000051575FFF78415410087FEAA10F7AE80000087BD55450855400BA002A",
INIT_34 => X"0000000000000000000000000000000000000000000002EAABFF0051400105D5",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000060000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(15),        -- Port A data input
DOA(0)   => data_read_a_lo_256(15),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(15),        -- Port B data input
DOB(0)   => data_read_b_lo_256(15),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_16_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"DA22C618B1000482B688B186588884862A400438255FC38381441205BA803003",
INIT_01 => X"8645A80028404C211203A952A90341080B173340412000E1005D628000820484",
INIT_02 => X"A101A9006DC1084833011850AAC55001349B10881802821808B4110007005E11",
INIT_03 => X"010108A802BB00080080006020020001A61036202800000D2410104200404550",
INIT_04 => X"8BFA58800005C40A46240252145148B38248030356415A4E62B6FC660F287240",
INIT_05 => X"0F05EA11E570000D610000000710296E542B6E3A825C15FB30A643695BFC2D56",
INIT_06 => X"00640044150C025A0000000901A054F2C0A8030140BCC0460050690A95C8383D",
INIT_07 => X"0288500102F85203E8010D0AA9BC4800015001219D0550077373CAA804000680",
INIT_08 => X"A2064193920A2004B51400001414091EAA14881C0002701881B120203B7A8012",
INIT_09 => X"C8204D02D965965200100104F2B0082251200000023153000C4400800000ACCA",
INIT_0A => X"000012C9000A0000D0A80000BF8028E87C1B9246002A8A562060410280081116",
INIT_0B => X"240014891801000495D40192D1000000000000A8A5AA80018120E00066000000",
INIT_0C => X"00088000880008800088000880008400044000400029011404008401CA809004",
INIT_0D => X"0140A80A5C8000102ED0044008004AD32400004001AB08C0031EDA7B08800088",
INIT_0E => X"04912AA28AA890BA00000024800480000000000000200802151025062C0BB400",
INIT_0F => X"1F554E11C596A64003195933741477264003195555B418687E35836020814004",
INIT_10 => X"0A499CF47DCB264003195933741597264003195555B4198843940076D296D003",
INIT_11 => X"00758486A556489347FE5F409CBC1362510695B6288743123C95251852041CD5",
INIT_12 => X"424EAE2992046EB70026486035600CEC45CBCA809654B48163CCC895E1E043D4",
INIT_13 => X"98E3A242DEA151848302BFD6D522B10C7EC71F6C1DB071D1216E078C4C1B1C74",
INIT_14 => X"037DAAABC982BE22267A2E2E4F44AA1DC5E37400C9EE1B7B638E8849D23C3832",
INIT_15 => X"2EE015998B28654565A003F0068E35352C1CAE48BFBF3A6C9B7B286B4DA8B93D",
INIT_16 => X"000009000040A8000452110A8442040D655602A102A0027E2C42320284086E6A",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"1451451451E96F2FC3C34F3CF3C2AC688AA263486D3260E34C0C3A7B451B0200",
INIT_1B => X"9F47A7D1E9F47A7D1E9F4D14D14D14D14D14D14D14D14D14D14D14D14D145145",
INIT_1C => X"F800007D3E9F4FA7D3E8F47A3D1E8F47A3D1E8F47A7D3E9F4FA7D3E9F4FA7D3E",
INIT_1D => X"FF00003FE005500000000000000000000000000000000000000000000000401F",
INIT_1E => X"4AA5D00001EFF78428AAA007BC2145F7843FFFFF7FBE8B45AAD568BFFFFAA975",
INIT_1F => X"8A105D2E974BAF7FBEAB45FFFFC00BAF780020005D2A95410FFFFC0000080415",
INIT_20 => X"821FFA2AAAAA00000417555FFD17DF45AAD157400007BEAAAAAAAE955555D556",
INIT_21 => X"BD74AAAAD17DF45F7D1421EF0055400AA007FC2000F78000010552E800AA002E",
INIT_22 => X"7BFDE00FFD140155F7AABDF55F7AE820AA08043FEBA5D55575FFF7AABFE00557",
INIT_23 => X"2FBE8B55FFFFD55FF557FC2000FF8015410FFD56AAAA5D043FFFFAAAABDEAA55",
INIT_24 => X"000000000007FFDF45FF84000BA552ABDFEF08517DF55A2FBEAB555D04154BAA",
INIT_25 => X"5B6DF6DBFFF7AA955C71C043FE10490000000000000000000000000000000000",
INIT_26 => X"38FFF1C7038140012482550E021C7EB8028A821C7BC516DFF8438FC7E3F1EAB5",
INIT_27 => X"A82AAA0955455D556DA00492490492F7FBE8B55FFF1C70BAF78A000005D20974",
INIT_28 => X"20285D2085092002A801FFB6AAA8A10080E1757DEBD17FF6DAADB504001C71ED",
INIT_29 => X"555FFE3AABFE005D71D5492BED17FF45E3DF471C70851400BA0071C5028FF840",
INIT_2A => X"A3FFD7AAA4B8E824971F8E38E3DF45155EBA4BAF6DE3AA8709208043FEBA555B",
INIT_2B => X"FBE8B555D04124BAB6FBE8B45E3FBD55D7557BC0028E38412428EBD16DA82410",
INIT_2C => X"000000000000000000000000000071FFF7DEB8000092552ABFFEF08517DF6DB6",
INIT_2D => X"F78428B55AAD168B55F7FFFDFEFFFAA9555555003DE000000000000000000000",
INIT_2E => X"AFFAE820105500154AAF7D5554BA5504000105D2A80145AA842AA00557BD75EF",
INIT_2F => X"FFAAFFC200055557DE00A2801554555557FE10000000010F7FBEAB45FFD1554A",
INIT_30 => X"0BA0055574BAF784000BA5D0017410082E801EFF7AEA8A10002E955FFA2D17DF",
INIT_31 => X"541000003DEBA557BD75EFA2AEBDE105D5557410F7D57DF55AAFBD5545005542",
INIT_32 => X"000AAAAD17FE00082EBDF45AA8428A10085568ABAA2FBD7545AA802ABEFA2AA9",
INIT_33 => X"ABDFFF08517FFFFF7FBEAB455D04020AAFFFBEAB45AAFFD55555D7FC20AAA280",
INIT_34 => X"000000000000000000000000000000000000000000000557FFEFA28402010552",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000020000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(16),        -- Port A data input
DOA(0)   => data_read_a_lo_256(16),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(16),        -- Port B data input
DOB(0)   => data_read_b_lo_256(16),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_17_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"5284CE4FB7BD2C8994A13392DBD02E14006B82AC7E800D44D3DD2FD5F9B961C0",
INIT_01 => X"F8ACD01F7E03FC6793F2199B39FC233C11D93AE6F3BB92B32091DBC339B24542",
INIT_02 => X"8F333007FD6808092A2AFA6667033DB50853379C10BFF70F1BD011110F205F18",
INIT_03 => X"294ADB4AFFCBF0DAD63ABF836B58EAFE060478202022234B2E0303FDC9E18339",
INIT_04 => X"DB7A40806FE4040840EBC563A0150A0926146FECB04196482236FC2005282AE1",
INIT_05 => X"0403DA0383200831C68206D7E6D0250834336D1E81500FDB306045255BFC2076",
INIT_06 => X"000A0E2D7D3EAFF15800100FBFB333C1CBC303163670497AFF00291B3C0E2015",
INIT_07 => X"451C581123AEE54DE8008B719E61C10BBA5DAAFA9DDA1194D51E067BB0000000",
INIT_08 => X"70320A9392083056C2270E004400091181168C4D14002A110C902481FC0B4212",
INIT_09 => X"0E28EFFC40C30E5F0182D0950190C0810BE00E9A76E4C7FD0E4700000B303806",
INIT_0A => X"C7DEF207000F00059D2ED56D7EED2ED3C9A86FB8013E7437823DF78CDB6CA60E",
INIT_0B => X"7C00319F8E853E64D73A08BFF0001D35682AC0CE8FCCC200A59BDD2FFE3F3EC7",
INIT_0C => X"7A7DE7A7DE7A7DE7A7DE7A7DE7A7DF3D3EF3D3C0030B889723782E816EC0A081",
INIT_0D => X"2D4CFEB69FF7A5F5AFFCCA787F7FE67C21800367451F8355EB9EDE7A7DE7A7DE",
INIT_0E => X"2C9F99FD0678B87A0003000D8D02E00000000000000040025D3C21463D6BFF25",
INIT_0F => X"232221ABD9CA854DFDD64A67D42C0F054DFDD64667D42C063E57A8F7B4594BB0",
INIT_10 => X"AEDAA504801F054DFDD64A67D42C0F054DFDD64667D42C07237DFE5865F6D2BF",
INIT_11 => X"FE58EAE7F5AB50D0806A9A2E0DFFF47DEDC496DA3181A0CC71440F9FBC3EFBB5",
INIT_12 => X"9C9C3FC95949AEFF556EF9C75E7DCF1EB1B6E6FCDC87CB35FC94B36AECF3A33D",
INIT_13 => X"382AF5B6AAAE594A4C0DBFDAD94AA669809809FEFAF4157ADB55572CA527056E",
INIT_14 => X"1AE33F32ADD543430808BABAF50E1A5EB4BAEA45A250202FE0ADD39387F92B29",
INIT_15 => X"669523E865D4B1293AB6B90BF2F0E30EDEFAFD0B3FBD72E9E90D20A003FBEBF4",
INIT_16 => X"00002F840000BCE0B6F67B3F845E017C833F6AAC02B002A2EFF22D4073DE83FB",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0600000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"9A69A69A6A4624C3434C0EBAEBA21B9001804F6E62029749701020B88A7CC0C0",
INIT_1B => X"41A0D46A341A0D46A341A69AEBA69A69AEBA69AEBA69A69AEBA69AEBA69A69A6",
INIT_1C => X"F8000046A351A8D46A351A8D46A351A8D46A351A8D068341A0D068341A0D0683",
INIT_1D => X"00F7D56ABFF55000000000000000000000000000000000000000000000007FFF",
INIT_1E => X"B45AAD568BFFFFAA975FF00003FE0055043FFFFFFFFFFFFFF7FBFDF55A284020",
INIT_1F => X"2145F7D568B45000002010552EBDF45A28028A00F7843FEBA55043FFFFF7FBE8",
INIT_20 => X"95410AAAEBFF55AAFFC00BAF7FFC00000804154AA5D00001EFF78428AAA007BC",
INIT_21 => X"E974BAF7FBEAB45FFFFC00BAF780020005D2A95410FFAE800105D2A95410002A",
INIT_22 => X"AE955555D5568A105D7FFFFEFA2D568BFFFFD57DE00F7AE800AAAAAABDFEF5D2",
INIT_23 => X"82A974105D003FF55F7802AAAAAAD168AAA5D517DF45AAD157400007BEAAAAAA",
INIT_24 => X"000000000000000010552E800AA002E821FFA2AAAAA00000417555FF8028B550",
INIT_25 => X"FE3F5FAF45AA8000038F7DB6FBD7490000000000000000000000000000000000",
INIT_26 => X"82490438FC7E3F1EAB55B6DF6DBFFF7AA955C71C043FE10490A3FFFFFFFFFDFE",
INIT_27 => X"1C7EB8028A821C7BC516DFFDF68B551C0E050384124BFF7DB68A28A38F7803DE",
INIT_28 => X"5000492495428082E95400AAA0BDF7DB6F5C70BAFFF1C7038140012482550E02",
INIT_29 => X"800BAB6AEBDFD75D2490492F7FBE8B55FFF1C70BAF78A000005D2097438FFAA8",
INIT_2A => X"B504001C71EDA82AAA0955455D556DA00497FFAFFFB6D56FBFFEBDB78E38F7AA",
INIT_2B => X"0E1757DEB8A2DB5514249243841003FF6DEB8028AAAB6D16FA8249517FF6DAAD",
INIT_2C => X"000000000000000000000000000004020285D2085092002A801FFB6AAA8A1008",
INIT_2D => X"002ABFFEFF7FBFDFFFAAD168B55AA80000BAF7FFFDF550000000000000000000",
INIT_2E => X"FFFAAA8AAAF7843FE10000428B55AAD168B55F7FFFDFEFFFAA9555555003DE00",
INIT_2F => X"BA5504000105D2A80145AA842AA00557BD75EFF7FBEAB45552E954BA08003DFF",
INIT_30 => X"0105500154AAF7AE974000800154AA002E95410AA843FFFFF7D5554BAF7D5554",
INIT_31 => X"FFEFAAFFE8ABAFFAA820BAF7AEBFF55550000010F7FBEAB45FFD1554AAFFAE82",
INIT_32 => X"7DE0000517DFFFAAFFC200055557DE00A2801554555557FE10007FEABEFFFD57",
INIT_33 => X"E801EFF7AEA8A10002E955FFA2AABFF455500020AA08003DFFFA28028AAAF7D1",
INIT_34 => X"00000000000000000000000000000000000000000000004000BA5D0017410082",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000067FFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(17),        -- Port A data input
DOA(0)   => data_read_a_lo_256(17),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(17),        -- Port B data input
DOB(0)   => data_read_b_lo_256(17),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_18_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"69844019080000A21A611406840014122A641074155FC28A2024001001801003",
INIT_01 => X"A643D920034004180005E9E3C90360C0041C0181002001602025800008440084",
INIT_02 => X"B7333980808408103F2000F81FC0FEDEAC2161B0B84D0002188011110C018041",
INIT_03 => X"0405D434003F2C020081587008020561E55116B0290000042B71240C800440F8",
INIT_04 => X"50805AC31007D6125724029216554A9847669903D640EC8E2001002604503004",
INIT_05 => X"07008000E0EA11803850C800010022660C1C0065003C0404002646DC20A02D40",
INIT_06 => X"8560000000022229A60B048048120FF040000000002C44D620F0228454C83810",
INIT_07 => X"058800A001D4033A004904087F9E3901218050018024110D6771C1F90C285682",
INIT_08 => X"F3020A82929A807B3731021400058C020000A9729400D10100420480202AC214",
INIT_09 => X"C820C802D86184A010180304307008025414204400220202F1A814A0080064C1",
INIT_0A => X"080003C32A10A19090C02010E10229440616900000022E0C6070000504102805",
INIT_0B => X"026226495446E2110AE44174112840880000060D7030C30B885200D274004008",
INIT_0C => X"840018400184001840018400184000C2000C200200301500C404C001B884B806",
INIT_0D => X"81010108003C000210020460801001FB3650D89888E06CAE1061018500184001",
INIT_0E => X"032007E281F840C00284A17210001060D8306C18360C1380A0260CB980840080",
INIT_0F => X"5D79BBEF8E50B041029075982BF3873041029079982BF39748AA0AC800014804",
INIT_10 => X"EA479BFD7F7F3041029075982BF3E73041029079982BF3F632C5F96D3C11555D",
INIT_11 => X"F96A595405FC7F1CFEBC7586C4100A53162B47FD7E39FFEECE1598702345156A",
INIT_12 => X"006FE037ACFB88083A99E06271BB0CA207DFDD5920057E0B001B0EBCC79932C5",
INIT_13 => X"5CA2A002DD51B6F7FC4A411D1E8D44517F14EAFE36E55150016EA8DB73E39464",
INIT_14 => X"953C30351452A13D55CFFA76E928E3891F148B30399F5FB7F28C800DFA06F5DF",
INIT_15 => X"5AC57DFEAEF1005475F1D1F608819CF0EE76E12C824ADD9089715F25FAF9DB84",
INIT_16 => X"0D834041A41A0000010180C02801680460FC900052FA10DC0006DA4881C11015",
INIT_17 => X"D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D836",
INIT_18 => X"8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360",
INIT_19 => X"00000000000000000000020D8360D8360D8360D8360D8360D8360D8360D8360D",
INIT_1A => X"8A28A28A2891182C8A82E0820825945DF675C0770B9E11807E54587BEF8B0000",
INIT_1B => X"44A2552A954AA5128944AAAA28A28A28AAAAAAA28A28A28AAAAAAA28A28A28A2",
INIT_1C => X"F80000128944A25128944A25128944A25128944A25128944A25128944A251289",
INIT_1D => X"BA5D04174AA0000000000000000000000000000000000000000000000000401F",
INIT_1E => X"FFFF7FBFDF55A28402000F7D56ABFF55043FFFFFFFFFFFFFFFFFFFFEFF7AE954",
INIT_1F => X"FE0055043FFFFFFFFFDFEFA2D56AB45AA8400145AA801741000043FFFFFFFFFF",
INIT_20 => X"FFFFFFF80021EF0855421EF00043FFFFF7FBE8B45AAD568BFFFFAA975FF00003",
INIT_21 => X"568B45000002010552EBDF45A28028A00F7843FEBA55557FFEFA2D168B55AAFB",
INIT_22 => X"8428AAA007BC2145F7D5400000004020AA5D2A82155F7AEBFEBAFFD56AA00A2D",
INIT_23 => X"82E954BA0004174AAAA8428B45082ABFEBAA2FFC00000804154AA5D00001EFF7",
INIT_24 => X"000000000002E800105D2A95410002A95410AAAEBFF55AAFFC00BAF7AE800100",
INIT_25 => X"FFFFBFDFEFFFAE954AA550415492140000000000000000000000000000000000",
INIT_26 => X"10140A3FFFFFFFFFDFEFE3F5FAF45AA8000038F7DB6FBD7490E3FFFFFFFFFFFF",
INIT_27 => X"BFFF7AA955C71C043FE1049043FFEFE3F1F8FD7AAD16FB6DBE8E00155BE80154",
INIT_28 => X"8FC7AAD56FB6DBEF1FAFD7E384001EF145B471C7140438FC7E3F1EAB55B6DF6D",
INIT_29 => X"BDE92FFD56FA28B6DF68B551C0E050384124BFF7DB68A28A38F7803DE82495B7",
INIT_2A => X"012482550E021C7EB8028A821C7BC516DFFD1420381C0A02082492A85155E3A4",
INIT_2B => X"F5C70BAFFAE870280024904BA1400174AABE8E28B7D1420BDEAAA2F1C7038140",
INIT_2C => X"00000000000000000000000000002A85000492495428082E95400AAA0BDF7DB6",
INIT_2D => X"002ABFFFFFFFFFFFEFF7FBFDFFFF7AA974BA5504154105500000000000000000",
INIT_2E => X"FF7AA82155F78015400552ABFFEFF7FBFDFFFAAD168B55AA80000BAF7FFFDF55",
INIT_2F => X"55AAD168B55F7FFFDFEFFFAA9555555003DE0000043DFEFA2D56AB45AAD57DFE",
INIT_30 => X"AAAF7843FE10007FEAB55A2D17FFEFFFD568B55A280021EF557FD7555550428B",
INIT_31 => X"2000002A95545A2843FE00F7D17FEAAF7FBEAB45552E954BA08003DFFFFFAAA8",
INIT_32 => X"3DEAAA2D5554BA5504000105D2A80145AA842AA00557BD75EFF7D1400AA5D2A8",
INIT_33 => X"E95410AA843FFFFF7D5554BAF7AE974BA0004020AA5D04154BAF7AEA8BEF5500",
INIT_34 => X"0000000000000000000000000000000000000000000002E974000800154AA002",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000020000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(18),        -- Port A data input
DOA(0)   => data_read_a_lo_256(18),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(18),        -- Port B data input
DOB(0)   => data_read_b_lo_256(18),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_19_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"042200000000000041088001001AA00000000000000000000000500802000003",
INIT_01 => X"200048000024000000000404000000000A22000800000800004A200000000001",
INIT_02 => X"032210008DEF00400060000001C008002489E0F0004037B00010101010000000",
INIT_03 => X"0000008128000000000000000000000024001620280000000000354200004008",
INIT_04 => X"000058800004C4024024001210001054B1C822009640000E2000002604003000",
INIT_05 => X"07008000E0200000000000000000200604000000001C04000026400000002C40",
INIT_06 => X"000000000000000100000000000001B040000000002C42010010200004C83810",
INIT_07 => X"0E0050A040041593104004500480090080A01120220140020420401800000000",
INIT_08 => X"130E409080188000021A0000100004082A140102B4020109801A4CE003710010",
INIT_09 => X"C80000005861840000000004301000B000000000001C1C0000000000000020C0",
INIT_0A => X"000002C30000000040500010301020400000000000022A040000000000000004",
INIT_0B => X"00000020001000022000000000000000000002F0001F00002024B20002000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"00108000EC000000000000000010004B20000000000000000000000000000000",
INIT_0E => X"0000006280180040000000000000000000000000000000000000000000000000",
INIT_0F => X"8084451B81A70AB3006BA0011400760AB3006BA0011400680F02096834820000",
INIT_10 => X"11204082248A0AB3006BA0011400160AB3006BA0011400084C780687DBA82800",
INIT_11 => X"068796E80A00802301BC0A7531EDD98E73B02800804620D030F873EB49F30B80",
INIT_12 => X"6B00000002044F091A860700FF9198AA115D5DA37F7A80C8A3604001C0664C78",
INIT_13 => X"98551AC9000000000314E01F9F30198600631448410A2A8D64800000081B0A93",
INIT_14 => X"2E00303842281C80A23004411AD661891F15148A4420804241526D6000000000",
INIT_15 => X"9D335F3D282000C6C5456C84850F61050C411AD6284FDA861682805A04A1046B",
INIT_16 => X"00000000000000000000000000000004600C0013800003088004202304366A4A",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"86186186186851046260A9A69A6039045DD1F863808633005010063A20C90000",
INIT_1B => X"D26930984C26130984C261861861869A61861861861869A61861861861861861",
INIT_1C => X"F800000984C26130984C26130984C26130984C26130984C26130984C26130984",
INIT_1D => X"BA5500020BA5D00000000000000000000000000000000000000000000000401F",
INIT_1E => X"FFFFFFFFFFEFF7AE954BA5D04174AA007BFFFFFFFFFFFFFFFFFFFFFFFFFAA954",
INIT_1F => X"ABFF557BFFFFFFFFFFFFFFFFFBFDFEFFFAA974BA5D517FFFF08043FFFFFFFFFF",
INIT_20 => X"6AB45AA8002000F7D5575455D043FFFFFFFFFFFFFF7FBFDF55A28402000F7D56",
INIT_21 => X"43FFFFFFFFFDFEFA2D56AB45AA8400145AA8017410007BFFFFFFFFFFFFEFF7D1",
INIT_22 => X"AA975FF00003FE00557BFFFFFFFFBFDF45AAD568B55F7AE955FFAA8402010080",
INIT_23 => X"7D168B55AAD17FFEFF7AE975FF00557FFFF5D043FFFFF7FBE8B45AAD568BFFFF",
INIT_24 => X"00000000000557FFEFA2D168B55AAFBFFFFFFF80021EF0855421EF002ABFFEFF",
INIT_25 => X"FFFFFFFFFFF7AA954BA550000082550000000000000000000000000000000000",
INIT_26 => X"C7080E3FFFFFFFFFFFFFFFFBFDFEFFFAE954AA5504154921471FFFFFFFFFFFFF",
INIT_27 => X"F45AA8000038F7DB6FBD74975FFFFFFFFFFFFEFF7FBFAFD7E3A4954BA555B7AF",
INIT_28 => X"FFFFF7FBF8FC7EBD568B55A28000000FFDF52545550A3FFFFFFFFFDFEFE3F5FA",
INIT_29 => X"955C7BE800000008043FFEFE3F1F8FD7AAD16FB6DBE8E00155BE8015410147FF",
INIT_2A => X"1EAB55B6DF6DBFFF7AA955C71C043FE10497BFDFC7E3F1FAF55A2DB6FB7DF7AE",
INIT_2B => X"5B471C71424B8FC7E3D56AB6DB6DF7AFC7EBA0955FF145B7AFC7410438FC7E3F",
INIT_2C => X"00000000000000000000000000005B78FC7AAD56FB6DBEF1FAFD7E384001EF14",
INIT_2D => X"55517FFFFFFFFFFFFFFFFFFFFEFF7AA974AA5500020005500000000000000000",
INIT_2E => X"5AA80154AA557BEAB45002ABFFFFFFFFFFFEFF7FBFDFFFF7AA974BA550415410",
INIT_2F => X"EFF7FBFDFFFAAD168B55AA80000BAF7FFFDF5500517FFFFFFFBFDFEFFFFFEAB4",
INIT_30 => X"155F78015400557BFDFEFF7FBEAB55A2D56AB55A28002000F7FFC2155552ABFF",
INIT_31 => X"8B45AAFBFFFFFFFAA95545F7840201000043DFEFA2D56AB45AAD57DFEFF7AA82",
INIT_32 => X"E8B55000428B55AAD168B55F7FFFDFEFFFAA9555555003DE00007FFDF45AAD56",
INIT_33 => X"568B55A280021EF557FD755555042AB55AAD16ABFFFFFBEAB45A280155EF557F",
INIT_34 => X"0000000000000000000000000000000000000000000007FEAB55A2D17FFEFFFD",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000040000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(19),        -- Port A data input
DOA(0)   => data_read_a_lo_256(19),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(19),        -- Port B data input
DOB(0)   => data_read_b_lo_256(19),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_20_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000003",
INIT_01 => X"A75FF80000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"14088080800008400F655001FFCFF80018FA8044000000000000011000000007",
INIT_03 => X"0000000000000000000000000000000024001660380000000000000000004FF8",
INIT_04 => X"000079800014CC02C034001600000000000000101EC0012EE0C0026E1E80F000",
INIT_05 => X"1F0FF433EFF0440C3902100002203F2EFC040388137C3E20C8EEC00284033CC0",
INIT_06 => X"00F00100002E22EB440012C809B2FFF7C8E8840155FDC0000010E40087D8787A",
INIT_07 => X"03B800000000000000008407FC800B0000000100600040000C205FF91C000F80",
INIT_08 => X"F28C0B0300020852000002101554021F00000000000000009049226020000200",
INIT_09 => X"D80000007BEFBC010002008FF7F00000000010018A81000041C401000004FFDF",
INIT_0A => X"00000ADF000000200000008000008028300100461003EAFE400000120000913F",
INIT_0B => X"0000000000000000000000000200200290000000000000000200000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000010001000000",
INIT_0D => X"00000100000010000002000080101FFB60000000000000000000000000000000",
INIT_0E => X"03007FE29FF800C00000001002040000000000000020480002E42429C0000080",
INIT_0F => X"0004D4E180010040000400000001E60040000400000001E6010003C000000000",
INIT_10 => X"000000094B1E0040000400000001E60040000400000001E60804000000400000",
INIT_11 => X"00002000000000033628000100100000004000000006170C0008001000004000",
INIT_12 => X"000000000295810000000A100020614148002000000000004307CC3CC0000804",
INIT_13 => X"5802000000000014AC000120200000000003F0D800020100000000000A4B0020",
INIT_14 => X"0020C0C00000000002E2D000001006204040000000005786C004000000000052",
INIT_15 => X"0100A0C0939BEE1810080200000E0CE0EC000010020000000000000AE8A00002",
INIT_16 => X"2008040400400C08080000000000049F6FFC0100000000000008008008000400",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0100000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0C30C30C320624C1090D0F3CF3CD038001801C10000804482A60D09008269020",
INIT_1B => X"90C86432190C86432190CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2C30C3",
INIT_1C => X"F80000432190C86432190C86432190C86432190C86432190C86432190C864321",
INIT_1D => X"AA5504020100800000000000000000000000000000000000000000000000401F",
INIT_1E => X"FFFFFFFFFFFFFFAA954BA5500020BA5D7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974",
INIT_1F => X"74AA00003FFFFFFFFFFFFFFFFFFFFFFF7AA974AA550002000007BFFFFFFFFFFF",
INIT_20 => X"FDFEFFFAE974AA5D003FE005D043FFFFFFFFFFFFFFFFFFFFEFF7AE954BA5D041",
INIT_21 => X"BFFFFFFFFFFFFFFFFFBFDFEFFFAA974BA5D517FFFF087FFFFFFFFFFFFFFFFFFF",
INIT_22 => X"8402000F7D56ABFF55003FFFFFFFFFFFFFF7FBFDFFFAA84000105D556AB55557",
INIT_23 => X"FFFFFFEFF7FBEAB55A28000010F7D16ABEF08043FFFFFFFFFFFFFF7FBFDF55A2",
INIT_24 => X"000000000007BFFFFFFFFFFFFEFF7D16AB45AA8002000F7D5575455D2EBFFFFF",
INIT_25 => X"FFFFFFFFFFFFAE974AA550400028000000000000000000000000000000000000",
INIT_26 => X"380071FFFFFFFFFFFFFFFFFFFFFFFF7AA954BA550000082557FFFFFFFFFFFFFF",
INIT_27 => X"FEFFFAE954AA55041549214043FFFFFFFFFFFFFFFFFFDFEFF7AE974BA5500050",
INIT_28 => X"FFFFFFFFFFFFFF7FBFDFFFFFAA974BA550038E285D0E3FFFFFFFFFFFFFFFFBFD",
INIT_29 => X"02028555F6FB7D5D75FFFFFFFFFFFFEFF7FBFAFD7E3A4954BA555B7AFC70871F",
INIT_2A => X"FFDFEFE3F5FAF45AA8000038F7DB6FBD7490E3FFFFFFFFFDFEFF7F1FAFC7A280",
INIT_2B => X"DF525455524BFFFFFFFBFDFC7E3F5E8B45A28402010FFDB6ABEF140A3FFFFFFF",
INIT_2C => X"00000000000000000000000000007FFFFFFF7FBF8FC7EBD568B55A28000000FF",
INIT_2D => X"557FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5504000BA0800000000000000000",
INIT_2E => X"FFFAE954BA5500174AA08517FFFFFFFFFFFFFFFFFFFFEFF7AA974AA550002000",
INIT_2F => X"FFFFFFFFFEFF7FBFDFFFF7AA974BA55041541055043FFFFFFFFFFFFFF7FBFDFE",
INIT_30 => X"4AA557BEAB4500557FFFFFFFFFDFEFF7FFFFFEFF7AE974AA550028AAA5D2ABFF",
INIT_31 => X"DFEFFFD568B55A284020BA557FFFFFF5D517FFFFFFFBFDFEFFFFFEAB45AA8015",
INIT_32 => X"EABEF5D2ABFFEFF7FBFDFFFAAD168B55AA80000BAF7FFFDF55002EBFFFFF7FBF",
INIT_33 => X"56AB55A28002000F7FFC215555043DFEFF7FBFFF55A2D16AB45AA8402000F7FB",
INIT_34 => X"0000000000000000000000000000000000000000000007BFDFEFF7FBEAB55A2D",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000007FFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(20),        -- Port A data input
DOA(0)   => data_read_a_lo_256(20),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(20),        -- Port B data input
DOB(0)   => data_read_b_lo_256(20),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_21_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"4A302428B824900A128C090A5C1800261500213C005FE812D10420054085A202",
INIT_01 => X"081FFE3440B609703B0427F801A40B8115BC4F655300340288A40D30040E4DD8",
INIT_02 => X"0109095C30C98809800000F9FFFFFFFF149FF1FCA4C0421B182E3490DF145FE4",
INIT_03 => X"084A76341244919000099486400026523C041660BA000100CC12701015007FF8",
INIT_04 => X"000079800014CC03C075161E001118653D2408041FC004AEF000816E1C11F541",
INIT_05 => X"3F0F807BFFE000240100004683103E7FFE02482553FC3C0204EFC25010143CC0",
INIT_06 => X"008808210996035A000006EC2E04FFFFC0A0000101FFE4036450E08247F87870",
INIT_07 => X"4003400812A156C002822987FC830F40134CC74D002016612DE87FFE00400804",
INIT_08 => X"F02348D2D00080C0C53400044114000000D022640B42406808790055043A8282",
INIT_09 => X"F84056387FEFBC110008420F7FF388B70A20389346FE9F26120200800008FDFF",
INIT_0A => X"4518DBFF00020004C0A6044901112A0908AA14601DE3EBFE0A812D8D5B742D3F",
INIT_0B => X"104032901CC63410ABD249C4B3007127080806FF917FC30010107688862A28C5",
INIT_0C => X"46C9146C9146C9146C9146C9146CC8A3648A3642003184822040D000D8C41807",
INIT_0D => X"201800500941044312000900D4621FFBE0008A94C822CA8919018206C9146C91",
INIT_0E => X"2029FFEADFF8050250010030165290008800440022201082401A002000C48000",
INIT_0F => X"18048A004A6C0D2820302C005A83480D1820302A009B02B101390C0CB2830816",
INIT_10 => X"1408904831400D1820302C005A83480D2820302A009B02B021A85C0941150013",
INIT_11 => X"5C08834600024D052C1051E0B92D400360520202682C19024B6164E300448510",
INIT_12 => X"6404093E22A2012418A9D1D44ADD9E0F174103820101C0B8160D5516259FA1A8",
INIT_13 => X"60D8AA288209E615100280DA0052000C5006402000206C55144104D510CC1B0D",
INIT_14 => X"0A0D50020C04023033C52009144231D902818100C90058010361AC808126C886",
INIT_15 => X"2202386454988140600C0181500A13E830011008B0374007000B4E0CD0002450",
INIT_16 => X"0080224004002000000703804008001F7FFF01B982B01258088C008CC41198A1",
INIT_17 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_18 => X"8020080200802008020080200802008020080200802008020080200802008020",
INIT_19 => X"0000000000000000000002008020080200802008020080200802008020080200",
INIT_1A => X"BEFBEFBEFBFF7FEFEFFFE79E79FFFF7CFF77FBFFEFBFF9F7E0FDF9EFEFBF0000",
INIT_1B => X"DFEFF7FBFDFEFF7FBFDFEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEF",
INIT_1C => X"F80000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"BA5D00020000800000000000000000000000000000000000000000000000401F",
INIT_1E => X"FFFFFFFFFFFFFFAE974AA550402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974",
INIT_1F => X"20BA5D7FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5D00020AA5D7FFFFFFFFFFFF",
INIT_20 => X"FFFFFF7AA974BA5D0402000557BFFFFFFFFFFFFFFFFFFFFFFFFFAA954BA55000",
INIT_21 => X"03FFFFFFFFFFFFFFFFFFFFFFF7AA974AA55000200000003FFFFFFFFFFFFFFFFF",
INIT_22 => X"AE954BA5D04174AA00003FFFFFFFFFFFFFFFFFFFFEFF7AE974BA5D00174BA000",
INIT_23 => X"FFFFFFFFFFFFFDFEFF7AE954AA5500174BA5D043FFFFFFFFFFFFFFFFFFFFEFF7",
INIT_24 => X"000000000007FFFFFFFFFFFFFFFFFFFFDFEFFFAE974AA5D003FE005D2EBFFFFF",
INIT_25 => X"FFFFFFFFFFFFAE974BA5D0000010000000000000000000000000000000000000",
INIT_26 => X"BA557FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550400028007FFFFFFFFFFFFFF",
INIT_27 => X"FFFF7AA954BA550000082557BFFFFFFFFFFFFFFFFFFFFFFFFFAA954BA5D00000",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFEFF7AA974AA5D04050005571FFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"954BA5D00154AA00043FFFFFFFFFFFFFFFFFFDFEFF7AE974BA55000503800003",
INIT_2A => X"FFFFFFFFFBFDFEFFFAE954AA550415492140E3FFFFFFFFFFFFFFFFFFDFEFF7AE",
INIT_2B => X"0038E285D2ABFFFFFFFFFFFFFFFFBFDFEFFFAA974BA5D00104925D0E3FFFFFFF",
INIT_2C => X"000000000000000000000000000071FFFFFFFFFFFFFFF7FBFDFFFFFAA974BA55",
INIT_2D => X"087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D00000100000000000000000000",
INIT_2E => X"FF7AA954BA5D00000BA5D7FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5504000BA",
INIT_2F => X"FFFFFFFFFFFFFFFFFFEFF7AA974AA550002000557BFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA5500174AA08043FFFFFFFFFFFFFFFFBFDFEFF7AE954AA5D041740055517FF",
INIT_31 => X"FFFFF7FBFDFFFFFAA974AA5D00174BA08043FFFFFFFFFFFFFF7FBFDFEFFFAE95",
INIT_32 => X"00010552ABFFFFFFFFFFFEFF7FBFDFFFF7AA974BA550415410552ABFFFFFFFFF",
INIT_33 => X"FFFFEFF7AE974AA550028AAA5D2EBFFFFFFFFFDFEFF7FBFFFFFF7AE954BA5D00",
INIT_34 => X"000000000000000000000000000000000000000000000557FFFFFFFFFDFEFF7F",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(21),        -- Port A data input
DOA(0)   => data_read_a_lo_256(21),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(21),        -- Port B data input
DOB(0)   => data_read_b_lo_256(21),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_22_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"5290F4CDE914905A14A43D33F488243E17122300F55FEB189B343A1140548380",
INIT_01 => X"A94007B259F6A975386262000C344BA9573C6FF57B18A5FB0ABFCD3C2C5F4F0C",
INIT_02 => X"877FE30EB378008D202551040030071869D0040180AC4B685F6E26FAA0810006",
INIT_03 => X"431965109E4481D6B5AAD6875AD6AB5A1815600802888808DEA83552954D3000",
INIT_04 => X"492C0020220001010E4916C884DCD607E5EC2A344103E48003D0800023D0072C",
INIT_05 => X"00107C441001100D620A06D683018001023D37E5088043620101179092540112",
INIT_06 => X"40111C2D50A46AE45281502E4A2200081ADA0E054402365774611E047020008E",
INIT_07 => X"680BD5AA4BF5C91F840C1710010344DB9A808FDFF3DE0313014A200754040180",
INIT_08 => X"0EA212D6D481ADF0CE47CA21544009007A64EBD64049D028B93D9561A48F6027",
INIT_09 => X"207246A80400015805060040080A2A0F4A82381B4000BFB65A0283800AA50020",
INIT_0A => X"4539C020E11810098D4067EFF9FF284D483E35602820110204804818CD280100",
INIT_0B => X"10081E9528963546278008AA800470370000A0004D0000002126F30C902A29C5",
INIT_0C => X"40E1540E1540E1540E1540E1540E4AA070AA07000A0000308000190168200281",
INIT_0D => X"6870A9CA0D458D131652A154D46B600085080B14009A2B2906504940E1540E15",
INIT_0E => X"448C00044000A1EC1C44140D101A54280A14050A028500A84F02842A24C594A0",
INIT_0F => X"38359E0C4E6C256690581800F1C3E82562B0581200F1C3F08145602280402080",
INIT_10 => X"100AB8581B602562B0581800F1C3E8256690581200F1C3F1238473F121000613",
INIT_11 => X"73F0E1050083750B3E4275F829547008600C030374361FA2CEE046D48122C438",
INIT_12 => X"C4CC012A66F61154C019511628756231018500C00203E1380615651607822384",
INIT_13 => X"608AA612C0096C37B00D1724801A0009C606D1221D104553096004B61BCC1128",
INIT_14 => X"12A41E0F0600035842E7601C2C4AC68A98810080AA825A890225189980254CDE",
INIT_15 => X"A89637E00D0A1080301401C390320188321C2C0B13890105800D520AF94870B0",
INIT_16 => X"88222F110111B281A54753AA004002601001918008C10912A4440B24E8B58234",
INIT_17 => X"8220882208822088220882208822088220882208822088220882208822088220",
INIT_18 => X"2008020080200802008020080200802008020080200802208822088220882208",
INIT_19 => X"1448000000001FFFFFFFFC802008020080200802008020080200802008020080",
INIT_1A => X"9E79E79E7BFF3FEFEBEEEFBEFBEFBEFDFEF7F47F8FBEF5EB7E6CFEFBEFBE8289",
INIT_1B => X"CFE7F3F9FCFE7F3F9FCFE79E79E79E79E79E79E79E79E79E79E79E79E79E79E7",
INIT_1C => X"F800003F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9F",
INIT_1D => X"BA5D04000000000000000000000000000000000000000000000000000000401F",
INIT_1E => X"FFFFFFFFFFFFFFAE974BA5D0002000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974",
INIT_1F => X"2010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA550000010007FFFFFFFFFFFF",
INIT_20 => X"FFFFFFFAE954AA5D00000AA007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA55040",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5D00020AA5D7FFFFFFFFFFFFFFFFFFF",
INIT_22 => X"AA954BA5500020BA5D7FFFFFFFFFFFFFFFFFFFFFFFFFFAA954BA5504000AA557",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFAA954BA5500000BA5D7BFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"00000000000003FFFFFFFFFFFFFFFFFFFFFFF7AA974BA5D040200055517FFFFF",
INIT_25 => X"FFFFFFFFFFFFAE974BA5D0402000080000000000000000000000000000000000",
INIT_26 => X"10087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0000010007FFFFFFFFFFFFFF",
INIT_27 => X"FFFFFAE974AA550400028007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA5500020",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFAE954AA5D00020BA087FFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"954BA5504020AA5D7BFFFFFFFFFFFFFFFFFFFFFFFFFAA954BA5D00000BA557FF",
INIT_2A => X"FFFFFFFFFFFFFFFF7AA954BA5500000825571FFFFFFFFFFFFFFFFFFFFFFFFFAA",
INIT_2B => X"040500055517FFFFFFFFFFFFFFFFFFFFFFF7AA974AA5D00070925D71FFFFFFFF",
INIT_2C => X"0000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFEFF7AA974AA5D",
INIT_2D => X"007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020000800000000000000000",
INIT_2E => X"FFFAE974AA550002000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0000010",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFAE954AA5504000BA087FFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA5D00000BA5D7BFFFFFFFFFFFFFFFFFFFFFFFFFAA954AA5D00020AA007FFFF",
INIT_31 => X"FFFFFFFFFFFEFF7AA974BA5504020BA557BFFFFFFFFFFFFFFFFFFFFFFFF7AA95",
INIT_32 => X"154105D517FFFFFFFFFFFFFFFFFFFFEFF7AA974AA55000200055517FFFFFFFFF",
INIT_33 => X"BFDFEFF7AE954AA5D041740055557FFFFFFFFFFFFFFFFFFDFEFF7AE974AA5D00",
INIT_34 => X"000000000000000000000000000000000000000000000043FFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000007FFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(22),        -- Port A data input
DOA(0)   => data_read_a_lo_256(22),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(22),        -- Port B data input
DOB(0)   => data_read_b_lo_256(22),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_23_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"EF20906D902424807BC8241BC81801B97D38AD3C0800103362A6741C80A12A02",
INIT_01 => X"001FFF8409F089003B4422000D80C80106804A7951C5B9D1C828043EA28838F9",
INIT_02 => X"073B8858218C2C50801000F9FFEFF8E72CA7F5FC2E048026496834D84721DFE0",
INIT_03 => X"2C4360101A4001001005080400401420350016E0BB222341C312000014006FF8",
INIT_04 => X"00017B810015DC03D034201E14000036486008101FC0002EE006297E1C05F561",
INIT_05 => X"BF0F817FFFE80100004044800080BEFFFC0248005FFC3C18A5FFC2444484BCC0",
INIT_06 => X"0400000409120338860900482404FFFFC000000001FFC0832050E00047F97870",
INIT_07 => X"200246801C41C3E81E872C8FFE900FC31348EFDF03BE15E22DA07FF92C204102",
INIT_08 => X"F6220280D2B025988311AB14155421006891A1089F6E200000022C140068EB90",
INIT_09 => X"F8001011FFEFBC80000000077FF184B03010004002FE000000201000000FFDFF",
INIT_0A => X"00001BFFA800808189A657EF81DD0C00079CD00837C3EBFD4201258112D4487F",
INIT_0B => X"24483890564084198AD249C433200180082A06FF907FC3081812048006000000",
INIT_0C => X"8608086080860808608086080860804304043042003184822150C000D8C41806",
INIT_0D => X"03000100200180480000095280001FFBF040C088CD20E0A21921828608086080",
INIT_0E => X"3821FFEAFFF805025E00853B92588000400020001000020A8018008002000014",
INIT_0F => X"486148484054395E27E428002A4200397E07E422002A420100382FCC30832A16",
INIT_10 => X"0C0788417000397E07E428002A4200395E27E422002A420110A51C01C0590401",
INIT_11 => X"1C01A2490040590C08120558C1759BE1C05A0400383808800DA1929F72864110",
INIT_12 => X"20000136006000215EA0A4833A32C8832050028603050014031B3950000C90A5",
INIT_13 => X"006658280009A2030108B14AC05C00112405222088B8332C140004D101800CE7",
INIT_14 => X"196B6808060201281004228996085F10020180C030880D11019CE4000026C00C",
INIT_15 => X"52A49DC7143F01C04240030720641E0A028996483A17204680410A04104A2659",
INIT_16 => X"0401000080080000000000002001201F7FFC0011C2F81A48080CA32800A01081",
INIT_17 => X"4010040100401004010040100401004010040100401004010040100401004010",
INIT_18 => X"0100401004010040100401004010040100401004010040100401004010040100",
INIT_19 => X"0000000000000000000000040100401004010040100401004010040100401004",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"F800000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"BA5D04020100000000000000000000000000000000000000000000000000401F",
INIT_1E => X"FFFFFFFFFFFFFFAE974BA5D0400000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974",
INIT_1F => X"2000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400010087FFFFFFFFFFFF",
INIT_20 => X"FFFFFFFAE974BA550002000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D000",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA550000010007FFFFFFFFFFFFFFFFFFF",
INIT_22 => X"AE974AA550402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550400000087",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFAE974AA550402000087FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5D00000AA007FFFFFFF",
INIT_25 => X"FFFFFFFFFFFFAE974BA5D0402010000000000000000000000000000000000000",
INIT_26 => X"10087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000087FFFFFFFFFFFFFF",
INIT_27 => X"FFFFFAE974BA5D0000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04000",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFAE974BA550002000007FFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974AA550400010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550002010087FF",
INIT_2A => X"FFFFFFFFFFFFFFFFFAE974AA550400028007FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_2B => X"00020BA087FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5D0402038007FFFFFFFFF",
INIT_2C => X"00000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5D",
INIT_2D => X"087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020100000000000000000000",
INIT_2E => X"FFFAE974BA5D0400000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D0000010007FFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4AA550002000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA550002010087FFFF",
INIT_31 => X"FFFFFFFFFFFFFFFAE954AA550400010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_32 => X"000AA087FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5504000BA087FFFFFFFFFFF",
INIT_33 => X"FFFFFFFFAA954AA5D00020AA007BFFFFFFFFFFFFFFFFFFFFFFFFFAA954AA5D04",
INIT_34 => X"0000000000000000000000000000000000000000000007BFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000007FFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(23),        -- Port A data input
DOA(0)   => data_read_a_lo_256(23),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(23),        -- Port B data input
DOB(0)   => data_read_b_lo_256(23),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_24_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100600007FFF000080108004000800020000840041000080808",
INIT_02 => X"172A00D000EF8210000000F9FFEFF8E7240FF1FC224087B1000639401D005FC0",
INIT_03 => X"00003A2E200811000000000400000000340016603A0000004860400014006FFF",
INIT_04 => X"000079800014CC03C034001E04010850300000101FC0002EE000006E1C00F500",
INIT_05 => X"1F0F8033FFE000000000000000003E2FFC024800137C3C0000EFC00000003CC0",
INIT_06 => X"0000000009120110020100002404FFFFC000000001FFC0000010E00007F87870",
INIT_07 => X"200102050840950002802C87FC800FCAA035400001B918600C207FF800000000",
INIT_08 => X"F6234AD280B02500063AC2840001610020408178B600C2400013649608730004",
INIT_09 => X"F80000007FEFBC00000000077FF000B00000000002FE0000000000000000FDFF",
INIT_0A => X"00001BFFA0000005501AA00000CE20000094000011C3EBFC020125811254083F",
INIT_0B => X"0040A040004000008012414433000100080806FD107FC3000000000006000000",
INIT_0C => X"0608006080060800608006080060800304003042003180822040C00090C41806",
INIT_0D => X"004800B0000000000000000000001FFBE0008080C820C0801801800608006080",
INIT_0E => X"2021FFEADFF80002080000000208800000000000000000020018000000000000",
INIT_0F => X"840009181008024A00043601100210024A00043C0110020901382CCCB28B0806",
INIT_10 => X"180040A03080024A00043601100210024A00043C01100209240C840C201D0210",
INIT_11 => X"840A604E0080820009908008341B000A8212070082002890010068320860C920",
INIT_12 => X"40600800082041205EC00044C1ACB66C37542082030281E0580001012811A40C",
INIT_13 => X"80B27A004300004103160DB3005E000618040C022000593D002180002090166B",
INIT_14 => X"2BBFF20406040084210C062000C2A2DDD00180C04504086002CD680C01000104",
INIT_15 => X"20804295C98F80400008040CC0582169022000C2876C40478002850016088001",
INIT_16 => X"0000000000000000000000000000001F7FFC001B823018F00880008805241060",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"9EF9EF9EFB263CC3090CABAEBAFF96857757B73E6089966B9EF9D5A220CC8000",
INIT_1B => X"C1E0F0783C1E0F0783C1EFBEFBEFBE79E79E79E79E79EFBEFBEFBEFBEFBEF9EF",
INIT_1C => X"F800000783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783",
INIT_1D => X"BA5D04020100800000000000000000000000000000000000000000000000401F",
INIT_1E => X"FFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974",
INIT_1F => X"0000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000087FFFFFFFFFFFF",
INIT_20 => X"FFFFFFFAE974BA5D0400000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400010087FFFFFFFFFFFFFFFFFFF",
INIT_22 => X"AE974BA5D0002000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0000010007",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFAE974BA5D0002000007FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA550002000007FFFFFFF",
INIT_25 => X"FFFFFFFFFFFFAE974BA5D0402010080000000000000000000000000000000000",
INIT_26 => X"00087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFF",
INIT_27 => X"FFFFFAE974BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000007FFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA5D0000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400010087FF",
INIT_2A => X"FFFFFFFFFFFFFFFFFAE974BA5D0000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_2B => X"0002000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA550002000087FFFFFFFFF",
INIT_2C => X"00000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA55",
INIT_2D => X"007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020100800000000000000000",
INIT_2E => X"FFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA5D0400000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000007FFFF",
INIT_31 => X"FFFFFFFFFFFFFFFAE974BA5D0000010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_32 => X"00010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0000010007FFFFFFFFFFF",
INIT_33 => X"FFFFFFFFAE974BA550002010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5500",
INIT_34 => X"0000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(24),        -- Port A data input
DOA(0)   => data_read_a_lo_256(24),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(24),        -- Port B data input
DOB(0)   => data_read_b_lo_256(24),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_25_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100200002000000080100004000000020000800041000080808",
INIT_02 => X"1000218000000800000000F9FFEFF8E738FFF1FC20400400000004455A375FE0",
INIT_03 => X"00002000000001000000000400000000340016623A0000004000000014006FFF",
INIT_04 => X"924279824C94CC1BE0B4001F20000000020380401FE0082EF000106E1C00F500",
INIT_05 => X"1F0F8033FFF048202582800100523E2FFE024820137C3C0040EFE02000003CE4",
INIT_06 => X"10DC00CC0992033A062116E82404FFFFC0E0801101FFC0000010E08A07FC7870",
INIT_07 => X"000000000000000002802C87FC800F8000000000019810600C207FFF3C410D84",
INIT_08 => X"FE8002000080281000008A0000014100200081000000000080480AE000000200",
INIT_09 => X"FC0020007FEFBE031018C31F7FFBAEBC0020008086FE0000100280800000FDFF",
INIT_0A => X"00001BFFE00301000000000000CC02000014000191C3EBFF4A7DF795965C6D3F",
INIT_0B => X"0040200000400000801243443B000100880806FD107FC3018000000006000000",
INIT_0C => X"0608006080060800608006080060800304003042003B99862444E61492C41806",
INIT_0D => X"00000000000000000000001280001FFBE0008080C820C4801801800608006080",
INIT_0E => X"3021FFEADFF805025C0304001E58906088304418222C108A009A090400000000",
INIT_0F => X"00000100100000480000200100000000480000200100000100380F0C30830A06",
INIT_10 => X"0000008000000048000020010000000048000020010000000004040000010000",
INIT_11 => X"0400004000000000008080000011000000020000000020000000001200000100",
INIT_12 => X"000000000800002018C010000020800000800122000000004004000008000004",
INIT_13 => X"0002080000000040000001020020000000000800200001040000000020000021",
INIT_14 => X"0021000008001000000800200000021000020100000000200004200000000100",
INIT_15 => X"0000008400000000605000000000200000200000020400000000000002008000",
INIT_16 => X"288226410410346010000000400A011F7FFE0031823010400800000800001840",
INIT_17 => X"8822088220882208822088220882208822088220882208822088220882208822",
INIT_18 => X"8220882208822088220882208822088220882208822088220882208822088220",
INIT_19 => X"00017FFFFFFFFFFFFFFFFE088220882208822088220882208822088220882208",
INIT_1A => X"2410492410A048029890AD34D35FDD144A50CB5462D14997BE09E760AED04040",
INIT_1B => X"8C46231188C46231188C49249249249249249249249241041041041041041049",
INIT_1C => X"F80000B158AC562B158AC562B158AC562B158AC562B158AC562B158AC562B158",
INIT_1D => X"BA5D040201000000000000000000000000000000000000000000000000007FFF",
INIT_1E => X"FFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974",
INIT_1F => X"2010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFF",
INIT_20 => X"FFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000087FFFFFFFFFFFFFFFFFFF",
INIT_22 => X"AE974BA5D0400000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000007",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFAE974BA5D0400000087FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000007FFFFFFF",
INIT_25 => X"FFFFFFFFFFFFAE974BA5D0402010000000000000000000000000000000000000",
INIT_26 => X"10087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFF",
INIT_27 => X"FFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA5D0402000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000087FF",
INIT_2A => X"FFFFFFFFFFFFFFFFFAE974BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_2B => X"0400000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000087FFFFFFFFF",
INIT_2C => X"00000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D",
INIT_2D => X"087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020100000000000000000000",
INIT_2E => X"FFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFF",
INIT_31 => X"FFFFFFFFFFFFFFFAE974BA5D0402000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_32 => X"02000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000087FFFFFFFFFFF",
INIT_33 => X"FFFFFFFFAE974BA5D0400000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_34 => X"0000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000007FFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(25),        -- Port A data input
DOA(0)   => data_read_a_lo_256(25),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(25),        -- Port B data input
DOB(0)   => data_read_b_lo_256(25),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_26_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"E9264EAB20190CA3BA4997AA9002AE9C001006B0778015CFA17E0811039879C7",
INIT_01 => X"F1FFF9BB1F773C7F9BB07DFFFDD863FC5FFF3FEFFBBF9FFB22FFFBC7B9F30686",
INIT_02 => X"1B33188302E708180F6FFBFFFFCFFFFF9C7FF7FC24350B99082400001D00DFD8",
INIT_03 => X"4A53D958C50000DCE7366303739CD98C27C57EF57980014F271807E3C9E9CFF8",
INIT_04 => X"DBFAFBD7FB1CDEBEF1BE17F7AC88042787FBFFF8FEE9FF7EE6F4C0EE1FFAF869",
INIT_05 => X"5F0FFEB3EFFEFFBDA7F7FED508707E2EFEBF6FFEB37C3FF302EEEDFF9B487CF6",
INIT_06 => X"AFBE564C71268F3BBF5FBFC2A427FFF7C3E3A74667FDDB7FB870FF30FFDEF87F",
INIT_07 => X"03BC18306396FBEC14489737FDC00B13BB79DFDB83BF4112AF205FFBDD3AFB93",
INIT_08 => X"F21E4391909B381B0B1F8E041051831FA3068D77E000030021324620C0B9C206",
INIT_09 => X"DE89ECC0FBEFBEBF30B8D79FF7F451F33CFD60FE8FFFDF58003B1D4223B4FFDF",
INIT_0A => X"8ED6BFDF3EB3EBF9DDBCE7FDC1DF8A760F3EB980580BFAFFF37DF7B9DF7DCB3F",
INIT_0B => X"6EE6F5E7FAC4C03DB856CD4CF73AC1FC98884FFF19FFC71FEFED7B251E35768E",
INIT_0C => X"06BC606BC606BC606BC606BC606BD3035E3035C62B7BB987666DEF8A90CCFA8F",
INIT_0D => X"CF6100C0E60FB9FC3A80EF69A04DFFFF7FF5F9A0DC33E9B41D01D207BC606BC6",
INIT_0E => X"7027FFFF9FF8FAFAA3ADEBFB9726BAF5FD7AFEBD7F7EFFD7ACDB7F947F0EA035",
INIT_0F => X"E020080A40403E8BD8002000FC02003E8BD8002000FC02010979AFFE36C36B86",
INIT_10 => X"000EE00034003E8BD8002000FC02003E8BD8002000FC020037B0040A00010003",
INIT_11 => X"040C00400003D80008160400FD81341C00020003B80008C00801EF0285380100",
INIT_12 => X"90981038406809677FA080468C46A81080581002000780C8001C8100201037B0",
INIT_13 => X"00F90D162001C803411FC0024080001F80040026C0807C868B1000E401A01F11",
INIT_14 => X"3F810503A00003E020042AC080CEB01228A80000F600080123E232130407080D",
INIT_15 => X"0087520750001064180807868000110C02C080CFA0042400000F8800105B0201",
INIT_16 => X"7FDFF7EFEEFF3EEC3FF7FBFFBCB7FFFFEFFE00BFF7FEBF420800EC0CBEE61F81",
INIT_17 => X"FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F",
INIT_18 => X"D7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5",
INIT_19 => X"43237FFFFFFFFFFFFFFFFF5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5F",
INIT_1A => X"A69A61861BAF15EAA6AFC38E38EA3AD8ADE7A48F0B366429F434AA9FC376DAE4",
INIT_1B => X"C26130984C26130984C261861861861861861861861861861861861861861869",
INIT_1C => X"F800000984C26130984C26130984C26130984C26130984C26130984C26130984",
INIT_1D => X"BA5D04020100000000000000000000000000000000000000000000000000401F",
INIT_1E => X"FFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974",
INIT_1F => X"2010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFF",
INIT_20 => X"FFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFF",
INIT_22 => X"AE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFF",
INIT_25 => X"FFFFFFFFFFFFAE974BA5D0402010000000000000000000000000000000000000",
INIT_26 => X"10007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFF",
INIT_27 => X"FFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FF",
INIT_2A => X"FFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_2B => X"0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFF",
INIT_2C => X"00000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D",
INIT_2D => X"007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020100000000000000000000",
INIT_2E => X"FFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFF",
INIT_31 => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_32 => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_33 => X"FFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_34 => X"0000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(26),        -- Port A data input
DOA(0)   => data_read_a_lo_256(26),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(26),        -- Port B data input
DOB(0)   => data_read_b_lo_256(26),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_27_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"00080A40000A41248002029000050A088000008242A0004404480002000A1155",
INIT_01 => X"F1FFF1C11F781C129C107DFFFE0860941E81258CA2B71C2220EC1B86E1A00002",
INIT_02 => X"4000002100000014400FF6FFFF0FFFFF8007F1FC211100014200800000887FC0",
INIT_03 => X"0842D85841000098C63061026318C18404C459757000015F00088BE3C0618FF8",
INIT_04 => X"DBEAE5D6D91C2EBCE1B21EA72C00000007FBE7C8F8E9EF79E6D440E91FDAE061",
INIT_05 => X"5C8FFCB38FF6B68984B5BCE408347E28FEBF6FEEB3723F7102E8EDBF8A4872F6",
INIT_06 => X"AB98420C71408D113956AFD0842FFFC7C3032646EFF1DB7FA868FE30EF1CE47E",
INIT_07 => X"10041830600640C415004637FC4003021259CFDB01BF80028E001FF8251AB9D1",
INIT_08 => X"F200822020842203000082050000110023068D03000002820000000840000005",
INIT_09 => X"1C852440E3DF7E2FB0B8E717C7F411F3BC6D60B60FFDDE480018AC4AA3B0FD1F",
INIT_0A => X"18109E1F16B16B71092CE7ED81CF403601229880400BE0FC137FF7A0FF75813F",
INIT_0B => X"86F7D5E382A440349816DD4C755AC16C1A884FFE18FFD757E7ED7A211E81C098",
INIT_0C => X"061A2061A2061A2061A2061A2061E1030D1030D6A37FB9872E65E6AA90CD5AAF",
INIT_0D => X"8FC10080A20ED1D41880CC61A044DFFC6EB5BCA0DE31F8B41C01E0071A2061A2",
INIT_0E => X"2023FFE91FF98AEAA1AC6AC9A3A4AAD5B56ADAB56D5AFD572C597B147506203E",
INIT_0F => X"E020000260403C8948002000EC0000BC8948002000EC00010878AC3CB8AB8857",
INIT_10 => X"000EE0000400BC8948002000EC0000BC8948002000EC000097B0040200010003",
INIT_11 => X"040400400003D80000070400DD81041400020003B80000410801AF0204180100",
INIT_12 => X"101010384008086378A080428C46A80080081002000780C800188000301017B0",
INIT_13 => X"02E909042001C800409FC0020080001F80000007C0807484821000E400205D11",
INIT_14 => X"3F810100A00003E020000BC0808EB01020280000F60000002BA2220204070801",
INIT_15 => X"0007520750000024080807868000100403C0808FA0040400000F8800001F0200",
INIT_16 => X"5B5EF3AF6AF6389C2FE128971AB2DDDF8FFE0031B776BF4208006C0C92621F81",
INIT_17 => X"B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D",
INIT_18 => X"56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5",
INIT_19 => X"43A3FFFFFFFFFFFFFFFFFD5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B",
INIT_1A => X"0000000001E0080397908000000A48710B4080240E543021B438A010825238B4",
INIT_1B => X"0804020100804020100800000000000000000000000000000000000000008200",
INIT_1C => X"F80000A05028140A05028140A05028140A05028140A05028140A05028140A050",
INIT_1D => X"BA5D04020100000000000000000000000000000000000000000000000000401F",
INIT_1E => X"FFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974",
INIT_1F => X"2010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFF",
INIT_20 => X"FFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFF",
INIT_22 => X"AE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFF",
INIT_25 => X"FFFFFFFFFFFFAE974BA5D0402010000000000000000000000000000000000000",
INIT_26 => X"10007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFF",
INIT_27 => X"FFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FF",
INIT_2A => X"FFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_2B => X"0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFF",
INIT_2C => X"00000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D",
INIT_2D => X"007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020100000000000000000000",
INIT_2E => X"FFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_31 => X"FFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_32 => X"02010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFF",
INIT_33 => X"FFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_34 => X"0000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000007FFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(27),        -- Port A data input
DOA(0)   => data_read_a_lo_256(27),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(27),        -- Port B data input
DOB(0)   => data_read_b_lo_256(27),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_28_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"02200AA400180030808802A900002A08001280A08A801044104A1000001818C3",
INIT_01 => X"50A00011460214428114180000882214413D0A71592A01D92213D28005210202",
INIT_02 => X"1444428102100884000AA30200000000C1000401041108404400022220800000",
INIT_03 => X"461080404900000C6314A900318C52A40051081000888806108802A141288001",
INIT_04 => X"00800040110102000902002000888400081045A8A00003C00000500000080008",
INIT_05 => X"0000000000024CA0A0101800032000400000000B800000014000000B08180000",
INIT_06 => X"814016012000C405280200008001000011110012220009A88800009A88000000",
INIT_07 => X"0004891224228810080010200040001020800000004000008200000240081400",
INIT_08 => X"00A010040401080308400821155540001122448142491008A004912040840221",
INIT_09 => X"0020405000000124058200408000880004440004080160C8100A858009940000",
INIT_0A => X"4D29400002002038104000000020003204000880082800010000000C0000E400",
INIT_0B => X"12220122A000416811040000400800081022C0000080000206CB0821082B694D",
INIT_0C => X"80B0280B0280B0280B0280B0280B01405814058009000421833010800A000200",
INIT_0D => X"C4210040860B188C0A8065302005A004039010280001001600200081B0280B02",
INIT_0E => X"500600010000280000802050010660001000080004004900204020105302A000",
INIT_0F => X"0000000A00000081480000001400000081480000001400000800C01082082210",
INIT_10 => X"0000000024000081480000001400000081480000001400000010000200000000",
INIT_11 => X"0004000000000000001400000080041400000000000000C00000010004180000",
INIT_12 => X"1010100000480802A40000000400000080081000000000000004800000000010",
INIT_13 => X"0001010420000002400040000080000000000024400000808210000001200010",
INIT_14 => X"04000100A0000000000028400004000020280000000000012002020204000009",
INIT_15 => X"0001000000000024080000000000010400400004000004000000000000510000",
INIT_16 => X"0108408420430E699AA42A1508104EA08000000810020000000044001AC20500",
INIT_17 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_18 => X"0040100401004010040100401004010040100401004010040100401004010040",
INIT_19 => X"1708000000000000000000010040100401004010040100401004010040100401",
INIT_1A => X"20820820800D41A8283AC618618EF1088160885001234B96061CCDEC4D205061",
INIT_1B => X"0C06030180C06030180C08208208208208208208208208208208208208208208",
INIT_1C => X"F80000B0582C160B0582C160B0582C160B0582C160B0582C160B0582C160B058",
INIT_1D => X"BA5D04020100000000000000000000000000000000000000000000000000401F",
INIT_1E => X"FFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974",
INIT_1F => X"2010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFF",
INIT_20 => X"FFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFF",
INIT_22 => X"AE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFF",
INIT_25 => X"FFFFFFFFFFFFAE974BA5D0402010000000000000000000000000000000000000",
INIT_26 => X"10007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFF",
INIT_27 => X"FFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FF",
INIT_2A => X"FFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_2B => X"0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFF",
INIT_2C => X"00000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D",
INIT_2D => X"007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020100000000000000000000",
INIT_2E => X"FFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_31 => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_32 => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_33 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_34 => X"0000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000007FFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(28),        -- Port A data input
DOA(0)   => data_read_a_lo_256(28),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(28),        -- Port B data input
DOB(0)   => data_read_b_lo_256(28),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_29_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"79964E4BA01DACAB9E659792D00AAE160002829C7FDFEFCEE97C2815039D70C3",
INIT_01 => X"50BFF9AB0775343F9AB01DF80D5821FC0FFF3FEFD1AF9FF1207FFBC7B9720586",
INIT_02 => X"0B33180300E700080F6AAA7BFFC007189C7FF2FC003503980A0000001D00DFD8",
INIT_03 => X"0401D940CD0000C8421A2B03210868AC23403E903900010E271006A148A0C000",
INIT_04 => X"49B87A417315D20A313E17F1800000058013DDF8BE21F36E02F0D06E03E8F800",
INIT_05 => X"1F007E33E01A4D9C87525E5101603E6E023D27DA937C03E340EE25CB9B483C12",
INIT_06 => X"85AA06002026872BAE0B1282A005FFF001E1870223FC3BFC98101F109FC6780F",
INIT_07 => X"03BC081023B233E804488527FDC008019968D74982C94110AF204001BC285A82",
INIT_08 => X"001E4191901A101B031F84000000831FA1028575A000110800124600C039C002",
INIT_09 => X"C60888D0782082B50080508FF00048B124D4005C8AFF4158102914800110FFC0",
INIT_0A => X"8AD6ABC02A02A0B0CCB463B4C0748A720B1EA980100BFA02E204D2154D28AA3F",
INIT_0B => X"6A22B126DA40C03531440800C22800B8900042FF0180000ABFEF89250815568A",
INIT_0C => X"803468034680346803468034680353401A340180010A0801422829800A00A001",
INIT_0D => X"87410080C60AB0F42A804628200DBFFF13D05928040329160520528134680346",
INIT_0E => X"2006FFFF8000F8F80281A16A1504302058102C0816244B82A0CA25907D0AA015",
INIT_0F => X"0000080A40000283D80000001402000283D80000001402010901A7D694494192",
INIT_10 => X"0000000034000283D80000001402000283D80000001402002010000A00000000",
INIT_11 => X"000C000000000000081600002080341C00000000000008C00000410085380000",
INIT_12 => X"90981000006809076B2000040400001080581000000000000004810020002010",
INIT_13 => X"0011051620000003410040004080000000040026C00008828B10000001A00210",
INIT_14 => X"04000503A000000000042AC00044000228A8000000000801204212130400000D",
INIT_15 => X"0081000000001064180000000000010C02C000440000240000000000105B0001",
INIT_16 => X"258964C4A44A0C689FF3F9FFEC5D6DBFE0020096528A0B000000CC043EC60780",
INIT_17 => X"5816058160581605816058160581605816058160581605816058160581605816",
INIT_18 => X"8160581605816058160581605816058160581605816058160581605816058160",
INIT_19 => X"03017FFFFFFFFFFFFFFFFE058160581605816058160581605816058160581605",
INIT_1A => X"AEBAEBAEBFFF7FEFCFDF7FFFFFF5DE7CFCB773FFEFBFF3C7E1E779FFEFFF5060",
INIT_1B => X"FEFF7FBFDFEFF7FBFDFEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEEBAEB",
INIT_1C => X"F80000FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFD",
INIT_1D => X"BA5D04020100000000000000000000000000000000000000000000000000401F",
INIT_1E => X"FFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974",
INIT_1F => X"2010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFF",
INIT_20 => X"FFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFF",
INIT_22 => X"AE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFF",
INIT_25 => X"FFFFFFFFFFFFAE974BA5D0402010000000000000000000000000000000000000",
INIT_26 => X"10007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFF",
INIT_27 => X"FFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FF",
INIT_2A => X"FFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_2B => X"0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFF",
INIT_2C => X"00000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D",
INIT_2D => X"007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020100000000000000000000",
INIT_2E => X"FFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_31 => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_32 => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_33 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_34 => X"0000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(29),        -- Port A data input
DOA(0)   => data_read_a_lo_256(29),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(29),        -- Port B data input
DOB(0)   => data_read_b_lo_256(29),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_30_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"9E79E79E7BAF7DEBAFAFEFBEFBFFBFFDFFF7FCFF0FBFFDFF7EFDDFFFEFFE8000",
INIT_1B => X"CFE7F3F9FCFE7F3F9FCFE79E79E79E79E79E79E79E79E79E79E79E79E79E79E7",
INIT_1C => X"F800003F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9F",
INIT_1D => X"BA5D04020100000000000000000000000000000000000000000000000000401F",
INIT_1E => X"FFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974",
INIT_1F => X"2010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFF",
INIT_20 => X"FFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFF",
INIT_22 => X"AE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFF",
INIT_25 => X"FFFFFFFFFFFFAE974BA5D0402010000000000000000000000000000000000000",
INIT_26 => X"10007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFF",
INIT_27 => X"FFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FF",
INIT_2A => X"FFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_2B => X"0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFF",
INIT_2C => X"00000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D",
INIT_2D => X"007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020100000000000000000000",
INIT_2E => X"FFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_31 => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_32 => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_33 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_34 => X"0000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(30),        -- Port A data input
DOA(0)   => data_read_a_lo_256(30),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(30),        -- Port B data input
DOB(0)   => data_read_b_lo_256(30),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_31_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"129000008004A00804A40000400800020000000C005FEA005800200400050100",
INIT_01 => X"A15FF18019700810180065FFFC0040801E80258CA2951C2200EC0906A0804140",
INIT_02 => X"0000000000000011000550FDFF0FFFFF0007F1FC200000011000000000205FC0",
INIT_03 => X"08425818000000908428C0024210A30004045060302223490002014280410FF8",
INIT_04 => X"DB6A618248140C18E0B016872400000007EBA24058E1ECA8E2D400681FD0E061",
INIT_05 => X"1C0FFC338FF01009048084C400103E28FE3F6FE513703F7000E8E5B4825030F6",
INIT_06 => X"0098000C51000910100006C00426FFC7C202060445F1F2572060FE82671C607E",
INIT_07 => X"40001020400440C41C000617FC0003021259CFDB01BF00020C001FF804000980",
INIT_08 => X"F200020000802000000082044000010022048902000002000000000000000004",
INIT_09 => X"1C002400E3CF3E0B1118C31747F000B33820209206FC9E80000000000220FD1F",
INIT_0A => X"00001A1F00110101092CE7ED81CF0004012290000023E0FC027DF780DF74013F",
INIT_0B => X"044094C1028400548812494C31004124080886FE187FC301B124F20016000000",
INIT_0C => X"0608006080060800608006080060C00304003042023B99862444E60090C41887",
INIT_0D => X"0B400080200481501000884080405FF864008880CC30E8A01C01C00608006080",
INIT_0E => X"2021FFE81FF880EA000400098200C04080204010200810020C18090424040034",
INIT_0F => X"E020000040403C0800002000E800003C0800002000E8000100780C2C30830806",
INIT_10 => X"000EE00000003C0800002000E800003C0800002000E8000017A0040000010003",
INIT_11 => X"040000400003D80000020400DD01000000020003B80000000801AE0200000100",
INIT_12 => X"000000384000006118A080428846A80000000002000780C800180000201017A0",
INIT_13 => X"00E808000001C800001F80020000001F8000000280807404000000E400001D01",
INIT_14 => X"3B810000000003E020000280808AB01000000000F600000003A0200000070800",
INIT_15 => X"000652075000000000080786800010000280808BA0040000000F8800000A0200",
INIT_16 => X"080223010010308025410082404A015F0FFE003182701B420800280C80201A81",
INIT_17 => X"8020080200802008020080200802008020080200802008020080200802008020",
INIT_18 => X"0200802008020080200802008020080200802008020080200802008020080200",
INIT_19 => X"04017FFFFFFFFFFFFFFFFC080200802008020080200802008020080200802008",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000080",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"F800000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"BA5D04020100000000000000000000000000000000000000000000000000401F",
INIT_1E => X"FFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974",
INIT_1F => X"2010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFF",
INIT_20 => X"FFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFF",
INIT_22 => X"AE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFF",
INIT_25 => X"FFFFFFFFFFFFAE974BA5D0402010000000000000000000000000000000000000",
INIT_26 => X"10007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFF",
INIT_27 => X"FFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FF",
INIT_2A => X"FFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_2B => X"0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFF",
INIT_2C => X"00000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D",
INIT_2D => X"007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020100000000000000000000",
INIT_2E => X"FFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_31 => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_32 => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_33 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_34 => X"0000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(31),        -- Port A data input
DOA(0)   => data_read_a_lo_256(31),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(31),        -- Port B data input
DOB(0)   => data_read_b_lo_256(31),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_0_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"ED39BA795990D275FB4A6E96ACC4731DEA4598B0AFB54867F6EE4618C3749803",
INIT_01 => X"58A0047D8607944AC7DA180001ECA2544042106208408208C20022E9173734B3",
INIT_02 => X"9F775E7CB273E6CCA7DAAF00001000000478020113C9C38E09FB7CCCDD9F203E",
INIT_03 => X"441406267B4CB04443163C91110C58F24A31000B8028A810A3D0F8B169A01006",
INIT_04 => X"0005802424830120024121209088809DF81454ACA01E03501D0A3B91E00F0A00",
INIT_05 => X"E0F001CC00012034C20B0232838F80D001C0100AEC83C008EF101A034C8CC300",
INIT_06 => X"582541A028D584E40CB0583CCA0100000161F84322000DA8C40F003C80030780",
INIT_07 => X"2BF70E1C3BBBB1138AF7F888025340C0888430047040FEE182CA00044BC5827C",
INIT_08 => X"0CAFC1F1F07F0FE1C94F65B11555EAFFC1C306758B24197ABCDA467F2C9CF9B3",
INIT_09 => X"027BDA3B0000011420A61080800B6E4C464258094101606E5A47A2A2098B0200",
INIT_0A => X"40198000D1281220444210123820B43B40804CE9AFC800017D82082E2081B6C0",
INIT_0B => X"CA2E0B32B01A752B078412A24844B01302A26900C4801854069B0C888890A081",
INIT_0C => X"C0F33C0F73C0F33C0F73C0F33C0E39E0319E0710A9402011C22908B56A21A020",
INIT_0D => X"8429A95E954868AD0E52273F542580000808061C0389161F027039C1F33C0F73",
INIT_0E => X"5C94001120055704FC4A1624485E2489024481224091282C4300942A19439481",
INIT_0F => X"1C55D65C3E3F01F52FFC1E0013C1F801F52FFC1E0013C1F8090423D38A18E3B1",
INIT_10 => X"1C0118796BE001F567FC1E0013C1F801F567FC1E0013C1F9085DFBF7E15C0610",
INIT_11 => X"FBF7E30F00C0270F3751F1FD00FECBF7E25C0700463E17B2C7F811FD7ADECC38",
INIT_12 => X"6474190626D6491063597F9177B956EF378D33E4030061341F077C571F8F885D",
INIT_13 => X"E207F328E3082636B2807FFD80FE00007E03F7207D3E03F9167184131B5C40FE",
INIT_14 => X"047EFA0CAE06101C53E3647D3F144FCDD22B81C0098E57D9081FCE8C8520C4DA",
INIT_15 => X"FF31ADF08DBF81846A540049707E0FE3307D3F141FFB45478040570EED41F4FE",
INIT_16 => X"902C189601208A1502B4AA5584B4068000019A80098120BCA4C617635C938574",
INIT_17 => X"0240902409024090240902409024090240902409024090240902409024090240",
INIT_18 => X"2409024090240902409024090240902409024090240902409024090240902409",
INIT_19 => X"424A800000000000000000902409024090240902409024090240902409024090",
INIT_1A => X"08208208208831042720EE38E38AAF9C4C704DAB63A6D58B3C10BAE8E789AA09",
INIT_1B => X"0F87C3E1F0F87C3E1F0F82082082082082082082082082082082082082082082",
INIT_1C => X"F800003E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F",
INIT_1D => X"55557BD75EF5D00000000000000000000000000000000000000000000018401F",
INIT_1E => X"FEFA28428B455D0017410A28428AAAA2FBD54BAF7FFD55EF007FD75EFFFAE975",
INIT_1F => X"0145F7AEBFFFF08002AA10A2AABFEAAA2FFC0000AA843FE00AAFBE8B45AA803D",
INIT_20 => X"974AA5D7BFFE000804000BAAAAAAAB45557FFFEBAA2D5401450051401555D7FC",
INIT_21 => X"FD7410557FC21555D51574AAA2FFE8B455D7BD755555517FFEFA280021FF082E",
INIT_22 => X"AEBFE00A2803FEBA002A820AA0800174BA5D2EA8B45005168A10AA8028A10087",
INIT_23 => X"7FFE8B45FFFBC00005D003FF45557FC01FFFFAE95410AA80000005D003FEAAFF",
INIT_24 => X"00000000000557DF5500003DFEFFF84175EFA2AEA8A10000417410A2FFE8BEFF",
INIT_25 => X"F0075D75EFEBAE9554540754717F1F8000000000000000000000000000000000",
INIT_26 => X"47E00A2DB45AA8A3AFD7B68E2AB78550E12555F524AFE38B780154BAFFF1D54A",
INIT_27 => X"1D500002A150038038E285D7F78FD7000B6AB50B6AABDE12BEA0AF010B7D1F8F",
INIT_28 => X"D5C7AA854008700249243A412EBFF5542A43FE9257F1E816D557095EAAA2D140",
INIT_29 => X"EDBC0B680900AAF52B474385D75C502D157545A87AAD178A8002D1D21C5E8257",
INIT_2A => X"F6A150012A2F02AFFDF40E85F475451D502D152A82000E3A5D2150AB8F401471",
INIT_2B => X"51EAFEDB52E3F1EFFFF485A2DA3D5D24BD417FD7E9541242FE920AD082E10A28",
INIT_2C => X"00000000000000000000000000005AAF555080550E87B7A405B52AAD152BD001",
INIT_2D => X"FA69574BAF7D5555AF0D79D55FFA2AC97445057F405458500000000000000000",
INIT_2E => X"0FF16565B2FA9075F4F7B3EBDF50FEAEAAB55F7AEAABFF5D2A81151FB8635A02",
INIT_2F => X"4D5D51F5E08A394003A908B8410E707EF34A08D46F6ABE7082AAAAF2FAC77FE0",
INIT_30 => X"FAE8C798A11A0EAEF75F7AA84001A7052C95256803CE3AEB038662E5D8140601",
INIT_31 => X"A05051023F9A9D57B63BFBF906CB45FABC0954AF0151555AF58794040077D774",
INIT_32 => X"FEE5555BE48AB2A2AE0A0F20C43EAC562245B4E1870108B11020AD4AA05542A0",
INIT_33 => X"D407A97F6F35F498B96BEB12DAAB77558ABD5F5F0DA6BC9525688C1A2A0C06E9",
INIT_34 => X"8000000FF8000000FF8000000FF8000000FF8000000FF80F55E25C00A0BA7FBE",
INIT_35 => X"F8000000FF8000000FF8000000FF8000000FF8000000FF8000000FF8000000FF",
INIT_36 => X"000000000000000000000000000000000000000000000000000000000000000F",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000008000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(0),        -- Port A data input
DOA(0)   => data_read_a_hi_256(0),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(0),        -- Port B data input
DOB(0)   => data_read_b_hi_256(0),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_1_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"212C001411984004084D000508C53810A03D1450E839B003342114428A000807",
INIT_01 => X"08000010400A0008010600000084004000400002000000000000000000140000",
INIT_02 => X"484DEBA0111800C004400D000000000028800001CC404E6008B4933336880010",
INIT_03 => X"650C00000848A0423183089008C604224200000100A200002C280810098C0001",
INIT_04 => X"00000004208B00200E010800006667BE7000102C00080000040012010000080C",
INIT_05 => X"0080000000002020600100208D04414000800000000200004800080000800200",
INIT_06 => X"0820196100006044401008100208000008082010000000800488000000020400",
INIT_07 => X"1210C18306788C00894098000011000820001000104050004108000001008250",
INIT_08 => X"00A48903121780004C6000311555521F183060AC564BF818B5EDFDE004460030",
INIT_09 => X"02AD881200100140A0223480000458400000480840002002184581A020000200",
INIT_0A => X"140040001020020410000010082080010400002001041001B102002E20013600",
INIT_0B => X"0895400004201001010884000000901100800800000004140002008280A8A815",
INIT_0C => X"C8D00C8D00C8D40C8D40C8D00C8D20642A06468400000030480808020F08E008",
INIT_0D => X"20BC417C16004C0B83822109040180000801000910000003203220C8C40C8D40",
INIT_0E => X"5C96000000010200200802100022008100408020401020040100142200E0E08A",
INIT_0F => X"0000021E300B000000781E00140018000000781E00140018000002430E30E061",
INIT_10 => X"1C00000024E0000000781E00140018000000781E0014001908400005E11C0610",
INIT_11 => X"0003C30F00C000000155800D00000003E21C0700000000F00118000000468C38",
INIT_12 => X"60640900004A400081401A0000004041218503E4030060000004804318008840",
INIT_13 => X"A0001208C30800025200003D807E000000000725201600090461840001340002",
INIT_14 => X"0000F00C0E06100000012D2005100409520381C00000005920004C0C81200009",
INIT_15 => X"25000120850B8180625400400000010711200510004B41478040000005548016",
INIT_16 => X"10040002002080040000804000A0000000011A000100208C008611430A000040",
INIT_17 => X"0040100401004010040100401004010040100401004010040100401004010040",
INIT_18 => X"0401004010040100401004010040100401004010040100401004010040100401",
INIT_19 => X"5000800000000000000000100401004010040100401004010040100401004010",
INIT_1A => X"8A28A28A2AC8090C69606492492C09945235D5F7E2A5040B80E1C863A2958000",
INIT_1B => X"5BADD6EB75BADD6EB75BAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA28A2",
INIT_1C => X"FC00002E974BA5D2E974BA5D2E974BA5D2E974BA5D2E974BA5D2E974BA5D2E97",
INIT_1D => X"BA55556AAAAAA800000000000000000000000000000000000000000000607FFF",
INIT_1E => X"F45A2FBD75EFA2AE97555F7FBFFF45FFAE80010AAAABFFFFFF803FE10F7D17FE",
INIT_1F => X"8AAAF7FBD54AA002A955555D7FE8ABA082EBFEBAFFD555400557BD54BA5D7FFD",
INIT_20 => X"17555AA8028BEFAAAE97555082A80000AA802ABEFA2D568A005D5157400AA802",
INIT_21 => X"EBDFEF5D7FEAA00AAAABFEAA007BC0145FFFFFDF55AAFBC00105555400105504",
INIT_22 => X"D5575555D7FC2155F7AEA8BEFAAAA954BA557BD7410550428ABA5D5168ABA552",
INIT_23 => X"FD57DF45F7D568ABAF7AABFFFF082ABFFFFFFFFEAB55557FFFEBAAAD568B45A2",
INIT_24 => X"000000000002EBFFEFA280021FF082E974AA5D7BD74000804154BA082ABFF55F",
INIT_25 => X"7F78A3FE28E3D17DEAA485FE8E02B50000000000000000000000000000000000",
INIT_26 => X"6D5D75D54BA5D7BFFF7DA2FFD55EFAAA495545E175EFF57BF8FC2000BEA4BAE9",
INIT_27 => X"A28550E10405F7A4AFE38EAA0924921C2FD55455571E8A2A087BF8EAAEB8E001",
INIT_28 => X"7A28415A001684104155C5B6DF6DBEFBFAA07157428145A00AA8A2FBD7B6DF6A",
INIT_29 => X"AAABF1FFBC7010FF8A38FEF557FEAB78B6AAB8E971471C7010B7D168F47400A0",
INIT_2A => X"495EAAA2D16D1FDBED56A55557A43DE385FD4BFBD7B6A0BF492415FC20105D24",
INIT_2B => X"F5D717FE2AAAA56DEBD17FE3DF7FB7FEBFE38017EBA4A8EB8F6FFD5FE8B7D557",
INIT_2C => X"00000000000000000000000000002A3D5C7AA854008700249243A417FFF41542",
INIT_2D => X"AF2A00010F78028B15F7823FEAAA2D57DFBA007DFCA127B80000000000000000",
INIT_2E => X"A0869AAAB8A7C19C55550E8574BA557BFFFEFAAFBD55FFAA8416545A6FB60F47",
INIT_2F => X"10A2AEBFF55F7BAAA8565DBAC1112FFAC21A022A38C20B2552E975F758516AAA",
INIT_30 => X"01E7AD1FFF5575841DE08007FC2048002895755FFEFBCEE5FBAACB10085EE5DE",
INIT_31 => X"D4000D7FC00FC5D062BBA05ED5034472A02EABEA097BEAAFAF2863FA00DD5742",
INIT_32 => X"62B0A2F7AE8B5D5D51F5E18ABD5EAFFF2AF9554FF57EFBFA18D4FBFFF40FF809",
INIT_33 => X"C95256807DC31AA8114DE55F5BED201FFFED17DFBFF6963FCAAA2283CF140500",
INIT_34 => X"0000000000000000000000000000000000000000000002CB75F7AA84001A7052",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000008000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(1),        -- Port A data input
DOA(0)   => data_read_a_hi_256(1),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(1),        -- Port B data input
DOB(0)   => data_read_b_hi_256(1),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_2_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10E44660018259B2843913100062C98004802322D3E030235201006009B2816",
INIT_01 => X"8005A188084900481C8024A542400340404000720885800802000906E4910204",
INIT_02 => X"5C010802020408040C640850AA055254090541A111240A104A0000000908B510",
INIT_03 => X"0C1101108800004481060A001204102803156020218808002440850008C80550",
INIT_04 => X"8840C08122050400582812C21C0804040968987810688899444090C10A124A69",
INIT_05 => X"4885109105400129210040010340086856B141212252142242A068A080106372",
INIT_06 => X"047450004062400090000202000054C28012204400908281302852A6710AA420",
INIT_07 => X"121810000230089008408402A800011012D41D518044411005000AA8A5004390",
INIT_08 => X"A214110514163218085008010141421F02000124000010880000442080810201",
INIT_09 => X"0A09E89041451581B53A739C42A0C9223000004881708D80100331CA8A848E0A",
INIT_0A => X"1009020A30020008096A06B8C1208A000A9C20004820B0573165541CD5482216",
INIT_0B => X"ACC084404A8000490152D100344001108AA88B1D007291402802B1041632A011",
INIT_0C => X"8696086860869608686086920868004309043414A2191C24485C4D2A9A0DF823",
INIT_0D => X"484000804201C1102080215900038AD030014588D200F0221821808682086820",
INIT_0E => X"00002AA00AA80240A001010026824040C000201030000200C8980080260C201E",
INIT_0F => X"0000000A20001602900020001400002A029000200014000100280E6694490312",
INIT_10 => X"0000000024002A02900020001400001602900020001400002700000800010000",
INIT_11 => X"0008004000000000001500006C00300800020000000000C100014A0081200100",
INIT_12 => X"8088000000480005188000440840081000500002000000000004800010003420",
INIT_13 => X"0070041200000002411280004000000000000026000038020900000001201300",
INIT_14 => X"2A0004030000000000002A00004A100208800000000000012260101100000009",
INIT_15 => X"0084420300001040100000000000010402000049800020000000000000580001",
INIT_16 => X"040111000008001505448340606B21090556002E00000000000080002A040A00",
INIT_17 => X"401004010040300C0300C0300C0100401004010040300C0300C0300C01004010",
INIT_18 => X"0200400004000040000C0200C0200C0200400004000040300C0300C0300C0100",
INIT_19 => X"14A97C0FC0FC1F81F81F800C0200C0200C0200400004000040000C0200C0200C",
INIT_1A => X"0410410411823A4301040B2CB2CBACB002009C6B860185AA1491B0E2863EA015",
INIT_1B => X"8944A25128944A25128941041041041041041041041041041041041041041041",
INIT_1C => X"FC703F25128944A25128944A25128944A25128944A25128944A25128944A2512",
INIT_1D => X"AA0004001550000000000000000000000000000000000000000000000078401F",
INIT_1E => X"5FF5D003FE10F7D17FEBAF7D5420AA0855420AAAA843DFFFAAD1554005D7FD74",
INIT_1F => X"FF45AAFBC20AAF7D1575EF55517DF555D2EBFF45AAAAA8A10A2AE80010A2AA97",
INIT_20 => X"AABEFAAD1575EFAAAE974AA5D51554BA5D7FFFF45A2AA975EFA2FFD7555FFFBF",
INIT_21 => X"5554AA555555555557FE8ABA082EBFFFFAAAE95555552E974105D517DF55AAAA",
INIT_22 => X"D540000AA802AABAF7FFC2010AAAE821EF552E82010F7AABFE10FFD542145FFD",
INIT_23 => X"02E800AA08042AB45007FC00BAFFD168BEFF7FBC0010AA802ABEFAAD540000FF",
INIT_24 => X"000000000002E80010555540010550417555AA8028BEFAAAE821550851420AA0",
INIT_25 => X"7A2DF55400557FD54AA1D04001C5150000000000000000000000000000000000",
INIT_26 => X"D5F7A482000BEAE905C755003FE28E3D17DEAAE95F40002157F470AABE803AE9",
INIT_27 => X"5EFAAA495545E3F5EFF57F7FE80082FFDE105EF55517DFC5552ABDF45B6AEAFF",
INIT_28 => X"24105D5B7FF7DB6AAAABC7BEDB505EFBEA4070BA5FD0154BA5D7BFAF7DA2AE95",
INIT_29 => X"38E00B6DF68FEF4871D24BA495B5556D5571E8AAF082AB8EAAEB8E0016D5D2A9",
INIT_2A => X"E2FBD7B6DF47A00EBDB50000A380AAE28E80495038AAAEAF1D7410E80000FF84",
INIT_2B => X"FBC703AE2DF42AAA002A851C214003FF680071ED1EFEAF1EFFFDEAD1C5010AA8",
INIT_2C => X"00000000000000000000000000002087A28415A001684104155C5B68E2DBEFBF",
INIT_2D => X"51FBD74BAF7802AB05AAFBD5400557BD54AA5500021555100000000000000000",
INIT_2E => X"55D2ABDF55F782BEB47AFAD00010F7AA8215555003FEAAAAD57DEBAA2FDDC010",
INIT_2F => X"BA557BEABEFAAEBD55FFAA1456547A2D360F47AF7FC20B2F7FBC015D58517FF5",
INIT_30 => X"AB4A78016545540400010557BFDFFFF7822A955FFFFC20FFF3AE544108410174",
INIT_31 => X"D545002A800A8FF862BA00F2F9E8F0050D4420BA547FD75FF58516AAAA0828AA",
INIT_32 => X"35B57AB5155400A2AEBFF45FFFB404007FFBD550AAFACAAA122AA8954BAA2AE9",
INIT_33 => X"895755FFAEBCFE57BBA57002DF3C4AAAA002E954505C417FFFF08555555BAAD3",
INIT_34 => X"000000000000000000000000000000000000000000000061DE08007FC2048002",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000010000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(2),        -- Port A data input
DOA(0)   => data_read_a_hi_256(2),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(2),        -- Port B data input
DOB(0)   => data_read_b_hi_256(2),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_3_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"210C44A20020248B08431120001604B8156023104C40771B3430400A02380206",
INIT_01 => X"014C9A4250B0296D3C2422C992100B49404040028804A0080A000416A8D90A0C",
INIT_02 => X"4809A900031800444460589C66E331352180D468B8040E600C0081110B802CD0",
INIT_03 => X"6D0B6110880001D23583480648D60520330066810A80881068A808029CC56330",
INIT_04 => X"48221A066A09D03B348C1C1928DD5A4402A13868070940842640902107002D24",
INIT_05 => X"058318035328202004C1C4E50B44644B30A86D01014A0D224063090082100E34",
INIT_06 => X"08381A010040200AC2190ED2002ACD99881822104C5A40942048288234629414",
INIT_07 => X"0218408142740E2C0948C3066400071913209CC8004640100D003999552083D2",
INIT_08 => X"900409231292A8080C2000110001521F0810A92E7402F08AB0016CA000C60011",
INIT_09 => X"620C889014D30E4A210214D5099058808010605A81A41480102130C020A43A39",
INIT_0A => X"512850E61822020C899046740121820004102000402079CCA037A02C68552A35",
INIT_0B => X"8895000026A00141015290040460C0B4828289AC1011954C0026A20400882914",
INIT_0C => X"80CA080DA080DA080CA080CE080DB0402F040654A2442834C0092E228A0DF2AB",
INIT_0D => X"289080600E04C50206808059000999C98840C508D220108200202080DA080CA0",
INIT_0E => X"300E6660599802602209021204A050E1C850C428521C208480821D842085A03E",
INIT_0F => X"0000010000003202900000010000000A02900000010000008038666920920A24",
INIT_10 => X"0000008000002202900000010000001E02900000010000002380000800000000",
INIT_11 => X"0008000000000000008000002D00300800000000000020010001620081200000",
INIT_12 => X"8088000008001021C88000048800281000500000000000004000000000003600",
INIT_13 => X"00B8041200000040011980004000000000000803000068020900000020001B00",
INIT_14 => X"29800403000000000008030000C83002088000000000002002E0101100000100",
INIT_15 => X"00841003100010401000000000002000030000C38000200000000000020C0001",
INIT_16 => X"108722420420A0100006D34A404800185CCE0128410820000008008021C40A00",
INIT_17 => X"0872108721085218852188521885218852188521887210872108721087210872",
INIT_18 => X"8721086214872108621C852188421C852188421C852188721087210872108721",
INIT_19 => X"54A2EAA555AAB554AAB5561C852188421C852188421C85218842148721086214",
INIT_1A => X"0410410412881D0B0000092492480A981E063C638321450A08899A62C314A014",
INIT_1B => X"9D4EA753A9D4EA753A9D49249249249249249249249249249249249249241041",
INIT_1C => X"FAABC4351A8D46A351A8D46A351A8D46A351A8D46A351A8D46A351A8D46A351A",
INIT_1D => X"5500002AA100000000000000000000000000000000000000000000000000401F",
INIT_1E => X"FFFAAD1554005D7FD74AAA284001550055421EFAAFFD54AAF7D168B45AAAABDF",
INIT_1F => X"20AA080400155AAD5554AAF7802AB4500043DF45FFD168AAA0855420AAAA843D",
INIT_20 => X"021550855555FFAA84001FFAAAE80010A2AA955FF5D003FE10F7803FEBAFFD54",
INIT_21 => X"BC20AAA284175EF55517DF555D2EBFE00AA8028B45A2AE82155A2FBFFEBA0800",
INIT_22 => X"7BD7555FFFBFDF55AAFBD55EF5D2EBFE10085168ABAFFFBD54BAAAAE97400A2F",
INIT_23 => X"D0015410F7AAAAAAA55043DE00FFFFD5555AAAA954AA5D7FFFF45AAAA975EF00",
INIT_24 => X"0000000000004174105D517DF55AAAAAABEFAAD1575EFAAAE974AA5D00175555",
INIT_25 => X"2EBD56DB7DBEAEBFF551C042AA101D0000000000000000000000000000000000",
INIT_26 => X"D75D5B470AABE8A3AFD7A2DF55400557FD54AABC04001C51551471D7AAF1D05D",
INIT_27 => X"E28E3D17DEAAEBDF40002550F47155AADB50492EB842FB5508043FF55EBD56AB",
INIT_28 => X"017DAAFFFAE821C0A0717D1C5B575FFB68E82557FD2082000BEAE905C755003F",
INIT_29 => X"D74BAE3AE85480FFFFC00AABE8E105C755517DF40552ABDF45B6AEAFFD5F7A48",
INIT_2A => X"FFAF7DA2AE905EF0075D5545E3F5EFF57F7D5C55D7492E90E3808756DA92EBFF",
INIT_2B => X"F5C7092FF801756D490A10438EBA4B8E9241043AE10EAF5C5547FF80954AA5D7",
INIT_2C => X"00000000000000000000000000000E124105D5B7FF7DB6AAAABC7BEDB505EFBE",
INIT_2D => X"515157555AAD142040A2D57FFFFFFAEBFF555D0028A005100000000000000000",
INIT_2E => X"500003FF55AAFD6AB455157D74BAF7AAA8B45AAFBD54005D7BD54AAF78002155",
INIT_2F => X"10F7AA8215555003FEAAAAC53DEB8A2FDDC01051AE955F7AAFBC0000AF843FF5",
INIT_30 => X"F51F782BCB47ABAE801FFAAFBEAA105D2E955FF557BD74EFFBACD41577B84000",
INIT_31 => X"0AAA00557FEA8A2FDD64BAAF8282012AFFEC20BAF7AA8015558517FF555D2ABD",
INIT_32 => X"48547AE04174BA557BEABEFA2AA951FF88554214FA2D3EAF57AFFDD7555082AA",
INIT_33 => X"22A955FFFFC21FFF3BE40412DE02955FF082A820AAAB842AA00000028AB0AAFF",
INIT_34 => X"0000000000000000000000000000000000000000000002A80010557BFDFFFF78",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000008000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(3),        -- Port A data input
DOA(0)   => data_read_a_hi_256(3),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(3),        -- Port B data input
DOB(0)   => data_read_b_hi_256(3),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_4_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10804002061080A284201081034809800A00230340007833522C82D04A16006",
INIT_01 => X"804399801838084C0420450E1E104348403008418984014902030006A0910204",
INIT_02 => X"480108A200000000446418E01E80F00A4104311868240200080000000988A390",
INIT_03 => X"065140108800004080064A0002001128270072E03000000030808D00888100F0",
INIT_04 => X"9100EB836A155C1AF0B81CD60433B944022AB8385AC0D4B8E02010E81C32E821",
INIT_05 => X"5C0F20B36F08000024C084C501441C4CF01C489533483C8042EAC190001074C4",
INIT_06 => X"0034420151620118120106902406C3C7800201448DD9D2871020F2AA375A6071",
INIT_07 => X"12181000023480040840C001E080030032009700024641000C00187A442007C2",
INIT_08 => X"8084830110160218004000001101121F220000260000108AA000440880000000",
INIT_09 => X"5A8C881063DF3E839008F29F407448F200B020DA841CA2001001008882046647",
INIT_0A => X"C61504C1380101801900439001FD8804041400001002003C230B6715A4786E0F",
INIT_0B => X"ACD1240522E000098100D104B26041348A088078116C105DA006D10416BE3002",
INIT_0C => X"8608086180860808608086180860A0434C0430D4A25F3182CC4D5D221A09E821",
INIT_0D => X"0BC28081080549504400A8080009B878184044881222D1821821A08628086180",
INIT_0E => X"20481E0E18790012820001100200D02048300418022C1282809A09040415002A",
INIT_0F => X"0000010020005E0090000001000000C6009000000100000000380E6C30830806",
INIT_10 => X"000000800000D20090000001000000EE0090000001000000A6A2000000000000",
INIT_11 => X"0000000000000000008100003B00200800000000000020010002EA0080200000",
INIT_12 => X"80800000080000211D80000C0044281000400000000000004000000010003282",
INIT_13 => X"03B00410000000400121800000000000000008020000B8020800000020006F00",
INIT_14 => X"59000402000000000008020000C9000200800000000000200FC0101000000100",
INIT_15 => X"008A500100001040000000000000200002000042E00000000000000002080001",
INIT_16 => X"08820440040802500104C34820E3031B63C20530C01800410009009821040A00",
INIT_17 => X"C832008020C812008220C81200802048320880204832008020C8320082204812",
INIT_18 => X"8120481208822008020C812048320880208802048320C8120882204812088020",
INIT_19 => X"10A3A5930C9A6CB261934E048320C81200822008220C81204832008020882204",
INIT_1A => X"8A28A28A2BD30264686668A28A2605145031C03F028000A1C2ED7831A2822250",
INIT_1B => X"51A8D46A351A8D46A351AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA28A2",
INIT_1C => X"F94304068341A0D068341A0D068341A0D068341A0D068341A0D068341A0D0683",
INIT_1D => X"BAAA84154005500000000000000000000000000000000000000000000000401F",
INIT_1E => X"4AAF7D168B45AAAABDF55A2802AA1000002ABFF087FFDF5508003FEBA087FD54",
INIT_1F => X"015500002AABA082E954005500021FF5D2EBFF5500003DF455555421EFAAFFD5",
INIT_20 => X"174BAA2AABDE0055517FF555555420AAAA843DFFFAAD1554005D7FD74AAAA840",
INIT_21 => X"400155AAD1554AAF7802AB4500043DF45FFD168BEF080028BFF0855555455500",
INIT_22 => X"803FEBAFFD5420BA085168A00007BFDE10085168ABA0055574BA5555554BA5D0",
INIT_23 => X"02A97545F7D1555EF55043DF5555517DEAA5D0400010A2AA955FF55003FE10F7",
INIT_24 => X"000000000002A82155A2FBFFEBA0800021550855555FFAA84001FFAAFBEAB450",
INIT_25 => X"5080A3AEAA007BD2482BE84124285C0000000000000000000000000000000000",
INIT_26 => X"381451471D7AAFBD0492EBD56DB7DBEAEBFF55BC042AA101D0A28BC7007FFDF4",
INIT_27 => X"400557FD54AABE84001C5550A28ABA1424974004100021FF492AB8F7D1C0438E",
INIT_28 => X"8BEF005557545490012482B6A0BAE2849557AFED1C5F470AABE8A3AFD7A2DF55",
INIT_29 => X"504924955524AA140E0717DAADB50492EB842FB5508043FF55EBD56ABD75D042",
INIT_2A => X"A905C755003FE28E3803DEAAEBDF40002557F6DA101475FDE10145F68A921C55",
INIT_2B => X"DF425575D7BEFB55002097555FFD5401EF5D043AF6D405F78E3A1C2002000BEA",
INIT_2C => X"0000000000000000000000000000208017DAAFFFAE821C0A0717D1C5B575FFB6",
INIT_2D => X"512EAAB45007FFFF55082EA8AAA087FC2010F784000AA5900000000000000000",
INIT_2E => X"F002EA8BEF5D0428ABA595557555AAFBC2000A2D57FFFFF7AEBFF55FF8028A00",
INIT_2F => X"BAF7AAA8B45AAFBD54005D7BD54AAF78002155512AAAA085D04174100800021F",
INIT_30 => X"F55AAFD6AB4551002ABEF005555555000402000FF802ABAA04552ABFF597FD74",
INIT_31 => X"DE005D7BE8AA85555400100879560AA592F955FFAAFBC0000AF843FF5500003F",
INIT_32 => X"FCABA598400010F7AA8215555003FEAAAA843DEB0A2FD5600051537DE005D557",
INIT_33 => X"E955FF557BD75EFFBBCD415521FBFDF45000417545FFD5421FF5D0428BEF0079",
INIT_34 => X"00000000000000000000000000000000000000000000004001FFAAFBEAA105D2",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000010000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(4),        -- Port A data input
DOA(0)   => data_read_a_hi_256(4),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(4),        -- Port B data input
DOB(0)   => data_read_b_hi_256(4),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_5_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50DB4A0791B1B4B694369283C81F9996A091832112004AB37B20E07C0C1E006",
INIT_01 => X"085FBC448000804C446A00000034826841280A00084000C8C212802EE2953235",
INIT_02 => X"C809AD5CB118E640A4D018FC011FF0002080000082C8C66609DB7DDDCB1F2036",
INIT_03 => X"250907263E4C90D210835C82484205720B20640A88800000B8E0F810A8C4500E",
INIT_04 => X"4005102126898100064D20001044429C7824382C0416C087198AB916E0551A24",
INIT_05 => X"A370C14CA0E101094008002389CFE2F20D7D7A114CB5C20AE514178054948912",
INIT_06 => X"547319A1499121D4C0A046FC4E06C030581859058C2404844437118630839B88",
INIT_07 => X"2A53468D1A758C038AFFEA9FE39348C9204C389672407EF120EA5806E6C543AC",
INIT_08 => X"8C05896372728FE0C420619000003AFF48D1222E5D26F06ABCC96CD72C463990",
INIT_09 => X"82DE9AB9182080C801041080300F6F0E42821809C2FEA0B65A212282002B029F",
INIT_0A => X"1688E480D10A90049026145B3830B64944904569E7E00A002C836D35B68D26C0",
INIT_0B => X"88990E14269AB54B078092E6BD4431138A00AEFDD567DA480816848C94180846",
INIT_0C => X"C0591C0791C0491C0791C0591C06A8E0248E03D68860A0106119883D6AE1A0A4",
INIT_0D => X"23D829FA654184533252095E542387F81008071C1BAAD68B027029C0491C0691",
INIT_0E => X"0CA7FE0227FC25847C4395166C5844480204011210A11028C380802A24C89494",
INIT_0F => X"1C55D65E3E3C017C37FC3E0017C1F8017C37FC3E0017C1F90005024108308061",
INIT_10 => X"1C0118796FE0017CA7FC3E0017C1F8017CA7FC3E0017C1F9100DFFF5E15D0610",
INIT_11 => X"FFF3E34F00C0270F3755F1F8007FCBEBE25E0700463E17F2C7E014FF7AE6CD38",
INIT_12 => X"64E4090626DE40100459759173BBD6EF37C523E6030061341F07FC571F8F800D",
INIT_13 => X"E0A6FE28C3082636F201BFFF807E00007E03F7243D38337D1C6184131B7C1DEF",
INIT_14 => X"397FFA0E0E06101C53E36C3D3E884FDDD28381C0098E57D923BDFC8C8120C4DB",
INIT_15 => X"FA36FDF58DBF81C062540049707E0FE7303D3E03BFFF41478040570EED50F4F8",
INIT_16 => X"88212B100901A2349004C26A624A21040FC190050A2110B8ACC40B204A119074",
INIT_17 => X"C20080230802108C2008C22080210882108C220842208821088210842208C200",
INIT_18 => X"20084220842208C2008823080230802108823084220842008821080230842008",
INIT_19 => X"54C1892596D34924B2DA6884220842008C20084220802108821080230802308C",
INIT_1A => X"BEFBEFBEFB7F7FE7EFEEE79E79EFAF2DDA73FBDCEDBFF9D3F0FDE0DB6DBF6218",
INIT_1B => X"DEEF77BBDDEEF77BBDDEEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEF",
INIT_1C => X"FAF3167BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBD",
INIT_1D => X"BA5D2ABFFEFFF80000000000000000000000000000000000000000000000401F",
INIT_1E => X"F5508003FEBA087FD54BA0804154005555574AAA2802AA10FFFFFDE0008556AA",
INIT_1F => X"AA1000003FEBA00002AABA5D2EBFEBAAAD16AABAF7AAA8BFFAA802ABFF087FFD",
INIT_20 => X"E8B45FF80001555D2E955FFFFD5421EFAAFFD54AAF7D168B45AAAABDF55AA802",
INIT_21 => X"02AABA082E954005500021FF5D2EBFF5500003DE005555575EFA2D142145A2FF",
INIT_22 => X"7FD74AAAA840014500517FFEF007BEABFF5D7FC00BA5D5568AAAF7AAAAAAAAA8",
INIT_23 => X"2FBEAA105D2E97410FFD16AAAA5D2ABDEBAFFD5420AAAA843DFFFAAD1554005D",
INIT_24 => X"000000000000028BFF0855555455500174BAA2AABDE0055517FF555504154BAA",
INIT_25 => X"0FFFFFFE38085F6FA92552AB8FEFF78000000000000000000000000000000000",
INIT_26 => X"C7B68A28BC70075FDF45080A3AEAA007BD24821E84124285C51574BAB68A2DA0",
INIT_27 => X"B7DBEAEBFF55BE842AA105D0A38EBA1C0428A925D2AB8EBABEDB6AA92F7AAA8B",
INIT_28 => X"75EFA2DB45145B6F5EFB6DF78E05145552A925FFFFD1471D7AAFBD0492EBD56D",
INIT_29 => X"68AAAF7AAAAA82BE8A28A921424974004100021FF492AB8F7D1C0438E38145B5",
INIT_2A => X"A3AFD7A2DF55400557FD54AABE84001C555517DFC70875EABC7557FC20AA415F",
INIT_2B => X"043AFED1C0E10492B6FFEFA105D2A95410FFDB6FABA542ABAE2AF7DF470AABE8",
INIT_2C => X"00000000000000000000000000000428BEF005557545490012482B6A0BAE2849",
INIT_2D => X"5955554BAFFAEBDE10F7FBFDEBA007BFDE005D2AAABEFFB80000000000000000",
INIT_2E => X"AF7FBE8A00FFAEAAB45F3AAAAB4500557FF55082EA8AAA087FC20105504000AA",
INIT_2F => X"55AAFBC2000A2D57FFFFF7AEBFF55FF8028A00512AA8AAA5D0028A005D2AA8AB",
INIT_30 => X"BEF5D0428ABA597FD55FFA2FFD5555FFD57FFEFFFAA97545552A821EFFBD5575",
INIT_31 => X"8B55557FC0012087FEAABAF7AAAAA10F3AAAAA005D04174100800021FF002EA8",
INIT_32 => X"A8ABAFBFFD74BAF7AAA8B45AAFBD54005D7BD54AAF7800015551517DF4500516",
INIT_33 => X"402000FF802AAAA04452ABFF592E80010FFFFFFE005D2A95410F7FFFFEBA5D2E",
INIT_34 => X"000000000000000000000000000000000000000000000002ABEF005555555000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000060000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(5),        -- Port A data input
DOA(0)   => data_read_a_hi_256(5),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(5),        -- Port B data input
DOB(0)   => data_read_b_hi_256(5),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_6_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10804B0061A010A2840012C030028180004003220200403302301C0381A0086",
INIT_01 => X"A70041CA3839684D18A160000C52424841000000090800090210080008110204",
INIT_02 => X"080108200C1000004465480400C0080100000000010432400800800009882050",
INIT_03 => X"040001008C2340D0842208624210802182800584488000103080014E08C10000",
INIT_04 => X"00101611A029B08410044800000000040088122A44281C040400900500001800",
INIT_05 => X"02800000400C820934E4A0002900404402820024000A00824004283011200A00",
INIT_06 => X"2632000004084804134DA7C011A83FC012122100C80812D00308010000829400",
INIT_07 => X"02181020423088002940C2401D0480112000100004404014602447F805326393",
INIT_08 => X"7004812130160008304000000000021F020408244000108A0000440003040000",
INIT_09 => X"020C889010104088A000348037F05840303902E814000010341108802020FF40",
INIT_0A => X"86C8B5DF1C83C9C8900000100220C244840021100017E2FD200000A40001223F",
INIT_0B => X"88D1804122A088018152D144317205502A880C00107FD75DE922005026A62A15",
INIT_0C => X"B6284B6284B6184B6184B6384B62825B0425B0568075A0826849C8229AC5F8AE",
INIT_0D => X"03C440C054048850A300A8480009A0020865A588DA20F1A2D92D82B6084B6084",
INIT_0E => X"031001E0800122100321C89214A01A742D3A168D1B4686D100234B442428C034",
INIT_0F => X"000008AB80030202800000001402068202800000001402067400026000000000",
INIT_10 => X"00000000341E8202100000001402068202100000001402062840000800000000",
INIT_11 => X"0008000000000000083C00052000300000000000000008CD0018400081000000",
INIT_12 => X"800800000069A48584000A0400000010001000000000000000048128C0002840",
INIT_13 => X"1A480012000000034C1E000040000000000400FE000644020100000001A34000",
INIT_14 => X"02800401000000000004BA000112B0020800000000000807E80000110000000D",
INIT_15 => X"0500020250001000100000000000010CCE000198000020000000000010F80006",
INIT_16 => X"62D18468CE8402440404D24A3081B020603E0A20640C8400010298432A002A00",
INIT_17 => X"ED3B4ED0B42D1B4ED3B42D0B42D1B4ED2B42D0B46D3B4ED2B42D1B46D3B4AD2B",
INIT_18 => X"D0B46D3B4AD0B46D1B4AD3B4ED0B42D1B4ED2B4ED1B42D0B4AD3B4ED0B42D0B4",
INIT_19 => X"002331C618E38E38C31C7346D3B4AD2B46D1B42D2B4ED2B42D1B46D2B4AD1B42",
INIT_1A => X"8E38E38E39DB3B676F66EFBEFBEFAFBC5E73FC7F87A7D4ABFE7CFAFBE7BF8040",
INIT_1B => X"CFE7F3F9FCFE7F3F9FCFE38E38E38E38E38E38E38E38E38E38E38E38E38E38E3",
INIT_1C => X"FF75A43F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9F",
INIT_1D => X"BA5D7BEAAAAFF80000000000000000000000000000000000000000000060401F",
INIT_1E => X"A10FFFFFDE0008556AABA5D2ABFFEFFF843DFEFA2FBD54BA5555554BAAAFBC20",
INIT_1F => X"5400550428AAAAA84021FF007BD54BAAAD17DEBA0855421455555574AAA2802A",
INIT_20 => X"17400AAFBE8ABAF7FFD54AAAA802ABFF087FFDF5508003FEBA087FD54BA00041",
INIT_21 => X"03FEBA00002AABA5D2EBFEBAAAD16AABAF7AAA8BFFAAD1554BA002A95555A284",
INIT_22 => X"AABDF55AA802AA100000001EF087FEAA00FFFBD5545080417555A2D17FE10000",
INIT_23 => X"2803DFEF0855401FF082EA8B555D7FC21FFFFD5421EFAAFFD54AAF7D168B45AA",
INIT_24 => X"0000000000055575EFA2D142145A2FFE8B45FF80001555D2E955FFFF843DEAAA",
INIT_25 => X"A415B52492B6F5C20825D7FE8A92FF8000000000000000000000000000000000",
INIT_26 => X"555551574BAB68A2DA00FFFFFFE38085F6FA92552AB8FEFF78E3DFFFAAFFD04A",
INIT_27 => X"EAA007BD24821C04124281C0E2DA82BE8E001EF147BD2482BED57AE921451421",
INIT_28 => X"24AA14209557DA28E15400BEF1EFA92FFFFD24BAB68A28BC70075FDF45080A3A",
INIT_29 => X"17545B6D178E281C0A38EBA1C0428A925D2AB8EBABEDB6AA92F7AAA8BC7B6D55",
INIT_2A => X"BD0492EBD56DB7DBEAEBFF55BE842AA105D0E071FF0071EDA38F7F1D55550004",
INIT_2B => X"2A925FFFF8E3DE82BE8E38FFF0851401C70824A8B555C7FC2147F7D1471D7AAF",
INIT_2C => X"00000000000000000000000000005B575EFA2DB45145B6F5EFB6DF78E0514555",
INIT_2D => X"FBAABDFEFAAFBC00BA007BC0000FFD542000557FE8A00F380000000000000000",
INIT_2E => X"0F7D168A105D55421455155554BAFFAEBDE10F7FBFDEBA007BFDE005D2AAABEF",
INIT_2F => X"4500557FF55082EA8AAA087FC20105504000AA592ABFE00F7AA821FF557FC001",
INIT_30 => X"A00FFAEAAB45F3D5400BA5504155EFAAAE95410F7D57DE00FFFBC00AAFBAAAAB",
INIT_31 => X"FEAAF7D157545080417545F7D56AAAA592AA8AAA5D0028A005D2AA8ABAF7FBE8",
INIT_32 => X"C2145F3D557555AAFBC2000A2D57FFFFF7AEBFF55FF8028A00512E975FF08557",
INIT_33 => X"57FFEFFFAA97545552A821EFFBAABDE00F7AAAABEF005542155000028B555D7F",
INIT_34 => X"0000000000000000000000000000000000000000000007FD55FFA2FFD5555FFD",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000048000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(6),        -- Port A data input
DOA(0)   => data_read_a_hi_256(6),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(6),        -- Port B data input
DOB(0)   => data_read_b_hi_256(6),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_7_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10840B0048225802842102C02450418800002300500030B313300C418992002",
INIT_01 => X"A34009C23838684D1C20E0000E11426840000000080000080200090000510200",
INIT_02 => X"4801082048100000446558040080000041000000000622400800000009000010",
INIT_03 => X"040001818CA144D0842248424210812102000400088000003080014688800000",
INIT_04 => X"000010002041800000048000000000040088322944200C850001940400301800",
INIT_05 => X"0200000040004100280040204104004402000025000800065004203030320800",
INIT_06 => X"0430060044084804900806D1112A002012120004440812D40120008200829001",
INIT_07 => X"02181020423408002940C24001A4A010200018920646C10C7035000244004380",
INIT_08 => X"008481213016020C204000000000121F020408264000100AA000440012040000",
INIT_09 => X"820C899410000000A100348020005902B1A0048825008091350100CAA0200280",
INIT_0A => X"50140A0010058188100004590331C9C4A400231200340C012100002400012200",
INIT_0B => X"1811C44D22A1884141600411800008104080890023000009A926801050001C00",
INIT_0C => X"9002C9002C9022C9022C9022C903064809648080204020004009080A0A00E088",
INIT_0D => X"0880144434A0010012280008031980036000014A0046206241A4069002C9002C",
INIT_0E => X"0216000200010000000081102080400040002000002010000004008080048A00",
INIT_0F => X"038A2881210382000000001E003E0582000000001E003E042283424000000000",
INIT_10 => X"60700706901982000000001E003E0582000000001E003E046840000000009864",
INIT_11 => X"00000000330C00F0C8210807200000000000581C01C1C809201C400000000001",
INIT_12 => X"0000C2419121028C00020A2400000000000080082C180603A0E003A090406840",
INIT_13 => X"14E8000004321189085F8000000061E001FC00C00207740000021908C4829D00",
INIT_14 => X"BB800000009864038C14800201BAB000000026130071A80613A0000018483224",
INIT_15 => X"0546520350000600812058100F81C018880201BBA0000008239020F110800806",
INIT_16 => X"24003300080022140444D268624B210040004A08000000044222900320C84008",
INIT_17 => X"4010040100402000000000000003004010040100000000000000100401004010",
INIT_18 => X"0000C01004010000000001004010040000000004010040300400000000000200",
INIT_19 => X"54A2C208200010410400000800000000040100C01000000000100C0100400000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000002A10",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FAF8800000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"55002E820AAAA80000000000000000000000000000000000000000000000401F",
INIT_1E => X"4BA5555554BAAAFBC20BA5D7BEAAAAFFFBC00AAF7D5575455D557DFEF002AAAB",
INIT_1F => X"FFEFFFAAAAAAAF7D57FFEFF7D555555A2AEAAB55007FD74AAAA843DFEFA2FBD5",
INIT_20 => X"FDF550000175555504175450055574AAA2802AA10FFFFFDE0008556AABA5D2AB",
INIT_21 => X"428AAAAA84021FF007BD54BAAAD17DEBA085542145552ABDFEFFFAA801EFFFFB",
INIT_22 => X"7FD54BA000415400557BD74BAFFD140000082A975EF00003DF55555168A00000",
INIT_23 => X"5557FEAAA2843FF55A2AEA8B55AAAABDEAAFF802ABFF087FFDF5508003FEBA08",
INIT_24 => X"0000000000051554BA002A95555A28417400AAFBE8ABAF7FFD54AAAAAEA8ABA5",
INIT_25 => X"5415178FD7082EAAB550820870BAAA8000000000000000000000000000000000",
INIT_26 => X"82AA8E3DFFFAAFFD04AA415B52492B6F5C20825D7FE8A92FFFFC70BAE3D15555",
INIT_27 => X"E38085F6FA92552AB8FEFF7A0ADABAEBD578FFFEBD55557DBEA4AFB550871D74",
INIT_28 => X"DFD7FFA4801D7F7F5FDF55000E17545410E175550051574BAB68A2DA00FFFFFF",
INIT_29 => X"3AF55415F6DA38080E2DA82BE8E001EF147BD2482BED57AE921451421555524B",
INIT_2A => X"5FDF45080A3AEAA007BD24821C04124281C7BD2482E3D1450381C20905EF0800",
INIT_2B => X"FFD24BAB6A4A8A82495F78E92AA843DF45BEAAAFB55ABA0BDE02EB8A28BC7007",
INIT_2C => X"000000000000000000000000000055524AA14209557DA28E15400BEF1EFA92FF",
INIT_2D => X"F3FFD54BAAAD15754508556AB45002AA8B450800174BAA680000000000000000",
INIT_2E => X"FF7803DF45085557410AEAABDFEFAAFBC00BA007BC0000FFD542000557FE8A00",
INIT_2F => X"BAFFAEBDE10F7FBFDEBA007BFDE005D2AAABEFFB803DEAAAAD56ABEFAAD5575E",
INIT_30 => X"A105D554214551003FF45FF8400145FFD57FF55082E97555002E955550C55554",
INIT_31 => X"54AA5500021EF000028B55087BFDEBA042ABFE00F7AA821FF557FC0010F7D168",
INIT_32 => X"3FE10AEAAAAB4500557FF55082EA8AAA087FC20105504000AA597FC2010A2D15",
INIT_33 => X"E95410F7D57DE00FFFBC00AAFB8028A00007FE8A00A2803FF45F7AABDF55AA84",
INIT_34 => X"00000000000000000000000000000000000000000000055400BA5504155EFAAA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000007FFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(7),        -- Port A data input
DOA(0)   => data_read_a_hi_256(7),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(7),        -- Port B data input
DOB(0)   => data_read_b_hi_256(7),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_8_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00000648E2840112C00000418000002700500030B3132000400812082",
INIT_01 => X"A14008420008204D042100000212026840000000180800080200090048510204",
INIT_02 => X"080108000090000004655C040080000051000000000402400800000009000010",
INIT_03 => X"00000100803008D0842240024210810002800584488000103080894288800000",
INIT_04 => X"00009610A028B084000440C0040000040088323244280C950400808500321800",
INIT_05 => X"42800080400C8A09306420202804400402800035200A00020204283001114A00",
INIT_06 => X"2230400041404B141345A7C20426FFC01292214444081254002801A200821400",
INIT_07 => X"021810204214080069408200008C1010200018920E06C0000020DFFA453223D3",
INIT_08 => X"0084010110120008024000000000021F02040826400000008000440000240000",
INIT_09 => X"828D8880100040898128768820045142B0B902E815008080A0B13848A2200280",
INIT_0A => X"9148A4801C81C9C8100004590711800414002004402008013000403084090200",
INIT_0B => X"BC95C44522A002410040940084720450220089000100104DE924800030821452",
INIT_0C => X"0000400004000040000400004000220010200114AA4020004009092A0009E0A8",
INIT_0D => X"0BC4028430108150900408590109A00209642500120230200100220020400004",
INIT_0E => X"0010000600002210A320C89000005A142D0A16850B6294D10023420124240114",
INIT_0F => X"00000800008100020003C1FE00020080020003C1FE0002004401426008208041",
INIT_10 => X"E3F00000100080020003C1FE00020080020003C1FE000200080000081EA2F9EC",
INIT_11 => X"00081CB0FF3C000008000201000010001DA1F8FC0000080110080000010132C7",
INIT_12 => X"0B0BE6C00020040580040200000001004832CC19FCF81E000000010000200800",
INIT_13 => X"020000C31CF60001008000007F01FFE00004000200420000618E7B0000804000",
INIT_14 => X"000000F151F9EC0000040200401000200D547E3F00000800080001617AD80004",
INIT_15 => X"0100000822406E1B95A3F83000000008020040100000BAB87FB0000010080102",
INIT_16 => X"66D1A368C68D26000544D26A504AB12040022220640484000110184300002A02",
INIT_17 => X"6D1B46D1B46D1B46D1B46D1B46D0B42D0B42D0B42D0B42D0B42D1B46D1B46D1B",
INIT_18 => X"D1B42D0B42D0B42D0B42D1B46D1B46D1B46D1B42D0B42D0B42D0B42D0B42D0B4",
INIT_19 => X"442200000000000000000346D1B46D1B42D0B42D0B42D0B42D1B46D1B46D1B46",
INIT_1A => X"9E79E79E7B7F11E66C6FAD96D96520145052A1F5E2BD085122ED48F3AEB20840",
INIT_1B => X"C3E1F0F87C3E1F0F87C3E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7",
INIT_1C => X"FA2A6D4F87D3E1F4F87D3E1F4F87D3E1F4F87D3E1F4F87D3E1F4F87D3E1F4F87",
INIT_1D => X"FFFF84000AAFF80000000000000000000000000000000000000000000000401F",
INIT_1E => X"5455D557DFEF002AAAB55002E820AAAA840000000043DF55087BC01EF007FD75",
INIT_1F => X"AAAAFFAA95545552ABFE00087BC00AA082EBFE10A28028AAAAAFBC00AAF7D557",
INIT_20 => X"E8BFFA2FBFFFFFAAD5400AAFF843DFEFA2FBD54BA5555554BAAAFBC20BA5D7BE",
INIT_21 => X"AAAAAAF7D57FFEFF7D555555A2AEAAB55007FD74AAAAD57FF45002A975FF007B",
INIT_22 => X"556AABA5D2ABFFEFFFAA82000555555545AAFBE8A00082A97410F7D5555EFAAA",
INIT_23 => X"87BC2010AAD54014500516ABFFA2AABDF450055574AAA2802AA10FFFFFDE0008",
INIT_24 => X"000000000002ABDFEFFFAA801EFFFFBFDF550000175555504175450000155450",
INIT_25 => X"50075C71FF087BD75D7FF84050BAEB8000000000000000000000000000000000",
INIT_26 => X"BABEFFC70BAE3D155555415178FD7082EAAB550820870BAAA8407000140038F4",
INIT_27 => X"492B6F5C20825D7FE8A92FFA497545552AB8E10007FC50BA002ABFE00AA8A2AA",
INIT_28 => X"DF451C24955EF0875EFBD7B6F1FFFC7BEDB45082EB8E3DFFFAAFFD04AA415B52",
INIT_29 => X"92410EBD5505EFB6A0ADABAEBD578FFFEBD55557DBEA4AFB550871D7482AAD17",
INIT_2A => X"A2DA00FFFFFFE38085F6FA92552AB8FEFF7AA87000415B5057DAAFBE8A100820",
INIT_2B => X"0E17555000E17545007BC0000BED14217D005B6ABC7B6AABFFED0051574BAB68",
INIT_2C => X"000000000000000000000000000024BDFD7FFA4801D7F7F5FDF55000E1754541",
INIT_2D => X"A684174105D042AB550055555FF007BD7555F784174AAA280000000000000000",
INIT_2E => X"A082EBDE10AAAEA8ABAF7FFD54BAAAD15754508556AB45002AA8B450800174BA",
INIT_2F => X"EFAAFBC00BA007BC0000FFD542000557FE8A00F384175555D2EA8A00087BD74B",
INIT_30 => X"F45085557410AED17FF455D04155FF00557DF55FFD57DF55FFFBD5400A2AABDF",
INIT_31 => X"21EFA2FFEAA00000002010A2D5421FFFF803DEAAAAD56ABEFAAD5575EFF7803D",
INIT_32 => X"BDFEF0855554BAFFAEBDE10F7FBFDEBA007BFDE005D2AAABEFFBAE97410087BC",
INIT_33 => X"57FF55082E97555002E955550C2E95555087BC0010FFD1401EF087FE8B55FFAE",
INIT_34 => X"000000000000000000000000000000000000000000000003FF45FF8400145FFD",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000020000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(8),        -- Port A data input
DOA(0)   => data_read_a_hi_256(8),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(8),        -- Port B data input
DOB(0)   => data_read_b_hi_256(8),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_9_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00018248A2840112C00002C18000002300500030B3132000400812006",
INIT_01 => X"A1400802000020490000000000000240413C0A61590001D90213C90008510204",
INIT_02 => X"680108200010000054655C040080000041000000010402400800800009082011",
INIT_03 => X"00040100800020D0842240124210810042800504488000103081894288800000",
INIT_04 => X"00001410A00AA084000400C0060000040088323044201C850020820400101880",
INIT_05 => X"0200020040048A09202420000C00410402000025000800020804203000100800",
INIT_06 => X"22320400404048041144A7D2003A002012120004DC08125400A0008300821000",
INIT_07 => X"06181020421C08000940820000800010200018B20206C00000200002441223C1",
INIT_08 => X"0184010110120008004000000000061F02040826400008118000440000040000",
INIT_09 => X"8208888210004009010852882000510230A900A8040080800055086002200280",
INIT_0A => X"1402008004814948100004590111C004040120000020080121024012A4081200",
INIT_0B => X"2C91844522A0004100488000801200D00000880001000415E1248002103C2294",
INIT_0C => X"080040820408004082040800408202040020410402000000400809080508A080",
INIT_0D => X"0B4000803200C150108008490809A00219246101100220202102020820408204",
INIT_0E => X"00160006000120002120499020A04A14650A328519629651900142002404201E",
INIT_0F => X"0000080A20010002100000001402008002100000001402000001426008208041",
INIT_10 => X"0000000034008002800000001402008002800000001402008800000800000000",
INIT_11 => X"0008000000000000081500010000100800000000000008C10008000001200000",
INIT_12 => X"0088000000680005800002000000000000500000000000000004810010000800",
INIT_13 => X"02E8040200000003401F80004000000000040027000274000900000001A05D00",
INIT_14 => X"3B8000030000000000042B00009AB00008800000000008012BA010010000000D",
INIT_15 => X"0106520350000040100000000000010C0300009BA000200000000000105C0002",
INIT_16 => X"6651B328CA8D26540544924272EB91004002022024048400000098030A000A00",
INIT_17 => X"2509425094250942509425094250942509425094250942509425194651946519",
INIT_18 => X"5094250942509425094251946519465194651946519465194651946519465194",
INIT_19 => X"0480800000000000000001465194651946519465194651946509425094250942",
INIT_1A => X"34D34D34D1285B080201C92410480AB9A26667A46F345448020082E1C712A054",
INIT_1B => X"8341A0D068341A0D06834514514514514514514514514514514514514514D34D",
INIT_1C => X"F8B2B60D069349A0D068341A4D268341A4D268341A0D069349A0D069349A0D06",
INIT_1D => X"EFA2FFFFF555D000000000000000000000000000000000000000000000007FFF",
INIT_1E => X"F55087BC01EF007FD75FFFF84000AAFFD57DF45A280154BA5555401EFFFD5421",
INIT_1F => X"20AAAA843DFEF00517DEBA007BFDFEFFFD1575EF00557DF555D040000000043D",
INIT_20 => X"68AAAF7802AA00FFFBD7555087BC00AAF7D5575455D557DFEF002AAAB55002E8",
INIT_21 => X"A95545552ABFE00087BC00AA082EBFE10A28028AAAAAAABDF45F7803FFEF5555",
INIT_22 => X"FBC20BA5D7BEAAAAFFFBC00AA552E95545087BD54BA550417400085155555082",
INIT_23 => X"2FFFDF555D7BE8BFF5D51575EFA280175555D043DFEFA2FBD54BA5555554BAAA",
INIT_24 => X"00000000000557FF45002A975FF007BE8BFFA2FBFFFFFAAD5400AAFF8402000A",
INIT_25 => X"2415B471C7E3DF451EFBEFBFAF45490000000000000000000000000000000000",
INIT_26 => X"45490407000140038F450075C71FF087BD75D7FF84050BAEBDF78F45B6801048",
INIT_27 => X"FD7082EAAB550820870BAAA8438FFF00517DE82007FFAFEFE3DB505EF1C5B7AF",
INIT_28 => X"8F45F78A3DFD741516DAAAE38E2DA28EBFFD55451C7FC70BAE3D155555415178",
INIT_29 => X"1543808515756D1C2497545552AB8E10007FC50BA002ABFE00AA8A2AABABEAEB",
INIT_2A => X"FD04AA415B52492B6F5C20825D7FE8A92FFFFC20BA5D2E905550071D54825D0A",
INIT_2B => X"DB45082EB8002000AAFFFDF6D417FEABEF5D55505FFBE801256D490E3DFFFAAF",
INIT_2C => X"0000000000000000000000000000517DF451C24955EF0875EFBD7B6F1FFFC7BE",
INIT_2D => X"A2FBEAB45F78402010007BD5545AAFFD55EFF7FBE8B550000000000000000000",
INIT_2E => X"FAAFFC01FF557FE8B550004174105D042AB550055555FF007BD7555F784174AA",
INIT_2F => X"BAAAD15754508556AB45002AA8B450800174BAA68028BEF00517FE10007BE8BF",
INIT_30 => X"E10AAAEA8ABAF7AAAAB45F7AEBFF4508557FEAAAAAEBFEAAAAFFD5545557FD54",
INIT_31 => X"0145005557400552A954BA0051575EF5504175555D2EA8A00087BD74BA082EBD",
INIT_32 => X"021FF002ABDFEFAAFBC00BA007BC0000FFD542000557FE8A00F3FFC00BA552E8",
INIT_33 => X"57DF55FFD57DF55FFFBD5400A28400010A2FBFDFFF007FE8BFF5551401EFF784",
INIT_34 => X"000000000000000000000000000000000000000000000517FF455D04155FF005",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000040000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(9),        -- Port A data input
DOA(0)   => data_read_a_hi_256(9),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(9),        -- Port B data input
DOB(0)   => data_read_b_hi_256(9),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_10_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000B0001800002840002C0000281800020030000000033022000000180006",
INIT_01 => X"0000098218302849180060000C00424040000000080000080200090008510200",
INIT_02 => X"0801080200100000044008000080000041000000002002400800000009008010",
INIT_03 => X"0001000004000040000202000000000802006400088000003080040008C10000",
INIT_04 => X"0000100022008000000C08C00C00000400201830040000040000000400001820",
INIT_05 => X"0200000040000000248080210044000400000000000800000004004010000800",
INIT_06 => X"0030040000404004000006D00008002010100000880800001000000030829000",
INIT_07 => X"02100000021008000940800001800010200018920206C01020200002440003C0",
INIT_08 => X"0084010110120010004000000000021F00000024400000008000440080040000",
INIT_09 => X"8288880010100001200852882004404000000008800000100001004202000280",
INIT_0A => X"0000008000020008100004590111824004000100000008012000401084080200",
INIT_0B => X"AC04400022808001200014000040001082800000000010500000010400808000",
INIT_0C => X"002200002000020002200022000020000100011082442000480909220001E020",
INIT_0D => X"0080000010044000000080080001800200000400020011000000200002000220",
INIT_0E => X"001000020001000020010010248000200010000800040000008009040000002A",
INIT_0F => X"0000000A00010200800000001400008200800000001400000000024008208041",
INIT_10 => X"0000000024008200100000001400008200100000001400002800000000000000",
INIT_11 => X"0000000000000000001400012000200000000000000000C10008400080000000",
INIT_12 => X"8000000000480000040002040000001000000000000000000004800000002800",
INIT_13 => X"0000001000000002408000000000000000000025000200020000000001200000",
INIT_14 => X"0000040000000000000029000010000200000000000000012000001000000009",
INIT_15 => X"0100000000001000000000000000010401000010000000000000000000540002",
INIT_16 => X"00001400080002100544924002A000004000020000080000000010032A000000",
INIT_17 => X"4010040100401004010040100401004010040100401004010040000000000000",
INIT_18 => X"0000000000000000000001004010040100401004010040100401004010040100",
INIT_19 => X"1080800000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"8A28A28A28D532A0CCC2A28A28A7AA344854A07F069CB8930AFD6A1AAA902A14",
INIT_1B => X"4CA6532994CA6532994CA28A28A28A28A28A28A28A28A28A28A28A28A28A28A2",
INIT_1C => X"FB3CC772B94CA6532994CA6572B95CAE532994CA6532995CAE572B94CA653299",
INIT_1D => X"55A2AABFFEF0800000000000000000000000000000000000000000000000401F",
INIT_1E => X"4BA5555401EFFFD5421EFA2FFFFF555D003FE10AAFBE8AAAA2D540000F7D57DF",
INIT_1F => X"00AAFF8002155AAFFE8B45AAD540000087FFDF45FFFBC2010AAD57DF45A28015",
INIT_20 => X"D5400FFD568B555D00155EF08040000000043DF55087BC01EF007FD75FFFF840",
INIT_21 => X"43DFEF00517DEBA007BFDFEFFFD1575EF00557DF555D517FEBA082A801EFF7FB",
INIT_22 => X"2AAAB55002E820AAAA803FEBA082AAAAAAF7FBFDE00A2FBC0145005168A10AA8",
INIT_23 => X"FAEAAB55AAD568B455D00154BAFFFBD75EF5D7BC00AAF7D5575455D557DFEF00",
INIT_24 => X"000000000002ABDF45F7803FFEF555568AAAF7802AA00FFFBD7555082E82155F",
INIT_25 => X"AAAD547038EBD57DF7DA2AEB8FC7000000000000000000000000000000000000",
INIT_26 => X"38A2DF78F45B68010482415B471C7E3DF451EFBEFBFAF4549003DE10BEF5EDAA",
INIT_27 => X"1FF087BD75D7FF84050BAEB8002155BEF5EDB6DAADF470280075FFF45E3F1C70",
INIT_28 => X"DEAA0824851EFEBFBD2410EBD168B7D410A175C7000407000140038F450075C7",
INIT_29 => X"C2155005F68A10A28438FFF00517DE82007FFAFEFE3DB505EF1C5B7AF45495B7",
INIT_2A => X"155555415178FD7082EAAB550820870BAAA8038EAA0824A8AAAEBF5FAE28AAF1",
INIT_2B => X"FFD55451C2087155EBA4A8B7DAADF68B7D4104104AAF7F1D75EF557FC70BAE3D",
INIT_2C => X"00000000000000000000000000002EB8F45F78A3DFD741516DAAAE38E2DA28EB",
INIT_2D => X"00043FE00F7D17FEBAA2D5574BAAAD17DFEFA2AEAAB550000000000000000000",
INIT_2E => X"A00557FF45A2D5554AAA2FBEAB45F78402010007BD5545AAFFD55EFF7FBE8B55",
INIT_2F => X"105D042AB550055555FF007BD7555F784174AAA28002155FFD17FFFFA2FBD74B",
INIT_30 => X"1FF557FE8B55007FFDEAA0004175FFA2FBC2000AAD16ABFF002A975450004174",
INIT_31 => X"AABAAAD56AABAAAD140155087FEAA10A28028BEF00517FE10007BE8BFFAAFFC0",
INIT_32 => X"555EF557FD54BAAAD15754508556AB45002AA8B450800174BAA68428AAA08042",
INIT_33 => X"57FEAAAAAEBFEAAAAFFD5545550015555A2842ABEFAAFBE8BFF0004020AAFFD5",
INIT_34 => X"0000000000000000000000000000000000000000000002AAAB45F7AEBFF45085",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000047FFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(10),        -- Port A data input
DOA(0)   => data_read_a_hi_256(10),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(10),        -- Port B data input
DOB(0)   => data_read_b_hi_256(10),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_11_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10180B05A0010402840602C2D001019000000300000000330A20080EC180002",
INIT_01 => X"AB400984B830084C1820E0000C36424840000000080000088200000802112220",
INIT_02 => X"8801081438106400A4F55800008000004100000040CCE24208005000C9060032",
INIT_03 => X"000406A492E6E440842254D002108153432004800880000030C0315688C00006",
INIT_04 => X"00001201200090001205400000000094108C322644240C840008030440111800",
INIT_05 => X"222000444008010028404002A002009402400025080880000C04223000170900",
INIT_06 => X"0431018040014804920906C74B32002012121004540816544522008200821100",
INIT_07 => X"3A5B1220421408004A56E840008B90D0200018B60A0650D450FC800644A0438A",
INIT_08 => X"0485816170760268E04000000000323F42C50826490640D28088445B0E041900",
INIT_09 => X"820F8B2C100000808120308020024002B3B01AC9540080A623213008800A0280",
INIT_0A => X"10000080D80381881000045B0511D28D94012671272008013002000220001240",
INIT_0B => X"8811865D22BB384100E010908060349322008000A1001C49A9348498B0808010",
INIT_0C => X"50639504395063950639504395062CA821CA8210A0040000480808214001A020",
INIT_0D => X"088812203360410110A40008553980021040465602023269400A202863950439",
INIT_0E => X"01160006000101004A01811064B050204810240812241280D00200A08044290A",
INIT_0F => X"1B0482A01AAEC3602330CD2A02952DC3502330CB4A0318B41400024008208041",
INIT_10 => X"1630144C0155C3502330CD2A02952DC3602330CB4A0318B5600C587149B6D014",
INIT_11 => X"587083B6A51005956308D1E8202C436375908AA840AD4513437640F15245B455",
INIT_12 => X"67062F47B2872400044959BC42B1060F0D036B80B548523136C158878D8FE04E",
INIT_13 => X"7010A2699AAA3794392000D81852B0A050C224180062085134CD1719564E020C",
INIT_14 => X"400C50500D94C8121713C02B555101C90705D71009604140C0418CE0C378F0B2",
INIT_15 => X"27C828E024D8C50965A40821568A06113801505010334AA73AA0666DAC20AD57",
INIT_16 => X"048123408C0822040004C248604B2100400100084008001D0113920060CDC06A",
INIT_17 => X"4812048120481204812048120481204812048120481204812048120481204812",
INIT_18 => X"8020080200802008020081204812048120481204812048120481204812048120",
INIT_19 => X"1420000000000000000002008020080200802008020080200802008020080200",
INIT_1A => X"2082082082815220A4A380000002A8313044020C0605885026853A1082100A00",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000008208",
INIT_1C => X"F83F070000000000000100800000000000000000004020000000000000000000",
INIT_1D => X"EF0855400005500000000000000000000000000000000000000000000000401F",
INIT_1E => X"AAAA2D540000F7D57DF55A2AABFFEF0804155EFAA842ABEFA280155EFFFFBC01",
INIT_1F => X"FF555D51575FFA2FFD75FF550015400FFFBFFF4508514000000003FE10AAFBE8",
INIT_20 => X"155EF0051555FF0804155FFF7D57DF45A280154BA5555401EFFFD5421EFA2FFF",
INIT_21 => X"002155AAFFE8B45AAD540000087FFDF45FFFBC2010AAD568AAAAAD142145FF80",
INIT_22 => X"7FD75FFFF84000AAFF802ABFFA2AABFE1008001540008514215555003DFFFA28",
INIT_23 => X"85142010FFAE800AA5D7BFDF45F7FFEAA0000040000000043DF55087BC01EF00",
INIT_24 => X"00000000000517FEBA082A801EFF7FBD5400FFD568B555D00155EF085168B450",
INIT_25 => X"7BE8A155EFE3FBC71FF145B42038550000000000000000000000000000000000",
INIT_26 => X"381C003DE10BEF5EDAAAAAD547038EBD57DF7DA2AEB8FC70000175EFB6802DBC",
INIT_27 => X"1C7E3DF451EFBEFBFAF45495F575FFBEF5D05EF550E15400E3F1FFF7D085B420",
INIT_28 => X"8ABAB6D145145FF84155D7085B555C71404105C7F7DF78F45B68010482415B47",
INIT_29 => X"4515549003FFC7BE8002155BEF5EDB6DAADF470280075FFF45E3F1C7038A2DB6",
INIT_2A => X"038F450075C71FF087BD75D7FF84050BAEB8428BEFBEA4BDE28140A154380051",
INIT_2B => X"0A175C7005B6DB55145140000FFAE85082417FFFF7DE3F1EFA10140407000140",
INIT_2C => X"00000000000000000000000000005B7DEAA0824851EFEBFBD2410EBD168B7D41",
INIT_2D => X"0004175FFF7803DF45FFAE955EFAAFBD55EF557BC20AA5D00000000000000000",
INIT_2E => X"0AAD17DFEF007FC20AA5D043FE00F7D17FEBAA2D5574BAAAD17DFEFA2AEAAB55",
INIT_2F => X"45F78402010007BD5545AAFFD55EFF7FBE8B55007FD75FFF7D5401EF5D2E9741",
INIT_30 => X"F45A2D5554AAA2FBEAAAAFFD555545FF8015555007FD5545550400145FFFBEAB",
INIT_31 => X"DEAA5D2E974AA00515754500003FF55FF8002155FFD17FFFFA2FBD74BA00557F",
INIT_32 => X"7FE105D04174105D042AB550055555FF007BD7555F784174AAA2842ABEFFF803",
INIT_33 => X"BC2000AAD16ABFF002A97545007FFFF45555540000FFAE97410007BFFFFFA2D5",
INIT_34 => X"0000000000000000000000000000000000000000000007FFDEAA0004175FFA2F",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000040000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(11),        -- Port A data input
DOA(0)   => data_read_a_hi_256(11),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(11),        -- Port B data input
DOB(0)   => data_read_b_hi_256(11),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_12_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50080B01BC002006940202C0DE041196A83183000000023322287E0FC000006",
INIT_01 => X"0E000C048000C048400380000007026040000000080000088200002802153231",
INIT_02 => X"2809AD0E7D180040945008040090000061800000C0E2F66009DA3D11CB148015",
INIT_03 => X"210D050012F6F8D2108216E24842005B8A20640008800000B8E0141C28851006",
INIT_04 => X"0080100022408000060DE0000066630C70241827041000040800820480001AA4",
INIT_05 => X"0240000C400000003C808003E0C8001401000000040900020904004000070800",
INIT_06 => X"00300D800C1960C4400006E10B90002018184000100804005784000130821200",
INIT_07 => X"0652428112180C03E8E5A2C800A3F018200418927E06686450FF8006460003A0",
INIT_08 => X"09840903525281D4F460409000000E3F08D1202C5C26A0719CC96CC7BF462990",
INIT_09 => X"82488BAE10000040000410802008600843001E09F00000276F81020000230280",
INIT_0A => X"00000080000C000C100204593F11A489F480067D04D40C012400080000800240",
INIT_0B => X"0800021826933E03662802B300003C13E0000000460000000000010CE0000000",
INIT_0C => X"78419784197861978419784197860CBC30CBC20000000010400808056500A080",
INIT_0D => X"201E7F3F01F40401C17E800C7F33800200000357008C0249E2DE0D7841978619",
INIT_0E => X"0F500002200004005002001408400000000000000000000053A4096F80705FA0",
INIT_0F => X"1B17B2C53F2FC16691DB587201EDDF4162B1DB527201EDDC4607024100100020",
INIT_10 => X"F2A01D5CC9794162B1DB587201EDDF416691DB527201EDDD884272592D6246FC",
INIT_11 => X"7258E995D5A825DBA569F9FF02547068618CD3CC45B7863AE7EC00D4B122A67D",
INIT_12 => X"C6CCA5C33717461C045B5B182019473D19D7CCD856106F31A683621BDFC28800",
INIT_13 => X"FB10A652CC8E3538BBA01624E51AA6C0469AC5493F5688532966471A9C5F6208",
INIT_14 => X"40041E1F5759001B4AA1853E6D5144AA9C914C8608D2724A4C4118D992B866E2",
INIT_15 => X"AD9825682D4A36C0B0B4B85112B2C4A05D3E6D5051893335EB0072AA85A4F9B7",
INIT_16 => X"000008000000821000048260020000004001DC0800000010E7F70171401DE07E",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0100401004010040100400000000000000000000000000000000000000000000",
INIT_19 => X"1080800000000000000000040100401004010040100401004010040100401004",
INIT_1A => X"249249249120780800016A28A288028DCA30444409B054A88C5890486582A210",
INIT_1B => X"86432190C86432190C8641041041041041041041041041041041041041049249",
INIT_1C => X"FBC007592C964B2592C964B2592C964B2592C964B2592C964B2592C964B2592C",
INIT_1D => X"FF55002ABEF0800000000000000000000000000000000000000000000000401F",
INIT_1E => X"BEFA280155EFFFFBC01EF0855400005555421FF00042ABEFFF8400010082EAAB",
INIT_1F => X"FFEF08556AA10000028AAAFFD15541000002ABEFFFFBD54000004155EFAA842A",
INIT_20 => X"001FF00041554555557FE005D003FE10AAFBE8AAAA2D540000F7D57DF55A2AAB",
INIT_21 => X"1575FFA2FFD75FF550015400FFFBFFF45085140000005168AAA087BFFFFF5D04",
INIT_22 => X"D5421EFA2FFFFF555D0000145082E955FF0851555FF082AA8B55F7AEA8BEF555",
INIT_23 => X"000020BAAA801541055042ABEFFFFBD5410AAD57DF45A280154BA5555401EFFF",
INIT_24 => X"000000000005568AAAAAD142145FF80155EF0051555FF0804155FFF7842AA100",
INIT_25 => X"7EB80000280824ADBD7490E28BEF080000000000000000000000000000000000",
INIT_26 => X"101C00175EFB6802DBC7BE8A155EFE3FBC71FF145B42038555F401D71C0A2DBC",
INIT_27 => X"038EBD57DF7DA2AEB8FC7005F6AA381C0A2DA82FFDB5243800002FBD7EBFBD24",
INIT_28 => X"AA82147FF8FEF410E001FF000E17555555B7AE1041003DE10BEF5EDAAAAAD547",
INIT_29 => X"ADB45F7AEA8BEF555F575FFBEF5D05EF550E15400E3F1FFF7D085B420381C5B6",
INIT_2A => X"010482415B471C7E3DF451EFBEFBFAF4549000017D142E905EF1451525C7082A",
INIT_2B => X"04105C7F7842FA381C0A00082AA8A1041041002FBEFEBFBD2410AADF78F45B68",
INIT_2C => X"00000000000000000000000000005B68ABAB6D145145FF84155D7085B555C714",
INIT_2D => X"5D7BC01555D2EBFF55A284000AA08003FF55002AA8BEF0000000000000000000",
INIT_2E => X"A08003FF55A2FBC00105D04175FFF7803DF45FFAE955EFAAFBD55EF557BC20AA",
INIT_2F => X"00F7D17FEBAA2D5574BAAAD17DFEFA2AEAAB55007BE8AAA5D2EBDE00FFFFC00A",
INIT_30 => X"FEF007FC20AA5D7BE8A005D7FEABFF002E821FF082A97555557FE8A0000043FE",
INIT_31 => X"01EF5D5142145082EBFF55F7AAAABEF5D7FD75FFF7D5401EF5D2E97410AAD17D",
INIT_32 => X"C2010A2FBEAB45F78402010007BD5545AAFFD55EFF7FBE8B550004001FF5D2A8",
INIT_33 => X"015555007FD5545550400145FF843DEAA552A82010A2AA8000008043FFFFA2FB",
INIT_34 => X"0000000000000000000000000000000000000000000007BEAAAAFFD555545FF8",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000007FFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(12),        -- Port A data input
DOA(0)   => data_read_a_hi_256(12),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(12),        -- Port B data input
DOB(0)   => data_read_b_hi_256(12),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_13_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10110A0441812402840402822007818000E00700000000330A3000000008042",
INIT_01 => X"A1400984B830C848180260000C0042404001000008220008A200100802110200",
INIT_02 => X"88010C02801040002475580400800000410000000064024608134C0CC9018034",
INIT_03 => X"00010100926220D084234212421085084300648A0880000630C0654288C10000",
INIT_04 => X"0004122122029100100C00001200009C40A83A2044360C84190BAC04E0101820",
INIT_05 => X"027000004009050064C8C00104C10184034010250089C00EB004327064B60900",
INIT_06 => X"543000004080480492A946CE1032002012125804440812541027008230821380",
INIT_07 => X"0A581424525408000AE2AA8002BC00D020003896020658FC4030000246E543AE",
INIT_08 => X"04840101107200B80040210000002ABF02450A264002C8008000441680041900",
INIT_09 => X"825A98801000008001041080200B660E30B200C8840080808065102000280280",
INIT_0A => X"00000080C90391881000145B0111A30404016003A56008012C80080200801280",
INIT_0B => X"08088C5D2288004120E80290882400908000A000A1000809A93485D610000000",
INIT_0C => X"002000000000000002000000000000001000000000000000400808154100A080",
INIT_0D => X"08000000360401021280800E400B800610C84100014224200000000020000000",
INIT_0E => X"0086000600040D045E4195104D5854284A14250A12A512A8808289840084A020",
INIT_0F => X"0949E07A80948354B6E68982167061037496E683821670620681024000000000",
INIT_10 => X"8E510B456587037496E689821670610354B6E6838216706220431961CA985D48",
INIT_11 => X"196186A91674011CE61403562274AA49CD594CF00039C7C414B6509DA2265213",
INIT_12 => X"A983014780CC8604040424A5323845932E620295879818170304B2F5002C2043",
INIT_13 => X"451654B9104A328665603148895D44E0251142B42A3D8B2A5C8825194328A2E6",
INIT_14 => X"C06A6C6A465AA0091482382B17614F2202858EE300991415B45CD5306028F019",
INIT_15 => X"52E08DC8047F17D1C7C3C02128E587D6A02B17605A130A4E8BF002258850AC5D",
INIT_16 => X"84A123508508220808048240604B2100C00022084809000D000393722A140000",
INIT_17 => X"4A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A12",
INIT_18 => X"A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A128",
INIT_19 => X"154000000000000000000284A1284A1284A1284A1284A1284A1284A1284A1284",
INIT_1A => X"BAEBAEBAEBFF6FEFEFEEEAAAAAAFBF7DDF77F9FBEFBFF9F3F0FDFCFBEFBF1228",
INIT_1B => X"5FAFD7EBF5FAFD7EBF5FAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAE",
INIT_1C => X"F800077EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF",
INIT_1D => X"00FFD140155F780000000000000000000000000000000000000000000000401F",
INIT_1E => X"BEFFF8400010082EAABFF55002ABEF08556AAAA5D043FFFFAAAABDEAA557BFDE",
INIT_1F => X"000055043DEBAF7843FFFFF7AABDF55A2AA97400AAD540155A2D5421FF00042A",
INIT_20 => X"E8B45557FD7410552EAAABAAA84155EFAA842ABEFA280155EFFFFBC01EF08554",
INIT_21 => X"56AA10000028AAAFFD15541000002ABEFFFFBD5400005568A1055043DEBAAAFF",
INIT_22 => X"D57DF55A2AABFFEF085557545FFD17DEBAA2FFE8ABAAA8428A00087BD7555FFD",
INIT_23 => X"57BEAABA5D2ABDF450851420AA5D7FD5555A2803FE10AAFBE8AAAA2D540000F7",
INIT_24 => X"000000000005168AAA087BFFFFF5D04001FF00041554555557FE005D00001555",
INIT_25 => X"7AAA4B8E824971F8E38E3DF45155EB8000000000000000000000000000000000",
INIT_26 => X"55A2DF401D71C0A2DBC7EB80000280824ADBD7490E28BEF08516DA82410A3FFD",
INIT_27 => X"5EFE3FBC71FF145B42038550E38E92EB803FFD7EBA4BDF45AAAA90410BEDF451",
INIT_28 => X"FA38490A3FE92BEFFEAB45417FD24385D2AAFA82B680175EFB6802DBC7BE8A15",
INIT_29 => X"28A10007FD557DFFDF6AA381C0A2DA82FFDB5243800002FBD7EBFBD24101C556",
INIT_2A => X"5EDAAAAAD547038EBD57DF7DA2AEB8FC700515056DE3D17FE92BEF1EFA92AA84",
INIT_2B => X"5B7AE10410E00155497FEFABA4120B8F55085B400925D7FD557DA2803DE10BEF",
INIT_2C => X"00000000000000000000000000005B6AA82147FF8FEF410E001FF000E1755555",
INIT_2D => X"00517FE00082EBDF45AA8428A10085568ABAA2FBD7545AA80000000000000000",
INIT_2E => X"5AAAE82000F7FBD5545AAFBC01555D2EBFF55A284000AA08003FF55002AA8BEF",
INIT_2F => X"FFF7803DF45FFAE955EFAAFBD55EF557BC20AA5D2EA8A00A2803DF45AA843DF5",
INIT_30 => X"F55A2FBC00105D517FEAA082EBFE10F7FFE8B55087FC00BA552ABFE10F784175",
INIT_31 => X"FE10F7D57DE00AA842AA00007FD75FFF7FBE8AAA5D2EBDE00FFFFC00AA08003F",
INIT_32 => X"D55FFAA843FE00F7D17FEBAA2D5574BAAAD17DFEFA2AEAAB550051401FFA2D57",
INIT_33 => X"E821FF082A97555557FE8A00002E82155007BFDEAA08042AB45087FC0010557F",
INIT_34 => X"0000000000000000000000000000000000000000000007BE8A005D7FEABFF002",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000067FFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(13),        -- Port A data input
DOA(0)   => data_read_a_hi_256(13),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(13),        -- Port B data input
DOB(0)   => data_read_b_hi_256(13),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_14_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10020A000180000284008280000281800000030000000033022000000580002",
INIT_01 => X"A140098018300848184860000C20C24040000000084000084200000000110200",
INIT_02 => X"88010C5A8010A600A4F558040080000041000000022C024008003CCCC9028030",
INIT_03 => X"000103A7A00904D0842242024210810803006480088000003081054288C10000",
INIT_04 => X"0000120122009000100C00000000000400A83A2044200C840000800400101820",
INIT_05 => X"020000004008010024C0C0010040000402000025000800020004207000100800",
INIT_06 => X"0430000040004804920906C20022002012120004440812541020008230821000",
INIT_07 => X"2A5A14285A15080008768A80008000D0200018B202067AF100A0000244204382",
INIT_08 => X"04850101105205380040000000000A7F42840A264920406080004400A0040900",
INIT_09 => X"8208888010000080010010802000400230B000C8840080800021100000200280",
INIT_0A => X"00000080C8038188100004590111B68404012000016008012000000000000200",
INIT_0B => X"080084452280004120400000802000908000800001000009A924810410000000",
INIT_0C => X"000000000000200000000000000200000000000000000000400808000000A080",
INIT_0D => X"080000002204010010808008000B800210404100000220200000000020000200",
INIT_0E => X"0000000600000000020181100400502048102408122412808082098400042020",
INIT_0F => X"0480040A100A42008000161C140000420080001C1C1400003201024000000000",
INIT_10 => X"39600022260042001000161C140000420010001C1C140001604E8084341CBA34",
INIT_11 => X"8082580E2B8802201014800C220A21829A302F1C024010C001124020C8C1A8A0",
INIT_12 => X"CA60CA000048228404401004418012787124648157780120B8678C000801E04E",
INIT_13 => X"001072D04730000241000CB1325E78E0186030240000083B602398000120024A",
INIT_14 => X"001EF6F4163C480481506800004000CFD55196CB012481812049495C19400009",
INIT_15 => X"248800108B8FB61A0401200845594965000000400568D0CFB780055060500001",
INIT_16 => X"048123408408220000048240604B210040000008400800B0000090022A140068",
INIT_17 => X"4812048120481204812048120481204812048120481204812048120481204812",
INIT_18 => X"8120481204812048120481204812048120481204812048120481204812048120",
INIT_19 => X"1400000000000000000002048120481204812048120481204812048120481204",
INIT_1A => X"9E79E79E79FF3BEEEEEFE79E79EFAABCDA72E47F87BDF4EBAE7CFAFBEFB28200",
INIT_1B => X"CFE7F3F9FCFE7F3F9FCFE79E79E79E79E79E79E79E79E79E79E79E79E79E79E7",
INIT_1C => X"FBFFF83F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9F",
INIT_1D => X"555D5568A105D00000000000000000000000000000000000000000000000401F",
INIT_1E => X"FFFAAAABDEAA557BFDE00FFD140155F7D17DF45AAD157400007BEAAAAAAAE955",
INIT_1F => X"ABEF085155400FFD1420100055574AAA2AA800AAF784020AAF7D56AAAA5D043F",
INIT_20 => X"FFE105D7BD7545A284020BA0055421FF00042ABEFFF8400010082EAABFF55002",
INIT_21 => X"43DEBAF7843FFFFF7AABDF55A2AA97400AAD540155A28028B550051574005D7F",
INIT_22 => X"FBC01EF08554000055002AB455D51420100851421FF5D7FFDEBA085168B45FF8",
INIT_23 => X"AD140000002EBFFEFA2AAA8BEFF780021FF5504155EFAA842ABEFA280155EFFF",
INIT_24 => X"000000000005568A1055043DEBAAAFFE8B45557FD7410552EAAABAAA8017400A",
INIT_25 => X"01C71EDA82AAA0955455D556DA00490000000000000000000000000000000000",
INIT_26 => X"BAEBD16DA82410A3FFD7AAA4B8E824971F8E38E3DF45155EBD17FF6DAADB5040",
INIT_27 => X"0280824ADBD7490E28BEF085157428FFDB420101C55554AAAAA480082FF84000",
INIT_28 => X"AB7D0051504005D71F8E004975D556DB68405092085F401D71C0A2DBC7EB8000",
INIT_29 => X"FAEAA08516AB45E38E38E92EB803FFD7EBA4BDF45AAAA90410BEDF45155A28E2",
INIT_2A => X"02DBC7BE8A155EFE3FBC71FF145B42038550028B6D5D51420101C5B401EF417B",
INIT_2B => X"2AAFA82B68015400AADB40000082EBFFC7A2AEAFBC7EB80071FF5500175EFB68",
INIT_2C => X"0000000000000000000000000000556FA38490A3FE92BEFFEAB45417FD24385D",
INIT_2D => X"AAD17DFFFAAFFC200055557DE00A2801554555557FE100000000000000000000",
INIT_2E => X"AA28400000F784020BAAAD17FE00082EBDF45AA8428A10085568ABAA2FBD7545",
INIT_2F => X"555D2EBFF55A284000AA08003FF55002AA8BEF0051554AAFFFFC00105D55554B",
INIT_30 => X"000F7FBD5545AAAEAABFF0051400105D5568A000051575FFF78415410087BC01",
INIT_31 => X"2000557FC01EF007FEAABA00556AB55A2AEA8A00A2803DF45AA843DF55AAAE82",
INIT_32 => X"175FF5D04175FFF7803DF45FFAE955EFAAFBD55EF557BC20AA5D042ABFF55514",
INIT_33 => X"FE8B55087FC00BA552ABFE10F78415400A2FBC0010082EBDF55A2AABDF45A284",
INIT_34 => X"000000000000000000000000000000000000000000000517FEAA082EBFE10F7F",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000007FFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(14),        -- Port A data input
DOA(0)   => data_read_a_hi_256(14),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(14),        -- Port B data input
DOB(0)   => data_read_b_hi_256(14),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_15_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000A000000000284000280000001800020030000000033022000000180002",
INIT_01 => X"A140098018300848180060000C00424040000000080000080200000000110200",
INIT_02 => X"080108000010E60004E55800008000004100000000040240080000C009170016",
INIT_03 => X"0000000080000040842240000210810002000400888000003080014288C00000",
INIT_04 => X"0001100024A0800000440000000000040088322044200C840000011400151800",
INIT_05 => X"A200014C4000000020000000000B8094020000254C8800000514203000108800",
INIT_06 => X"0031042040804804100006EE4032002012120005540812540020008600831000",
INIT_07 => X"021912244A14080008408880008000D020001892020656300020000244000380",
INIT_08 => X"048501415032000800406180000002DF02440826400000008000440000043080",
INIT_09 => X"8208880110000000010010802000400230A000880400808000450200000B0280",
INIT_0A => X"00000080C003010810000459011182040400200003E0080120000000000002C0",
INIT_0B => X"080084452280004100400000800000100000800001000001A124800010000000",
INIT_0C => X"002000020000000000000000000200001000010000000000400808000020A000",
INIT_0D => X"08000000260001001280000C400B000200000000000220200000000020000200",
INIT_0E => X"008400060000000000010010040040000000000000201000000000000004A000",
INIT_0F => X"0000000000000202100000000000000202100000000000004600024000000000",
INIT_10 => X"0000000000000202800000000000000202800000000000002000000800000000",
INIT_11 => X"0008000000000000000000002000100800000000000000000000400001200000",
INIT_12 => X"00880000000006000400080C0000000000D08120280000000000000000002000",
INIT_13 => X"0010040200000000010000004020010000000000000008000900000000000200",
INIT_14 => X"0000000308801400000000000040000008822110000000000040100100000000",
INIT_15 => X"0080000000004840717050000000000000000040000020000000000000000001",
INIT_16 => X"000023000000220000048240404A010040000008000000000000000020C40000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"1400000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000200",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"F800000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"AA007BC2145F780000000000000000000000000000000000000000000000401F",
INIT_1E => X"400007BEAAAAAAAE955555D5568A105D7FC00000804154AA5D00001EFF78428A",
INIT_1F => X"0155F7FBD74AAAAD17DF45F7D1421EF0055400AA007FC2000F7D17DF45AAD157",
INIT_20 => X"BDFEF08517DF55A2FBEAB555D556AAAA5D043FFFFAAAABDEAA557BFDE00FFD14",
INIT_21 => X"155400FFD1420100055574AAA2AA800AAF784020AAF7FFFDF45FF84000BA552A",
INIT_22 => X"2EAABFF55002ABEF087BE8ABA555168B55AAFFEAB45F7843FF45082A801FF005",
INIT_23 => X"284000AA0055401550055574005D2E800AAA2D5421FF00042ABEFFF840001008",
INIT_24 => X"000000000000028B550051574005D7FFFE105D7BD7545A284020BA007FFFE10A",
INIT_25 => X"2550E021C7EB8028A821C7BC516DFF8000000000000000000000000000000000",
INIT_26 => X"28FFD17FF6DAADB504001C71EDA82AAA0955455D556DA004971C703814001248",
INIT_27 => X"E824971F8E38E3DF45155EBF1D5492BED17FF45E3DF471C70851400BA0071C50",
INIT_28 => X"FF7DEB8000092552ABFFEF08517DF6DB6FBE8B555D516DA82410A3FFD7AAA4B8",
INIT_29 => X"3DF551C20801C71C5157428FFDB420101C55554AAAAA480082FF84000BAEBF1F",
INIT_2A => X"A2DBC7EB80000280824ADBD7490E28BEF087FEFA8241516DB55A2FFEAB6DEB84",
INIT_2B => X"8405092087FF8E00BE8A02082005F47145085550428412A85082BEDF401D71C0",
INIT_2C => X"00000000000000000000000000000E2AB7D0051504005D71F8E004975D556DB6",
INIT_2D => X"0055554BA5504000105D2A80145AA842AA00557BD75EFF780000000000000000",
INIT_2E => X"50055420BA0055574BAF7D17DFFFAAFFC200055557DE00A2801554555557FE10",
INIT_2F => X"00082EBDF45AA8428A10085568ABAA2FBD7545AAD557410F7D57DF55AAFBD554",
INIT_30 => X"000F784020BAAAD57FFEFA28402010552ABDFFF08517FFFFF7FBEAB455D517FE",
INIT_31 => X"DF45AAFBE8BEFA2803FF455504001555551554AAFFFFC00105D55554BAA28400",
INIT_32 => X"95400F7FBC01555D2EBFF55A284000AA08003FF55002AA8BEF007FFDE1000557",
INIT_33 => X"568A000051575FFF78415410087FEAA10F7AE80000087BD55450855400BA002A",
INIT_34 => X"0000000000000000000000000000000000000000000002EAABFF0051400105D5",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000060000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(15),        -- Port A data input
DOA(0)   => data_read_a_hi_256(15),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(15),        -- Port B data input
DOB(0)   => data_read_b_hi_256(15),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_16_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"DA22C618B1000482B688B186588884862A400438255FC38381441205BA803003",
INIT_01 => X"8645A80028404C211203A952A90341080B173340412000E1005D628000820484",
INIT_02 => X"A101A9006DC1084833011850AAC55001349B10881802821808B4110007005E11",
INIT_03 => X"010108A802BB00080080006020020001A61036202800000D2410104200404550",
INIT_04 => X"8BFA58800005C40A46240252145148B38248030356415A4E62B6FC660F287240",
INIT_05 => X"0F05EA11E570000D610000000710296E542B6E3A825C15FB30A643695BFC2D56",
INIT_06 => X"00640044150C025A0000000901A054F2C0A8030140BCC0460050690A95C8383D",
INIT_07 => X"0288500102F85203E8010D0AA9BC4800015001219D0550077373CAA804000680",
INIT_08 => X"A2064193920A2004B51400001414091EAA14881C0002701881B120203B7A8012",
INIT_09 => X"C8204D02D965965200100104F2B0082251200000023153000C4400800000ACCA",
INIT_0A => X"000012C9000A0000D0A80000BF8028E87C1B9246002A8A562060410280081116",
INIT_0B => X"240014891801000495D40192D1000000000000A8A5AA80018120E00066000000",
INIT_0C => X"00088000880008800088000880008400044000400029011404008401CA809004",
INIT_0D => X"0140A80A5C8000102ED0044008004AD32400004001AB08C0031EDA7B08800088",
INIT_0E => X"04912AA28AA890BA00000024800480000000000000200802151025062C0BB400",
INIT_0F => X"1F554E11C596A64003195933741477264003195555B418687E35836020814004",
INIT_10 => X"0A499CF47DCB264003195933741597264003195555B4198843940076D296D003",
INIT_11 => X"00758486A556489347FE5F409CBC1362510695B6288743123C95251852041CD5",
INIT_12 => X"424EAE2992046EB70026486035600CEC45CBCA809654B48163CCC895E1E043D4",
INIT_13 => X"98E3A242DEA151848302BFD6D522B10C7EC71F6C1DB071D1216E078C4C1B1C74",
INIT_14 => X"037DAAABC982BE22267A2E2E4F44AA1DC5E37400C9EE1B7B638E8849D23C3832",
INIT_15 => X"2EE015998B28654565A003F0068E35352C1CAE48BFBF3A6C9B7B286B4DA8B93D",
INIT_16 => X"000009000040A8000452110A8442040D655602A102A0027E2C42320284086E6A",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"1451451451E96F2FC3C34F3CF3C2AC688AA263486D3260E34C0C3A7B451B0200",
INIT_1B => X"9F47A7D1E9F47A7D1E9F4D14D14D14D14D14D14D14D14D14D14D14D14D145145",
INIT_1C => X"F800007D3E9F4FA7D3E8F47A3D1E8F47A3D1E8F47A7D3E9F4FA7D3E9F4FA7D3E",
INIT_1D => X"FF00003FE005500000000000000000000000000000000000000000000000401F",
INIT_1E => X"4AA5D00001EFF78428AAA007BC2145F7843FFFFF7FBE8B45AAD568BFFFFAA975",
INIT_1F => X"8A105D2E974BAF7FBEAB45FFFFC00BAF780020005D2A95410FFFFC0000080415",
INIT_20 => X"821FFA2AAAAA00000417555FFD17DF45AAD157400007BEAAAAAAAE955555D556",
INIT_21 => X"BD74AAAAD17DF45F7D1421EF0055400AA007FC2000F78000010552E800AA002E",
INIT_22 => X"7BFDE00FFD140155F7AABDF55F7AE820AA08043FEBA5D55575FFF7AABFE00557",
INIT_23 => X"2FBE8B55FFFFD55FF557FC2000FF8015410FFD56AAAA5D043FFFFAAAABDEAA55",
INIT_24 => X"000000000007FFDF45FF84000BA552ABDFEF08517DF55A2FBEAB555D04154BAA",
INIT_25 => X"5B6DF6DBFFF7AA955C71C043FE10490000000000000000000000000000000000",
INIT_26 => X"38FFF1C7038140012482550E021C7EB8028A821C7BC516DFF8438FC7E3F1EAB5",
INIT_27 => X"A82AAA0955455D556DA00492490492F7FBE8B55FFF1C70BAF78A000005D20974",
INIT_28 => X"20285D2085092002A801FFB6AAA8A10080E1757DEBD17FF6DAADB504001C71ED",
INIT_29 => X"555FFE3AABFE005D71D5492BED17FF45E3DF471C70851400BA0071C5028FF840",
INIT_2A => X"A3FFD7AAA4B8E824971F8E38E3DF45155EBA4BAF6DE3AA8709208043FEBA555B",
INIT_2B => X"FBE8B555D04124BAB6FBE8B45E3FBD55D7557BC0028E38412428EBD16DA82410",
INIT_2C => X"000000000000000000000000000071FFF7DEB8000092552ABFFEF08517DF6DB6",
INIT_2D => X"F78428B55AAD168B55F7FFFDFEFFFAA9555555003DE000000000000000000000",
INIT_2E => X"AFFAE820105500154AAF7D5554BA5504000105D2A80145AA842AA00557BD75EF",
INIT_2F => X"FFAAFFC200055557DE00A2801554555557FE10000000010F7FBEAB45FFD1554A",
INIT_30 => X"0BA0055574BAF784000BA5D0017410082E801EFF7AEA8A10002E955FFA2D17DF",
INIT_31 => X"541000003DEBA557BD75EFA2AEBDE105D5557410F7D57DF55AAFBD5545005542",
INIT_32 => X"000AAAAD17FE00082EBDF45AA8428A10085568ABAA2FBD7545AA802ABEFA2AA9",
INIT_33 => X"ABDFFF08517FFFFF7FBEAB455D04020AAFFFBEAB45AAFFD55555D7FC20AAA280",
INIT_34 => X"000000000000000000000000000000000000000000000557FFEFA28402010552",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000020000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(16),        -- Port A data input
DOA(0)   => data_read_a_hi_256(16),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(16),        -- Port B data input
DOB(0)   => data_read_b_hi_256(16),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_17_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"5284CE4FB7BD2C8994A13392DBD02E14006B82AC7E800D44D3DD2FD5F9B961C0",
INIT_01 => X"F8ACD01F7E03FC6793F2199B39FC233C11D93AE6F3BB92B32091DBC339B24542",
INIT_02 => X"8F333007FD6808092A2AFA6667033DB50853379C10BFF70F1BD011110F205F18",
INIT_03 => X"294ADB4AFFCBF0DAD63ABF836B58EAFE060478202022234B2E0303FDC9E18339",
INIT_04 => X"DB7A40806FE4040840EBC563A0150A0926146FECB04196482236FC2005282AE1",
INIT_05 => X"0403DA0383200831C68206D7E6D0250834336D1E81500FDB306045255BFC2076",
INIT_06 => X"000A0E2D7D3EAFF15800100FBFB333C1CBC303163670497AFF00291B3C0E2015",
INIT_07 => X"451C581123AEE54DE8008B719E61C10BBA5DAAFA9DDA1194D51E067BB0000000",
INIT_08 => X"70320A9392083056C2270E004400091181168C4D14002A110C902481FC0B4212",
INIT_09 => X"0E28EFFC40C30E5F0182D0950190C0810BE00E9A76E4C7FD0E4700000B303806",
INIT_0A => X"C7DEF207000F00059D2ED56D7EED2ED3C9A86FB8013E7437823DF78CDB6CA60E",
INIT_0B => X"7C00319F8E853E64D73A08BFF0001D35682AC0CE8FCCC200A59BDD2FFE3F3EC7",
INIT_0C => X"7A7DE7A7DE7A7DE7A7DE7A7DE7A7DF3D3EF3D3C0030B889723782E816EC0A081",
INIT_0D => X"2D4CFEB69FF7A5F5AFFCCA787F7FE67C21800367451F8355EB9EDE7A7DE7A7DE",
INIT_0E => X"2C9F99FD0678B87A0003000D8D02E00000000000000040025D3C21463D6BFF25",
INIT_0F => X"232221ABD9CA854DFDD64A67D42C0F054DFDD64667D42C063E57A8F7B4594BB0",
INIT_10 => X"AEDAA504801F054DFDD64A67D42C0F054DFDD64667D42C07237DFE5865F6D2BF",
INIT_11 => X"FE58EAE7F5AB50D0806A9A2E0DFFF47DEDC496DA3181A0CC71440F9FBC3EFBB5",
INIT_12 => X"9C9C3FC95949AEFF556EF9C75E7DCF1EB1B6E6FCDC87CB35FC94B36AECF3A33D",
INIT_13 => X"382AF5B6AAAE594A4C0DBFDAD94AA669809809FEFAF4157ADB55572CA527056E",
INIT_14 => X"1AE33F32ADD543430808BABAF50E1A5EB4BAEA45A250202FE0ADD39387F92B29",
INIT_15 => X"669523E865D4B1293AB6B90BF2F0E30EDEFAFD0B3FBD72E9E90D20A003FBEBF4",
INIT_16 => X"00002F840000BCE0B6F67B3F845E017C833F6AAC02B002A2EFF22D4073DE83FB",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0600000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"9A69A69A6A4624C3434C0EBAEBA21B9001804F6E62029749701020B88A7CC0C0",
INIT_1B => X"41A0D46A341A0D46A341A69AEBA69A69AEBA69AEBA69A69AEBA69AEBA69A69A6",
INIT_1C => X"F8000046A351A8D46A351A8D46A351A8D46A351A8D068341A0D068341A0D0683",
INIT_1D => X"00F7D56ABFF55000000000000000000000000000000000000000000000007FFF",
INIT_1E => X"B45AAD568BFFFFAA975FF00003FE0055043FFFFFFFFFFFFFF7FBFDF55A284020",
INIT_1F => X"2145F7D568B45000002010552EBDF45A28028A00F7843FEBA55043FFFFF7FBE8",
INIT_20 => X"95410AAAEBFF55AAFFC00BAF7FFC00000804154AA5D00001EFF78428AAA007BC",
INIT_21 => X"E974BAF7FBEAB45FFFFC00BAF780020005D2A95410FFAE800105D2A95410002A",
INIT_22 => X"AE955555D5568A105D7FFFFEFA2D568BFFFFD57DE00F7AE800AAAAAABDFEF5D2",
INIT_23 => X"82A974105D003FF55F7802AAAAAAD168AAA5D517DF45AAD157400007BEAAAAAA",
INIT_24 => X"000000000000000010552E800AA002E821FFA2AAAAA00000417555FF8028B550",
INIT_25 => X"FE3F5FAF45AA8000038F7DB6FBD7490000000000000000000000000000000000",
INIT_26 => X"82490438FC7E3F1EAB55B6DF6DBFFF7AA955C71C043FE10490A3FFFFFFFFFDFE",
INIT_27 => X"1C7EB8028A821C7BC516DFFDF68B551C0E050384124BFF7DB68A28A38F7803DE",
INIT_28 => X"5000492495428082E95400AAA0BDF7DB6F5C70BAFFF1C7038140012482550E02",
INIT_29 => X"800BAB6AEBDFD75D2490492F7FBE8B55FFF1C70BAF78A000005D2097438FFAA8",
INIT_2A => X"B504001C71EDA82AAA0955455D556DA00497FFAFFFB6D56FBFFEBDB78E38F7AA",
INIT_2B => X"0E1757DEB8A2DB5514249243841003FF6DEB8028AAAB6D16FA8249517FF6DAAD",
INIT_2C => X"000000000000000000000000000004020285D2085092002A801FFB6AAA8A1008",
INIT_2D => X"002ABFFEFF7FBFDFFFAAD168B55AA80000BAF7FFFDF550000000000000000000",
INIT_2E => X"FFFAAA8AAAF7843FE10000428B55AAD168B55F7FFFDFEFFFAA9555555003DE00",
INIT_2F => X"BA5504000105D2A80145AA842AA00557BD75EFF7FBEAB45552E954BA08003DFF",
INIT_30 => X"0105500154AAF7AE974000800154AA002E95410AA843FFFFF7D5554BAF7D5554",
INIT_31 => X"FFEFAAFFE8ABAFFAA820BAF7AEBFF55550000010F7FBEAB45FFD1554AAFFAE82",
INIT_32 => X"7DE0000517DFFFAAFFC200055557DE00A2801554555557FE10007FEABEFFFD57",
INIT_33 => X"E801EFF7AEA8A10002E955FFA2AABFF455500020AA08003DFFFA28028AAAF7D1",
INIT_34 => X"00000000000000000000000000000000000000000000004000BA5D0017410082",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000067FFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(17),        -- Port A data input
DOA(0)   => data_read_a_hi_256(17),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(17),        -- Port B data input
DOB(0)   => data_read_b_hi_256(17),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_18_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"69844019080000A21A611406840014122A641074155FC28A2024001001801003",
INIT_01 => X"A643D920034004180005E9E3C90360C0041C0181002001602025800008440084",
INIT_02 => X"B7333980808408103F2000F81FC0FEDEAC2161B0B84D0002188011110C018041",
INIT_03 => X"0405D434003F2C020081587008020561E55116B0290000042B71240C800440F8",
INIT_04 => X"50805AC31007D6125724029216554A9847669903D640EC8E2001002604503004",
INIT_05 => X"07008000E0EA11803850C800010022660C1C0065003C0404002646DC20A02D40",
INIT_06 => X"8560000000022229A60B048048120FF040000000002C44D620F0228454C83810",
INIT_07 => X"058800A001D4033A004904087F9E3901218050018024110D6771C1F90C285682",
INIT_08 => X"F3020A82929A807B3731021400058C020000A9729400D10100420480202AC214",
INIT_09 => X"C820C802D86184A010180304307008025414204400220202F1A814A0080064C1",
INIT_0A => X"080003C32A10A19090C02010E10229440616900000022E0C6070000504102805",
INIT_0B => X"026226495446E2110AE44174112840880000060D7030C30B885200D274004008",
INIT_0C => X"840018400184001840018400184000C2000C200200301500C404C001B884B806",
INIT_0D => X"81010108003C000210020460801001FB3650D89888E06CAE1061018500184001",
INIT_0E => X"032007E281F840C00284A17210001060D8306C18360C1380A0260CB980840080",
INIT_0F => X"5D79BBEF8E50B041029075982BF3873041029079982BF39748AA0AC800014804",
INIT_10 => X"EA479BFD7F7F3041029075982BF3E73041029079982BF3F632C5F96D3C11555D",
INIT_11 => X"F96A595405FC7F1CFEBC7586C4100A53162B47FD7E39FFEECE1598702345156A",
INIT_12 => X"006FE037ACFB88083A99E06271BB0CA207DFDD5920057E0B001B0EBCC79932C5",
INIT_13 => X"5CA2A002DD51B6F7FC4A411D1E8D44517F14EAFE36E55150016EA8DB73E39464",
INIT_14 => X"953C30351452A13D55CFFA76E928E3891F148B30399F5FB7F28C800DFA06F5DF",
INIT_15 => X"5AC57DFEAEF1005475F1D1F608819CF0EE76E12C824ADD9089715F25FAF9DB84",
INIT_16 => X"0D834041A41A0000010180C02801680460FC900052FA10DC0006DA4881C11015",
INIT_17 => X"D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D836",
INIT_18 => X"8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360",
INIT_19 => X"00000000000000000000020D8360D8360D8360D8360D8360D8360D8360D8360D",
INIT_1A => X"8A28A28A2891182C8A82E0820825945DF675C0770B9E11807E54587BEF8B0000",
INIT_1B => X"44A2552A954AA5128944AAAA28A28A28AAAAAAA28A28A28AAAAAAA28A28A28A2",
INIT_1C => X"F80000128944A25128944A25128944A25128944A25128944A25128944A251289",
INIT_1D => X"BA5D04174AA0000000000000000000000000000000000000000000000000401F",
INIT_1E => X"FFFF7FBFDF55A28402000F7D56ABFF55043FFFFFFFFFFFFFFFFFFFFEFF7AE954",
INIT_1F => X"FE0055043FFFFFFFFFDFEFA2D56AB45AA8400145AA801741000043FFFFFFFFFF",
INIT_20 => X"FFFFFFF80021EF0855421EF00043FFFFF7FBE8B45AAD568BFFFFAA975FF00003",
INIT_21 => X"568B45000002010552EBDF45A28028A00F7843FEBA55557FFEFA2D168B55AAFB",
INIT_22 => X"8428AAA007BC2145F7D5400000004020AA5D2A82155F7AEBFEBAFFD56AA00A2D",
INIT_23 => X"82E954BA0004174AAAA8428B45082ABFEBAA2FFC00000804154AA5D00001EFF7",
INIT_24 => X"000000000002E800105D2A95410002A95410AAAEBFF55AAFFC00BAF7AE800100",
INIT_25 => X"FFFFBFDFEFFFAE954AA550415492140000000000000000000000000000000000",
INIT_26 => X"10140A3FFFFFFFFFDFEFE3F5FAF45AA8000038F7DB6FBD7490E3FFFFFFFFFFFF",
INIT_27 => X"BFFF7AA955C71C043FE1049043FFEFE3F1F8FD7AAD16FB6DBE8E00155BE80154",
INIT_28 => X"8FC7AAD56FB6DBEF1FAFD7E384001EF145B471C7140438FC7E3F1EAB55B6DF6D",
INIT_29 => X"BDE92FFD56FA28B6DF68B551C0E050384124BFF7DB68A28A38F7803DE82495B7",
INIT_2A => X"012482550E021C7EB8028A821C7BC516DFFD1420381C0A02082492A85155E3A4",
INIT_2B => X"F5C70BAFFAE870280024904BA1400174AABE8E28B7D1420BDEAAA2F1C7038140",
INIT_2C => X"00000000000000000000000000002A85000492495428082E95400AAA0BDF7DB6",
INIT_2D => X"002ABFFFFFFFFFFFEFF7FBFDFFFF7AA974BA5504154105500000000000000000",
INIT_2E => X"FF7AA82155F78015400552ABFFEFF7FBFDFFFAAD168B55AA80000BAF7FFFDF55",
INIT_2F => X"55AAD168B55F7FFFDFEFFFAA9555555003DE0000043DFEFA2D56AB45AAD57DFE",
INIT_30 => X"AAAF7843FE10007FEAB55A2D17FFEFFFD568B55A280021EF557FD7555550428B",
INIT_31 => X"2000002A95545A2843FE00F7D17FEAAF7FBEAB45552E954BA08003DFFFFFAAA8",
INIT_32 => X"3DEAAA2D5554BA5504000105D2A80145AA842AA00557BD75EFF7D1400AA5D2A8",
INIT_33 => X"E95410AA843FFFFF7D5554BAF7AE974BA0004020AA5D04154BAF7AEA8BEF5500",
INIT_34 => X"0000000000000000000000000000000000000000000002E974000800154AA002",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000020000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(18),        -- Port A data input
DOA(0)   => data_read_a_hi_256(18),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(18),        -- Port B data input
DOB(0)   => data_read_b_hi_256(18),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_19_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"042200000000000041088001001AA00000000000000000000000500802000003",
INIT_01 => X"200048000024000000000404000000000A22000800000800004A200000000001",
INIT_02 => X"032210008DEF00400060000001C008002489E0F0004037B00010101010000000",
INIT_03 => X"0000008128000000000000000000000024001620280000000000354200004008",
INIT_04 => X"000058800004C4024024001210001054B1C822009640000E2000002604003000",
INIT_05 => X"07008000E0200000000000000000200604000000001C04000026400000002C40",
INIT_06 => X"000000000000000100000000000001B040000000002C42010010200004C83810",
INIT_07 => X"0E0050A040041593104004500480090080A01120220140020420401800000000",
INIT_08 => X"130E409080188000021A0000100004082A140102B4020109801A4CE003710010",
INIT_09 => X"C80000005861840000000004301000B000000000001C1C0000000000000020C0",
INIT_0A => X"000002C30000000040500010301020400000000000022A040000000000000004",
INIT_0B => X"00000020001000022000000000000000000002F0001F00002024B20002000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"00108000EC000000000000000010004B20000000000000000000000000000000",
INIT_0E => X"0000006280180040000000000000000000000000000000000000000000000000",
INIT_0F => X"8084451B81A70AB3006BA0011400760AB3006BA0011400680F02096834820000",
INIT_10 => X"11204082248A0AB3006BA0011400160AB3006BA0011400084C780687DBA82800",
INIT_11 => X"068796E80A00802301BC0A7531EDD98E73B02800804620D030F873EB49F30B80",
INIT_12 => X"6B00000002044F091A860700FF9198AA115D5DA37F7A80C8A3604001C0664C78",
INIT_13 => X"98551AC9000000000314E01F9F30198600631448410A2A8D64800000081B0A93",
INIT_14 => X"2E00303842281C80A23004411AD661891F15148A4420804241526D6000000000",
INIT_15 => X"9D335F3D282000C6C5456C84850F61050C411AD6284FDA861682805A04A1046B",
INIT_16 => X"00000000000000000000000000000004600C0013800003088004202304366A4A",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"86186186186851046260A9A69A6039045DD1F863808633005010063A20C90000",
INIT_1B => X"D26930984C26130984C261861861869A61861861861869A61861861861861861",
INIT_1C => X"F800000984C26130984C26130984C26130984C26130984C26130984C26130984",
INIT_1D => X"BA5500020BA5D00000000000000000000000000000000000000000000000401F",
INIT_1E => X"FFFFFFFFFFEFF7AE954BA5D04174AA007BFFFFFFFFFFFFFFFFFFFFFFFFFAA954",
INIT_1F => X"ABFF557BFFFFFFFFFFFFFFFFFBFDFEFFFAA974BA5D517FFFF08043FFFFFFFFFF",
INIT_20 => X"6AB45AA8002000F7D5575455D043FFFFFFFFFFFFFF7FBFDF55A28402000F7D56",
INIT_21 => X"43FFFFFFFFFDFEFA2D56AB45AA8400145AA8017410007BFFFFFFFFFFFFEFF7D1",
INIT_22 => X"AA975FF00003FE00557BFFFFFFFFBFDF45AAD568B55F7AE955FFAA8402010080",
INIT_23 => X"7D168B55AAD17FFEFF7AE975FF00557FFFF5D043FFFFF7FBE8B45AAD568BFFFF",
INIT_24 => X"00000000000557FFEFA2D168B55AAFBFFFFFFF80021EF0855421EF002ABFFEFF",
INIT_25 => X"FFFFFFFFFFF7AA954BA550000082550000000000000000000000000000000000",
INIT_26 => X"C7080E3FFFFFFFFFFFFFFFFBFDFEFFFAE954AA5504154921471FFFFFFFFFFFFF",
INIT_27 => X"F45AA8000038F7DB6FBD74975FFFFFFFFFFFFEFF7FBFAFD7E3A4954BA555B7AF",
INIT_28 => X"FFFFF7FBF8FC7EBD568B55A28000000FFDF52545550A3FFFFFFFFFDFEFE3F5FA",
INIT_29 => X"955C7BE800000008043FFEFE3F1F8FD7AAD16FB6DBE8E00155BE8015410147FF",
INIT_2A => X"1EAB55B6DF6DBFFF7AA955C71C043FE10497BFDFC7E3F1FAF55A2DB6FB7DF7AE",
INIT_2B => X"5B471C71424B8FC7E3D56AB6DB6DF7AFC7EBA0955FF145B7AFC7410438FC7E3F",
INIT_2C => X"00000000000000000000000000005B78FC7AAD56FB6DBEF1FAFD7E384001EF14",
INIT_2D => X"55517FFFFFFFFFFFFFFFFFFFFEFF7AA974AA5500020005500000000000000000",
INIT_2E => X"5AA80154AA557BEAB45002ABFFFFFFFFFFFEFF7FBFDFFFF7AA974BA550415410",
INIT_2F => X"EFF7FBFDFFFAAD168B55AA80000BAF7FFFDF5500517FFFFFFFBFDFEFFFFFEAB4",
INIT_30 => X"155F78015400557BFDFEFF7FBEAB55A2D56AB55A28002000F7FFC2155552ABFF",
INIT_31 => X"8B45AAFBFFFFFFFAA95545F7840201000043DFEFA2D56AB45AAD57DFEFF7AA82",
INIT_32 => X"E8B55000428B55AAD168B55F7FFFDFEFFFAA9555555003DE00007FFDF45AAD56",
INIT_33 => X"568B55A280021EF557FD755555042AB55AAD16ABFFFFFBEAB45A280155EF557F",
INIT_34 => X"0000000000000000000000000000000000000000000007FEAB55A2D17FFEFFFD",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000040000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(19),        -- Port A data input
DOA(0)   => data_read_a_hi_256(19),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(19),        -- Port B data input
DOB(0)   => data_read_b_hi_256(19),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_20_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000003",
INIT_01 => X"A75FF80000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"14088080800008400F655001FFCFF80018FA8044000000000000011000000007",
INIT_03 => X"0000000000000000000000000000000024001660380000000000000000004FF8",
INIT_04 => X"000079800014CC02C034001600000000000000101EC0012EE0C0026E1E80F000",
INIT_05 => X"1F0FF433EFF0440C3902100002203F2EFC040388137C3E20C8EEC00284033CC0",
INIT_06 => X"00F00100002E22EB440012C809B2FFF7C8E8840155FDC0000010E40087D8787A",
INIT_07 => X"03B800000000000000008407FC800B0000000100600040000C205FF91C000F80",
INIT_08 => X"F28C0B0300020852000002101554021F00000000000000009049226020000200",
INIT_09 => X"D80000007BEFBC010002008FF7F00000000010018A81000041C401000004FFDF",
INIT_0A => X"00000ADF000000200000008000008028300100461003EAFE400000120000913F",
INIT_0B => X"0000000000000000000000000200200290000000000000000200000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000010001000000",
INIT_0D => X"00000100000010000002000080101FFB60000000000000000000000000000000",
INIT_0E => X"03007FE29FF800C00000001002040000000000000020480002E42429C0000080",
INIT_0F => X"0004D4E180010040000400000001E60040000400000001E6010003C000000000",
INIT_10 => X"000000094B1E0040000400000001E60040000400000001E60804000000400000",
INIT_11 => X"00002000000000033628000100100000004000000006170C0008001000004000",
INIT_12 => X"000000000295810000000A100020614148002000000000004307CC3CC0000804",
INIT_13 => X"5802000000000014AC000120200000000003F0D800020100000000000A4B0020",
INIT_14 => X"0020C0C00000000002E2D000001006204040000000005786C004000000000052",
INIT_15 => X"0100A0C0939BEE1810080200000E0CE0EC000010020000000000000AE8A00002",
INIT_16 => X"2008040400400C08080000000000049F6FFC0100000000000008008008000400",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0100000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0C30C30C320624C1090D0F3CF3CD038001801C10000804482A60D09008269020",
INIT_1B => X"90C86432190C86432190CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2C30C3",
INIT_1C => X"F80000432190C86432190C86432190C86432190C86432190C86432190C864321",
INIT_1D => X"AA5504020100800000000000000000000000000000000000000000000000401F",
INIT_1E => X"FFFFFFFFFFFFFFAA954BA5500020BA5D7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974",
INIT_1F => X"74AA00003FFFFFFFFFFFFFFFFFFFFFFF7AA974AA550002000007BFFFFFFFFFFF",
INIT_20 => X"FDFEFFFAE974AA5D003FE005D043FFFFFFFFFFFFFFFFFFFFEFF7AE954BA5D041",
INIT_21 => X"BFFFFFFFFFFFFFFFFFBFDFEFFFAA974BA5D517FFFF087FFFFFFFFFFFFFFFFFFF",
INIT_22 => X"8402000F7D56ABFF55003FFFFFFFFFFFFFF7FBFDFFFAA84000105D556AB55557",
INIT_23 => X"FFFFFFEFF7FBEAB55A28000010F7D16ABEF08043FFFFFFFFFFFFFF7FBFDF55A2",
INIT_24 => X"000000000007BFFFFFFFFFFFFEFF7D16AB45AA8002000F7D5575455D2EBFFFFF",
INIT_25 => X"FFFFFFFFFFFFAE974AA550400028000000000000000000000000000000000000",
INIT_26 => X"380071FFFFFFFFFFFFFFFFFFFFFFFF7AA954BA550000082557FFFFFFFFFFFFFF",
INIT_27 => X"FEFFFAE954AA55041549214043FFFFFFFFFFFFFFFFFFDFEFF7AE974BA5500050",
INIT_28 => X"FFFFFFFFFFFFFF7FBFDFFFFFAA974BA550038E285D0E3FFFFFFFFFFFFFFFFBFD",
INIT_29 => X"02028555F6FB7D5D75FFFFFFFFFFFFEFF7FBFAFD7E3A4954BA555B7AFC70871F",
INIT_2A => X"FFDFEFE3F5FAF45AA8000038F7DB6FBD7490E3FFFFFFFFFDFEFF7F1FAFC7A280",
INIT_2B => X"DF525455524BFFFFFFFBFDFC7E3F5E8B45A28402010FFDB6ABEF140A3FFFFFFF",
INIT_2C => X"00000000000000000000000000007FFFFFFF7FBF8FC7EBD568B55A28000000FF",
INIT_2D => X"557FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5504000BA0800000000000000000",
INIT_2E => X"FFFAE954BA5500174AA08517FFFFFFFFFFFFFFFFFFFFEFF7AA974AA550002000",
INIT_2F => X"FFFFFFFFFEFF7FBFDFFFF7AA974BA55041541055043FFFFFFFFFFFFFF7FBFDFE",
INIT_30 => X"4AA557BEAB4500557FFFFFFFFFDFEFF7FFFFFEFF7AE974AA550028AAA5D2ABFF",
INIT_31 => X"DFEFFFD568B55A284020BA557FFFFFF5D517FFFFFFFBFDFEFFFFFEAB45AA8015",
INIT_32 => X"EABEF5D2ABFFEFF7FBFDFFFAAD168B55AA80000BAF7FFFDF55002EBFFFFF7FBF",
INIT_33 => X"56AB55A28002000F7FFC215555043DFEFF7FBFFF55A2D16AB45AA8402000F7FB",
INIT_34 => X"0000000000000000000000000000000000000000000007BFDFEFF7FBEAB55A2D",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000007FFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(20),        -- Port A data input
DOA(0)   => data_read_a_hi_256(20),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(20),        -- Port B data input
DOB(0)   => data_read_b_hi_256(20),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_21_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"4A302428B824900A128C090A5C1800261500213C005FE812D10420054085A202",
INIT_01 => X"081FFE3440B609703B0427F801A40B8115BC4F655300340288A40D30040E4DD8",
INIT_02 => X"0109095C30C98809800000F9FFFFFFFF149FF1FCA4C0421B182E3490DF145FE4",
INIT_03 => X"084A76341244919000099486400026523C041660BA000100CC12701015007FF8",
INIT_04 => X"000079800014CC03C075161E001118653D2408041FC004AEF000816E1C11F541",
INIT_05 => X"3F0F807BFFE000240100004683103E7FFE02482553FC3C0204EFC25010143CC0",
INIT_06 => X"008808210996035A000006EC2E04FFFFC0A0000101FFE4036450E08247F87870",
INIT_07 => X"4003400812A156C002822987FC830F40134CC74D002016612DE87FFE00400804",
INIT_08 => X"F02348D2D00080C0C53400044114000000D022640B42406808790055043A8282",
INIT_09 => X"F84056387FEFBC110008420F7FF388B70A20389346FE9F26120200800008FDFF",
INIT_0A => X"4518DBFF00020004C0A6044901112A0908AA14601DE3EBFE0A812D8D5B742D3F",
INIT_0B => X"104032901CC63410ABD249C4B3007127080806FF917FC30010107688862A28C5",
INIT_0C => X"46C9146C9146C9146C9146C9146CC8A3648A3642003184822040D000D8C41807",
INIT_0D => X"201800500941044312000900D4621FFBE0008A94C822CA8919018206C9146C91",
INIT_0E => X"2029FFEADFF8050250010030165290008800440022201082401A002000C48000",
INIT_0F => X"18048A004A6C0D2820302C005A83480D1820302A009B02B101390C0CB2830816",
INIT_10 => X"1408904831400D1820302C005A83480D2820302A009B02B021A85C0941150013",
INIT_11 => X"5C08834600024D052C1051E0B92D400360520202682C19024B6164E300448510",
INIT_12 => X"6404093E22A2012418A9D1D44ADD9E0F174103820101C0B8160D5516259FA1A8",
INIT_13 => X"60D8AA288209E615100280DA0052000C5006402000206C55144104D510CC1B0D",
INIT_14 => X"0A0D50020C04023033C52009144231D902818100C90058010361AC808126C886",
INIT_15 => X"2202386454988140600C0181500A13E830011008B0374007000B4E0CD0002450",
INIT_16 => X"0080224004002000000703804008001F7FFF01B982B01258088C008CC41198A1",
INIT_17 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_18 => X"8020080200802008020080200802008020080200802008020080200802008020",
INIT_19 => X"0000000000000000000002008020080200802008020080200802008020080200",
INIT_1A => X"BEFBEFBEFBFF7FEFEFFFE79E79FFFF7CFF77FBFFEFBFF9F7E0FDF9EFEFBF0000",
INIT_1B => X"DFEFF7FBFDFEFF7FBFDFEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEF",
INIT_1C => X"F80000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"BA5D00020000800000000000000000000000000000000000000000000000401F",
INIT_1E => X"FFFFFFFFFFFFFFAE974AA550402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974",
INIT_1F => X"20BA5D7FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5D00020AA5D7FFFFFFFFFFFF",
INIT_20 => X"FFFFFF7AA974BA5D0402000557BFFFFFFFFFFFFFFFFFFFFFFFFFAA954BA55000",
INIT_21 => X"03FFFFFFFFFFFFFFFFFFFFFFF7AA974AA55000200000003FFFFFFFFFFFFFFFFF",
INIT_22 => X"AE954BA5D04174AA00003FFFFFFFFFFFFFFFFFFFFEFF7AE974BA5D00174BA000",
INIT_23 => X"FFFFFFFFFFFFFDFEFF7AE954AA5500174BA5D043FFFFFFFFFFFFFFFFFFFFEFF7",
INIT_24 => X"000000000007FFFFFFFFFFFFFFFFFFFFDFEFFFAE974AA5D003FE005D2EBFFFFF",
INIT_25 => X"FFFFFFFFFFFFAE974BA5D0000010000000000000000000000000000000000000",
INIT_26 => X"BA557FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550400028007FFFFFFFFFFFFFF",
INIT_27 => X"FFFF7AA954BA550000082557BFFFFFFFFFFFFFFFFFFFFFFFFFAA954BA5D00000",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFEFF7AA974AA5D04050005571FFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"954BA5D00154AA00043FFFFFFFFFFFFFFFFFFDFEFF7AE974BA55000503800003",
INIT_2A => X"FFFFFFFFFBFDFEFFFAE954AA550415492140E3FFFFFFFFFFFFFFFFFFDFEFF7AE",
INIT_2B => X"0038E285D2ABFFFFFFFFFFFFFFFFBFDFEFFFAA974BA5D00104925D0E3FFFFFFF",
INIT_2C => X"000000000000000000000000000071FFFFFFFFFFFFFFF7FBFDFFFFFAA974BA55",
INIT_2D => X"087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D00000100000000000000000000",
INIT_2E => X"FF7AA954BA5D00000BA5D7FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5504000BA",
INIT_2F => X"FFFFFFFFFFFFFFFFFFEFF7AA974AA550002000557BFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA5500174AA08043FFFFFFFFFFFFFFFFBFDFEFF7AE954AA5D041740055517FF",
INIT_31 => X"FFFFF7FBFDFFFFFAA974AA5D00174BA08043FFFFFFFFFFFFFF7FBFDFEFFFAE95",
INIT_32 => X"00010552ABFFFFFFFFFFFEFF7FBFDFFFF7AA974BA550415410552ABFFFFFFFFF",
INIT_33 => X"FFFFEFF7AE974AA550028AAA5D2EBFFFFFFFFFDFEFF7FBFFFFFF7AE954BA5D00",
INIT_34 => X"000000000000000000000000000000000000000000000557FFFFFFFFFDFEFF7F",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(21),        -- Port A data input
DOA(0)   => data_read_a_hi_256(21),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(21),        -- Port B data input
DOB(0)   => data_read_b_hi_256(21),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_22_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"5290F4CDE914905A14A43D33F488243E17122300F55FEB189B343A1140548380",
INIT_01 => X"A94007B259F6A975386262000C344BA9573C6FF57B18A5FB0ABFCD3C2C5F4F0C",
INIT_02 => X"877FE30EB378008D202551040030071869D0040180AC4B685F6E26FAA0810006",
INIT_03 => X"431965109E4481D6B5AAD6875AD6AB5A1815600802888808DEA83552954D3000",
INIT_04 => X"492C0020220001010E4916C884DCD607E5EC2A344103E48003D0800023D0072C",
INIT_05 => X"00107C441001100D620A06D683018001023D37E5088043620101179092540112",
INIT_06 => X"40111C2D50A46AE45281502E4A2200081ADA0E054402365774611E047020008E",
INIT_07 => X"680BD5AA4BF5C91F840C1710010344DB9A808FDFF3DE0313014A200754040180",
INIT_08 => X"0EA212D6D481ADF0CE47CA21544009007A64EBD64049D028B93D9561A48F6027",
INIT_09 => X"207246A80400015805060040080A2A0F4A82381B4000BFB65A0283800AA50020",
INIT_0A => X"4539C020E11810098D4067EFF9FF284D483E35602820110204804818CD280100",
INIT_0B => X"10081E9528963546278008AA800470370000A0004D0000002126F30C902A29C5",
INIT_0C => X"40E1540E1540E1540E1540E1540E4AA070AA07000A0000308000190168200281",
INIT_0D => X"6870A9CA0D458D131652A154D46B600085080B14009A2B2906504940E1540E15",
INIT_0E => X"448C00044000A1EC1C44140D101A54280A14050A028500A84F02842A24C594A0",
INIT_0F => X"38359E0C4E6C256690581800F1C3E82562B0581200F1C3F08145602280402080",
INIT_10 => X"100AB8581B602562B0581800F1C3E8256690581200F1C3F1238473F121000613",
INIT_11 => X"73F0E1050083750B3E4275F829547008600C030374361FA2CEE046D48122C438",
INIT_12 => X"C4CC012A66F61154C019511628756231018500C00203E1380615651607822384",
INIT_13 => X"608AA612C0096C37B00D1724801A0009C606D1221D104553096004B61BCC1128",
INIT_14 => X"12A41E0F0600035842E7601C2C4AC68A98810080AA825A890225189980254CDE",
INIT_15 => X"A89637E00D0A1080301401C390320188321C2C0B13890105800D520AF94870B0",
INIT_16 => X"88222F110111B281A54753AA004002601001918008C10912A4440B24E8B58234",
INIT_17 => X"8220882208822088220882208822088220882208822088220882208822088220",
INIT_18 => X"2008020080200802008020080200802008020080200802208822088220882208",
INIT_19 => X"1448000000001FFFFFFFFC802008020080200802008020080200802008020080",
INIT_1A => X"9E79E79E7BFF3FEFEBEEEFBEFBEFBEFDFEF7F47F8FBEF5EB7E6CFEFBEFBE8289",
INIT_1B => X"CFE7F3F9FCFE7F3F9FCFE79E79E79E79E79E79E79E79E79E79E79E79E79E79E7",
INIT_1C => X"F800003F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9F",
INIT_1D => X"BA5D04000000000000000000000000000000000000000000000000000000401F",
INIT_1E => X"FFFFFFFFFFFFFFAE974BA5D0002000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974",
INIT_1F => X"2010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA550000010007FFFFFFFFFFFF",
INIT_20 => X"FFFFFFFAE954AA5D00000AA007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA55040",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5D00020AA5D7FFFFFFFFFFFFFFFFFFF",
INIT_22 => X"AA954BA5500020BA5D7FFFFFFFFFFFFFFFFFFFFFFFFFFAA954BA5504000AA557",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFAA954BA5500000BA5D7BFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"00000000000003FFFFFFFFFFFFFFFFFFFFFFF7AA974BA5D040200055517FFFFF",
INIT_25 => X"FFFFFFFFFFFFAE974BA5D0402000080000000000000000000000000000000000",
INIT_26 => X"10087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0000010007FFFFFFFFFFFFFF",
INIT_27 => X"FFFFFAE974AA550400028007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA5500020",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFAE954AA5D00020BA087FFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"954BA5504020AA5D7BFFFFFFFFFFFFFFFFFFFFFFFFFAA954BA5D00000BA557FF",
INIT_2A => X"FFFFFFFFFFFFFFFF7AA954BA5500000825571FFFFFFFFFFFFFFFFFFFFFFFFFAA",
INIT_2B => X"040500055517FFFFFFFFFFFFFFFFFFFFFFF7AA974AA5D00070925D71FFFFFFFF",
INIT_2C => X"0000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFEFF7AA974AA5D",
INIT_2D => X"007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020000800000000000000000",
INIT_2E => X"FFFAE974AA550002000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0000010",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFAE954AA5504000BA087FFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA5D00000BA5D7BFFFFFFFFFFFFFFFFFFFFFFFFFAA954AA5D00020AA007FFFF",
INIT_31 => X"FFFFFFFFFFFEFF7AA974BA5504020BA557BFFFFFFFFFFFFFFFFFFFFFFFF7AA95",
INIT_32 => X"154105D517FFFFFFFFFFFFFFFFFFFFEFF7AA974AA55000200055517FFFFFFFFF",
INIT_33 => X"BFDFEFF7AE954AA5D041740055557FFFFFFFFFFFFFFFFFFDFEFF7AE974AA5D00",
INIT_34 => X"000000000000000000000000000000000000000000000043FFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000007FFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(22),        -- Port A data input
DOA(0)   => data_read_a_hi_256(22),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(22),        -- Port B data input
DOB(0)   => data_read_b_hi_256(22),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_23_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"EF20906D902424807BC8241BC81801B97D38AD3C0800103362A6741C80A12A02",
INIT_01 => X"001FFF8409F089003B4422000D80C80106804A7951C5B9D1C828043EA28838F9",
INIT_02 => X"073B8858218C2C50801000F9FFEFF8E72CA7F5FC2E048026496834D84721DFE0",
INIT_03 => X"2C4360101A4001001005080400401420350016E0BB222341C312000014006FF8",
INIT_04 => X"00017B810015DC03D034201E14000036486008101FC0002EE006297E1C05F561",
INIT_05 => X"BF0F817FFFE80100004044800080BEFFFC0248005FFC3C18A5FFC2444484BCC0",
INIT_06 => X"0400000409120338860900482404FFFFC000000001FFC0832050E00047F97870",
INIT_07 => X"200246801C41C3E81E872C8FFE900FC31348EFDF03BE15E22DA07FF92C204102",
INIT_08 => X"F6220280D2B025988311AB14155421006891A1089F6E200000022C140068EB90",
INIT_09 => X"F8001011FFEFBC80000000077FF184B03010004002FE000000201000000FFDFF",
INIT_0A => X"00001BFFA800808189A657EF81DD0C00079CD00837C3EBFD4201258112D4487F",
INIT_0B => X"24483890564084198AD249C433200180082A06FF907FC3081812048006000000",
INIT_0C => X"8608086080860808608086080860804304043042003184822150C000D8C41806",
INIT_0D => X"03000100200180480000095280001FFBF040C088CD20E0A21921828608086080",
INIT_0E => X"3821FFEAFFF805025E00853B92588000400020001000020A8018008002000014",
INIT_0F => X"486148484054395E27E428002A4200397E07E422002A420100382FCC30832A16",
INIT_10 => X"0C0788417000397E07E428002A4200395E27E422002A420110A51C01C0590401",
INIT_11 => X"1C01A2490040590C08120558C1759BE1C05A0400383808800DA1929F72864110",
INIT_12 => X"20000136006000215EA0A4833A32C8832050028603050014031B3950000C90A5",
INIT_13 => X"006658280009A2030108B14AC05C00112405222088B8332C140004D101800CE7",
INIT_14 => X"196B6808060201281004228996085F10020180C030880D11019CE4000026C00C",
INIT_15 => X"52A49DC7143F01C04240030720641E0A028996483A17204680410A04104A2659",
INIT_16 => X"0401000080080000000000002001201F7FFC0011C2F81A48080CA32800A01081",
INIT_17 => X"4010040100401004010040100401004010040100401004010040100401004010",
INIT_18 => X"0100401004010040100401004010040100401004010040100401004010040100",
INIT_19 => X"0000000000000000000000040100401004010040100401004010040100401004",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"F800000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"BA5D04020100000000000000000000000000000000000000000000000000401F",
INIT_1E => X"FFFFFFFFFFFFFFAE974BA5D0400000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974",
INIT_1F => X"2000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400010087FFFFFFFFFFFF",
INIT_20 => X"FFFFFFFAE974BA550002000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D000",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA550000010007FFFFFFFFFFFFFFFFFFF",
INIT_22 => X"AE974AA550402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550400000087",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFAE974AA550402000087FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5D00000AA007FFFFFFF",
INIT_25 => X"FFFFFFFFFFFFAE974BA5D0402010000000000000000000000000000000000000",
INIT_26 => X"10087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000087FFFFFFFFFFFFFF",
INIT_27 => X"FFFFFAE974BA5D0000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04000",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFAE974BA550002000007FFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974AA550400010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550002010087FF",
INIT_2A => X"FFFFFFFFFFFFFFFFFAE974AA550400028007FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_2B => X"00020BA087FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5D0402038007FFFFFFFFF",
INIT_2C => X"00000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5D",
INIT_2D => X"087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020100000000000000000000",
INIT_2E => X"FFFAE974BA5D0400000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D0000010007FFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4AA550002000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA550002010087FFFF",
INIT_31 => X"FFFFFFFFFFFFFFFAE954AA550400010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_32 => X"000AA087FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5504000BA087FFFFFFFFFFF",
INIT_33 => X"FFFFFFFFAA954AA5D00020AA007BFFFFFFFFFFFFFFFFFFFFFFFFFAA954AA5D04",
INIT_34 => X"0000000000000000000000000000000000000000000007BFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000007FFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(23),        -- Port A data input
DOA(0)   => data_read_a_hi_256(23),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(23),        -- Port B data input
DOB(0)   => data_read_b_hi_256(23),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_24_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100600007FFF000080108004000800020000840041000080808",
INIT_02 => X"172A00D000EF8210000000F9FFEFF8E7240FF1FC224087B1000639401D005FC0",
INIT_03 => X"00003A2E200811000000000400000000340016603A0000004860400014006FFF",
INIT_04 => X"000079800014CC03C034001E04010850300000101FC0002EE000006E1C00F500",
INIT_05 => X"1F0F8033FFE000000000000000003E2FFC024800137C3C0000EFC00000003CC0",
INIT_06 => X"0000000009120110020100002404FFFFC000000001FFC0000010E00007F87870",
INIT_07 => X"200102050840950002802C87FC800FCAA035400001B918600C207FF800000000",
INIT_08 => X"F6234AD280B02500063AC2840001610020408178B600C2400013649608730004",
INIT_09 => X"F80000007FEFBC00000000077FF000B00000000002FE0000000000000000FDFF",
INIT_0A => X"00001BFFA0000005501AA00000CE20000094000011C3EBFC020125811254083F",
INIT_0B => X"0040A040004000008012414433000100080806FD107FC3000000000006000000",
INIT_0C => X"0608006080060800608006080060800304003042003180822040C00090C41806",
INIT_0D => X"004800B0000000000000000000001FFBE0008080C820C0801801800608006080",
INIT_0E => X"2021FFEADFF80002080000000208800000000000000000020018000000000000",
INIT_0F => X"840009181008024A00043601100210024A00043C0110020901382CCCB28B0806",
INIT_10 => X"180040A03080024A00043601100210024A00043C01100209240C840C201D0210",
INIT_11 => X"840A604E0080820009908008341B000A8212070082002890010068320860C920",
INIT_12 => X"40600800082041205EC00044C1ACB66C37542082030281E0580001012811A40C",
INIT_13 => X"80B27A004300004103160DB3005E000618040C022000593D002180002090166B",
INIT_14 => X"2BBFF20406040084210C062000C2A2DDD00180C04504086002CD680C01000104",
INIT_15 => X"20804295C98F80400008040CC0582169022000C2876C40478002850016088001",
INIT_16 => X"0000000000000000000000000000001F7FFC001B823018F00880008805241060",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"9EF9EF9EFB263CC3090CABAEBAFF96857757B73E6089966B9EF9D5A220CC8000",
INIT_1B => X"C1E0F0783C1E0F0783C1EFBEFBEFBE79E79E79E79E79EFBEFBEFBEFBEFBEF9EF",
INIT_1C => X"F800000783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783",
INIT_1D => X"BA5D04020100800000000000000000000000000000000000000000000000401F",
INIT_1E => X"FFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974",
INIT_1F => X"0000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000087FFFFFFFFFFFF",
INIT_20 => X"FFFFFFFAE974BA5D0400000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400010087FFFFFFFFFFFFFFFFFFF",
INIT_22 => X"AE974BA5D0002000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0000010007",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFAE974BA5D0002000007FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA550002000007FFFFFFF",
INIT_25 => X"FFFFFFFFFFFFAE974BA5D0402010080000000000000000000000000000000000",
INIT_26 => X"00087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFF",
INIT_27 => X"FFFFFAE974BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000007FFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA5D0000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400010087FF",
INIT_2A => X"FFFFFFFFFFFFFFFFFAE974BA5D0000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_2B => X"0002000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA550002000087FFFFFFFFF",
INIT_2C => X"00000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA55",
INIT_2D => X"007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020100800000000000000000",
INIT_2E => X"FFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA5D0400000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000007FFFF",
INIT_31 => X"FFFFFFFFFFFFFFFAE974BA5D0000010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_32 => X"00010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0000010007FFFFFFFFFFF",
INIT_33 => X"FFFFFFFFAE974BA550002010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5500",
INIT_34 => X"0000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(24),        -- Port A data input
DOA(0)   => data_read_a_hi_256(24),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(24),        -- Port B data input
DOB(0)   => data_read_b_hi_256(24),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_25_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100200002000000080100004000000020000800041000080808",
INIT_02 => X"1000218000000800000000F9FFEFF8E738FFF1FC20400400000004455A375FE0",
INIT_03 => X"00002000000001000000000400000000340016623A0000004000000014006FFF",
INIT_04 => X"924279824C94CC1BE0B4001F20000000020380401FE0082EF000106E1C00F500",
INIT_05 => X"1F0F8033FFF048202582800100523E2FFE024820137C3C0040EFE02000003CE4",
INIT_06 => X"10DC00CC0992033A062116E82404FFFFC0E0801101FFC0000010E08A07FC7870",
INIT_07 => X"000000000000000002802C87FC800F8000000000019810600C207FFF3C410D84",
INIT_08 => X"FE8002000080281000008A0000014100200081000000000080480AE000000200",
INIT_09 => X"FC0020007FEFBE031018C31F7FFBAEBC0020008086FE0000100280800000FDFF",
INIT_0A => X"00001BFFE00301000000000000CC02000014000191C3EBFF4A7DF795965C6D3F",
INIT_0B => X"0040200000400000801243443B000100880806FD107FC3018000000006000000",
INIT_0C => X"0608006080060800608006080060800304003042003B99862444E61492C41806",
INIT_0D => X"00000000000000000000001280001FFBE0008080C820C4801801800608006080",
INIT_0E => X"3021FFEADFF805025C0304001E58906088304418222C108A009A090400000000",
INIT_0F => X"00000100100000480000200100000000480000200100000100380F0C30830A06",
INIT_10 => X"0000008000000048000020010000000048000020010000000004040000010000",
INIT_11 => X"0400004000000000008080000011000000020000000020000000001200000100",
INIT_12 => X"000000000800002018C010000020800000800122000000004004000008000004",
INIT_13 => X"0002080000000040000001020020000000000800200001040000000020000021",
INIT_14 => X"0021000008001000000800200000021000020100000000200004200000000100",
INIT_15 => X"0000008400000000605000000000200000200000020400000000000002008000",
INIT_16 => X"288226410410346010000000400A011F7FFE0031823010400800000800001840",
INIT_17 => X"8822088220882208822088220882208822088220882208822088220882208822",
INIT_18 => X"8220882208822088220882208822088220882208822088220882208822088220",
INIT_19 => X"00017FFFFFFFFFFFFFFFFE088220882208822088220882208822088220882208",
INIT_1A => X"2410492410A048029890AD34D35FDD144A50CB5462D14997BE09E760AED04040",
INIT_1B => X"8C46231188C46231188C49249249249249249249249241041041041041041049",
INIT_1C => X"F80000B158AC562B158AC562B158AC562B158AC562B158AC562B158AC562B158",
INIT_1D => X"BA5D040201000000000000000000000000000000000000000000000000007FFF",
INIT_1E => X"FFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974",
INIT_1F => X"2010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFF",
INIT_20 => X"FFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000087FFFFFFFFFFFFFFFFFFF",
INIT_22 => X"AE974BA5D0400000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000007",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFAE974BA5D0400000087FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000007FFFFFFF",
INIT_25 => X"FFFFFFFFFFFFAE974BA5D0402010000000000000000000000000000000000000",
INIT_26 => X"10087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFF",
INIT_27 => X"FFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA5D0402000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000087FF",
INIT_2A => X"FFFFFFFFFFFFFFFFFAE974BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_2B => X"0400000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000087FFFFFFFFF",
INIT_2C => X"00000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D",
INIT_2D => X"087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020100000000000000000000",
INIT_2E => X"FFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFF",
INIT_31 => X"FFFFFFFFFFFFFFFAE974BA5D0402000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_32 => X"02000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000087FFFFFFFFFFF",
INIT_33 => X"FFFFFFFFAE974BA5D0400000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_34 => X"0000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000007FFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(25),        -- Port A data input
DOA(0)   => data_read_a_hi_256(25),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(25),        -- Port B data input
DOB(0)   => data_read_b_hi_256(25),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_26_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"E9264EAB20190CA3BA4997AA9002AE9C001006B0778015CFA17E0811039879C7",
INIT_01 => X"F1FFF9BB1F773C7F9BB07DFFFDD863FC5FFF3FEFFBBF9FFB22FFFBC7B9F30686",
INIT_02 => X"1B33188302E708180F6FFBFFFFCFFFFF9C7FF7FC24350B99082400001D00DFD8",
INIT_03 => X"4A53D958C50000DCE7366303739CD98C27C57EF57980014F271807E3C9E9CFF8",
INIT_04 => X"DBFAFBD7FB1CDEBEF1BE17F7AC88042787FBFFF8FEE9FF7EE6F4C0EE1FFAF869",
INIT_05 => X"5F0FFEB3EFFEFFBDA7F7FED508707E2EFEBF6FFEB37C3FF302EEEDFF9B487CF6",
INIT_06 => X"AFBE564C71268F3BBF5FBFC2A427FFF7C3E3A74667FDDB7FB870FF30FFDEF87F",
INIT_07 => X"03BC18306396FBEC14489737FDC00B13BB79DFDB83BF4112AF205FFBDD3AFB93",
INIT_08 => X"F21E4391909B381B0B1F8E041051831FA3068D77E000030021324620C0B9C206",
INIT_09 => X"DE89ECC0FBEFBEBF30B8D79FF7F451F33CFD60FE8FFFDF58003B1D4223B4FFDF",
INIT_0A => X"8ED6BFDF3EB3EBF9DDBCE7FDC1DF8A760F3EB980580BFAFFF37DF7B9DF7DCB3F",
INIT_0B => X"6EE6F5E7FAC4C03DB856CD4CF73AC1FC98884FFF19FFC71FEFED7B251E35768E",
INIT_0C => X"06BC606BC606BC606BC606BC606BD3035E3035C62B7BB987666DEF8A90CCFA8F",
INIT_0D => X"CF6100C0E60FB9FC3A80EF69A04DFFFF7FF5F9A0DC33E9B41D01D207BC606BC6",
INIT_0E => X"7027FFFF9FF8FAFAA3ADEBFB9726BAF5FD7AFEBD7F7EFFD7ACDB7F947F0EA035",
INIT_0F => X"E020080A40403E8BD8002000FC02003E8BD8002000FC02010979AFFE36C36B86",
INIT_10 => X"000EE00034003E8BD8002000FC02003E8BD8002000FC020037B0040A00010003",
INIT_11 => X"040C00400003D80008160400FD81341C00020003B80008C00801EF0285380100",
INIT_12 => X"90981038406809677FA080468C46A81080581002000780C8001C8100201037B0",
INIT_13 => X"00F90D162001C803411FC0024080001F80040026C0807C868B1000E401A01F11",
INIT_14 => X"3F810503A00003E020042AC080CEB01228A80000F600080123E232130407080D",
INIT_15 => X"0087520750001064180807868000110C02C080CFA0042400000F8800105B0201",
INIT_16 => X"7FDFF7EFEEFF3EEC3FF7FBFFBCB7FFFFEFFE00BFF7FEBF420800EC0CBEE61F81",
INIT_17 => X"FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F",
INIT_18 => X"D7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5",
INIT_19 => X"43237FFFFFFFFFFFFFFFFF5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5F",
INIT_1A => X"A69A61861BAF15EAA6AFC38E38EA3AD8ADE7A48F0B366429F434AA9FC376DAE4",
INIT_1B => X"C26130984C26130984C261861861861861861861861861861861861861861869",
INIT_1C => X"F800000984C26130984C26130984C26130984C26130984C26130984C26130984",
INIT_1D => X"BA5D04020100000000000000000000000000000000000000000000000000401F",
INIT_1E => X"FFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974",
INIT_1F => X"2010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFF",
INIT_20 => X"FFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFF",
INIT_22 => X"AE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFF",
INIT_25 => X"FFFFFFFFFFFFAE974BA5D0402010000000000000000000000000000000000000",
INIT_26 => X"10007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFF",
INIT_27 => X"FFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FF",
INIT_2A => X"FFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_2B => X"0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFF",
INIT_2C => X"00000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D",
INIT_2D => X"007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020100000000000000000000",
INIT_2E => X"FFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFF",
INIT_31 => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_32 => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_33 => X"FFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_34 => X"0000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(26),        -- Port A data input
DOA(0)   => data_read_a_hi_256(26),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(26),        -- Port B data input
DOB(0)   => data_read_b_hi_256(26),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_27_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"00080A40000A41248002029000050A088000008242A0004404480002000A1155",
INIT_01 => X"F1FFF1C11F781C129C107DFFFE0860941E81258CA2B71C2220EC1B86E1A00002",
INIT_02 => X"4000002100000014400FF6FFFF0FFFFF8007F1FC211100014200800000887FC0",
INIT_03 => X"0842D85841000098C63061026318C18404C459757000015F00088BE3C0618FF8",
INIT_04 => X"DBEAE5D6D91C2EBCE1B21EA72C00000007FBE7C8F8E9EF79E6D440E91FDAE061",
INIT_05 => X"5C8FFCB38FF6B68984B5BCE408347E28FEBF6FEEB3723F7102E8EDBF8A4872F6",
INIT_06 => X"AB98420C71408D113956AFD0842FFFC7C3032646EFF1DB7FA868FE30EF1CE47E",
INIT_07 => X"10041830600640C415004637FC4003021259CFDB01BF80028E001FF8251AB9D1",
INIT_08 => X"F200822020842203000082050000110023068D03000002820000000840000005",
INIT_09 => X"1C852440E3DF7E2FB0B8E717C7F411F3BC6D60B60FFDDE480018AC4AA3B0FD1F",
INIT_0A => X"18109E1F16B16B71092CE7ED81CF403601229880400BE0FC137FF7A0FF75813F",
INIT_0B => X"86F7D5E382A440349816DD4C755AC16C1A884FFE18FFD757E7ED7A211E81C098",
INIT_0C => X"061A2061A2061A2061A2061A2061E1030D1030D6A37FB9872E65E6AA90CD5AAF",
INIT_0D => X"8FC10080A20ED1D41880CC61A044DFFC6EB5BCA0DE31F8B41C01E0071A2061A2",
INIT_0E => X"2023FFE91FF98AEAA1AC6AC9A3A4AAD5B56ADAB56D5AFD572C597B147506203E",
INIT_0F => X"E020000260403C8948002000EC0000BC8948002000EC00010878AC3CB8AB8857",
INIT_10 => X"000EE0000400BC8948002000EC0000BC8948002000EC000097B0040200010003",
INIT_11 => X"040400400003D80000070400DD81041400020003B80000410801AF0204180100",
INIT_12 => X"101010384008086378A080428C46A80080081002000780C800188000301017B0",
INIT_13 => X"02E909042001C800409FC0020080001F80000007C0807484821000E400205D11",
INIT_14 => X"3F810100A00003E020000BC0808EB01020280000F60000002BA2220204070801",
INIT_15 => X"0007520750000024080807868000100403C0808FA0040400000F8800001F0200",
INIT_16 => X"5B5EF3AF6AF6389C2FE128971AB2DDDF8FFE0031B776BF4208006C0C92621F81",
INIT_17 => X"B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D",
INIT_18 => X"56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5",
INIT_19 => X"43A3FFFFFFFFFFFFFFFFFD5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B",
INIT_1A => X"0000000001E0080397908000000A48710B4080240E543021B438A010825238B4",
INIT_1B => X"0804020100804020100800000000000000000000000000000000000000008200",
INIT_1C => X"F80000A05028140A05028140A05028140A05028140A05028140A05028140A050",
INIT_1D => X"BA5D04020100000000000000000000000000000000000000000000000000401F",
INIT_1E => X"FFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974",
INIT_1F => X"2010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFF",
INIT_20 => X"FFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFF",
INIT_22 => X"AE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFF",
INIT_25 => X"FFFFFFFFFFFFAE974BA5D0402010000000000000000000000000000000000000",
INIT_26 => X"10007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFF",
INIT_27 => X"FFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FF",
INIT_2A => X"FFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_2B => X"0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFF",
INIT_2C => X"00000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D",
INIT_2D => X"007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020100000000000000000000",
INIT_2E => X"FFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_31 => X"FFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_32 => X"02010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFF",
INIT_33 => X"FFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_34 => X"0000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000007FFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(27),        -- Port A data input
DOA(0)   => data_read_a_hi_256(27),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(27),        -- Port B data input
DOB(0)   => data_read_b_hi_256(27),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_28_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"02200AA400180030808802A900002A08001280A08A801044104A1000001818C3",
INIT_01 => X"50A00011460214428114180000882214413D0A71592A01D92213D28005210202",
INIT_02 => X"1444428102100884000AA30200000000C1000401041108404400022220800000",
INIT_03 => X"461080404900000C6314A900318C52A40051081000888806108802A141288001",
INIT_04 => X"00800040110102000902002000888400081045A8A00003C00000500000080008",
INIT_05 => X"0000000000024CA0A0101800032000400000000B800000014000000B08180000",
INIT_06 => X"814016012000C405280200008001000011110012220009A88800009A88000000",
INIT_07 => X"0004891224228810080010200040001020800000004000008200000240081400",
INIT_08 => X"00A010040401080308400821155540001122448142491008A004912040840221",
INIT_09 => X"0020405000000124058200408000880004440004080160C8100A858009940000",
INIT_0A => X"4D29400002002038104000000020003204000880082800010000000C0000E400",
INIT_0B => X"12220122A000416811040000400800081022C0000080000206CB0821082B694D",
INIT_0C => X"80B0280B0280B0280B0280B0280B01405814058009000421833010800A000200",
INIT_0D => X"C4210040860B188C0A8065302005A004039010280001001600200081B0280B02",
INIT_0E => X"500600010000280000802050010660001000080004004900204020105302A000",
INIT_0F => X"0000000A00000081480000001400000081480000001400000800C01082082210",
INIT_10 => X"0000000024000081480000001400000081480000001400000010000200000000",
INIT_11 => X"0004000000000000001400000080041400000000000000C00000010004180000",
INIT_12 => X"1010100000480802A40000000400000080081000000000000004800000000010",
INIT_13 => X"0001010420000002400040000080000000000024400000808210000001200010",
INIT_14 => X"04000100A0000000000028400004000020280000000000012002020204000009",
INIT_15 => X"0001000000000024080000000000010400400004000004000000000000510000",
INIT_16 => X"0108408420430E699AA42A1508104EA08000000810020000000044001AC20500",
INIT_17 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_18 => X"0040100401004010040100401004010040100401004010040100401004010040",
INIT_19 => X"1708000000000000000000010040100401004010040100401004010040100401",
INIT_1A => X"20820820800D41A8283AC618618EF1088160885001234B96061CCDEC4D205061",
INIT_1B => X"0C06030180C06030180C08208208208208208208208208208208208208208208",
INIT_1C => X"F80000B0582C160B0582C160B0582C160B0582C160B0582C160B0582C160B058",
INIT_1D => X"BA5D04020100000000000000000000000000000000000000000000000000401F",
INIT_1E => X"FFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974",
INIT_1F => X"2010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFF",
INIT_20 => X"FFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFF",
INIT_22 => X"AE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFF",
INIT_25 => X"FFFFFFFFFFFFAE974BA5D0402010000000000000000000000000000000000000",
INIT_26 => X"10007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFF",
INIT_27 => X"FFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FF",
INIT_2A => X"FFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_2B => X"0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFF",
INIT_2C => X"00000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D",
INIT_2D => X"007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020100000000000000000000",
INIT_2E => X"FFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_31 => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_32 => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_33 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_34 => X"0000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000007FFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(28),        -- Port A data input
DOA(0)   => data_read_a_hi_256(28),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(28),        -- Port B data input
DOB(0)   => data_read_b_hi_256(28),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_29_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"79964E4BA01DACAB9E659792D00AAE160002829C7FDFEFCEE97C2815039D70C3",
INIT_01 => X"50BFF9AB0775343F9AB01DF80D5821FC0FFF3FEFD1AF9FF1207FFBC7B9720586",
INIT_02 => X"0B33180300E700080F6AAA7BFFC007189C7FF2FC003503980A0000001D00DFD8",
INIT_03 => X"0401D940CD0000C8421A2B03210868AC23403E903900010E271006A148A0C000",
INIT_04 => X"49B87A417315D20A313E17F1800000058013DDF8BE21F36E02F0D06E03E8F800",
INIT_05 => X"1F007E33E01A4D9C87525E5101603E6E023D27DA937C03E340EE25CB9B483C12",
INIT_06 => X"85AA06002026872BAE0B1282A005FFF001E1870223FC3BFC98101F109FC6780F",
INIT_07 => X"03BC081023B233E804488527FDC008019968D74982C94110AF204001BC285A82",
INIT_08 => X"001E4191901A101B031F84000000831FA1028575A000110800124600C039C002",
INIT_09 => X"C60888D0782082B50080508FF00048B124D4005C8AFF4158102914800110FFC0",
INIT_0A => X"8AD6ABC02A02A0B0CCB463B4C0748A720B1EA980100BFA02E204D2154D28AA3F",
INIT_0B => X"6A22B126DA40C03531440800C22800B8900042FF0180000ABFEF89250815568A",
INIT_0C => X"803468034680346803468034680353401A340180010A0801422829800A00A001",
INIT_0D => X"87410080C60AB0F42A804628200DBFFF13D05928040329160520528134680346",
INIT_0E => X"2006FFFF8000F8F80281A16A1504302058102C0816244B82A0CA25907D0AA015",
INIT_0F => X"0000080A40000283D80000001402000283D80000001402010901A7D694494192",
INIT_10 => X"0000000034000283D80000001402000283D80000001402002010000A00000000",
INIT_11 => X"000C000000000000081600002080341C00000000000008C00000410085380000",
INIT_12 => X"90981000006809076B2000040400001080581000000000000004810020002010",
INIT_13 => X"0011051620000003410040004080000000040026C00008828B10000001A00210",
INIT_14 => X"04000503A000000000042AC00044000228A8000000000801204212130400000D",
INIT_15 => X"0081000000001064180000000000010C02C000440000240000000000105B0001",
INIT_16 => X"258964C4A44A0C689FF3F9FFEC5D6DBFE0020096528A0B000000CC043EC60780",
INIT_17 => X"5816058160581605816058160581605816058160581605816058160581605816",
INIT_18 => X"8160581605816058160581605816058160581605816058160581605816058160",
INIT_19 => X"03017FFFFFFFFFFFFFFFFE058160581605816058160581605816058160581605",
INIT_1A => X"AEBAEBAEBFFF7FEFCFDF7FFFFFF5DE7CFCB773FFEFBFF3C7E1E779FFEFFF5060",
INIT_1B => X"FEFF7FBFDFEFF7FBFDFEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEEBAEB",
INIT_1C => X"F80000FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFD",
INIT_1D => X"BA5D04020100000000000000000000000000000000000000000000000000401F",
INIT_1E => X"FFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974",
INIT_1F => X"2010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFF",
INIT_20 => X"FFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFF",
INIT_22 => X"AE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFF",
INIT_25 => X"FFFFFFFFFFFFAE974BA5D0402010000000000000000000000000000000000000",
INIT_26 => X"10007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFF",
INIT_27 => X"FFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FF",
INIT_2A => X"FFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_2B => X"0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFF",
INIT_2C => X"00000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D",
INIT_2D => X"007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020100000000000000000000",
INIT_2E => X"FFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_31 => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_32 => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_33 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_34 => X"0000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(29),        -- Port A data input
DOA(0)   => data_read_a_hi_256(29),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(29),        -- Port B data input
DOB(0)   => data_read_b_hi_256(29),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_30_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"9E79E79E7BAF7DEBAFAFEFBEFBFFBFFDFFF7FCFF0FBFFDFF7EFDDFFFEFFE8000",
INIT_1B => X"CFE7F3F9FCFE7F3F9FCFE79E79E79E79E79E79E79E79E79E79E79E79E79E79E7",
INIT_1C => X"F800003F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9F",
INIT_1D => X"BA5D04020100000000000000000000000000000000000000000000000000401F",
INIT_1E => X"FFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974",
INIT_1F => X"2010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFF",
INIT_20 => X"FFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFF",
INIT_22 => X"AE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFF",
INIT_25 => X"FFFFFFFFFFFFAE974BA5D0402010000000000000000000000000000000000000",
INIT_26 => X"10007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFF",
INIT_27 => X"FFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FF",
INIT_2A => X"FFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_2B => X"0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFF",
INIT_2C => X"00000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D",
INIT_2D => X"007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020100000000000000000000",
INIT_2E => X"FFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_31 => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_32 => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_33 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_34 => X"0000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(30),        -- Port A data input
DOA(0)   => data_read_a_hi_256(30),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(30),        -- Port B data input
DOB(0)   => data_read_b_hi_256(30),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_31_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"129000008004A00804A40000400800020000000C005FEA005800200400050100",
INIT_01 => X"A15FF18019700810180065FFFC0040801E80258CA2951C2200EC0906A0804140",
INIT_02 => X"0000000000000011000550FDFF0FFFFF0007F1FC200000011000000000205FC0",
INIT_03 => X"08425818000000908428C0024210A30004045060302223490002014280410FF8",
INIT_04 => X"DB6A618248140C18E0B016872400000007EBA24058E1ECA8E2D400681FD0E061",
INIT_05 => X"1C0FFC338FF01009048084C400103E28FE3F6FE513703F7000E8E5B4825030F6",
INIT_06 => X"0098000C51000910100006C00426FFC7C202060445F1F2572060FE82671C607E",
INIT_07 => X"40001020400440C41C000617FC0003021259CFDB01BF00020C001FF804000980",
INIT_08 => X"F200020000802000000082044000010022048902000002000000000000000004",
INIT_09 => X"1C002400E3CF3E0B1118C31747F000B33820209206FC9E80000000000220FD1F",
INIT_0A => X"00001A1F00110101092CE7ED81CF0004012290000023E0FC027DF780DF74013F",
INIT_0B => X"044094C1028400548812494C31004124080886FE187FC301B124F20016000000",
INIT_0C => X"0608006080060800608006080060C00304003042023B99862444E60090C41887",
INIT_0D => X"0B400080200481501000884080405FF864008880CC30E8A01C01C00608006080",
INIT_0E => X"2021FFE81FF880EA000400098200C04080204010200810020C18090424040034",
INIT_0F => X"E020000040403C0800002000E800003C0800002000E8000100780C2C30830806",
INIT_10 => X"000EE00000003C0800002000E800003C0800002000E8000017A0040000010003",
INIT_11 => X"040000400003D80000020400DD01000000020003B80000000801AE0200000100",
INIT_12 => X"000000384000006118A080428846A80000000002000780C800180000201017A0",
INIT_13 => X"00E808000001C800001F80020000001F8000000280807404000000E400001D01",
INIT_14 => X"3B810000000003E020000280808AB01000000000F600000003A0200000070800",
INIT_15 => X"000652075000000000080786800010000280808BA0040000000F8800000A0200",
INIT_16 => X"080223010010308025410082404A015F0FFE003182701B420800280C80201A81",
INIT_17 => X"8020080200802008020080200802008020080200802008020080200802008020",
INIT_18 => X"0200802008020080200802008020080200802008020080200802008020080200",
INIT_19 => X"04017FFFFFFFFFFFFFFFFC080200802008020080200802008020080200802008",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000080",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"F800000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"BA5D04020100000000000000000000000000000000000000000000000000401F",
INIT_1E => X"FFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974",
INIT_1F => X"2010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFF",
INIT_20 => X"FFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFF",
INIT_22 => X"AE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFF",
INIT_25 => X"FFFFFFFFFFFFAE974BA5D0402010000000000000000000000000000000000000",
INIT_26 => X"10007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFF",
INIT_27 => X"FFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FF",
INIT_2A => X"FFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_2B => X"0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFF",
INIT_2C => X"00000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D",
INIT_2D => X"007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020100000000000000000000",
INIT_2E => X"FFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFF",
INIT_31 => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_32 => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_33 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_34 => X"0000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(31),        -- Port A data input
DOA(0)   => data_read_a_hi_256(31),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(31),        -- Port B data input
DOB(0)   => data_read_b_hi_256(31),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


end;