library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_misc.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library UNISIM;
use UNISIM.vcomponents.all;

entity ram_plasma is
	port(clk             : in  std_logic;
        address_a       : in  std_logic_vector(31 downto 2);
        enable_a        : in  std_logic;
        wbe_a           : in  std_logic_vector(3 downto 0);
        data_write_a    : in  std_logic_vector(31 downto 0);
        data_read_a     : out std_logic_vector(31 downto 0);

        address_b       : in  std_logic_vector(31 downto 2);
        enable_b        : in  std_logic;
        wbe_b           : in  std_logic_vector(3 downto 0);
        data_write_b    : in  std_logic_vector(31 downto 0);
        data_read_b     : out std_logic_vector(31 downto 0));
end; --entity ram     

architecture ram_plasma of ram_plasma is
signal enable_a_lo       : std_logic;
signal wbe_a_lo          : std_logic_vector(3 downto 0);
signal data_write_a_lo   : std_logic_vector(31 downto 0);
signal data_read_a_lo    : std_logic_vector(31 downto 0);
signal enable_b_lo       : std_logic;
signal wbe_b_lo          : std_logic_vector(3 downto 0);
signal data_read_b_lo    : std_logic_vector(31 downto 0);
signal enable_a_hi       : std_logic;
signal wbe_a_hi          : std_logic_vector(3 downto 0);
signal data_read_a_hi   : std_logic_vector(31 downto 0);
signal enable_b_hi       : std_logic;
signal wbe_b_hi          : std_logic_vector(3 downto 0);
signal data_read_b_hi    : std_logic_vector(31 downto 0);
signal address_a_reg     : std_logic_vector(31 downto 2);
signal address_b_reg     : std_logic_vector(31 downto 2);
signal enable_a_lo_256       : std_logic;
signal wbe_a_lo_256          : std_logic_vector(3 downto 0);
signal data_write_a_lo_256   : std_logic_vector(31 downto 0);
signal data_read_a_lo_256    : std_logic_vector(31 downto 0);
signal enable_b_lo_256       : std_logic;
signal wbe_b_lo_256          : std_logic_vector(3 downto 0);
signal data_read_b_lo_256    : std_logic_vector(31 downto 0);
signal enable_a_hi_256       : std_logic;
signal wbe_a_hi_256          : std_logic_vector(3 downto 0);
signal data_read_a_hi_256   : std_logic_vector(31 downto 0);
signal enable_b_hi_256       : std_logic;
signal wbe_b_hi_256          : std_logic_vector(3 downto 0);
signal data_read_b_hi_256    : std_logic_vector(31 downto 0);
begin
process(clk)
begin
if rising_edge(clk) then
	address_a_reg <= address_a;
	address_b_reg <= address_b;
	end if;
end process;
data_read_a <= data_read_a_lo when (address_a_reg < x"0001000"&"00") else
data_read_a_hi when ((address_a_reg >= x"0001000"&"00") and (address_a_reg < x"0002000"&"00")) else 
data_read_a_lo_256 when ((address_a_reg >= x"0002000"&"00") and (address_a_reg < x"0003000"&"00")) else 
data_read_a_hi_256 when ((address_a_reg >= x"0003000"&"00") and (address_a_reg < x"0004000"&"00"));
data_read_b <= data_read_b_lo when (address_b_reg < x"0001000"&"00") else
data_read_b_hi when ((address_b_reg >= x"0001000"&"00") and (address_b_reg < x"0002000"&"00")) else
data_read_b_lo_256 when ((address_b_reg >= x"0002000"&"00") and (address_a_reg < x"0003000"&"00")) else 
data_read_b_hi_256 when ((address_b_reg >= x"0003000"&"00") and (address_b_reg< x"0004000"&"00"));
enable_a_lo <= enable_a when (address_a < x"0001000"&"00") else '0';
enable_b_lo <= enable_b when (address_b < x"0001000"&"00") else '0';
enable_a_hi <= enable_a when ((address_a >= x"0001000"&"00") and (address_a < x"0002000"&"00")) else '0';
enable_b_hi <= enable_b when ((address_b >= x"0001000"&"00") and (address_b < x"0002000"&"00")) else '0';
enable_a_lo_256 <= enable_a when ((address_a >= x"0002000"&"00") and (address_a < x"0003000"&"00")) else '0';
enable_b_lo_256 <= enable_b when ((address_b >= x"0002000"&"00") and (address_b < x"0003000"&"00")) else '0';
enable_a_hi_256 <= enable_a when ((address_a >= x"0003000"&"00") and (address_a < x"0004000"&"00")) else '0';
enable_b_hi_256 <= enable_b when ((address_b >= x"0003000"&"00") and (address_b < x"0004000"&"00")) else '0';
wbe_a_lo <= wbe_a when  enable_a_lo='1' else x"0";
wbe_a_hi <= wbe_a when  enable_a_hi='1' else x"0";
wbe_b_lo <= wbe_b when  enable_b_lo='1' else x"0";
wbe_b_hi <= wbe_b when  enable_b_hi='1' else x"0";
wbe_a_lo_256 <= wbe_a when  enable_a_lo_256='1' else x"0";
wbe_a_hi_256 <= wbe_a when  enable_a_hi_256='1' else x"0";
wbe_b_lo_256 <= wbe_b when  enable_b_lo_256='1' else x"0";
wbe_b_hi_256 <= wbe_b when  enable_b_hi_256='1' else x"0";



ram_bit_0_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"DA9918630DD2200000000000012800000040002000A106001180000000008007",
INIT_01 => X"80202100005CD2C7B4E6C1E566434955ED29B05AB311C477A91660C2B4D5208F",
INIT_02 => X"11840040D2AC24048604810082640D046B24CC461E01332121AD800087828206",
INIT_03 => X"080029800001E5202400B85242009129400A2A042000F22200808420C4108104",
INIT_04 => X"000FFF9D8F603C21282300100003000404F0100838008ED10C280E44011DA811",
INIT_05 => X"5000032408000000808000349D2934800010180000802B000060040012120000",
INIT_06 => X"40261C93C1345120821204AE0A41780DC6D01980827218422A0C004092B00A14",
INIT_07 => X"400AF9C0A003557C605D491DA48448900A020810000202AAEA922236141141A2",
INIT_08 => X"9030DA025E0900002300040002000840C204C2C131209008137028AD0779C23B",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF80C11F1127D082",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(0),        -- Port A data input
DOA(0)   => data_read_a_lo(0),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(0),        -- Port B data input
DOB(0)   => data_read_b_lo(0),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_1_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"C08451022808200000000000002000000000000010000C001108000000028002",
INIT_01 => X"22402100005000008490005046680400213C00142300E04080F4514BA066C00C",
INIT_02 => X"00000000000020044400010000C28410230CC4480000024000A1800182C12400",
INIT_03 => X"00001000000000000810440001002000802880040000A2020000800004000000",
INIT_04 => X"00006D858F602400280300100001400452000008000004A0000004A002090008",
INIT_05 => X"501000209000000080000020010008000090900090000B000000000048484000",
INIT_06 => X"09000900010410A082084002000002000012000214208008A890001284200000",
INIT_07 => X"4005010C10002000042028092400884080000000080A08222A22000200004009",
INIT_08 => X"947022015EA802000108121004000000090A458294C24001820004404205F012",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF81809307840190",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(1),        -- Port A data input
DOA(0)   => data_read_a_lo(1),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(1),        -- Port B data input
DOB(0)   => data_read_b_lo(1),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_2_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"C4804010026CA010101010110092D555550554161001447431116AAAAA820012",
INIT_01 => X"0A141D0A80440812841911980061967CA10E44C4000CB262012008C8B4780C08",
INIT_02 => X"100400000DD9AA5D050335002951264102C1C141491444444A90028282604143",
INIT_03 => X"82921220A28088500A92560801202412F06202040082080840808000E4110B00",
INIT_04 => X"42200020000040044004010208896AA03288101802A0242A0104843012480048",
INIT_05 => X"861A5082908814018000830A041400220C909115E12C4A02A00AA8054ACAD020",
INIT_06 => X"59510860140403E86A0AC8101AA88502590A401A542022AAAA0210378C24000B",
INIT_07 => X"010500130C048045913A20488481D851900022D048080090A2A0220280044209",
INIT_08 => X"B5013F1C742852CE43805274B40340150B9A8D46B4AE500242A910405294C091",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFFC8A0193716CC3A",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(2),        -- Port A data input
DOA(0)   => data_read_a_lo(2),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(2),        -- Port B data input
DOB(0)   => data_read_b_lo(2),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_3_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"C0C1002008E008110011001024C366666619989C00A105460141B33333020006",
INIT_01 => X"0004B50C84642830841112880080922C210C4480004812E055808C413181DC6C",
INIT_02 => X"1014001A2DD1BAA94D09640318C2C44822849440480EA80482208882C2050048",
INIT_03 => X"3183106A69989A5449B854A8102C241814A02200110008980280808005100940",
INIT_04 => X"02800040000040804084000020A9599012A1404041B024261084A4284A48426A",
INIT_05 => X"084C60828481CC880890A0020404028281A09081C02081418386630DCACBE422",
INIT_06 => X"5B410840148C02BA740ACA8100A00A283828400A542820800A90A6342866C040",
INIT_07 => X"0005020D0480604185022048040010518011018520110A2A2C208A1040220019",
INIT_08 => X"B000220C748E346521C072F0A541C38C199A8D46B4AE50018A0C004810148090",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF8D4015050C05A8",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(3),        -- Port A data input
DOA(0)   => data_read_a_lo(3),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(3),        -- Port B data input
DOB(0)   => data_read_b_lo(3),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_4_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"C0CB20AC108100111100001100FC78787806181894884518995E3C3C3C128002",
INIT_01 => X"081425AA60440802840100008184B200A108402040C21260028000C0C400122C",
INIT_02 => X"920406000DC124110442042878C2002022409101485E64140010200892014143",
INIT_03 => X"87840669E7D0189253BE47000009280008000000012E28805080601083130802",
INIT_04 => X"C800000000004084410000002A09B8651202020207C8240E8380941A3A480026",
INIT_05 => X"14308401842A3C60A30184200440000613808401C0020003971E190CC8C94422",
INIT_06 => X"1B750810100D02FD0008C2A0402D080011410A909028432604AB74B20028904A",
INIT_07 => X"0420400900004001142AA0480610B04390803784EC884A00090F984AC90E0119",
INIT_08 => X"044015114600F6E44900731CA503C63C19AA150A8C824001020B024202848090",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFFB5208A0F988902",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(4),        -- Port A data input
DOA(0)   => data_read_a_lo(4),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(4),        -- Port B data input
DOB(0)   => data_read_b_lo(4),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_5_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"CAC8380F010300111111110000D7807F8048181E94A84D60A555C03FC0120002",
INIT_01 => X"082025234054C8C69416C281E46C6D05A50DA0A0F217E665A82468C854801EAC",
INIT_02 => X"918425025D5524110746040A8752890040A491061F213021492C800087230206",
INIT_03 => X"6860699410016D322440A8DA0620950314200004212C10A25082501400108001",
INIT_04 => X"000FFFFD8F703C2168230012AAA207E424011018B8028E516C681E45831CB911",
INIT_05 => X"041007240429826183011006880D1004421104108202B1405161FD051010B800",
INIT_06 => X"02429C80C53D41A8DE1006824B604A05D690D122917A18678266086280B6004A",
INIT_07 => X"0406B3CD3480653D617FE11C8680A882100228620C804220481000302CD14002",
INIT_08 => X"0FB5FF3F7A550B6269C0046C8500294342B41A0D190C8001837B0AED157C8239",
INIT_09 => X"00000000000000000000000000000000000005FFFFFFFFFFFFC1E3BE7EA3DDBF",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(5),        -- Port A data input
DOA(0)   => data_read_a_lo(5),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(5),        -- Port B data input
DOB(0)   => data_read_b_lo(5),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_6_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"C0CC0708E06000111111111100D7FF80000FE01E10200D600155FFC000000002",
INIT_01 => X"0800250C41440812842112C018619238A10844B00C14B062001008C094001C2C",
INIT_02 => X"1204201000902411040204000042000008809100000220000020000080010002",
INIT_03 => X"400010080000000208585481800020D004200004000208080082000000121000",
INIT_04 => X"000000005086000044000A02AAA8401432890000000024204000842102480108",
INIT_05 => X"0010008180010020889110006000C2A441A090040200000012000068CA4B4400",
INIT_06 => X"5901080010040128000A428008200800101000008020002D2B89083200220000",
INIT_07 => X"0020410910004041000220480490005080810006E888081880A80040C9000219",
INIT_08 => X"B541FF1F3E2802610100721081840200198A8542A4A250010008000000048090",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF9CE19F3B9FDCBA",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(6),        -- Port A data input
DOA(0)   => data_read_a_lo(6),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(6),        -- Port B data input
DOB(0)   => data_read_b_lo(6),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_7_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"C48C031862648011111111110000000000000000840844008100000000100006",
INIT_01 => X"0804258020440802842002C012090410A10000B009000060000000C00000000C",
INIT_02 => X"100400100090A4110402042001D2040000809100410220144820000090210042",
INIT_03 => X"40001008001210084840108880600C4034200000000000098080000000100000",
INIT_04 => X"00000000208000484200860AAAA9401100810000000065204001852102CA0428",
INIT_05 => X"00100099010100408384820A241440920A310501C10AC0400200000802830600",
INIT_06 => X"40014A20340D27F32203201048088808011040028029002A8802082200220000",
INIT_07 => X"15010709148C40401108A0CA0E83B81A1001A00404204000000800000080C000",
INIT_08 => X"00000000000000990980406C748102002030D86C382C10850003920010048194",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF94000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(7),        -- Port A data input
DOA(0)   => data_read_a_lo(7),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(7),        -- Port B data input
DOB(0)   => data_read_b_lo(7),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_8_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"D08800000008001111111111000000000000000084884C009100000000100002",
INIT_01 => X"081025A001440802842002C000090410A10800B000140062000001C80080000C",
INIT_02 => X"100400120000A4110542042801520000008011010102200048200000C0210102",
INIT_03 => X"50000008080202000050448984202CD214200004000208088080000000301000",
INIT_04 => X"800000021000010244405806AAA8001032010000400000005000000102004000",
INIT_05 => X"0010009180010048838000026404C08002B38480800290500280000848CD4600",
INIT_06 => X"09240010048900A0024840A14009080001504880800800040000083200260000",
INIT_07 => X"04000309148040401100A0000600A9429800300404094A0888A8001000804909",
INIT_08 => X"2A303F1F5850050749C052F804C40200092A150A948A44210003020010048000",
INIT_09 => X"00000000000000000000000000000000000005FFFFFFFFFFFFF52080369848B3",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(8),        -- Port A data input
DOA(0)   => data_read_a_lo(8),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(8),        -- Port B data input
DOB(0)   => data_read_b_lo(8),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_9_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"C4C800100204810000000000000000000000000000000C001100000000000002",
INIT_01 => X"000025AAA0440812840112C000609228A10044B00000B060000008C014000C2C",
INIT_02 => X"B20427920090A4110542042800C2046008C000000002641002302002D2014003",
INIT_03 => X"5000100808000A10085044800000281004200004012E088850827814C2B20003",
INIT_04 => X"CAA0006000104084018401400000401032090000400000A0500010A102014008",
INIT_05 => X"0410008384290028881100000000022400B38084800000101280006548CCFA22",
INIT_06 => X"09640110008011A0024840A10809080801500A8000008221202008328026004B",
INIT_07 => X"C0204309148040401008200164108940808000040089083888A1005008804B09",
INIT_08 => X"97F13F36608800010140121004400200090A058284C244210000000200848002",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF98813550204088",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(9),        -- Port A data input
DOA(0)   => data_read_a_lo(9),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(9),        -- Port B data input
DOB(0)   => data_read_b_lo(9),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_10_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"C4C800100264811111111111000000000000000084884C009100000000100002",
INIT_01 => X"081025A360440812840112C000609228A10044B00000B060000808C014000C2C",
INIT_02 => X"100400120010A411054204280152000000801101010220104820000090210102",
INIT_03 => X"4000000800000810004800880020040014200000052C00885080000000100000",
INIT_04 => X"4AA000600010408441840142AAA8001400090000000020004000800102400000",
INIT_05 => X"04100082042900408B900002040402A0030004048002C0400200002D8001BC22",
INIT_06 => X"12650010140900A0040080204001080800404AA010080020200008028026014B",
INIT_07 => X"040000091000404001008040060030031001200404084A3880A8000000808310",
INIT_08 => X"3B0568176850000109C0206C040002001030180C180C00010003024210008080",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF9DC39405BE0525",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(10),        -- Port A data input
DOA(0)   => data_read_a_lo(10),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(10),        -- Port B data input
DOB(0)   => data_read_b_lo(10),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_11_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"C2880203B0600020202020200000000000400000000004000100000000000006",
INIT_01 => X"0824250C40448882840602C168004100A10180B0B4004064000000C00000000C",
INIT_02 => X"1104000010042411060204000042010000801104540220240024000080010042",
INIT_03 => X"4000088800004100204000930200018104200000000000028080000000100000",
INIT_04 => X"000355134A4410692C6086140000001000010000100000C0402000C103962001",
INIT_05 => X"001002300001000080000000C801900000000000800000000220000000000000",
INIT_06 => X"00025600802060A0000000020000080084000000005300000004080200B20000",
INIT_07 => X"0004248920084018401441960402000000000004000000000000000004800000",
INIT_08 => X"0181683650100000010000000400020020000000000000850300808C0518832D",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF9CE13045200411",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(11),        -- Port A data input
DOA(0)   => data_read_a_lo(11),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(11),        -- Port B data input
DOB(0)   => data_read_b_lo(11),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_12_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"C88A1F83F000020022002200020000000040004000000480012A000000000002",
INIT_01 => X"081025A00054C8C6940202C06F000801A50080B037810465AA0C60C00000008C",
INIT_02 => X"110400125014A4110746042880428100008411010603302100248000C0030106",
INIT_03 => X"4000018800010400044000DB822095C1142000002000102B8080000000100000",
INIT_04 => X"000F9B1B4E8208012E6294080002001000011010200000904800008103978000",
INIT_05 => X"001003BC0101000980000006E80DD00000000080800021000240000000000000",
INIT_06 => X"0002568081A070A08000000300004A04C0801100005380400000084200B60000",
INIT_07 => X"C000820D24806530004001976400000000028004000100000000000000910000",
INIT_08 => X"A4C48D264409000101C0000004C002400000000000000001806000000400832E",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF9C0025401700A6",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(12),        -- Port A data input
DOA(0)   => data_read_a_lo(12),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(12),        -- Port B data input
DOB(0)   => data_read_b_lo(12),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_13_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"C6CC00100206811133331111580000000000010084084480A320000000100002",
INIT_01 => X"083425A020C40812840552811060DB28A10144A08801F060003809C014000C2C",
INIT_02 => X"114400321014A4110742042803520800408011054102201449240000D4210342",
INIT_03 => X"4800000800016D300048A0880020041014200001832C10A85080020000104400",
INIT_04 => X"5AACE2ED56765C846DC75B56AAAA0010A40901093800EB004C298B010240A800",
INIT_05 => X"04100381042900489B100086080C122003214484800290400A60042D9091BE22",
INIT_06 => X"12410180759900A00430800142004804868051000008004010000822003600CA",
INIT_07 => X"0412B2C9048040306145C0400608308310412804044140104010002006818612",
INIT_08 => X"0FB5F7397E30000109C0246C04401A0052341A8D194C821101530AA515688080",
INIT_09 => X"00000000000000000000000000000000000005FFFFFFFFFFFFE0E7BE7F83DDBF",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(13),        -- Port A data input
DOA(0)   => data_read_a_lo(13),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(13),        -- Port B data input
DOB(0)   => data_read_b_lo(13),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_14_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"C088000001600222000000005A0000000040014000000480012A000000000002",
INIT_01 => X"08002500004408028400828000600000A10020A00000A060000000C00000000C",
INIT_02 => X"1084000000002411040204000042000000801100000220000028000081010002",
INIT_03 => X"4000000800000000004000800000000004200000000000000080000000108000",
INIT_04 => X"00000D8731063940000210140002001000010000000000004000000102000000",
INIT_05 => X"0010000000010000800000000000000000000000000000000200000000000000",
INIT_06 => X"0000000000000020000000000000080100000000000000000000080200220000",
INIT_07 => X"000000090000400C000000000400000000000004000000000000000000800000",
INIT_08 => X"BF45FF1F3CC80000110000000000020000000000000000010000000000008000",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF81E39533BF4DBE",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(14),        -- Port A data input
DOA(0)   => data_read_a_lo(14),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(14),        -- Port B data input
DOB(0)   => data_read_b_lo(14),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_15_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"C08800000060022222222222000000000040000000000400010A000000000002",
INIT_01 => X"08002500004408028400028000000000A10000A000000060000800C00000000C",
INIT_02 => X"1004000000002411040204000042000000A01102160220000020000080010002",
INIT_03 => X"4000298800000000244008800000000004200000000000000080000000100000",
INIT_04 => X"000000008000042B242188000002001000010000000000514000004502000011",
INIT_05 => X"0010000000010000800000000000000000000000000010000200000000000000",
INIT_06 => X"0000000000000020000004000040080000000000000010000004080200220000",
INIT_07 => X"0000000900004000001000008400000000000804000000000000000000800000",
INIT_08 => X"0000000000000000010000000000020000000000000000010000000000008001",
INIT_09 => X"00000000000000000000000000000000000005FFFFFFFFFFFF80000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(15),        -- Port A data input
DOA(0)   => data_read_a_lo(15),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(15),        -- Port B data input
DOB(0)   => data_read_b_lo(15),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_16_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"05104816EA00C199999999998B82D55555055577C0000675C3816AAAAAB80003",
INIT_01 => X"8014102000081213688B1862C400120ADA22C61962221218A90010E0957F0E0E",
INIT_02 => X"C200BAC50001061C8901300A2C0980A50085C801003641100400A00980206443",
INIT_03 => X"E2D5423CB284889002E20281C02900E8CC00000340A9401040162E6680824001",
INIT_04 => X"2FDAC651494D654F010FCA0208282AB240330303829FBF0A61DAFF19988017A2",
INIT_05 => X"252A5018058B9611A81110887160E2205004010210480142D30AA9290000198B",
INIT_06 => X"0050400484141401508000004500050248210008000041000000BC86424A9650",
INIT_07 => X"0208023485003A048820088005000200124342D66130400000008809D0C62220",
INIT_08 => X"1D75310E66E4584AA2AC002B005A631500000000001000005485220000000102",
INIT_09 => X"00000000000000000000000000000000000005FFFFFFFFFFFF80C3183DBECD8E",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(16),        -- Port A data input
DOA(0)   => data_read_a_lo(16),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(16),        -- Port B data input
DOB(0)   => data_read_b_lo(16),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_17_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"4F74BF57E6E587FFFFFFFFFF92D71999998E665DC000E1D9E8758CCCCCF80000",
INIT_01 => X"2ADE30F033C915094A13393EDEF4B2265284CE4B6F40B85001AE0AB1FA003513",
INIT_02 => X"664123B786736A3991E3A47C1D59727F83855D59A1AC21CA6C30AAA2F8F149E3",
INIT_03 => X"01EF407061DE98DF4182021FC45117E22A0888D2C6F8E0FE6823B275CDE77725",
INIT_04 => X"EDD90A855E9396159B5AEBFD777C19EBC03E272701DDBF0600D8FF080FE617A2",
INIT_05 => X"79639AE01E360FDFCF3BEBFFF17FEE5BBC021EE7D7EDBD79F0067A7300009CCD",
INIT_06 => X"005379675FEBE2F7E860285FE282B5A25822E00003FF001F9FEBA08437291FFC",
INIT_07 => X"D2780225C3B59F058DB28BFEEC394102168741D823F3F0040443B8C558020EE0",
INIT_08 => X"EAB0400D64A8399B47F1000937F4E00D0020100800010630ECAF77105801B3FD",
INIT_09 => X"00000000000000000000000000000000000005FFFFFFFFFFFF80203778BE0864",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(17),        -- Port A data input
DOA(0)   => data_read_a_lo(17),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(17),        -- Port B data input
DOB(0)   => data_read_b_lo(17),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_18_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"80900040060040000000000040039E1E1E0F80060E1C067E2F81CF0F0F000003",
INIT_01 => X"82500F0000100211A6110064200002886984501A10005048A99041D0557F0A28",
INIT_02 => X"C0404B0000108804C04211220424A28000C0804940226454001080009001A502",
INIT_03 => X"6078001C3080000000EB02801129001CDC40000100810011D008380302004002",
INIT_04 => X"40A662F955E7094500A5D54008A007F028431018808040026081000988000002",
INIT_05 => X"862CE019418B82203B5414007000E000436D2000000200044301F98CA1A12F12",
INIT_06 => X"36888606A41514081581900415241410202980184100E18000002CA9620A9000",
INIT_07 => X"04000A360D029582000000008204360921008066240000000104000060C2B094",
INIT_08 => X"274051317664099AEB04286408082303969048A41A4C084AD080000050000001",
INIT_09 => X"00000000000000000000000000000000000005FFFFFFFFFFFF8026A81B2A5022",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(18),        -- Port A data input
DOA(0)   => data_read_a_lo(18),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(18),        -- Port B data input
DOB(0)   => data_read_b_lo(18),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_19_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"00014020080007FFFFFFFFFF82D7E01FE008005FC000E7E1C1F5F00FF0380003",
INIT_01 => X"0000000000000004108800000000000104220004006A80000000000000000000",
INIT_02 => X"00009440000005400C0000020400000000000000002200000020000940000000",
INIT_03 => X"6040001C3080000000E20280000900000C000000000000000014440010000010",
INIT_04 => X"40018F03201F7C056400DE0C82A8007000030000808000026080000988000002",
INIT_05 => X"0090040000038200000000000000000000000000000000004300180000003022",
INIT_06 => X"00000000000000000000000000000200000000000000000000002C820C6E9000",
INIT_07 => X"0000000000002000000000000000000000000046200000000000000040C20000",
INIT_08 => X"520020232E240844100800000000230100000000000000000000000000000000",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF80A1321EAA8140",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(19),        -- Port A data input
DOA(0)   => data_read_a_lo(19),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(19),        -- Port B data input
DOB(0)   => data_read_b_lo(19),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_20_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"00000000000007FFFFFFFFFF82D7FFE0000FF85FC000E7E1C1F5FFF000380003",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000027C00000180004400007E00000000000000000000",
INIT_03 => X"E7C6867DF780000093E60380000900000C000000000000000000000000000000",
INIT_04 => X"1AA01182938901EA66400042A800BFF00003000087E2008EE386009BB8190046",
INIT_05 => X"000000000003BE0000000000000000240000430200400003CF1FF80000040140",
INIT_06 => X"00000000000000000000000000000000000000000000000000007C80000A9000",
INIT_07 => X"5200000000000000002008012D000000404007E6E000000000000008C3CE0000",
INIT_08 => X"80800812380CF801004001031202F73F00000000001120000000000000000402",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF810487600C0004",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(20),        -- Port A data input
DOA(0)   => data_read_a_lo(20),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(20),        -- Port B data input
DOB(0)   => data_read_b_lo(20),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_21_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"4410801502168D555555555520D7FFFFFF90001F8000057F8D55FFFFFFF00002",
INIT_01 => X"8880BE000439376128C090A2E09240284A30242970600098540084F0017FA04B",
INIT_02 => X"0511481A600817F8800B64437D11428202208800047EF900C80488000085480F",
INIT_03 => X"E7D80EFFF7CC20E513E60BF2044D11000C800040108C0022022B789ECAA60068",
INIT_04 => X"4AA339708A60102128A000100000BFF0000366668780201EE380801FFD140436",
INIT_05 => X"E82F02201003FE424043142491092829200010042020200BC71FF8010000B822",
INIT_06 => X"200A944880344004D8000806010285A00A09801841D2610A8A8A7E87620AD004",
INIT_07 => X"0400821589B43102800083140200010000811FE7E02200000516A82CC1EE0000",
INIT_08 => X"0F35FF3F5E36FDFE78800068F142E7BF0020100800000000F056102100480638",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF80E7BE7F83FDBF",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(21),        -- Port A data input
DOA(0)   => data_read_a_lo(21),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(21),        -- Port B data input
DOB(0)   => data_read_b_lo(21),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_22_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"6CD0E84501520D555555555524FFFFFFFF90009F8001C17F8055FFFFFFF00000",
INIT_01 => X"0A94BEAFE77D3C314A43D337A45241685290F4CFD22090F85C488C03D57FAC62",
INIT_02 => X"F6157F9A78589FFDD14B756901537001E028C4415900AB14E83DA22A50A5694B",
INIT_03 => X"0827A802001090086000807A1124150890A222023DA002AA52AE78DFEAF6314B",
INIT_04 => X"4AAFBB390A30488569A60142AAAA000304287676087620400446A00045541AC0",
INIT_05 => X"AB7FFAA014A840490B55B62E915D2A21A204059434223328000007AC10111C26",
INIT_06 => X"004B1C0A95B9400000D0060740E01FB25402400206DA180A8A9A020766044540",
INIT_07 => X"0561124C8480FA0545630B5480B002881117300105A340926202228100302A02",
INIT_08 => X"BFC5793F7CEA05FF48C00408F1C800800084422111088C6164DF1284170066A9",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF81E7BD7BBEDDAE",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(22),        -- Port A data input
DOA(0)   => data_read_a_lo(22),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(22),        -- Port B data input
DOB(0)   => data_read_b_lo(22),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_23_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"8A99D0720284A800000000006A000000005FFF400C1804002D00000000000002",
INIT_01 => X"A00080000420E3E7BC8241B640909201EF20906F206006E5F4E2B4F0200040CD",
INIT_02 => X"A39050087D451C8190084003FC04B16802C11910167EDC8180382AA20006800C",
INIT_03 => X"E7C02FFFF780000017EE0BA0044D00122CC888D0700CC010020D0094F2A38B73",
INIT_04 => X"000CCAAD86201C00280300100000BFF02003404087818A5FE3980A5FF8000017",
INIT_05 => X"EB7FFD010003FF226006CA081110001A0921000141088043C71FFF8180809200",
INIT_06 => X"121000064104000084008000160696210A020000002000800004FEA2020AD004",
INIT_07 => X"100002134014B008841000000801100108000FF7E00000000504880EE5FE8010",
INIT_08 => X"000000000006F800200020040002E7FF1200000008000002F834000000000000",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF80000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(23),        -- Port A data input
DOA(0)   => data_read_a_lo(23),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(23),        -- Port B data input
DOB(0)   => data_read_b_lo(23),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_24_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000D555555555524FFFFFFFF90009F8001C57F8155FFFFFFF00002",
INIT_01 => X"0000800004202020000000000000000000000000000000805400840000000040",
INIT_02 => X"0010800820001080000840037C00000000000000007E88008380000000040008",
INIT_03 => X"E7C0067FF780000013E603A0000D00000C800000100000000210008001000040",
INIT_04 => X"000065E581003800000200100000BFF0000340408780000EE380001BF8000006",
INIT_05 => X"040000000003FE0000000000000000000000000000000003C71FFF8000003000",
INIT_06 => X"00000000000000000000000000000000000000000000000000007E80098AD00A",
INIT_07 => X"00000000000004800000000000000000000007E7E000000001048808C1EE0000",
INIT_08 => X"8EB2CEAF580EF800100000000002E7BF00000000000000000000000000000000",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF806D2D66331814",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(24),        -- Port A data input
DOA(0)   => data_read_a_lo(24),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(24),        -- Port B data input
DOB(0)   => data_read_b_lo(24),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_25_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000D555555555524FFFFFFFF90009F8001C57F8155FFFFFFF00002",
INIT_01 => X"0000800004202020000000000000000000000000000000805400840000000040",
INIT_02 => X"0010000820001080000840037C00028600040000007E88008000000000040008",
INIT_03 => X"E7D8067FF7DC38FD53E623A0000D00000C800000100000000200008000000040",
INIT_04 => X"800000600C600421202100000000BFF0000340408780040EE380041BF8080426",
INIT_05 => X"000000000003FE0000000000000000645202140402000013D71FFF890105B400",
INIT_06 => X"200080600000065F7801285001000000A02980184100610000007E80000AD000",
INIT_07 => X"0400B0C0092001022015C00802002102008007E7E000000001148868C9EE0000",
INIT_08 => X"14B3C80EA076F800880701680006E7BF0230180C100C0000002200A541491010",
INIT_09 => X"00000000000000000000000000000000000003FFFFFFFFFFFF80883A7B42C803",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(25),        -- Port A data input
DOA(0)   => data_read_a_lo(25),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(25),        -- Port B data input
DOB(0)   => data_read_b_lo(25),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_26_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"85F820440E61E5DDDDDDDDDD81D7FFFFFF8FFE3FDEBCEF7FDFD5FFFFFFF80007",
INIT_01 => X"AA5E3FF033CC1A1BA4993AAC8064328EE9265EAA400ABA7000401AC1DE00573E",
INIT_02 => X"F645FFF78F73EF7DDDE3B57E7C6F72BF89C15D49E0FE675E24302AA9F8D1E5E3",
INIT_03 => X"E7FFD67DF7DE1ADFDBEF578C5479263E7E600053CEFDE25C78BFFE7FDFF77F3F",
INIT_04 => X"FFF000600019C294D19C21E3FFFDFFFBFAFF272787FF302EE3D6F03BBE6057EE",
INIT_05 => X"FFFFFCC1DABFBFFEFF7FFFFB1136267FFFFFFFE7D7EFDE7FFF1FFBFFEBEFFFFF",
INIT_06 => X"7FD9A0671ECB87FF7FEBFADDFDAEBDB23939E23AD10C6B9D1D69FCBF7F6F9FBE",
INIT_07 => X"17794B3BCFB7DA839D8AAA600FBDFF5BFFC567FEEFF3F234094F98D9DBCEFEFD",
INIT_08 => X"D082EF0B3EACFFFFFFFF7BFFFFFFF73F9DBA9D6EAEBF7E7B7C8F77525A85B4C0",
INIT_09 => X"00000000000000000000000000000000000003FFFFFFFFFFFF800B354D1138DC",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(26),        -- Port A data input
DOA(0)   => data_read_a_lo(26),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(26),        -- Port B data input
DOB(0)   => data_read_b_lo(26),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_27_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"11200008002844CCCCCCCCCC80D7FFFFFF8FFE1F5AB4AB7F5ED5FFFFFFEA8015",
INIT_01 => X"080A0E5012800008002029000029049200080A4000142822000002090A800110",
INIT_02 => X"4441D8370DC3416110A004547C8854AB88011100A0FC000A040022202A1000A0",
INIT_03 => X"97EF9671EFDC1ADDDB97570404512A062A000057CA7F0844783D024B19456E38",
INIT_04 => X"7FF000600019C294D19C21E3FFFDFFEE9A8E252547F7102E93D6603A3C2056EE",
INIT_05 => X"AFCF7842C23E3FD65FFECAC9041202FB2ADCE767554BCC6FEC9FFBBF6B6BFDFF",
INIT_06 => X"6DFCA0760E43875F7BAB7AF4EDAF80B83959EAB8D10463B03008F099E10914AB",
INIT_07 => X"1654452153BC0AC3998AA2200B2BAE5AF54467F8EF78FA3C88E88891D30E774D",
INIT_08 => X"4A825C88A220FFFFCC7F5AFBF93BF43F2DAA956AA6BB7AD42E0FD35A18942440",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF80F91049E10840",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(27),        -- Port A data input
DOA(0)   => data_read_a_lo(27),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(27),        -- Port B data input
DOB(0)   => data_read_b_lo(27),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_28_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"4128400000606088888888888000000000000000420526004380000000080003",
INIT_01 => X"220A20501184080808802A90006000C202200AA40000A820004A02822A004110",
INIT_02 => X"B24427A5000A440440A21114001A00002288C440A980220A0CA1088828B120A2",
INIT_03 => X"0000000000008000800100041110020C8222220186D182D428827A14E2B25403",
INIT_04 => X"B550000000098210901820A15554000988240303000014000000440000280000",
INIT_05 => X"40900040569400B4342934E101420804D04A727222611E1438000012202401D9",
INIT_06 => X"048028000A46800001601000A00008000002200206A4081A9A92000A040101A0",
INIT_07 => X"03310028020040000CA00828019805006CC0500802D2B086264222463A001C44",
INIT_08 => X"0501710016D0000034380903083410000400400012112631000041104A014050",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF809A223208608B",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(28),        -- Port A data input
DOA(0)   => data_read_a_lo(28),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(28),        -- Port B data input
DOB(0)   => data_read_b_lo(28),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_29_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A5F0A0540E75C5DDDDDDDDDD81000000000FFE20C60C677EC3D5FFFFFFD80003",
INIT_01 => X"805E1FFFF1C81619E659392E8076B2AE79965E4B402AB858000A0A71FF7FBF3B",
INIT_02 => X"E240FFF78F72EB588DE1A03E016D627D81408809E0FE455E66100001F850C5E1",
INIT_03 => X"E037C67C104E00C793E9038C403806345E4000438F5D604C281FFE7FDFA35F3F",
INIT_04 => X"FFF0000000098210901820A15554BFFBE8572323807E340EE046F41B866813C6",
INIT_05 => X"B8AF84C14A1781FEBF7B77D31026246DDD6B6EE3D3C59C1FFF0003F2A0A4BFFB",
INIT_06 => X"16C9282F1ACE82F32560B25DB402B59200202000022C001515697C2D7A6F8FFE",
INIT_07 => X"02380A338E97988008800068051D550176C167FE03D1B0140545104DFBC09EF4",
INIT_08 => X"2E77BF3F7E2405FFF7FA292FFFF6F700941008040A15263A748175100800B0D0",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF83D7BC7787BF7E",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(29),        -- Port A data input
DOA(0)   => data_read_a_lo(29),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(29),        -- Port B data input
DOB(0)   => data_read_b_lo(29),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_30_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000222222222225A00000000000140000000800020000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"DF83FF2F7CF80000000000000000000000000000000000000000000000000000",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF80FF3F7F3BF8DF",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(30),        -- Port A data input
DOA(0)   => data_read_a_lo(30),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(30),        -- Port B data input
DOB(0)   => data_read_b_lo(30),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_31_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"60008010001404444444444400D7FFFFFF8FFE1F0810817F0C55FFFFFFE00000",
INIT_01 => X"08800E0FC20105004A40000200128020129000010020000800000030017FA801",
INIT_02 => X"4401D8120D410161100004407D1050EB80011110017C00804A00222200200800",
INIT_03 => X"87EF8671E7DC18DD5386030004410002280888D2492C0080503D004B19452A38",
INIT_04 => X"4AA000600010408441840142AAA8BFE2000A242407F7000E83D6201A3C0016E6",
INIT_05 => X"AF4F7800042A3F424B56CA080010027B2A040505450A806BC41FFBAD0101BC26",
INIT_06 => X"2058806C0401065F78812A5045A680B03809C018418061800000F0816108144A",
INIT_07 => X"1440000141B40A83810282000A21220A110427E0E520401000008881C10E2200",
INIT_08 => X"000000000000FDFFC8470068F10AE43F00A05028100808402C0F120010000400",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF80000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(31),        -- Port A data input
DOA(0)   => data_read_a_lo(31),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(31),        -- Port B data input
DOB(0)   => data_read_b_lo(31),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_0_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"DA9918630DD2200000000000012800000040002000A106001180000000008007",
INIT_01 => X"80202100005CD2C7B4E6C1E566434955ED29B05AB311C477A91660C2B4D5208F",
INIT_02 => X"11840040D2AC24048604810082640D046B24CC461E01332121AD800087828206",
INIT_03 => X"080029800001E5202400B85242009129400A2A042000F22200808420C4108104",
INIT_04 => X"000FFF9D8F603C21282300100003000404F0100838008ED10C280E44011DA811",
INIT_05 => X"5000032408000000808000349D2934800010180000802B000060040012120000",
INIT_06 => X"40261C93C1345120821204AE0A41780DC6D01980827218422A0C004092B00A14",
INIT_07 => X"400AF9C0A003557C605D491DA48448900A020810000202AAEA922236141141A2",
INIT_08 => X"9030DA025E0900002300040002000840C204C2C131209008137028AD0779C23B",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF80C11F1127D082",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(0),        -- Port A data input
DOA(0)   => data_read_a_hi(0),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(0),        -- Port B data input
DOB(0)   => data_read_b_hi(0),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_1_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"C08451022808200000000000002000000000000010000C001108000000028002",
INIT_01 => X"22402100005000008490005046680400213C00142300E04080F4514BA066C00C",
INIT_02 => X"00000000000020044400010000C28410230CC4480000024000A1800182C12400",
INIT_03 => X"00001000000000000810440001002000802880040000A2020000800004000000",
INIT_04 => X"00006D858F602400280300100001400452000008000004A0000004A002090008",
INIT_05 => X"501000209000000080000020010008000090900090000B000000000048484000",
INIT_06 => X"09000900010410A082084002000002000012000214208008A890001284200000",
INIT_07 => X"4005010C10002000042028092400884080000000080A08222A22000200004009",
INIT_08 => X"947022015EA802000108121004000000090A458294C24001820004404205F012",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF81809307840190",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(1),        -- Port A data input
DOA(0)   => data_read_a_hi(1),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(1),        -- Port B data input
DOB(0)   => data_read_b_hi(1),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_2_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"C4804010026CA010101010110092D555550554161001447431116AAAAA820012",
INIT_01 => X"0A141D0A80440812841911980061967CA10E44C4000CB262012008C8B4780C08",
INIT_02 => X"100400000DD9AA5D050335002951264102C1C141491444444A90028282604143",
INIT_03 => X"82921220A28088500A92560801202412F06202040082080840808000E4110B00",
INIT_04 => X"42200020000040044004010208896AA03288101802A0242A0104843012480048",
INIT_05 => X"861A5082908814018000830A041400220C909115E12C4A02A00AA8054ACAD020",
INIT_06 => X"59510860140403E86A0AC8101AA88502590A401A542022AAAA0210378C24000B",
INIT_07 => X"010500130C048045913A20488481D851900022D048080090A2A0220280044209",
INIT_08 => X"B5013F1C742852CE43805274B40340150B9A8D46B4AE500242A910405294C091",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFFC8A0193716CC3A",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(2),        -- Port A data input
DOA(0)   => data_read_a_hi(2),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(2),        -- Port B data input
DOB(0)   => data_read_b_hi(2),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_3_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"C0C1002008E008110011001024C366666619989C00A105460141B33333020006",
INIT_01 => X"0004B50C84642830841112880080922C210C4480004812E055808C413181DC6C",
INIT_02 => X"1014001A2DD1BAA94D09640318C2C44822849440480EA80482208882C2050048",
INIT_03 => X"3183106A69989A5449B854A8102C241814A02200110008980280808005100940",
INIT_04 => X"02800040000040804084000020A9599012A1404041B024261084A4284A48426A",
INIT_05 => X"084C60828481CC880890A0020404028281A09081C02081418386630DCACBE422",
INIT_06 => X"5B410840148C02BA740ACA8100A00A283828400A542820800A90A6342866C040",
INIT_07 => X"0005020D0480604185022048040010518011018520110A2A2C208A1040220019",
INIT_08 => X"B000220C748E346521C072F0A541C38C199A8D46B4AE50018A0C004810148090",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF8D4015050C05A8",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(3),        -- Port A data input
DOA(0)   => data_read_a_hi(3),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(3),        -- Port B data input
DOB(0)   => data_read_b_hi(3),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_4_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"C0CB20AC108100111100001100FC78787806181894884518995E3C3C3C128002",
INIT_01 => X"081425AA60440802840100008184B200A108402040C21260028000C0C400122C",
INIT_02 => X"920406000DC124110442042878C2002022409101485E64140010200892014143",
INIT_03 => X"87840669E7D0189253BE47000009280008000000012E28805080601083130802",
INIT_04 => X"C800000000004084410000002A09B8651202020207C8240E8380941A3A480026",
INIT_05 => X"14308401842A3C60A30184200440000613808401C0020003971E190CC8C94422",
INIT_06 => X"1B750810100D02FD0008C2A0402D080011410A909028432604AB74B20028904A",
INIT_07 => X"0420400900004001142AA0480610B04390803784EC884A00090F984AC90E0119",
INIT_08 => X"044015114600F6E44900731CA503C63C19AA150A8C824001020B024202848090",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFFB5208A0F988902",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(4),        -- Port A data input
DOA(0)   => data_read_a_hi(4),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(4),        -- Port B data input
DOB(0)   => data_read_b_hi(4),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_5_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"CAC8380F010300111111110000D7807F8048181E94A84D60A555C03FC0120002",
INIT_01 => X"082025234054C8C69416C281E46C6D05A50DA0A0F217E665A82468C854801EAC",
INIT_02 => X"918425025D5524110746040A8752890040A491061F213021492C800087230206",
INIT_03 => X"6860699410016D322440A8DA0620950314200004212C10A25082501400108001",
INIT_04 => X"000FFFFD8F703C2168230012AAA207E424011018B8028E516C681E45831CB911",
INIT_05 => X"041007240429826183011006880D1004421104108202B1405161FD051010B800",
INIT_06 => X"02429C80C53D41A8DE1006824B604A05D690D122917A18678266086280B6004A",
INIT_07 => X"0406B3CD3480653D617FE11C8680A882100228620C804220481000302CD14002",
INIT_08 => X"0FB5FF3F7A550B6269C0046C8500294342B41A0D190C8001837B0AED157C8239",
INIT_09 => X"00000000000000000000000000000000000005FFFFFFFFFFFFC1E3BE7EA3DDBF",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(5),        -- Port A data input
DOA(0)   => data_read_a_hi(5),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(5),        -- Port B data input
DOB(0)   => data_read_b_hi(5),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_6_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"C0CC0708E06000111111111100D7FF80000FE01E10200D600155FFC000000002",
INIT_01 => X"0800250C41440812842112C018619238A10844B00C14B062001008C094001C2C",
INIT_02 => X"1204201000902411040204000042000008809100000220000020000080010002",
INIT_03 => X"400010080000000208585481800020D004200004000208080082000000121000",
INIT_04 => X"000000005086000044000A02AAA8401432890000000024204000842102480108",
INIT_05 => X"0010008180010020889110006000C2A441A090040200000012000068CA4B4400",
INIT_06 => X"5901080010040128000A428008200800101000008020002D2B89083200220000",
INIT_07 => X"0020410910004041000220480490005080810006E888081880A80040C9000219",
INIT_08 => X"B541FF1F3E2802610100721081840200198A8542A4A250010008000000048090",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF9CE19F3B9FDCBA",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(6),        -- Port A data input
DOA(0)   => data_read_a_hi(6),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(6),        -- Port B data input
DOB(0)   => data_read_b_hi(6),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_7_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"C48C031862648011111111110000000000000000840844008100000000100006",
INIT_01 => X"0804258020440802842002C012090410A10000B009000060000000C00000000C",
INIT_02 => X"100400100090A4110402042001D2040000809100410220144820000090210042",
INIT_03 => X"40001008001210084840108880600C4034200000000000098080000000100000",
INIT_04 => X"00000000208000484200860AAAA9401100810000000065204001852102CA0428",
INIT_05 => X"00100099010100408384820A241440920A310501C10AC0400200000802830600",
INIT_06 => X"40014A20340D27F32203201048088808011040028029002A8802082200220000",
INIT_07 => X"15010709148C40401108A0CA0E83B81A1001A00404204000000800000080C000",
INIT_08 => X"00000000000000990980406C748102002030D86C382C10850003920010048194",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF94000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(7),        -- Port A data input
DOA(0)   => data_read_a_hi(7),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(7),        -- Port B data input
DOB(0)   => data_read_b_hi(7),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_8_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"D08800000008001111111111000000000000000084884C009100000000100002",
INIT_01 => X"081025A001440802842002C000090410A10800B000140062000001C80080000C",
INIT_02 => X"100400120000A4110542042801520000008011010102200048200000C0210102",
INIT_03 => X"50000008080202000050448984202CD214200004000208088080000000301000",
INIT_04 => X"800000021000010244405806AAA8001032010000400000005000000102004000",
INIT_05 => X"0010009180010048838000026404C08002B38480800290500280000848CD4600",
INIT_06 => X"09240010048900A0024840A14009080001504880800800040000083200260000",
INIT_07 => X"04000309148040401100A0000600A9429800300404094A0888A8001000804909",
INIT_08 => X"2A303F1F5850050749C052F804C40200092A150A948A44210003020010048000",
INIT_09 => X"00000000000000000000000000000000000005FFFFFFFFFFFFF52080369848B3",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(8),        -- Port A data input
DOA(0)   => data_read_a_hi(8),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(8),        -- Port B data input
DOB(0)   => data_read_b_hi(8),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_9_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"C4C800100204810000000000000000000000000000000C001100000000000002",
INIT_01 => X"000025AAA0440812840112C000609228A10044B00000B060000008C014000C2C",
INIT_02 => X"B20427920090A4110542042800C2046008C000000002641002302002D2014003",
INIT_03 => X"5000100808000A10085044800000281004200004012E088850827814C2B20003",
INIT_04 => X"CAA0006000104084018401400000401032090000400000A0500010A102014008",
INIT_05 => X"0410008384290028881100000000022400B38084800000101280006548CCFA22",
INIT_06 => X"09640110008011A0024840A10809080801500A8000008221202008328026004B",
INIT_07 => X"C0204309148040401008200164108940808000040089083888A1005008804B09",
INIT_08 => X"97F13F36608800010140121004400200090A058284C244210000000200848002",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF98813550204088",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(9),        -- Port A data input
DOA(0)   => data_read_a_hi(9),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(9),        -- Port B data input
DOB(0)   => data_read_b_hi(9),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_10_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"C4C800100264811111111111000000000000000084884C009100000000100002",
INIT_01 => X"081025A360440812840112C000609228A10044B00000B060000808C014000C2C",
INIT_02 => X"100400120010A411054204280152000000801101010220104820000090210102",
INIT_03 => X"4000000800000810004800880020040014200000052C00885080000000100000",
INIT_04 => X"4AA000600010408441840142AAA8001400090000000020004000800102400000",
INIT_05 => X"04100082042900408B900002040402A0030004048002C0400200002D8001BC22",
INIT_06 => X"12650010140900A0040080204001080800404AA010080020200008028026014B",
INIT_07 => X"040000091000404001008040060030031001200404084A3880A8000000808310",
INIT_08 => X"3B0568176850000109C0206C040002001030180C180C00010003024210008080",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF9DC39405BE0525",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(10),        -- Port A data input
DOA(0)   => data_read_a_hi(10),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(10),        -- Port B data input
DOB(0)   => data_read_b_hi(10),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_11_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"C2880203B0600020202020200000000000400000000004000100000000000006",
INIT_01 => X"0824250C40448882840602C168004100A10180B0B4004064000000C00000000C",
INIT_02 => X"1104000010042411060204000042010000801104540220240024000080010042",
INIT_03 => X"4000088800004100204000930200018104200000000000028080000000100000",
INIT_04 => X"000355134A4410692C6086140000001000010000100000C0402000C103962001",
INIT_05 => X"001002300001000080000000C801900000000000800000000220000000000000",
INIT_06 => X"00025600802060A0000000020000080084000000005300000004080200B20000",
INIT_07 => X"0004248920084018401441960402000000000004000000000000000004800000",
INIT_08 => X"0181683650100000010000000400020020000000000000850300808C0518832D",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF9CE13045200411",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(11),        -- Port A data input
DOA(0)   => data_read_a_hi(11),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(11),        -- Port B data input
DOB(0)   => data_read_b_hi(11),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_12_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"C88A1F83F000020022002200020000000040004000000480012A000000000002",
INIT_01 => X"081025A00054C8C6940202C06F000801A50080B037810465AA0C60C00000008C",
INIT_02 => X"110400125014A4110746042880428100008411010603302100248000C0030106",
INIT_03 => X"4000018800010400044000DB822095C1142000002000102B8080000000100000",
INIT_04 => X"000F9B1B4E8208012E6294080002001000011010200000904800008103978000",
INIT_05 => X"001003BC0101000980000006E80DD00000000080800021000240000000000000",
INIT_06 => X"0002568081A070A08000000300004A04C0801100005380400000084200B60000",
INIT_07 => X"C000820D24806530004001976400000000028004000100000000000000910000",
INIT_08 => X"A4C48D264409000101C0000004C002400000000000000001806000000400832E",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF9C0025401700A6",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(12),        -- Port A data input
DOA(0)   => data_read_a_hi(12),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(12),        -- Port B data input
DOB(0)   => data_read_b_hi(12),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_13_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"C6CC00100206811133331111580000000000010084084480A320000000100002",
INIT_01 => X"083425A020C40812840552811060DB28A10144A08801F060003809C014000C2C",
INIT_02 => X"114400321014A4110742042803520800408011054102201449240000D4210342",
INIT_03 => X"4800000800016D300048A0880020041014200001832C10A85080020000104400",
INIT_04 => X"5AACE2ED56765C846DC75B56AAAA0010A40901093800EB004C298B010240A800",
INIT_05 => X"04100381042900489B100086080C122003214484800290400A60042D9091BE22",
INIT_06 => X"12410180759900A00430800142004804868051000008004010000822003600CA",
INIT_07 => X"0412B2C9048040306145C0400608308310412804044140104010002006818612",
INIT_08 => X"0FB5F7397E30000109C0246C04401A0052341A8D194C821101530AA515688080",
INIT_09 => X"00000000000000000000000000000000000005FFFFFFFFFFFFE0E7BE7F83DDBF",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(13),        -- Port A data input
DOA(0)   => data_read_a_hi(13),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(13),        -- Port B data input
DOB(0)   => data_read_b_hi(13),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_14_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"C088000001600222000000005A0000000040014000000480012A000000000002",
INIT_01 => X"08002500004408028400828000600000A10020A00000A060000000C00000000C",
INIT_02 => X"1084000000002411040204000042000000801100000220000028000081010002",
INIT_03 => X"4000000800000000004000800000000004200000000000000080000000108000",
INIT_04 => X"00000D8731063940000210140002001000010000000000004000000102000000",
INIT_05 => X"0010000000010000800000000000000000000000000000000200000000000000",
INIT_06 => X"0000000000000020000000000000080100000000000000000000080200220000",
INIT_07 => X"000000090000400C000000000400000000000004000000000000000000800000",
INIT_08 => X"BF45FF1F3CC80000110000000000020000000000000000010000000000008000",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF81E39533BF4DBE",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(14),        -- Port A data input
DOA(0)   => data_read_a_hi(14),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(14),        -- Port B data input
DOB(0)   => data_read_b_hi(14),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_15_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"C08800000060022222222222000000000040000000000400010A000000000002",
INIT_01 => X"08002500004408028400028000000000A10000A000000060000800C00000000C",
INIT_02 => X"1004000000002411040204000042000000A01102160220000020000080010002",
INIT_03 => X"4000298800000000244008800000000004200000000000000080000000100000",
INIT_04 => X"000000008000042B242188000002001000010000000000514000004502000011",
INIT_05 => X"0010000000010000800000000000000000000000000010000200000000000000",
INIT_06 => X"0000000000000020000004000040080000000000000010000004080200220000",
INIT_07 => X"0000000900004000001000008400000000000804000000000000000000800000",
INIT_08 => X"0000000000000000010000000000020000000000000000010000000000008001",
INIT_09 => X"00000000000000000000000000000000000005FFFFFFFFFFFF80000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(15),        -- Port A data input
DOA(0)   => data_read_a_hi(15),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(15),        -- Port B data input
DOB(0)   => data_read_b_hi(15),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_16_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"05104816EA00C199999999998B82D55555055577C0000675C3816AAAAAB80003",
INIT_01 => X"8014102000081213688B1862C400120ADA22C61962221218A90010E0957F0E0E",
INIT_02 => X"C200BAC50001061C8901300A2C0980A50085C801003641100400A00980206443",
INIT_03 => X"E2D5423CB284889002E20281C02900E8CC00000340A9401040162E6680824001",
INIT_04 => X"2FDAC651494D654F010FCA0208282AB240330303829FBF0A61DAFF19988017A2",
INIT_05 => X"252A5018058B9611A81110887160E2205004010210480142D30AA9290000198B",
INIT_06 => X"0050400484141401508000004500050248210008000041000000BC86424A9650",
INIT_07 => X"0208023485003A048820088005000200124342D66130400000008809D0C62220",
INIT_08 => X"1D75310E66E4584AA2AC002B005A631500000000001000005485220000000102",
INIT_09 => X"00000000000000000000000000000000000005FFFFFFFFFFFF80C3183DBECD8E",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(16),        -- Port A data input
DOA(0)   => data_read_a_hi(16),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(16),        -- Port B data input
DOB(0)   => data_read_b_hi(16),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_17_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"4F74BF57E6E587FFFFFFFFFF92D71999998E665DC000E1D9E8758CCCCCF80000",
INIT_01 => X"2ADE30F033C915094A13393EDEF4B2265284CE4B6F40B85001AE0AB1FA003513",
INIT_02 => X"664123B786736A3991E3A47C1D59727F83855D59A1AC21CA6C30AAA2F8F149E3",
INIT_03 => X"01EF407061DE98DF4182021FC45117E22A0888D2C6F8E0FE6823B275CDE77725",
INIT_04 => X"EDD90A855E9396159B5AEBFD777C19EBC03E272701DDBF0600D8FF080FE617A2",
INIT_05 => X"79639AE01E360FDFCF3BEBFFF17FEE5BBC021EE7D7EDBD79F0067A7300009CCD",
INIT_06 => X"005379675FEBE2F7E860285FE282B5A25822E00003FF001F9FEBA08437291FFC",
INIT_07 => X"D2780225C3B59F058DB28BFEEC394102168741D823F3F0040443B8C558020EE0",
INIT_08 => X"EAB0400D64A8399B47F1000937F4E00D0020100800010630ECAF77105801B3FD",
INIT_09 => X"00000000000000000000000000000000000005FFFFFFFFFFFF80203778BE0864",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(17),        -- Port A data input
DOA(0)   => data_read_a_hi(17),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(17),        -- Port B data input
DOB(0)   => data_read_b_hi(17),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_18_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"80900040060040000000000040039E1E1E0F80060E1C067E2F81CF0F0F000003",
INIT_01 => X"82500F0000100211A6110064200002886984501A10005048A99041D0557F0A28",
INIT_02 => X"C0404B0000108804C04211220424A28000C0804940226454001080009001A502",
INIT_03 => X"6078001C3080000000EB02801129001CDC40000100810011D008380302004002",
INIT_04 => X"40A662F955E7094500A5D54008A007F028431018808040026081000988000002",
INIT_05 => X"862CE019418B82203B5414007000E000436D2000000200044301F98CA1A12F12",
INIT_06 => X"36888606A41514081581900415241410202980184100E18000002CA9620A9000",
INIT_07 => X"04000A360D029582000000008204360921008066240000000104000060C2B094",
INIT_08 => X"274051317664099AEB04286408082303969048A41A4C084AD080000050000001",
INIT_09 => X"00000000000000000000000000000000000005FFFFFFFFFFFF8026A81B2A5022",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(18),        -- Port A data input
DOA(0)   => data_read_a_hi(18),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(18),        -- Port B data input
DOB(0)   => data_read_b_hi(18),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_19_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"00014020080007FFFFFFFFFF82D7E01FE008005FC000E7E1C1F5F00FF0380003",
INIT_01 => X"0000000000000004108800000000000104220004006A80000000000000000000",
INIT_02 => X"00009440000005400C0000020400000000000000002200000020000940000000",
INIT_03 => X"6040001C3080000000E20280000900000C000000000000000014440010000010",
INIT_04 => X"40018F03201F7C056400DE0C82A8007000030000808000026080000988000002",
INIT_05 => X"0090040000038200000000000000000000000000000000004300180000003022",
INIT_06 => X"00000000000000000000000000000200000000000000000000002C820C6E9000",
INIT_07 => X"0000000000002000000000000000000000000046200000000000000040C20000",
INIT_08 => X"520020232E240844100800000000230100000000000000000000000000000000",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF80A1321EAA8140",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(19),        -- Port A data input
DOA(0)   => data_read_a_hi(19),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(19),        -- Port B data input
DOB(0)   => data_read_b_hi(19),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_20_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"00000000000007FFFFFFFFFF82D7FFE0000FF85FC000E7E1C1F5FFF000380003",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000027C00000180004400007E00000000000000000000",
INIT_03 => X"E7C6867DF780000093E60380000900000C000000000000000000000000000000",
INIT_04 => X"1AA01182938901EA66400042A800BFF00003000087E2008EE386009BB8190046",
INIT_05 => X"000000000003BE0000000000000000240000430200400003CF1FF80000040140",
INIT_06 => X"00000000000000000000000000000000000000000000000000007C80000A9000",
INIT_07 => X"5200000000000000002008012D000000404007E6E000000000000008C3CE0000",
INIT_08 => X"80800812380CF801004001031202F73F00000000001120000000000000000402",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF810487600C0004",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(20),        -- Port A data input
DOA(0)   => data_read_a_hi(20),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(20),        -- Port B data input
DOB(0)   => data_read_b_hi(20),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_21_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"4410801502168D555555555520D7FFFFFF90001F8000057F8D55FFFFFFF00002",
INIT_01 => X"8880BE000439376128C090A2E09240284A30242970600098540084F0017FA04B",
INIT_02 => X"0511481A600817F8800B64437D11428202208800047EF900C80488000085480F",
INIT_03 => X"E7D80EFFF7CC20E513E60BF2044D11000C800040108C0022022B789ECAA60068",
INIT_04 => X"4AA339708A60102128A000100000BFF0000366668780201EE380801FFD140436",
INIT_05 => X"E82F02201003FE424043142491092829200010042020200BC71FF8010000B822",
INIT_06 => X"200A944880344004D8000806010285A00A09801841D2610A8A8A7E87620AD004",
INIT_07 => X"0400821589B43102800083140200010000811FE7E02200000516A82CC1EE0000",
INIT_08 => X"0F35FF3F5E36FDFE78800068F142E7BF0020100800000000F056102100480638",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF80E7BE7F83FDBF",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(21),        -- Port A data input
DOA(0)   => data_read_a_hi(21),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(21),        -- Port B data input
DOB(0)   => data_read_b_hi(21),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_22_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"6CD0E84501520D555555555524FFFFFFFF90009F8001C17F8055FFFFFFF00000",
INIT_01 => X"0A94BEAFE77D3C314A43D337A45241685290F4CFD22090F85C488C03D57FAC62",
INIT_02 => X"F6157F9A78589FFDD14B756901537001E028C4415900AB14E83DA22A50A5694B",
INIT_03 => X"0827A802001090086000807A1124150890A222023DA002AA52AE78DFEAF6314B",
INIT_04 => X"4AAFBB390A30488569A60142AAAA000304287676087620400446A00045541AC0",
INIT_05 => X"AB7FFAA014A840490B55B62E915D2A21A204059434223328000007AC10111C26",
INIT_06 => X"004B1C0A95B9400000D0060740E01FB25402400206DA180A8A9A020766044540",
INIT_07 => X"0561124C8480FA0545630B5480B002881117300105A340926202228100302A02",
INIT_08 => X"BFC5793F7CEA05FF48C00408F1C800800084422111088C6164DF1284170066A9",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF81E7BD7BBEDDAE",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(22),        -- Port A data input
DOA(0)   => data_read_a_hi(22),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(22),        -- Port B data input
DOB(0)   => data_read_b_hi(22),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_23_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"8A99D0720284A800000000006A000000005FFF400C1804002D00000000000002",
INIT_01 => X"A00080000420E3E7BC8241B640909201EF20906F206006E5F4E2B4F0200040CD",
INIT_02 => X"A39050087D451C8190084003FC04B16802C11910167EDC8180382AA20006800C",
INIT_03 => X"E7C02FFFF780000017EE0BA0044D00122CC888D0700CC010020D0094F2A38B73",
INIT_04 => X"000CCAAD86201C00280300100000BFF02003404087818A5FE3980A5FF8000017",
INIT_05 => X"EB7FFD010003FF226006CA081110001A0921000141088043C71FFF8180809200",
INIT_06 => X"121000064104000084008000160696210A020000002000800004FEA2020AD004",
INIT_07 => X"100002134014B008841000000801100108000FF7E00000000504880EE5FE8010",
INIT_08 => X"000000000006F800200020040002E7FF1200000008000002F834000000000000",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF80000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(23),        -- Port A data input
DOA(0)   => data_read_a_hi(23),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(23),        -- Port B data input
DOB(0)   => data_read_b_hi(23),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_24_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000D555555555524FFFFFFFF90009F8001C57F8155FFFFFFF00002",
INIT_01 => X"0000800004202020000000000000000000000000000000805400840000000040",
INIT_02 => X"0010800820001080000840037C00000000000000007E88008380000000040008",
INIT_03 => X"E7C0067FF780000013E603A0000D00000C800000100000000210008001000040",
INIT_04 => X"000065E581003800000200100000BFF0000340408780000EE380001BF8000006",
INIT_05 => X"040000000003FE0000000000000000000000000000000003C71FFF8000003000",
INIT_06 => X"00000000000000000000000000000000000000000000000000007E80098AD00A",
INIT_07 => X"00000000000004800000000000000000000007E7E000000001048808C1EE0000",
INIT_08 => X"8EB2CEAF580EF800100000000002E7BF00000000000000000000000000000000",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF806D2D66331814",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(24),        -- Port A data input
DOA(0)   => data_read_a_hi(24),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(24),        -- Port B data input
DOB(0)   => data_read_b_hi(24),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_25_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000D555555555524FFFFFFFF90009F8001C57F8155FFFFFFF00002",
INIT_01 => X"0000800004202020000000000000000000000000000000805400840000000040",
INIT_02 => X"0010000820001080000840037C00028600040000007E88008000000000040008",
INIT_03 => X"E7D8067FF7DC38FD53E623A0000D00000C800000100000000200008000000040",
INIT_04 => X"800000600C600421202100000000BFF0000340408780040EE380041BF8080426",
INIT_05 => X"000000000003FE0000000000000000645202140402000013D71FFF890105B400",
INIT_06 => X"200080600000065F7801285001000000A02980184100610000007E80000AD000",
INIT_07 => X"0400B0C0092001022015C00802002102008007E7E000000001148868C9EE0000",
INIT_08 => X"14B3C80EA076F800880701680006E7BF0230180C100C0000002200A541491010",
INIT_09 => X"00000000000000000000000000000000000003FFFFFFFFFFFF80883A7B42C803",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(25),        -- Port A data input
DOA(0)   => data_read_a_hi(25),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(25),        -- Port B data input
DOB(0)   => data_read_b_hi(25),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_26_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"85F820440E61E5DDDDDDDDDD81D7FFFFFF8FFE3FDEBCEF7FDFD5FFFFFFF80007",
INIT_01 => X"AA5E3FF033CC1A1BA4993AAC8064328EE9265EAA400ABA7000401AC1DE00573E",
INIT_02 => X"F645FFF78F73EF7DDDE3B57E7C6F72BF89C15D49E0FE675E24302AA9F8D1E5E3",
INIT_03 => X"E7FFD67DF7DE1ADFDBEF578C5479263E7E600053CEFDE25C78BFFE7FDFF77F3F",
INIT_04 => X"FFF000600019C294D19C21E3FFFDFFFBFAFF272787FF302EE3D6F03BBE6057EE",
INIT_05 => X"FFFFFCC1DABFBFFEFF7FFFFB1136267FFFFFFFE7D7EFDE7FFF1FFBFFEBEFFFFF",
INIT_06 => X"7FD9A0671ECB87FF7FEBFADDFDAEBDB23939E23AD10C6B9D1D69FCBF7F6F9FBE",
INIT_07 => X"17794B3BCFB7DA839D8AAA600FBDFF5BFFC567FEEFF3F234094F98D9DBCEFEFD",
INIT_08 => X"D082EF0B3EACFFFFFFFF7BFFFFFFF73F9DBA9D6EAEBF7E7B7C8F77525A85B4C0",
INIT_09 => X"00000000000000000000000000000000000003FFFFFFFFFFFF800B354D1138DC",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(26),        -- Port A data input
DOA(0)   => data_read_a_hi(26),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(26),        -- Port B data input
DOB(0)   => data_read_b_hi(26),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_27_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"11200008002844CCCCCCCCCC80D7FFFFFF8FFE1F5AB4AB7F5ED5FFFFFFEA8015",
INIT_01 => X"080A0E5012800008002029000029049200080A4000142822000002090A800110",
INIT_02 => X"4441D8370DC3416110A004547C8854AB88011100A0FC000A040022202A1000A0",
INIT_03 => X"97EF9671EFDC1ADDDB97570404512A062A000057CA7F0844783D024B19456E38",
INIT_04 => X"7FF000600019C294D19C21E3FFFDFFEE9A8E252547F7102E93D6603A3C2056EE",
INIT_05 => X"AFCF7842C23E3FD65FFECAC9041202FB2ADCE767554BCC6FEC9FFBBF6B6BFDFF",
INIT_06 => X"6DFCA0760E43875F7BAB7AF4EDAF80B83959EAB8D10463B03008F099E10914AB",
INIT_07 => X"1654452153BC0AC3998AA2200B2BAE5AF54467F8EF78FA3C88E88891D30E774D",
INIT_08 => X"4A825C88A220FFFFCC7F5AFBF93BF43F2DAA956AA6BB7AD42E0FD35A18942440",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF80F91049E10840",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(27),        -- Port A data input
DOA(0)   => data_read_a_hi(27),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(27),        -- Port B data input
DOB(0)   => data_read_b_hi(27),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_28_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"4128400000606088888888888000000000000000420526004380000000080003",
INIT_01 => X"220A20501184080808802A90006000C202200AA40000A820004A02822A004110",
INIT_02 => X"B24427A5000A440440A21114001A00002288C440A980220A0CA1088828B120A2",
INIT_03 => X"0000000000008000800100041110020C8222220186D182D428827A14E2B25403",
INIT_04 => X"B550000000098210901820A15554000988240303000014000000440000280000",
INIT_05 => X"40900040569400B4342934E101420804D04A727222611E1438000012202401D9",
INIT_06 => X"048028000A46800001601000A00008000002200206A4081A9A92000A040101A0",
INIT_07 => X"03310028020040000CA00828019805006CC0500802D2B086264222463A001C44",
INIT_08 => X"0501710016D0000034380903083410000400400012112631000041104A014050",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF809A223208608B",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(28),        -- Port A data input
DOA(0)   => data_read_a_hi(28),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(28),        -- Port B data input
DOB(0)   => data_read_b_hi(28),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_29_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A5F0A0540E75C5DDDDDDDDDD81000000000FFE20C60C677EC3D5FFFFFFD80003",
INIT_01 => X"805E1FFFF1C81619E659392E8076B2AE79965E4B402AB858000A0A71FF7FBF3B",
INIT_02 => X"E240FFF78F72EB588DE1A03E016D627D81408809E0FE455E66100001F850C5E1",
INIT_03 => X"E037C67C104E00C793E9038C403806345E4000438F5D604C281FFE7FDFA35F3F",
INIT_04 => X"FFF0000000098210901820A15554BFFBE8572323807E340EE046F41B866813C6",
INIT_05 => X"B8AF84C14A1781FEBF7B77D31026246DDD6B6EE3D3C59C1FFF0003F2A0A4BFFB",
INIT_06 => X"16C9282F1ACE82F32560B25DB402B59200202000022C001515697C2D7A6F8FFE",
INIT_07 => X"02380A338E97988008800068051D550176C167FE03D1B0140545104DFBC09EF4",
INIT_08 => X"2E77BF3F7E2405FFF7FA292FFFF6F700941008040A15263A748175100800B0D0",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF83D7BC7787BF7E",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(29),        -- Port A data input
DOA(0)   => data_read_a_hi(29),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(29),        -- Port B data input
DOB(0)   => data_read_b_hi(29),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_30_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000222222222225A00000000000140000000800020000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"DF83FF2F7CF80000000000000000000000000000000000000000000000000000",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF80FF3F7F3BF8DF",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(30),        -- Port A data input
DOA(0)   => data_read_a_hi(30),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(30),        -- Port B data input
DOB(0)   => data_read_b_hi(30),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_31_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"60008010001404444444444400D7FFFFFF8FFE1F0810817F0C55FFFFFFE00000",
INIT_01 => X"08800E0FC20105004A40000200128020129000010020000800000030017FA801",
INIT_02 => X"4401D8120D410161100004407D1050EB80011110017C00804A00222200200800",
INIT_03 => X"87EF8671E7DC18DD5386030004410002280888D2492C0080503D004B19452A38",
INIT_04 => X"4AA000600010408441840142AAA8BFE2000A242407F7000E83D6201A3C0016E6",
INIT_05 => X"AF4F7800042A3F424B56CA080010027B2A040505450A806BC41FFBAD0101BC26",
INIT_06 => X"2058806C0401065F78812A5045A680B03809C018418061800000F0816108144A",
INIT_07 => X"1440000141B40A83810282000A21220A110427E0E520401000008881C10E2200",
INIT_08 => X"000000000000FDFFC8470068F10AE43F00A05028100808402C0F120010000400",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF80000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(31),        -- Port A data input
DOA(0)   => data_read_a_hi(31),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(31),        -- Port B data input
DOB(0)   => data_read_b_hi(31),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_0_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"DA9918630DD2200000000000012800000040002000A106001180000000008007",
INIT_01 => X"80202100005CD2C7B4E6C1E566434955ED29B05AB311C477A91660C2B4D5208F",
INIT_02 => X"11840040D2AC24048604810082640D046B24CC461E01332121AD800087828206",
INIT_03 => X"080029800001E5202400B85242009129400A2A042000F22200808420C4108104",
INIT_04 => X"000FFF9D8F603C21282300100003000404F0100838008ED10C280E44011DA811",
INIT_05 => X"5000032408000000808000349D2934800010180000802B000060040012120000",
INIT_06 => X"40261C93C1345120821204AE0A41780DC6D01980827218422A0C004092B00A14",
INIT_07 => X"400AF9C0A003557C605D491DA48448900A020810000202AAEA922236141141A2",
INIT_08 => X"9030DA025E0900002300040002000840C204C2C131209008137028AD0779C23B",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF80C11F1127D082",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(0),        -- Port A data input
DOA(0)   => data_read_a_lo_256(0),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(0),        -- Port B data input
DOB(0)   => data_read_b_lo_256(0),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_1_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"C08451022808200000000000002000000000000010000C001108000000028002",
INIT_01 => X"22402100005000008490005046680400213C00142300E04080F4514BA066C00C",
INIT_02 => X"00000000000020044400010000C28410230CC4480000024000A1800182C12400",
INIT_03 => X"00001000000000000810440001002000802880040000A2020000800004000000",
INIT_04 => X"00006D858F602400280300100001400452000008000004A0000004A002090008",
INIT_05 => X"501000209000000080000020010008000090900090000B000000000048484000",
INIT_06 => X"09000900010410A082084002000002000012000214208008A890001284200000",
INIT_07 => X"4005010C10002000042028092400884080000000080A08222A22000200004009",
INIT_08 => X"947022015EA802000108121004000000090A458294C24001820004404205F012",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF81809307840190",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(1),        -- Port A data input
DOA(0)   => data_read_a_lo_256(1),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(1),        -- Port B data input
DOB(0)   => data_read_b_lo_256(1),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_2_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"C4804010026CA010101010110092D555550554161001447431116AAAAA820012",
INIT_01 => X"0A141D0A80440812841911980061967CA10E44C4000CB262012008C8B4780C08",
INIT_02 => X"100400000DD9AA5D050335002951264102C1C141491444444A90028282604143",
INIT_03 => X"82921220A28088500A92560801202412F06202040082080840808000E4110B00",
INIT_04 => X"42200020000040044004010208896AA03288101802A0242A0104843012480048",
INIT_05 => X"861A5082908814018000830A041400220C909115E12C4A02A00AA8054ACAD020",
INIT_06 => X"59510860140403E86A0AC8101AA88502590A401A542022AAAA0210378C24000B",
INIT_07 => X"010500130C048045913A20488481D851900022D048080090A2A0220280044209",
INIT_08 => X"B5013F1C742852CE43805274B40340150B9A8D46B4AE500242A910405294C091",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFFC8A0193716CC3A",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(2),        -- Port A data input
DOA(0)   => data_read_a_lo_256(2),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(2),        -- Port B data input
DOB(0)   => data_read_b_lo_256(2),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_3_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"C0C1002008E008110011001024C366666619989C00A105460141B33333020006",
INIT_01 => X"0004B50C84642830841112880080922C210C4480004812E055808C413181DC6C",
INIT_02 => X"1014001A2DD1BAA94D09640318C2C44822849440480EA80482208882C2050048",
INIT_03 => X"3183106A69989A5449B854A8102C241814A02200110008980280808005100940",
INIT_04 => X"02800040000040804084000020A9599012A1404041B024261084A4284A48426A",
INIT_05 => X"084C60828481CC880890A0020404028281A09081C02081418386630DCACBE422",
INIT_06 => X"5B410840148C02BA740ACA8100A00A283828400A542820800A90A6342866C040",
INIT_07 => X"0005020D0480604185022048040010518011018520110A2A2C208A1040220019",
INIT_08 => X"B000220C748E346521C072F0A541C38C199A8D46B4AE50018A0C004810148090",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF8D4015050C05A8",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(3),        -- Port A data input
DOA(0)   => data_read_a_lo_256(3),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(3),        -- Port B data input
DOB(0)   => data_read_b_lo_256(3),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_4_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"C0CB20AC108100111100001100FC78787806181894884518995E3C3C3C128002",
INIT_01 => X"081425AA60440802840100008184B200A108402040C21260028000C0C400122C",
INIT_02 => X"920406000DC124110442042878C2002022409101485E64140010200892014143",
INIT_03 => X"87840669E7D0189253BE47000009280008000000012E28805080601083130802",
INIT_04 => X"C800000000004084410000002A09B8651202020207C8240E8380941A3A480026",
INIT_05 => X"14308401842A3C60A30184200440000613808401C0020003971E190CC8C94422",
INIT_06 => X"1B750810100D02FD0008C2A0402D080011410A909028432604AB74B20028904A",
INIT_07 => X"0420400900004001142AA0480610B04390803784EC884A00090F984AC90E0119",
INIT_08 => X"044015114600F6E44900731CA503C63C19AA150A8C824001020B024202848090",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFFB5208A0F988902",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(4),        -- Port A data input
DOA(0)   => data_read_a_lo_256(4),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(4),        -- Port B data input
DOB(0)   => data_read_b_lo_256(4),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_5_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"CAC8380F010300111111110000D7807F8048181E94A84D60A555C03FC0120002",
INIT_01 => X"082025234054C8C69416C281E46C6D05A50DA0A0F217E665A82468C854801EAC",
INIT_02 => X"918425025D5524110746040A8752890040A491061F213021492C800087230206",
INIT_03 => X"6860699410016D322440A8DA0620950314200004212C10A25082501400108001",
INIT_04 => X"000FFFFD8F703C2168230012AAA207E424011018B8028E516C681E45831CB911",
INIT_05 => X"041007240429826183011006880D1004421104108202B1405161FD051010B800",
INIT_06 => X"02429C80C53D41A8DE1006824B604A05D690D122917A18678266086280B6004A",
INIT_07 => X"0406B3CD3480653D617FE11C8680A882100228620C804220481000302CD14002",
INIT_08 => X"0FB5FF3F7A550B6269C0046C8500294342B41A0D190C8001837B0AED157C8239",
INIT_09 => X"00000000000000000000000000000000000005FFFFFFFFFFFFC1E3BE7EA3DDBF",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(5),        -- Port A data input
DOA(0)   => data_read_a_lo_256(5),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(5),        -- Port B data input
DOB(0)   => data_read_b_lo_256(5),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_6_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"C0CC0708E06000111111111100D7FF80000FE01E10200D600155FFC000000002",
INIT_01 => X"0800250C41440812842112C018619238A10844B00C14B062001008C094001C2C",
INIT_02 => X"1204201000902411040204000042000008809100000220000020000080010002",
INIT_03 => X"400010080000000208585481800020D004200004000208080082000000121000",
INIT_04 => X"000000005086000044000A02AAA8401432890000000024204000842102480108",
INIT_05 => X"0010008180010020889110006000C2A441A090040200000012000068CA4B4400",
INIT_06 => X"5901080010040128000A428008200800101000008020002D2B89083200220000",
INIT_07 => X"0020410910004041000220480490005080810006E888081880A80040C9000219",
INIT_08 => X"B541FF1F3E2802610100721081840200198A8542A4A250010008000000048090",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF9CE19F3B9FDCBA",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(6),        -- Port A data input
DOA(0)   => data_read_a_lo_256(6),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(6),        -- Port B data input
DOB(0)   => data_read_b_lo_256(6),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_7_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"C48C031862648011111111110000000000000000840844008100000000100006",
INIT_01 => X"0804258020440802842002C012090410A10000B009000060000000C00000000C",
INIT_02 => X"100400100090A4110402042001D2040000809100410220144820000090210042",
INIT_03 => X"40001008001210084840108880600C4034200000000000098080000000100000",
INIT_04 => X"00000000208000484200860AAAA9401100810000000065204001852102CA0428",
INIT_05 => X"00100099010100408384820A241440920A310501C10AC0400200000802830600",
INIT_06 => X"40014A20340D27F32203201048088808011040028029002A8802082200220000",
INIT_07 => X"15010709148C40401108A0CA0E83B81A1001A00404204000000800000080C000",
INIT_08 => X"00000000000000990980406C748102002030D86C382C10850003920010048194",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF94000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(7),        -- Port A data input
DOA(0)   => data_read_a_lo_256(7),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(7),        -- Port B data input
DOB(0)   => data_read_b_lo_256(7),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_8_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"D08800000008001111111111000000000000000084884C009100000000100002",
INIT_01 => X"081025A001440802842002C000090410A10800B000140062000001C80080000C",
INIT_02 => X"100400120000A4110542042801520000008011010102200048200000C0210102",
INIT_03 => X"50000008080202000050448984202CD214200004000208088080000000301000",
INIT_04 => X"800000021000010244405806AAA8001032010000400000005000000102004000",
INIT_05 => X"0010009180010048838000026404C08002B38480800290500280000848CD4600",
INIT_06 => X"09240010048900A0024840A14009080001504880800800040000083200260000",
INIT_07 => X"04000309148040401100A0000600A9429800300404094A0888A8001000804909",
INIT_08 => X"2A303F1F5850050749C052F804C40200092A150A948A44210003020010048000",
INIT_09 => X"00000000000000000000000000000000000005FFFFFFFFFFFFF52080369848B3",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(8),        -- Port A data input
DOA(0)   => data_read_a_lo_256(8),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(8),        -- Port B data input
DOB(0)   => data_read_b_lo_256(8),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_9_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"C4C800100204810000000000000000000000000000000C001100000000000002",
INIT_01 => X"000025AAA0440812840112C000609228A10044B00000B060000008C014000C2C",
INIT_02 => X"B20427920090A4110542042800C2046008C000000002641002302002D2014003",
INIT_03 => X"5000100808000A10085044800000281004200004012E088850827814C2B20003",
INIT_04 => X"CAA0006000104084018401400000401032090000400000A0500010A102014008",
INIT_05 => X"0410008384290028881100000000022400B38084800000101280006548CCFA22",
INIT_06 => X"09640110008011A0024840A10809080801500A8000008221202008328026004B",
INIT_07 => X"C0204309148040401008200164108940808000040089083888A1005008804B09",
INIT_08 => X"97F13F36608800010140121004400200090A058284C244210000000200848002",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF98813550204088",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(9),        -- Port A data input
DOA(0)   => data_read_a_lo_256(9),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(9),        -- Port B data input
DOB(0)   => data_read_b_lo_256(9),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_10_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"C4C800100264811111111111000000000000000084884C009100000000100002",
INIT_01 => X"081025A360440812840112C000609228A10044B00000B060000808C014000C2C",
INIT_02 => X"100400120010A411054204280152000000801101010220104820000090210102",
INIT_03 => X"4000000800000810004800880020040014200000052C00885080000000100000",
INIT_04 => X"4AA000600010408441840142AAA8001400090000000020004000800102400000",
INIT_05 => X"04100082042900408B900002040402A0030004048002C0400200002D8001BC22",
INIT_06 => X"12650010140900A0040080204001080800404AA010080020200008028026014B",
INIT_07 => X"040000091000404001008040060030031001200404084A3880A8000000808310",
INIT_08 => X"3B0568176850000109C0206C040002001030180C180C00010003024210008080",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF9DC39405BE0525",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(10),        -- Port A data input
DOA(0)   => data_read_a_lo_256(10),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(10),        -- Port B data input
DOB(0)   => data_read_b_lo_256(10),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_11_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"C2880203B0600020202020200000000000400000000004000100000000000006",
INIT_01 => X"0824250C40448882840602C168004100A10180B0B4004064000000C00000000C",
INIT_02 => X"1104000010042411060204000042010000801104540220240024000080010042",
INIT_03 => X"4000088800004100204000930200018104200000000000028080000000100000",
INIT_04 => X"000355134A4410692C6086140000001000010000100000C0402000C103962001",
INIT_05 => X"001002300001000080000000C801900000000000800000000220000000000000",
INIT_06 => X"00025600802060A0000000020000080084000000005300000004080200B20000",
INIT_07 => X"0004248920084018401441960402000000000004000000000000000004800000",
INIT_08 => X"0181683650100000010000000400020020000000000000850300808C0518832D",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF9CE13045200411",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(11),        -- Port A data input
DOA(0)   => data_read_a_lo_256(11),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(11),        -- Port B data input
DOB(0)   => data_read_b_lo_256(11),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_12_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"C88A1F83F000020022002200020000000040004000000480012A000000000002",
INIT_01 => X"081025A00054C8C6940202C06F000801A50080B037810465AA0C60C00000008C",
INIT_02 => X"110400125014A4110746042880428100008411010603302100248000C0030106",
INIT_03 => X"4000018800010400044000DB822095C1142000002000102B8080000000100000",
INIT_04 => X"000F9B1B4E8208012E6294080002001000011010200000904800008103978000",
INIT_05 => X"001003BC0101000980000006E80DD00000000080800021000240000000000000",
INIT_06 => X"0002568081A070A08000000300004A04C0801100005380400000084200B60000",
INIT_07 => X"C000820D24806530004001976400000000028004000100000000000000910000",
INIT_08 => X"A4C48D264409000101C0000004C002400000000000000001806000000400832E",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF9C0025401700A6",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(12),        -- Port A data input
DOA(0)   => data_read_a_lo_256(12),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(12),        -- Port B data input
DOB(0)   => data_read_b_lo_256(12),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_13_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"C6CC00100206811133331111580000000000010084084480A320000000100002",
INIT_01 => X"083425A020C40812840552811060DB28A10144A08801F060003809C014000C2C",
INIT_02 => X"114400321014A4110742042803520800408011054102201449240000D4210342",
INIT_03 => X"4800000800016D300048A0880020041014200001832C10A85080020000104400",
INIT_04 => X"5AACE2ED56765C846DC75B56AAAA0010A40901093800EB004C298B010240A800",
INIT_05 => X"04100381042900489B100086080C122003214484800290400A60042D9091BE22",
INIT_06 => X"12410180759900A00430800142004804868051000008004010000822003600CA",
INIT_07 => X"0412B2C9048040306145C0400608308310412804044140104010002006818612",
INIT_08 => X"0FB5F7397E30000109C0246C04401A0052341A8D194C821101530AA515688080",
INIT_09 => X"00000000000000000000000000000000000005FFFFFFFFFFFFE0E7BE7F83DDBF",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(13),        -- Port A data input
DOA(0)   => data_read_a_lo_256(13),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(13),        -- Port B data input
DOB(0)   => data_read_b_lo_256(13),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_14_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"C088000001600222000000005A0000000040014000000480012A000000000002",
INIT_01 => X"08002500004408028400828000600000A10020A00000A060000000C00000000C",
INIT_02 => X"1084000000002411040204000042000000801100000220000028000081010002",
INIT_03 => X"4000000800000000004000800000000004200000000000000080000000108000",
INIT_04 => X"00000D8731063940000210140002001000010000000000004000000102000000",
INIT_05 => X"0010000000010000800000000000000000000000000000000200000000000000",
INIT_06 => X"0000000000000020000000000000080100000000000000000000080200220000",
INIT_07 => X"000000090000400C000000000400000000000004000000000000000000800000",
INIT_08 => X"BF45FF1F3CC80000110000000000020000000000000000010000000000008000",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF81E39533BF4DBE",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(14),        -- Port A data input
DOA(0)   => data_read_a_lo_256(14),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(14),        -- Port B data input
DOB(0)   => data_read_b_lo_256(14),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_15_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"C08800000060022222222222000000000040000000000400010A000000000002",
INIT_01 => X"08002500004408028400028000000000A10000A000000060000800C00000000C",
INIT_02 => X"1004000000002411040204000042000000A01102160220000020000080010002",
INIT_03 => X"4000298800000000244008800000000004200000000000000080000000100000",
INIT_04 => X"000000008000042B242188000002001000010000000000514000004502000011",
INIT_05 => X"0010000000010000800000000000000000000000000010000200000000000000",
INIT_06 => X"0000000000000020000004000040080000000000000010000004080200220000",
INIT_07 => X"0000000900004000001000008400000000000804000000000000000000800000",
INIT_08 => X"0000000000000000010000000000020000000000000000010000000000008001",
INIT_09 => X"00000000000000000000000000000000000005FFFFFFFFFFFF80000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(15),        -- Port A data input
DOA(0)   => data_read_a_lo_256(15),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(15),        -- Port B data input
DOB(0)   => data_read_b_lo_256(15),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_16_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"05104816EA00C199999999998B82D55555055577C0000675C3816AAAAAB80003",
INIT_01 => X"8014102000081213688B1862C400120ADA22C61962221218A90010E0957F0E0E",
INIT_02 => X"C200BAC50001061C8901300A2C0980A50085C801003641100400A00980206443",
INIT_03 => X"E2D5423CB284889002E20281C02900E8CC00000340A9401040162E6680824001",
INIT_04 => X"2FDAC651494D654F010FCA0208282AB240330303829FBF0A61DAFF19988017A2",
INIT_05 => X"252A5018058B9611A81110887160E2205004010210480142D30AA9290000198B",
INIT_06 => X"0050400484141401508000004500050248210008000041000000BC86424A9650",
INIT_07 => X"0208023485003A048820088005000200124342D66130400000008809D0C62220",
INIT_08 => X"1D75310E66E4584AA2AC002B005A631500000000001000005485220000000102",
INIT_09 => X"00000000000000000000000000000000000005FFFFFFFFFFFF80C3183DBECD8E",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(16),        -- Port A data input
DOA(0)   => data_read_a_lo_256(16),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(16),        -- Port B data input
DOB(0)   => data_read_b_lo_256(16),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_17_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"4F74BF57E6E587FFFFFFFFFF92D71999998E665DC000E1D9E8758CCCCCF80000",
INIT_01 => X"2ADE30F033C915094A13393EDEF4B2265284CE4B6F40B85001AE0AB1FA003513",
INIT_02 => X"664123B786736A3991E3A47C1D59727F83855D59A1AC21CA6C30AAA2F8F149E3",
INIT_03 => X"01EF407061DE98DF4182021FC45117E22A0888D2C6F8E0FE6823B275CDE77725",
INIT_04 => X"EDD90A855E9396159B5AEBFD777C19EBC03E272701DDBF0600D8FF080FE617A2",
INIT_05 => X"79639AE01E360FDFCF3BEBFFF17FEE5BBC021EE7D7EDBD79F0067A7300009CCD",
INIT_06 => X"005379675FEBE2F7E860285FE282B5A25822E00003FF001F9FEBA08437291FFC",
INIT_07 => X"D2780225C3B59F058DB28BFEEC394102168741D823F3F0040443B8C558020EE0",
INIT_08 => X"EAB0400D64A8399B47F1000937F4E00D0020100800010630ECAF77105801B3FD",
INIT_09 => X"00000000000000000000000000000000000005FFFFFFFFFFFF80203778BE0864",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(17),        -- Port A data input
DOA(0)   => data_read_a_lo_256(17),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(17),        -- Port B data input
DOB(0)   => data_read_b_lo_256(17),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_18_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"80900040060040000000000040039E1E1E0F80060E1C067E2F81CF0F0F000003",
INIT_01 => X"82500F0000100211A6110064200002886984501A10005048A99041D0557F0A28",
INIT_02 => X"C0404B0000108804C04211220424A28000C0804940226454001080009001A502",
INIT_03 => X"6078001C3080000000EB02801129001CDC40000100810011D008380302004002",
INIT_04 => X"40A662F955E7094500A5D54008A007F028431018808040026081000988000002",
INIT_05 => X"862CE019418B82203B5414007000E000436D2000000200044301F98CA1A12F12",
INIT_06 => X"36888606A41514081581900415241410202980184100E18000002CA9620A9000",
INIT_07 => X"04000A360D029582000000008204360921008066240000000104000060C2B094",
INIT_08 => X"274051317664099AEB04286408082303969048A41A4C084AD080000050000001",
INIT_09 => X"00000000000000000000000000000000000005FFFFFFFFFFFF8026A81B2A5022",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(18),        -- Port A data input
DOA(0)   => data_read_a_lo_256(18),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(18),        -- Port B data input
DOB(0)   => data_read_b_lo_256(18),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_19_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"00014020080007FFFFFFFFFF82D7E01FE008005FC000E7E1C1F5F00FF0380003",
INIT_01 => X"0000000000000004108800000000000104220004006A80000000000000000000",
INIT_02 => X"00009440000005400C0000020400000000000000002200000020000940000000",
INIT_03 => X"6040001C3080000000E20280000900000C000000000000000014440010000010",
INIT_04 => X"40018F03201F7C056400DE0C82A8007000030000808000026080000988000002",
INIT_05 => X"0090040000038200000000000000000000000000000000004300180000003022",
INIT_06 => X"00000000000000000000000000000200000000000000000000002C820C6E9000",
INIT_07 => X"0000000000002000000000000000000000000046200000000000000040C20000",
INIT_08 => X"520020232E240844100800000000230100000000000000000000000000000000",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF80A1321EAA8140",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(19),        -- Port A data input
DOA(0)   => data_read_a_lo_256(19),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(19),        -- Port B data input
DOB(0)   => data_read_b_lo_256(19),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_20_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"00000000000007FFFFFFFFFF82D7FFE0000FF85FC000E7E1C1F5FFF000380003",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000027C00000180004400007E00000000000000000000",
INIT_03 => X"E7C6867DF780000093E60380000900000C000000000000000000000000000000",
INIT_04 => X"1AA01182938901EA66400042A800BFF00003000087E2008EE386009BB8190046",
INIT_05 => X"000000000003BE0000000000000000240000430200400003CF1FF80000040140",
INIT_06 => X"00000000000000000000000000000000000000000000000000007C80000A9000",
INIT_07 => X"5200000000000000002008012D000000404007E6E000000000000008C3CE0000",
INIT_08 => X"80800812380CF801004001031202F73F00000000001120000000000000000402",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF810487600C0004",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(20),        -- Port A data input
DOA(0)   => data_read_a_lo_256(20),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(20),        -- Port B data input
DOB(0)   => data_read_b_lo_256(20),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_21_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"4410801502168D555555555520D7FFFFFF90001F8000057F8D55FFFFFFF00002",
INIT_01 => X"8880BE000439376128C090A2E09240284A30242970600098540084F0017FA04B",
INIT_02 => X"0511481A600817F8800B64437D11428202208800047EF900C80488000085480F",
INIT_03 => X"E7D80EFFF7CC20E513E60BF2044D11000C800040108C0022022B789ECAA60068",
INIT_04 => X"4AA339708A60102128A000100000BFF0000366668780201EE380801FFD140436",
INIT_05 => X"E82F02201003FE424043142491092829200010042020200BC71FF8010000B822",
INIT_06 => X"200A944880344004D8000806010285A00A09801841D2610A8A8A7E87620AD004",
INIT_07 => X"0400821589B43102800083140200010000811FE7E02200000516A82CC1EE0000",
INIT_08 => X"0F35FF3F5E36FDFE78800068F142E7BF0020100800000000F056102100480638",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF80E7BE7F83FDBF",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(21),        -- Port A data input
DOA(0)   => data_read_a_lo_256(21),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(21),        -- Port B data input
DOB(0)   => data_read_b_lo_256(21),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_22_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"6CD0E84501520D555555555524FFFFFFFF90009F8001C17F8055FFFFFFF00000",
INIT_01 => X"0A94BEAFE77D3C314A43D337A45241685290F4CFD22090F85C488C03D57FAC62",
INIT_02 => X"F6157F9A78589FFDD14B756901537001E028C4415900AB14E83DA22A50A5694B",
INIT_03 => X"0827A802001090086000807A1124150890A222023DA002AA52AE78DFEAF6314B",
INIT_04 => X"4AAFBB390A30488569A60142AAAA000304287676087620400446A00045541AC0",
INIT_05 => X"AB7FFAA014A840490B55B62E915D2A21A204059434223328000007AC10111C26",
INIT_06 => X"004B1C0A95B9400000D0060740E01FB25402400206DA180A8A9A020766044540",
INIT_07 => X"0561124C8480FA0545630B5480B002881117300105A340926202228100302A02",
INIT_08 => X"BFC5793F7CEA05FF48C00408F1C800800084422111088C6164DF1284170066A9",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF81E7BD7BBEDDAE",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(22),        -- Port A data input
DOA(0)   => data_read_a_lo_256(22),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(22),        -- Port B data input
DOB(0)   => data_read_b_lo_256(22),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_23_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"8A99D0720284A800000000006A000000005FFF400C1804002D00000000000002",
INIT_01 => X"A00080000420E3E7BC8241B640909201EF20906F206006E5F4E2B4F0200040CD",
INIT_02 => X"A39050087D451C8190084003FC04B16802C11910167EDC8180382AA20006800C",
INIT_03 => X"E7C02FFFF780000017EE0BA0044D00122CC888D0700CC010020D0094F2A38B73",
INIT_04 => X"000CCAAD86201C00280300100000BFF02003404087818A5FE3980A5FF8000017",
INIT_05 => X"EB7FFD010003FF226006CA081110001A0921000141088043C71FFF8180809200",
INIT_06 => X"121000064104000084008000160696210A020000002000800004FEA2020AD004",
INIT_07 => X"100002134014B008841000000801100108000FF7E00000000504880EE5FE8010",
INIT_08 => X"000000000006F800200020040002E7FF1200000008000002F834000000000000",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF80000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(23),        -- Port A data input
DOA(0)   => data_read_a_lo_256(23),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(23),        -- Port B data input
DOB(0)   => data_read_b_lo_256(23),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_24_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000D555555555524FFFFFFFF90009F8001C57F8155FFFFFFF00002",
INIT_01 => X"0000800004202020000000000000000000000000000000805400840000000040",
INIT_02 => X"0010800820001080000840037C00000000000000007E88008380000000040008",
INIT_03 => X"E7C0067FF780000013E603A0000D00000C800000100000000210008001000040",
INIT_04 => X"000065E581003800000200100000BFF0000340408780000EE380001BF8000006",
INIT_05 => X"040000000003FE0000000000000000000000000000000003C71FFF8000003000",
INIT_06 => X"00000000000000000000000000000000000000000000000000007E80098AD00A",
INIT_07 => X"00000000000004800000000000000000000007E7E000000001048808C1EE0000",
INIT_08 => X"8EB2CEAF580EF800100000000002E7BF00000000000000000000000000000000",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF806D2D66331814",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(24),        -- Port A data input
DOA(0)   => data_read_a_lo_256(24),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(24),        -- Port B data input
DOB(0)   => data_read_b_lo_256(24),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_25_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000D555555555524FFFFFFFF90009F8001C57F8155FFFFFFF00002",
INIT_01 => X"0000800004202020000000000000000000000000000000805400840000000040",
INIT_02 => X"0010000820001080000840037C00028600040000007E88008000000000040008",
INIT_03 => X"E7D8067FF7DC38FD53E623A0000D00000C800000100000000200008000000040",
INIT_04 => X"800000600C600421202100000000BFF0000340408780040EE380041BF8080426",
INIT_05 => X"000000000003FE0000000000000000645202140402000013D71FFF890105B400",
INIT_06 => X"200080600000065F7801285001000000A02980184100610000007E80000AD000",
INIT_07 => X"0400B0C0092001022015C00802002102008007E7E000000001148868C9EE0000",
INIT_08 => X"14B3C80EA076F800880701680006E7BF0230180C100C0000002200A541491010",
INIT_09 => X"00000000000000000000000000000000000003FFFFFFFFFFFF80883A7B42C803",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(25),        -- Port A data input
DOA(0)   => data_read_a_lo_256(25),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(25),        -- Port B data input
DOB(0)   => data_read_b_lo_256(25),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_26_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"85F820440E61E5DDDDDDDDDD81D7FFFFFF8FFE3FDEBCEF7FDFD5FFFFFFF80007",
INIT_01 => X"AA5E3FF033CC1A1BA4993AAC8064328EE9265EAA400ABA7000401AC1DE00573E",
INIT_02 => X"F645FFF78F73EF7DDDE3B57E7C6F72BF89C15D49E0FE675E24302AA9F8D1E5E3",
INIT_03 => X"E7FFD67DF7DE1ADFDBEF578C5479263E7E600053CEFDE25C78BFFE7FDFF77F3F",
INIT_04 => X"FFF000600019C294D19C21E3FFFDFFFBFAFF272787FF302EE3D6F03BBE6057EE",
INIT_05 => X"FFFFFCC1DABFBFFEFF7FFFFB1136267FFFFFFFE7D7EFDE7FFF1FFBFFEBEFFFFF",
INIT_06 => X"7FD9A0671ECB87FF7FEBFADDFDAEBDB23939E23AD10C6B9D1D69FCBF7F6F9FBE",
INIT_07 => X"17794B3BCFB7DA839D8AAA600FBDFF5BFFC567FEEFF3F234094F98D9DBCEFEFD",
INIT_08 => X"D082EF0B3EACFFFFFFFF7BFFFFFFF73F9DBA9D6EAEBF7E7B7C8F77525A85B4C0",
INIT_09 => X"00000000000000000000000000000000000003FFFFFFFFFFFF800B354D1138DC",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(26),        -- Port A data input
DOA(0)   => data_read_a_lo_256(26),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(26),        -- Port B data input
DOB(0)   => data_read_b_lo_256(26),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_27_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"11200008002844CCCCCCCCCC80D7FFFFFF8FFE1F5AB4AB7F5ED5FFFFFFEA8015",
INIT_01 => X"080A0E5012800008002029000029049200080A4000142822000002090A800110",
INIT_02 => X"4441D8370DC3416110A004547C8854AB88011100A0FC000A040022202A1000A0",
INIT_03 => X"97EF9671EFDC1ADDDB97570404512A062A000057CA7F0844783D024B19456E38",
INIT_04 => X"7FF000600019C294D19C21E3FFFDFFEE9A8E252547F7102E93D6603A3C2056EE",
INIT_05 => X"AFCF7842C23E3FD65FFECAC9041202FB2ADCE767554BCC6FEC9FFBBF6B6BFDFF",
INIT_06 => X"6DFCA0760E43875F7BAB7AF4EDAF80B83959EAB8D10463B03008F099E10914AB",
INIT_07 => X"1654452153BC0AC3998AA2200B2BAE5AF54467F8EF78FA3C88E88891D30E774D",
INIT_08 => X"4A825C88A220FFFFCC7F5AFBF93BF43F2DAA956AA6BB7AD42E0FD35A18942440",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF80F91049E10840",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(27),        -- Port A data input
DOA(0)   => data_read_a_lo_256(27),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(27),        -- Port B data input
DOB(0)   => data_read_b_lo_256(27),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_28_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"4128400000606088888888888000000000000000420526004380000000080003",
INIT_01 => X"220A20501184080808802A90006000C202200AA40000A820004A02822A004110",
INIT_02 => X"B24427A5000A440440A21114001A00002288C440A980220A0CA1088828B120A2",
INIT_03 => X"0000000000008000800100041110020C8222220186D182D428827A14E2B25403",
INIT_04 => X"B550000000098210901820A15554000988240303000014000000440000280000",
INIT_05 => X"40900040569400B4342934E101420804D04A727222611E1438000012202401D9",
INIT_06 => X"048028000A46800001601000A00008000002200206A4081A9A92000A040101A0",
INIT_07 => X"03310028020040000CA00828019805006CC0500802D2B086264222463A001C44",
INIT_08 => X"0501710016D0000034380903083410000400400012112631000041104A014050",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF809A223208608B",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(28),        -- Port A data input
DOA(0)   => data_read_a_lo_256(28),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(28),        -- Port B data input
DOB(0)   => data_read_b_lo_256(28),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_29_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A5F0A0540E75C5DDDDDDDDDD81000000000FFE20C60C677EC3D5FFFFFFD80003",
INIT_01 => X"805E1FFFF1C81619E659392E8076B2AE79965E4B402AB858000A0A71FF7FBF3B",
INIT_02 => X"E240FFF78F72EB588DE1A03E016D627D81408809E0FE455E66100001F850C5E1",
INIT_03 => X"E037C67C104E00C793E9038C403806345E4000438F5D604C281FFE7FDFA35F3F",
INIT_04 => X"FFF0000000098210901820A15554BFFBE8572323807E340EE046F41B866813C6",
INIT_05 => X"B8AF84C14A1781FEBF7B77D31026246DDD6B6EE3D3C59C1FFF0003F2A0A4BFFB",
INIT_06 => X"16C9282F1ACE82F32560B25DB402B59200202000022C001515697C2D7A6F8FFE",
INIT_07 => X"02380A338E97988008800068051D550176C167FE03D1B0140545104DFBC09EF4",
INIT_08 => X"2E77BF3F7E2405FFF7FA292FFFF6F700941008040A15263A748175100800B0D0",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF83D7BC7787BF7E",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(29),        -- Port A data input
DOA(0)   => data_read_a_lo_256(29),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(29),        -- Port B data input
DOB(0)   => data_read_b_lo_256(29),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_30_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000222222222225A00000000000140000000800020000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"DF83FF2F7CF80000000000000000000000000000000000000000000000000000",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF80FF3F7F3BF8DF",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(30),        -- Port A data input
DOA(0)   => data_read_a_lo_256(30),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(30),        -- Port B data input
DOB(0)   => data_read_b_lo_256(30),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_31_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"60008010001404444444444400D7FFFFFF8FFE1F0810817F0C55FFFFFFE00000",
INIT_01 => X"08800E0FC20105004A40000200128020129000010020000800000030017FA801",
INIT_02 => X"4401D8120D410161100004407D1050EB80011110017C00804A00222200200800",
INIT_03 => X"87EF8671E7DC18DD5386030004410002280888D2492C0080503D004B19452A38",
INIT_04 => X"4AA000600010408441840142AAA8BFE2000A242407F7000E83D6201A3C0016E6",
INIT_05 => X"AF4F7800042A3F424B56CA080010027B2A040505450A806BC41FFBAD0101BC26",
INIT_06 => X"2058806C0401065F78812A5045A680B03809C018418061800000F0816108144A",
INIT_07 => X"1440000141B40A83810282000A21220A110427E0E520401000008881C10E2200",
INIT_08 => X"000000000000FDFFC8470068F10AE43F00A05028100808402C0F120010000400",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF80000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(31),        -- Port A data input
DOA(0)   => data_read_a_lo_256(31),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(31),        -- Port B data input
DOB(0)   => data_read_b_lo_256(31),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_0_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"DA9918630DD2200000000000012800000040002000A106001180000000008007",
INIT_01 => X"80202100005CD2C7B4E6C1E566434955ED29B05AB311C477A91660C2B4D5208F",
INIT_02 => X"11840040D2AC24048604810082640D046B24CC461E01332121AD800087828206",
INIT_03 => X"080029800001E5202400B85242009129400A2A042000F22200808420C4108104",
INIT_04 => X"000FFF9D8F603C21282300100003000404F0100838008ED10C280E44011DA811",
INIT_05 => X"5000032408000000808000349D2934800010180000802B000060040012120000",
INIT_06 => X"40261C93C1345120821204AE0A41780DC6D01980827218422A0C004092B00A14",
INIT_07 => X"400AF9C0A003557C605D491DA48448900A020810000202AAEA922236141141A2",
INIT_08 => X"9030DA025E0900002300040002000840C204C2C131209008137028AD0779C23B",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF80C11F1127D082",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(0),        -- Port A data input
DOA(0)   => data_read_a_hi_256(0),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(0),        -- Port B data input
DOB(0)   => data_read_b_hi_256(0),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_1_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"C08451022808200000000000002000000000000010000C001108000000028002",
INIT_01 => X"22402100005000008490005046680400213C00142300E04080F4514BA066C00C",
INIT_02 => X"00000000000020044400010000C28410230CC4480000024000A1800182C12400",
INIT_03 => X"00001000000000000810440001002000802880040000A2020000800004000000",
INIT_04 => X"00006D858F602400280300100001400452000008000004A0000004A002090008",
INIT_05 => X"501000209000000080000020010008000090900090000B000000000048484000",
INIT_06 => X"09000900010410A082084002000002000012000214208008A890001284200000",
INIT_07 => X"4005010C10002000042028092400884080000000080A08222A22000200004009",
INIT_08 => X"947022015EA802000108121004000000090A458294C24001820004404205F012",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF81809307840190",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(1),        -- Port A data input
DOA(0)   => data_read_a_hi_256(1),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(1),        -- Port B data input
DOB(0)   => data_read_b_hi_256(1),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_2_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"C4804010026CA010101010110092D555550554161001447431116AAAAA820012",
INIT_01 => X"0A141D0A80440812841911980061967CA10E44C4000CB262012008C8B4780C08",
INIT_02 => X"100400000DD9AA5D050335002951264102C1C141491444444A90028282604143",
INIT_03 => X"82921220A28088500A92560801202412F06202040082080840808000E4110B00",
INIT_04 => X"42200020000040044004010208896AA03288101802A0242A0104843012480048",
INIT_05 => X"861A5082908814018000830A041400220C909115E12C4A02A00AA8054ACAD020",
INIT_06 => X"59510860140403E86A0AC8101AA88502590A401A542022AAAA0210378C24000B",
INIT_07 => X"010500130C048045913A20488481D851900022D048080090A2A0220280044209",
INIT_08 => X"B5013F1C742852CE43805274B40340150B9A8D46B4AE500242A910405294C091",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFFC8A0193716CC3A",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(2),        -- Port A data input
DOA(0)   => data_read_a_hi_256(2),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(2),        -- Port B data input
DOB(0)   => data_read_b_hi_256(2),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_3_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"C0C1002008E008110011001024C366666619989C00A105460141B33333020006",
INIT_01 => X"0004B50C84642830841112880080922C210C4480004812E055808C413181DC6C",
INIT_02 => X"1014001A2DD1BAA94D09640318C2C44822849440480EA80482208882C2050048",
INIT_03 => X"3183106A69989A5449B854A8102C241814A02200110008980280808005100940",
INIT_04 => X"02800040000040804084000020A9599012A1404041B024261084A4284A48426A",
INIT_05 => X"084C60828481CC880890A0020404028281A09081C02081418386630DCACBE422",
INIT_06 => X"5B410840148C02BA740ACA8100A00A283828400A542820800A90A6342866C040",
INIT_07 => X"0005020D0480604185022048040010518011018520110A2A2C208A1040220019",
INIT_08 => X"B000220C748E346521C072F0A541C38C199A8D46B4AE50018A0C004810148090",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF8D4015050C05A8",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(3),        -- Port A data input
DOA(0)   => data_read_a_hi_256(3),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(3),        -- Port B data input
DOB(0)   => data_read_b_hi_256(3),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_4_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"C0CB20AC108100111100001100FC78787806181894884518995E3C3C3C128002",
INIT_01 => X"081425AA60440802840100008184B200A108402040C21260028000C0C400122C",
INIT_02 => X"920406000DC124110442042878C2002022409101485E64140010200892014143",
INIT_03 => X"87840669E7D0189253BE47000009280008000000012E28805080601083130802",
INIT_04 => X"C800000000004084410000002A09B8651202020207C8240E8380941A3A480026",
INIT_05 => X"14308401842A3C60A30184200440000613808401C0020003971E190CC8C94422",
INIT_06 => X"1B750810100D02FD0008C2A0402D080011410A909028432604AB74B20028904A",
INIT_07 => X"0420400900004001142AA0480610B04390803784EC884A00090F984AC90E0119",
INIT_08 => X"044015114600F6E44900731CA503C63C19AA150A8C824001020B024202848090",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFFB5208A0F988902",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(4),        -- Port A data input
DOA(0)   => data_read_a_hi_256(4),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(4),        -- Port B data input
DOB(0)   => data_read_b_hi_256(4),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_5_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"CAC8380F010300111111110000D7807F8048181E94A84D60A555C03FC0120002",
INIT_01 => X"082025234054C8C69416C281E46C6D05A50DA0A0F217E665A82468C854801EAC",
INIT_02 => X"918425025D5524110746040A8752890040A491061F213021492C800087230206",
INIT_03 => X"6860699410016D322440A8DA0620950314200004212C10A25082501400108001",
INIT_04 => X"000FFFFD8F703C2168230012AAA207E424011018B8028E516C681E45831CB911",
INIT_05 => X"041007240429826183011006880D1004421104108202B1405161FD051010B800",
INIT_06 => X"02429C80C53D41A8DE1006824B604A05D690D122917A18678266086280B6004A",
INIT_07 => X"0406B3CD3480653D617FE11C8680A882100228620C804220481000302CD14002",
INIT_08 => X"0FB5FF3F7A550B6269C0046C8500294342B41A0D190C8001837B0AED157C8239",
INIT_09 => X"00000000000000000000000000000000000005FFFFFFFFFFFFC1E3BE7EA3DDBF",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(5),        -- Port A data input
DOA(0)   => data_read_a_hi_256(5),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(5),        -- Port B data input
DOB(0)   => data_read_b_hi_256(5),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_6_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"C0CC0708E06000111111111100D7FF80000FE01E10200D600155FFC000000002",
INIT_01 => X"0800250C41440812842112C018619238A10844B00C14B062001008C094001C2C",
INIT_02 => X"1204201000902411040204000042000008809100000220000020000080010002",
INIT_03 => X"400010080000000208585481800020D004200004000208080082000000121000",
INIT_04 => X"000000005086000044000A02AAA8401432890000000024204000842102480108",
INIT_05 => X"0010008180010020889110006000C2A441A090040200000012000068CA4B4400",
INIT_06 => X"5901080010040128000A428008200800101000008020002D2B89083200220000",
INIT_07 => X"0020410910004041000220480490005080810006E888081880A80040C9000219",
INIT_08 => X"B541FF1F3E2802610100721081840200198A8542A4A250010008000000048090",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF9CE19F3B9FDCBA",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(6),        -- Port A data input
DOA(0)   => data_read_a_hi_256(6),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(6),        -- Port B data input
DOB(0)   => data_read_b_hi_256(6),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_7_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"C48C031862648011111111110000000000000000840844008100000000100006",
INIT_01 => X"0804258020440802842002C012090410A10000B009000060000000C00000000C",
INIT_02 => X"100400100090A4110402042001D2040000809100410220144820000090210042",
INIT_03 => X"40001008001210084840108880600C4034200000000000098080000000100000",
INIT_04 => X"00000000208000484200860AAAA9401100810000000065204001852102CA0428",
INIT_05 => X"00100099010100408384820A241440920A310501C10AC0400200000802830600",
INIT_06 => X"40014A20340D27F32203201048088808011040028029002A8802082200220000",
INIT_07 => X"15010709148C40401108A0CA0E83B81A1001A00404204000000800000080C000",
INIT_08 => X"00000000000000990980406C748102002030D86C382C10850003920010048194",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF94000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(7),        -- Port A data input
DOA(0)   => data_read_a_hi_256(7),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(7),        -- Port B data input
DOB(0)   => data_read_b_hi_256(7),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_8_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"D08800000008001111111111000000000000000084884C009100000000100002",
INIT_01 => X"081025A001440802842002C000090410A10800B000140062000001C80080000C",
INIT_02 => X"100400120000A4110542042801520000008011010102200048200000C0210102",
INIT_03 => X"50000008080202000050448984202CD214200004000208088080000000301000",
INIT_04 => X"800000021000010244405806AAA8001032010000400000005000000102004000",
INIT_05 => X"0010009180010048838000026404C08002B38480800290500280000848CD4600",
INIT_06 => X"09240010048900A0024840A14009080001504880800800040000083200260000",
INIT_07 => X"04000309148040401100A0000600A9429800300404094A0888A8001000804909",
INIT_08 => X"2A303F1F5850050749C052F804C40200092A150A948A44210003020010048000",
INIT_09 => X"00000000000000000000000000000000000005FFFFFFFFFFFFF52080369848B3",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(8),        -- Port A data input
DOA(0)   => data_read_a_hi_256(8),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(8),        -- Port B data input
DOB(0)   => data_read_b_hi_256(8),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_9_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"C4C800100204810000000000000000000000000000000C001100000000000002",
INIT_01 => X"000025AAA0440812840112C000609228A10044B00000B060000008C014000C2C",
INIT_02 => X"B20427920090A4110542042800C2046008C000000002641002302002D2014003",
INIT_03 => X"5000100808000A10085044800000281004200004012E088850827814C2B20003",
INIT_04 => X"CAA0006000104084018401400000401032090000400000A0500010A102014008",
INIT_05 => X"0410008384290028881100000000022400B38084800000101280006548CCFA22",
INIT_06 => X"09640110008011A0024840A10809080801500A8000008221202008328026004B",
INIT_07 => X"C0204309148040401008200164108940808000040089083888A1005008804B09",
INIT_08 => X"97F13F36608800010140121004400200090A058284C244210000000200848002",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF98813550204088",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(9),        -- Port A data input
DOA(0)   => data_read_a_hi_256(9),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(9),        -- Port B data input
DOB(0)   => data_read_b_hi_256(9),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_10_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"C4C800100264811111111111000000000000000084884C009100000000100002",
INIT_01 => X"081025A360440812840112C000609228A10044B00000B060000808C014000C2C",
INIT_02 => X"100400120010A411054204280152000000801101010220104820000090210102",
INIT_03 => X"4000000800000810004800880020040014200000052C00885080000000100000",
INIT_04 => X"4AA000600010408441840142AAA8001400090000000020004000800102400000",
INIT_05 => X"04100082042900408B900002040402A0030004048002C0400200002D8001BC22",
INIT_06 => X"12650010140900A0040080204001080800404AA010080020200008028026014B",
INIT_07 => X"040000091000404001008040060030031001200404084A3880A8000000808310",
INIT_08 => X"3B0568176850000109C0206C040002001030180C180C00010003024210008080",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF9DC39405BE0525",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(10),        -- Port A data input
DOA(0)   => data_read_a_hi_256(10),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(10),        -- Port B data input
DOB(0)   => data_read_b_hi_256(10),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_11_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"C2880203B0600020202020200000000000400000000004000100000000000006",
INIT_01 => X"0824250C40448882840602C168004100A10180B0B4004064000000C00000000C",
INIT_02 => X"1104000010042411060204000042010000801104540220240024000080010042",
INIT_03 => X"4000088800004100204000930200018104200000000000028080000000100000",
INIT_04 => X"000355134A4410692C6086140000001000010000100000C0402000C103962001",
INIT_05 => X"001002300001000080000000C801900000000000800000000220000000000000",
INIT_06 => X"00025600802060A0000000020000080084000000005300000004080200B20000",
INIT_07 => X"0004248920084018401441960402000000000004000000000000000004800000",
INIT_08 => X"0181683650100000010000000400020020000000000000850300808C0518832D",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF9CE13045200411",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(11),        -- Port A data input
DOA(0)   => data_read_a_hi_256(11),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(11),        -- Port B data input
DOB(0)   => data_read_b_hi_256(11),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_12_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"C88A1F83F000020022002200020000000040004000000480012A000000000002",
INIT_01 => X"081025A00054C8C6940202C06F000801A50080B037810465AA0C60C00000008C",
INIT_02 => X"110400125014A4110746042880428100008411010603302100248000C0030106",
INIT_03 => X"4000018800010400044000DB822095C1142000002000102B8080000000100000",
INIT_04 => X"000F9B1B4E8208012E6294080002001000011010200000904800008103978000",
INIT_05 => X"001003BC0101000980000006E80DD00000000080800021000240000000000000",
INIT_06 => X"0002568081A070A08000000300004A04C0801100005380400000084200B60000",
INIT_07 => X"C000820D24806530004001976400000000028004000100000000000000910000",
INIT_08 => X"A4C48D264409000101C0000004C002400000000000000001806000000400832E",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF9C0025401700A6",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(12),        -- Port A data input
DOA(0)   => data_read_a_hi_256(12),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(12),        -- Port B data input
DOB(0)   => data_read_b_hi_256(12),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_13_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"C6CC00100206811133331111580000000000010084084480A320000000100002",
INIT_01 => X"083425A020C40812840552811060DB28A10144A08801F060003809C014000C2C",
INIT_02 => X"114400321014A4110742042803520800408011054102201449240000D4210342",
INIT_03 => X"4800000800016D300048A0880020041014200001832C10A85080020000104400",
INIT_04 => X"5AACE2ED56765C846DC75B56AAAA0010A40901093800EB004C298B010240A800",
INIT_05 => X"04100381042900489B100086080C122003214484800290400A60042D9091BE22",
INIT_06 => X"12410180759900A00430800142004804868051000008004010000822003600CA",
INIT_07 => X"0412B2C9048040306145C0400608308310412804044140104010002006818612",
INIT_08 => X"0FB5F7397E30000109C0246C04401A0052341A8D194C821101530AA515688080",
INIT_09 => X"00000000000000000000000000000000000005FFFFFFFFFFFFE0E7BE7F83DDBF",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(13),        -- Port A data input
DOA(0)   => data_read_a_hi_256(13),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(13),        -- Port B data input
DOB(0)   => data_read_b_hi_256(13),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_14_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"C088000001600222000000005A0000000040014000000480012A000000000002",
INIT_01 => X"08002500004408028400828000600000A10020A00000A060000000C00000000C",
INIT_02 => X"1084000000002411040204000042000000801100000220000028000081010002",
INIT_03 => X"4000000800000000004000800000000004200000000000000080000000108000",
INIT_04 => X"00000D8731063940000210140002001000010000000000004000000102000000",
INIT_05 => X"0010000000010000800000000000000000000000000000000200000000000000",
INIT_06 => X"0000000000000020000000000000080100000000000000000000080200220000",
INIT_07 => X"000000090000400C000000000400000000000004000000000000000000800000",
INIT_08 => X"BF45FF1F3CC80000110000000000020000000000000000010000000000008000",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF81E39533BF4DBE",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(14),        -- Port A data input
DOA(0)   => data_read_a_hi_256(14),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(14),        -- Port B data input
DOB(0)   => data_read_b_hi_256(14),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_15_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"C08800000060022222222222000000000040000000000400010A000000000002",
INIT_01 => X"08002500004408028400028000000000A10000A000000060000800C00000000C",
INIT_02 => X"1004000000002411040204000042000000A01102160220000020000080010002",
INIT_03 => X"4000298800000000244008800000000004200000000000000080000000100000",
INIT_04 => X"000000008000042B242188000002001000010000000000514000004502000011",
INIT_05 => X"0010000000010000800000000000000000000000000010000200000000000000",
INIT_06 => X"0000000000000020000004000040080000000000000010000004080200220000",
INIT_07 => X"0000000900004000001000008400000000000804000000000000000000800000",
INIT_08 => X"0000000000000000010000000000020000000000000000010000000000008001",
INIT_09 => X"00000000000000000000000000000000000005FFFFFFFFFFFF80000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(15),        -- Port A data input
DOA(0)   => data_read_a_hi_256(15),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(15),        -- Port B data input
DOB(0)   => data_read_b_hi_256(15),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_16_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"05104816EA00C199999999998B82D55555055577C0000675C3816AAAAAB80003",
INIT_01 => X"8014102000081213688B1862C400120ADA22C61962221218A90010E0957F0E0E",
INIT_02 => X"C200BAC50001061C8901300A2C0980A50085C801003641100400A00980206443",
INIT_03 => X"E2D5423CB284889002E20281C02900E8CC00000340A9401040162E6680824001",
INIT_04 => X"2FDAC651494D654F010FCA0208282AB240330303829FBF0A61DAFF19988017A2",
INIT_05 => X"252A5018058B9611A81110887160E2205004010210480142D30AA9290000198B",
INIT_06 => X"0050400484141401508000004500050248210008000041000000BC86424A9650",
INIT_07 => X"0208023485003A048820088005000200124342D66130400000008809D0C62220",
INIT_08 => X"1D75310E66E4584AA2AC002B005A631500000000001000005485220000000102",
INIT_09 => X"00000000000000000000000000000000000005FFFFFFFFFFFF80C3183DBECD8E",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(16),        -- Port A data input
DOA(0)   => data_read_a_hi_256(16),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(16),        -- Port B data input
DOB(0)   => data_read_b_hi_256(16),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_17_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"4F74BF57E6E587FFFFFFFFFF92D71999998E665DC000E1D9E8758CCCCCF80000",
INIT_01 => X"2ADE30F033C915094A13393EDEF4B2265284CE4B6F40B85001AE0AB1FA003513",
INIT_02 => X"664123B786736A3991E3A47C1D59727F83855D59A1AC21CA6C30AAA2F8F149E3",
INIT_03 => X"01EF407061DE98DF4182021FC45117E22A0888D2C6F8E0FE6823B275CDE77725",
INIT_04 => X"EDD90A855E9396159B5AEBFD777C19EBC03E272701DDBF0600D8FF080FE617A2",
INIT_05 => X"79639AE01E360FDFCF3BEBFFF17FEE5BBC021EE7D7EDBD79F0067A7300009CCD",
INIT_06 => X"005379675FEBE2F7E860285FE282B5A25822E00003FF001F9FEBA08437291FFC",
INIT_07 => X"D2780225C3B59F058DB28BFEEC394102168741D823F3F0040443B8C558020EE0",
INIT_08 => X"EAB0400D64A8399B47F1000937F4E00D0020100800010630ECAF77105801B3FD",
INIT_09 => X"00000000000000000000000000000000000005FFFFFFFFFFFF80203778BE0864",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(17),        -- Port A data input
DOA(0)   => data_read_a_hi_256(17),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(17),        -- Port B data input
DOB(0)   => data_read_b_hi_256(17),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_18_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"80900040060040000000000040039E1E1E0F80060E1C067E2F81CF0F0F000003",
INIT_01 => X"82500F0000100211A6110064200002886984501A10005048A99041D0557F0A28",
INIT_02 => X"C0404B0000108804C04211220424A28000C0804940226454001080009001A502",
INIT_03 => X"6078001C3080000000EB02801129001CDC40000100810011D008380302004002",
INIT_04 => X"40A662F955E7094500A5D54008A007F028431018808040026081000988000002",
INIT_05 => X"862CE019418B82203B5414007000E000436D2000000200044301F98CA1A12F12",
INIT_06 => X"36888606A41514081581900415241410202980184100E18000002CA9620A9000",
INIT_07 => X"04000A360D029582000000008204360921008066240000000104000060C2B094",
INIT_08 => X"274051317664099AEB04286408082303969048A41A4C084AD080000050000001",
INIT_09 => X"00000000000000000000000000000000000005FFFFFFFFFFFF8026A81B2A5022",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(18),        -- Port A data input
DOA(0)   => data_read_a_hi_256(18),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(18),        -- Port B data input
DOB(0)   => data_read_b_hi_256(18),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_19_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"00014020080007FFFFFFFFFF82D7E01FE008005FC000E7E1C1F5F00FF0380003",
INIT_01 => X"0000000000000004108800000000000104220004006A80000000000000000000",
INIT_02 => X"00009440000005400C0000020400000000000000002200000020000940000000",
INIT_03 => X"6040001C3080000000E20280000900000C000000000000000014440010000010",
INIT_04 => X"40018F03201F7C056400DE0C82A8007000030000808000026080000988000002",
INIT_05 => X"0090040000038200000000000000000000000000000000004300180000003022",
INIT_06 => X"00000000000000000000000000000200000000000000000000002C820C6E9000",
INIT_07 => X"0000000000002000000000000000000000000046200000000000000040C20000",
INIT_08 => X"520020232E240844100800000000230100000000000000000000000000000000",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF80A1321EAA8140",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(19),        -- Port A data input
DOA(0)   => data_read_a_hi_256(19),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(19),        -- Port B data input
DOB(0)   => data_read_b_hi_256(19),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_20_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"00000000000007FFFFFFFFFF82D7FFE0000FF85FC000E7E1C1F5FFF000380003",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000027C00000180004400007E00000000000000000000",
INIT_03 => X"E7C6867DF780000093E60380000900000C000000000000000000000000000000",
INIT_04 => X"1AA01182938901EA66400042A800BFF00003000087E2008EE386009BB8190046",
INIT_05 => X"000000000003BE0000000000000000240000430200400003CF1FF80000040140",
INIT_06 => X"00000000000000000000000000000000000000000000000000007C80000A9000",
INIT_07 => X"5200000000000000002008012D000000404007E6E000000000000008C3CE0000",
INIT_08 => X"80800812380CF801004001031202F73F00000000001120000000000000000402",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF810487600C0004",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(20),        -- Port A data input
DOA(0)   => data_read_a_hi_256(20),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(20),        -- Port B data input
DOB(0)   => data_read_b_hi_256(20),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_21_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"4410801502168D555555555520D7FFFFFF90001F8000057F8D55FFFFFFF00002",
INIT_01 => X"8880BE000439376128C090A2E09240284A30242970600098540084F0017FA04B",
INIT_02 => X"0511481A600817F8800B64437D11428202208800047EF900C80488000085480F",
INIT_03 => X"E7D80EFFF7CC20E513E60BF2044D11000C800040108C0022022B789ECAA60068",
INIT_04 => X"4AA339708A60102128A000100000BFF0000366668780201EE380801FFD140436",
INIT_05 => X"E82F02201003FE424043142491092829200010042020200BC71FF8010000B822",
INIT_06 => X"200A944880344004D8000806010285A00A09801841D2610A8A8A7E87620AD004",
INIT_07 => X"0400821589B43102800083140200010000811FE7E02200000516A82CC1EE0000",
INIT_08 => X"0F35FF3F5E36FDFE78800068F142E7BF0020100800000000F056102100480638",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF80E7BE7F83FDBF",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(21),        -- Port A data input
DOA(0)   => data_read_a_hi_256(21),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(21),        -- Port B data input
DOB(0)   => data_read_b_hi_256(21),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_22_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"6CD0E84501520D555555555524FFFFFFFF90009F8001C17F8055FFFFFFF00000",
INIT_01 => X"0A94BEAFE77D3C314A43D337A45241685290F4CFD22090F85C488C03D57FAC62",
INIT_02 => X"F6157F9A78589FFDD14B756901537001E028C4415900AB14E83DA22A50A5694B",
INIT_03 => X"0827A802001090086000807A1124150890A222023DA002AA52AE78DFEAF6314B",
INIT_04 => X"4AAFBB390A30488569A60142AAAA000304287676087620400446A00045541AC0",
INIT_05 => X"AB7FFAA014A840490B55B62E915D2A21A204059434223328000007AC10111C26",
INIT_06 => X"004B1C0A95B9400000D0060740E01FB25402400206DA180A8A9A020766044540",
INIT_07 => X"0561124C8480FA0545630B5480B002881117300105A340926202228100302A02",
INIT_08 => X"BFC5793F7CEA05FF48C00408F1C800800084422111088C6164DF1284170066A9",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF81E7BD7BBEDDAE",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(22),        -- Port A data input
DOA(0)   => data_read_a_hi_256(22),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(22),        -- Port B data input
DOB(0)   => data_read_b_hi_256(22),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_23_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"8A99D0720284A800000000006A000000005FFF400C1804002D00000000000002",
INIT_01 => X"A00080000420E3E7BC8241B640909201EF20906F206006E5F4E2B4F0200040CD",
INIT_02 => X"A39050087D451C8190084003FC04B16802C11910167EDC8180382AA20006800C",
INIT_03 => X"E7C02FFFF780000017EE0BA0044D00122CC888D0700CC010020D0094F2A38B73",
INIT_04 => X"000CCAAD86201C00280300100000BFF02003404087818A5FE3980A5FF8000017",
INIT_05 => X"EB7FFD010003FF226006CA081110001A0921000141088043C71FFF8180809200",
INIT_06 => X"121000064104000084008000160696210A020000002000800004FEA2020AD004",
INIT_07 => X"100002134014B008841000000801100108000FF7E00000000504880EE5FE8010",
INIT_08 => X"000000000006F800200020040002E7FF1200000008000002F834000000000000",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF80000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(23),        -- Port A data input
DOA(0)   => data_read_a_hi_256(23),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(23),        -- Port B data input
DOB(0)   => data_read_b_hi_256(23),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_24_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000D555555555524FFFFFFFF90009F8001C57F8155FFFFFFF00002",
INIT_01 => X"0000800004202020000000000000000000000000000000805400840000000040",
INIT_02 => X"0010800820001080000840037C00000000000000007E88008380000000040008",
INIT_03 => X"E7C0067FF780000013E603A0000D00000C800000100000000210008001000040",
INIT_04 => X"000065E581003800000200100000BFF0000340408780000EE380001BF8000006",
INIT_05 => X"040000000003FE0000000000000000000000000000000003C71FFF8000003000",
INIT_06 => X"00000000000000000000000000000000000000000000000000007E80098AD00A",
INIT_07 => X"00000000000004800000000000000000000007E7E000000001048808C1EE0000",
INIT_08 => X"8EB2CEAF580EF800100000000002E7BF00000000000000000000000000000000",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF806D2D66331814",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(24),        -- Port A data input
DOA(0)   => data_read_a_hi_256(24),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(24),        -- Port B data input
DOB(0)   => data_read_b_hi_256(24),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_25_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000D555555555524FFFFFFFF90009F8001C57F8155FFFFFFF00002",
INIT_01 => X"0000800004202020000000000000000000000000000000805400840000000040",
INIT_02 => X"0010000820001080000840037C00028600040000007E88008000000000040008",
INIT_03 => X"E7D8067FF7DC38FD53E623A0000D00000C800000100000000200008000000040",
INIT_04 => X"800000600C600421202100000000BFF0000340408780040EE380041BF8080426",
INIT_05 => X"000000000003FE0000000000000000645202140402000013D71FFF890105B400",
INIT_06 => X"200080600000065F7801285001000000A02980184100610000007E80000AD000",
INIT_07 => X"0400B0C0092001022015C00802002102008007E7E000000001148868C9EE0000",
INIT_08 => X"14B3C80EA076F800880701680006E7BF0230180C100C0000002200A541491010",
INIT_09 => X"00000000000000000000000000000000000003FFFFFFFFFFFF80883A7B42C803",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(25),        -- Port A data input
DOA(0)   => data_read_a_hi_256(25),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(25),        -- Port B data input
DOB(0)   => data_read_b_hi_256(25),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_26_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"85F820440E61E5DDDDDDDDDD81D7FFFFFF8FFE3FDEBCEF7FDFD5FFFFFFF80007",
INIT_01 => X"AA5E3FF033CC1A1BA4993AAC8064328EE9265EAA400ABA7000401AC1DE00573E",
INIT_02 => X"F645FFF78F73EF7DDDE3B57E7C6F72BF89C15D49E0FE675E24302AA9F8D1E5E3",
INIT_03 => X"E7FFD67DF7DE1ADFDBEF578C5479263E7E600053CEFDE25C78BFFE7FDFF77F3F",
INIT_04 => X"FFF000600019C294D19C21E3FFFDFFFBFAFF272787FF302EE3D6F03BBE6057EE",
INIT_05 => X"FFFFFCC1DABFBFFEFF7FFFFB1136267FFFFFFFE7D7EFDE7FFF1FFBFFEBEFFFFF",
INIT_06 => X"7FD9A0671ECB87FF7FEBFADDFDAEBDB23939E23AD10C6B9D1D69FCBF7F6F9FBE",
INIT_07 => X"17794B3BCFB7DA839D8AAA600FBDFF5BFFC567FEEFF3F234094F98D9DBCEFEFD",
INIT_08 => X"D082EF0B3EACFFFFFFFF7BFFFFFFF73F9DBA9D6EAEBF7E7B7C8F77525A85B4C0",
INIT_09 => X"00000000000000000000000000000000000003FFFFFFFFFFFF800B354D1138DC",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(26),        -- Port A data input
DOA(0)   => data_read_a_hi_256(26),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(26),        -- Port B data input
DOB(0)   => data_read_b_hi_256(26),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_27_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"11200008002844CCCCCCCCCC80D7FFFFFF8FFE1F5AB4AB7F5ED5FFFFFFEA8015",
INIT_01 => X"080A0E5012800008002029000029049200080A4000142822000002090A800110",
INIT_02 => X"4441D8370DC3416110A004547C8854AB88011100A0FC000A040022202A1000A0",
INIT_03 => X"97EF9671EFDC1ADDDB97570404512A062A000057CA7F0844783D024B19456E38",
INIT_04 => X"7FF000600019C294D19C21E3FFFDFFEE9A8E252547F7102E93D6603A3C2056EE",
INIT_05 => X"AFCF7842C23E3FD65FFECAC9041202FB2ADCE767554BCC6FEC9FFBBF6B6BFDFF",
INIT_06 => X"6DFCA0760E43875F7BAB7AF4EDAF80B83959EAB8D10463B03008F099E10914AB",
INIT_07 => X"1654452153BC0AC3998AA2200B2BAE5AF54467F8EF78FA3C88E88891D30E774D",
INIT_08 => X"4A825C88A220FFFFCC7F5AFBF93BF43F2DAA956AA6BB7AD42E0FD35A18942440",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF80F91049E10840",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(27),        -- Port A data input
DOA(0)   => data_read_a_hi_256(27),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(27),        -- Port B data input
DOB(0)   => data_read_b_hi_256(27),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_28_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"4128400000606088888888888000000000000000420526004380000000080003",
INIT_01 => X"220A20501184080808802A90006000C202200AA40000A820004A02822A004110",
INIT_02 => X"B24427A5000A440440A21114001A00002288C440A980220A0CA1088828B120A2",
INIT_03 => X"0000000000008000800100041110020C8222220186D182D428827A14E2B25403",
INIT_04 => X"B550000000098210901820A15554000988240303000014000000440000280000",
INIT_05 => X"40900040569400B4342934E101420804D04A727222611E1438000012202401D9",
INIT_06 => X"048028000A46800001601000A00008000002200206A4081A9A92000A040101A0",
INIT_07 => X"03310028020040000CA00828019805006CC0500802D2B086264222463A001C44",
INIT_08 => X"0501710016D0000034380903083410000400400012112631000041104A014050",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF809A223208608B",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(28),        -- Port A data input
DOA(0)   => data_read_a_hi_256(28),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(28),        -- Port B data input
DOB(0)   => data_read_b_hi_256(28),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_29_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A5F0A0540E75C5DDDDDDDDDD81000000000FFE20C60C677EC3D5FFFFFFD80003",
INIT_01 => X"805E1FFFF1C81619E659392E8076B2AE79965E4B402AB858000A0A71FF7FBF3B",
INIT_02 => X"E240FFF78F72EB588DE1A03E016D627D81408809E0FE455E66100001F850C5E1",
INIT_03 => X"E037C67C104E00C793E9038C403806345E4000438F5D604C281FFE7FDFA35F3F",
INIT_04 => X"FFF0000000098210901820A15554BFFBE8572323807E340EE046F41B866813C6",
INIT_05 => X"B8AF84C14A1781FEBF7B77D31026246DDD6B6EE3D3C59C1FFF0003F2A0A4BFFB",
INIT_06 => X"16C9282F1ACE82F32560B25DB402B59200202000022C001515697C2D7A6F8FFE",
INIT_07 => X"02380A338E97988008800068051D550176C167FE03D1B0140545104DFBC09EF4",
INIT_08 => X"2E77BF3F7E2405FFF7FA292FFFF6F700941008040A15263A748175100800B0D0",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF83D7BC7787BF7E",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(29),        -- Port A data input
DOA(0)   => data_read_a_hi_256(29),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(29),        -- Port B data input
DOB(0)   => data_read_b_hi_256(29),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_30_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000222222222225A00000000000140000000800020000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"DF83FF2F7CF80000000000000000000000000000000000000000000000000000",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF80FF3F7F3BF8DF",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(30),        -- Port A data input
DOA(0)   => data_read_a_hi_256(30),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(30),        -- Port B data input
DOB(0)   => data_read_b_hi_256(30),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_31_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"60008010001404444444444400D7FFFFFF8FFE1F0810817F0C55FFFFFFE00000",
INIT_01 => X"08800E0FC20105004A40000200128020129000010020000800000030017FA801",
INIT_02 => X"4401D8120D410161100004407D1050EB80011110017C00804A00222200200800",
INIT_03 => X"87EF8671E7DC18DD5386030004410002280888D2492C0080503D004B19452A38",
INIT_04 => X"4AA000600010408441840142AAA8BFE2000A242407F7000E83D6201A3C0016E6",
INIT_05 => X"AF4F7800042A3F424B56CA080010027B2A040505450A806BC41FFBAD0101BC26",
INIT_06 => X"2058806C0401065F78812A5045A680B03809C018418061800000F0816108144A",
INIT_07 => X"1440000141B40A83810282000A21220A110427E0E520401000008881C10E2200",
INIT_08 => X"000000000000FDFFC8470068F10AE43F00A05028100808402C0F120010000400",
INIT_09 => X"00000000000000000000000000000000000001FFFFFFFFFFFF80000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(31),        -- Port A data input
DOA(0)   => data_read_a_hi_256(31),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(31),        -- Port B data input
DOB(0)   => data_read_b_hi_256(31),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


end;