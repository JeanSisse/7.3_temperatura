library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_misc.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library UNISIM;
use UNISIM.vcomponents.all;

entity ram_master is
	port(clk             : in  std_logic;
        address_a       : in  std_logic_vector(31 downto 2);
        enable_a        : in  std_logic;
        wbe_a           : in  std_logic_vector(3 downto 0);
        data_write_a    : in  std_logic_vector(31 downto 0);
        data_read_a     : out std_logic_vector(31 downto 0);

        address_b       : in  std_logic_vector(31 downto 2);
        enable_b        : in  std_logic;
        wbe_b           : in  std_logic_vector(3 downto 0);
        data_write_b    : in  std_logic_vector(31 downto 0);
        data_read_b     : out std_logic_vector(31 downto 0));
end; --entity ram     

architecture ram_master of ram_master is
signal enable_a_lo       : std_logic;
signal wbe_a_lo          : std_logic_vector(3 downto 0);
signal data_write_a_lo   : std_logic_vector(31 downto 0);
signal data_read_a_lo    : std_logic_vector(31 downto 0);
signal enable_b_lo       : std_logic;
signal wbe_b_lo          : std_logic_vector(3 downto 0);
signal data_read_b_lo    : std_logic_vector(31 downto 0);
signal enable_a_hi       : std_logic;
signal wbe_a_hi          : std_logic_vector(3 downto 0);
signal data_read_a_hi   : std_logic_vector(31 downto 0);
signal enable_b_hi       : std_logic;
signal wbe_b_hi          : std_logic_vector(3 downto 0);
signal data_read_b_hi    : std_logic_vector(31 downto 0);
signal address_a_reg     : std_logic_vector(31 downto 2);
signal address_b_reg     : std_logic_vector(31 downto 2);
signal enable_a_lo_256       : std_logic;
signal wbe_a_lo_256          : std_logic_vector(3 downto 0);
signal data_write_a_lo_256   : std_logic_vector(31 downto 0);
signal data_read_a_lo_256    : std_logic_vector(31 downto 0);
signal enable_b_lo_256       : std_logic;
signal wbe_b_lo_256          : std_logic_vector(3 downto 0);
signal data_read_b_lo_256    : std_logic_vector(31 downto 0);
signal enable_a_hi_256       : std_logic;
signal wbe_a_hi_256          : std_logic_vector(3 downto 0);
signal data_read_a_hi_256   : std_logic_vector(31 downto 0);
signal enable_b_hi_256       : std_logic;
signal wbe_b_hi_256          : std_logic_vector(3 downto 0);
signal data_read_b_hi_256    : std_logic_vector(31 downto 0);
signal enable_a_lo_512       : std_logic;
signal wbe_a_lo_512          : std_logic_vector(3 downto 0);
signal data_write_a_lo_512   : std_logic_vector(31 downto 0);
signal data_read_a_lo_512    : std_logic_vector(31 downto 0);
signal enable_b_lo_512       : std_logic;
signal wbe_b_lo_512          : std_logic_vector(3 downto 0);
signal data_read_b_lo_512    : std_logic_vector(31 downto 0);
signal enable_a_hi_512       : std_logic;
signal wbe_a_hi_512          : std_logic_vector(3 downto 0);
signal data_read_a_hi_512   : std_logic_vector(31 downto 0);
signal enable_b_hi_512       : std_logic;
signal wbe_b_hi_512          : std_logic_vector(3 downto 0);
signal data_read_b_hi_512    : std_logic_vector(31 downto 0);
signal enable_a_lo_512_2       : std_logic;
signal wbe_a_lo_512_2          : std_logic_vector(3 downto 0);
signal data_write_a_lo_512_2   : std_logic_vector(31 downto 0);
signal data_read_a_lo_512_2    : std_logic_vector(31 downto 0);
signal enable_b_lo_512_2       : std_logic;
signal wbe_b_lo_512_2          : std_logic_vector(3 downto 0);
signal data_read_b_lo_512_2    : std_logic_vector(31 downto 0);
signal enable_a_hi_512_2       : std_logic;
signal wbe_a_hi_512_2          : std_logic_vector(3 downto 0);
signal data_read_a_hi_512_2   : std_logic_vector(31 downto 0);
signal enable_b_hi_512_2       : std_logic;
signal wbe_b_hi_512_2          : std_logic_vector(3 downto 0);
signal data_read_b_hi_512_2    : std_logic_vector(31 downto 0);
signal enable_a_lo_1024       : std_logic;
signal wbe_a_lo_1024          : std_logic_vector(3 downto 0);
signal data_write_a_lo_1024   : std_logic_vector(31 downto 0);
signal data_read_a_lo_1024    : std_logic_vector(31 downto 0);
signal enable_b_lo_1024       : std_logic;
signal wbe_b_lo_1024          : std_logic_vector(3 downto 0);
signal data_read_b_lo_1024    : std_logic_vector(31 downto 0);
signal enable_a_hi_1024       : std_logic;
signal wbe_a_hi_1024          : std_logic_vector(3 downto 0);
signal data_read_a_hi_1024   : std_logic_vector(31 downto 0);
signal enable_b_hi_1024       : std_logic;
signal wbe_b_hi_1024          : std_logic_vector(3 downto 0);
signal data_read_b_hi_1024    : std_logic_vector(31 downto 0);
signal enable_a_lo_1024_2       : std_logic;
signal wbe_a_lo_1024_2          : std_logic_vector(3 downto 0);
signal data_write_a_lo_1024_2   : std_logic_vector(31 downto 0);
signal data_read_a_lo_1024_2    : std_logic_vector(31 downto 0);
signal enable_b_lo_1024_2       : std_logic;
signal wbe_b_lo_1024_2          : std_logic_vector(3 downto 0);
signal data_read_b_lo_1024_2    : std_logic_vector(31 downto 0);
signal enable_a_hi_1024_2       : std_logic;
signal wbe_a_hi_1024_2          : std_logic_vector(3 downto 0);
signal data_read_a_hi_1024_2   : std_logic_vector(31 downto 0);
signal enable_b_hi_1024_2       : std_logic;
signal wbe_b_hi_1024_2          : std_logic_vector(3 downto 0);
signal data_read_b_hi_1024_2    : std_logic_vector(31 downto 0);
signal enable_a_lo_1024_3       : std_logic;
signal wbe_a_lo_1024_3          : std_logic_vector(3 downto 0);
signal data_write_a_lo_1024_3   : std_logic_vector(31 downto 0);
signal data_read_a_lo_1024_3    : std_logic_vector(31 downto 0);
signal enable_b_lo_1024_3       : std_logic;
signal wbe_b_lo_1024_3          : std_logic_vector(3 downto 0);
signal data_read_b_lo_1024_3    : std_logic_vector(31 downto 0);
signal enable_a_hi_1024_3       : std_logic;
signal wbe_a_hi_1024_3          : std_logic_vector(3 downto 0);
signal data_read_a_hi_1024_3   : std_logic_vector(31 downto 0);
signal enable_b_hi_1024_3       : std_logic;
signal wbe_b_hi_1024_3          : std_logic_vector(3 downto 0);
signal data_read_b_hi_1024_3    : std_logic_vector(31 downto 0);
signal enable_a_lo_1024_4       : std_logic;
signal wbe_a_lo_1024_4          : std_logic_vector(3 downto 0);
signal data_write_a_lo_1024_4   : std_logic_vector(31 downto 0);
signal data_read_a_lo_1024_4    : std_logic_vector(31 downto 0);
signal enable_b_lo_1024_4       : std_logic;
signal wbe_b_lo_1024_4          : std_logic_vector(3 downto 0);
signal data_read_b_lo_1024_4    : std_logic_vector(31 downto 0);
signal enable_a_hi_1024_4       : std_logic;
signal wbe_a_hi_1024_4          : std_logic_vector(3 downto 0);
signal data_read_a_hi_1024_4   : std_logic_vector(31 downto 0);
signal enable_b_hi_1024_4       : std_logic;
signal wbe_b_hi_1024_4          : std_logic_vector(3 downto 0);
signal data_read_b_hi_1024_4    : std_logic_vector(31 downto 0);
begin
process(clk)
begin
if rising_edge(clk) then
	address_a_reg <= address_a;
	address_b_reg <= address_b;
	end if;
end process;
data_read_a <= data_read_a_lo when (address_a_reg < x"0001000"&"00") else
data_read_a_hi when ((address_a_reg >= x"0001000"&"00") and (address_a_reg < x"0002000"&"00")) else 
data_read_a_lo_256 when ((address_a_reg >= x"0002000"&"00") and (address_a_reg < x"0003000"&"00")) else 
data_read_a_hi_256 when ((address_a_reg >= x"0003000"&"00") and (address_a_reg < x"0004000"&"00")) else 
data_read_a_lo_512 when ((address_a_reg >= x"0004000"&"00") and (address_a_reg < x"0005000"&"00")) else 
data_read_a_hi_512 when ((address_a_reg >= x"0005000"&"00") and (address_a_reg < x"0006000"&"00")) else 
data_read_a_lo_512_2 when ((address_a_reg >= x"0006000"&"00") and (address_a_reg < x"0007000"&"00")) else 
data_read_a_hi_512_2 when ((address_a_reg >= x"0007000"&"00") and (address_a_reg < x"0008000"&"00")) else 
data_read_a_lo_1024 when ((address_a_reg >= x"0008000"&"00") and (address_a_reg < x"0009000"&"00")) else 
data_read_a_hi_1024 when ((address_a_reg >= x"0009000"&"00") and (address_a_reg < x"000A000"&"00")) else 
data_read_a_lo_1024_2 when ((address_a_reg >= x"000A000"&"00") and (address_a_reg < x"000B000"&"00")) else 
data_read_a_hi_1024_2 when ((address_a_reg >= x"000B000"&"00") and (address_a_reg < x"000C000"&"00")) else 
data_read_a_lo_1024_3 when ((address_a_reg >= x"000C000"&"00") and (address_a_reg < x"000D000"&"00")) else 
data_read_a_hi_1024_3 when ((address_a_reg >= x"000D000"&"00") and (address_a_reg < x"000E000"&"00")) else 
data_read_a_lo_1024_4 when ((address_a_reg >= x"000E000"&"00") and (address_a_reg < x"000F000"&"00")) else 
data_read_a_hi_1024_4 when ((address_a_reg >= x"000F000"&"00") and (address_a_reg < x"0010000"&"00")); 
data_read_b <= data_read_b_lo when (address_b_reg < x"0001000"&"00") else
data_read_b_hi when ((address_b_reg >= x"0001000"&"00") and (address_b_reg < x"0002000"&"00")) else
data_read_b_lo_256 when ((address_b_reg >= x"0002000"&"00") and (address_a_reg < x"0003000"&"00")) else 
data_read_b_hi_256 when ((address_b_reg >= x"0003000"&"00") and (address_b_reg< x"0004000"&"00")) else 
data_read_b_lo_512 when ((address_b_reg >= x"0004000"&"00") and (address_b_reg< x"0005000"&"00")) else 
data_read_b_hi_512 when ((address_b_reg >= x"0005000"&"00") and (address_b_reg< x"0006000"&"00")) else 
data_read_b_lo_512_2 when ((address_b_reg >= x"0006000"&"00") and (address_b_reg< x"0007000"&"00")) else 
data_read_b_hi_512_2 when ((address_b_reg >= x"0007000"&"00") and (address_b_reg< x"0008000"&"00")) else 
data_read_b_lo_1024 when ((address_b_reg >= x"0008000"&"00") and (address_b_reg< x"0009000"&"00")) else 
data_read_b_hi_1024 when ((address_b_reg >= x"0009000"&"00") and (address_b_reg< x"000A000"&"00")) else 
data_read_b_lo_1024_2 when ((address_b_reg >= x"000A000"&"00") and (address_b_reg< x"000B000"&"00")) else 
data_read_b_hi_1024_2 when ((address_b_reg >= x"000B000"&"00") and (address_b_reg< x"000C000"&"00")) else 
data_read_b_lo_1024_3 when ((address_b_reg >= x"000C000"&"00") and (address_b_reg< x"000D000"&"00")) else 
data_read_b_hi_1024_3 when ((address_b_reg >= x"000D000"&"00") and (address_b_reg< x"000E000"&"00")) else 
data_read_b_lo_1024_4 when ((address_b_reg >= x"000E000"&"00") and (address_b_reg< x"000F000"&"00")) else 
data_read_b_hi_1024_4 when ((address_b_reg >= x"000F000"&"00") and (address_b_reg< x"0010000"&"00")); 
enable_a_lo <= enable_a when (address_a < x"0001000"&"00") else '0';
enable_b_lo <= enable_b when (address_b < x"0001000"&"00") else '0';
enable_a_hi <= enable_a when ((address_a >= x"0001000"&"00") and (address_a < x"0002000"&"00")) else '0';
enable_b_hi <= enable_b when ((address_b >= x"0001000"&"00") and (address_b < x"0002000"&"00")) else '0';
enable_a_lo_256 <= enable_a when ((address_a >= x"0002000"&"00") and (address_a < x"0003000"&"00")) else '0';
enable_b_lo_256 <= enable_b when ((address_b >= x"0002000"&"00") and (address_b < x"0003000"&"00")) else '0';
enable_a_hi_256 <= enable_a when ((address_a >= x"0003000"&"00") and (address_a < x"0004000"&"00")) else '0';
enable_b_hi_256 <= enable_b when ((address_b >= x"0003000"&"00") and (address_b < x"0004000"&"00")) else '0';
enable_a_lo_512 <= enable_a when ((address_a >= x"0004000"&"00") and (address_a < x"0005000"&"00")) else '0';
enable_b_lo_512 <= enable_b when ((address_b >= x"0004000"&"00") and (address_b < x"0005000"&"00")) else '0';
enable_a_hi_512 <= enable_a when ((address_a >= x"0005000"&"00") and (address_a < x"0006000"&"00")) else '0';
enable_b_hi_512 <= enable_b when ((address_b >= x"0005000"&"00") and (address_b < x"0006000"&"00")) else '0';
enable_a_lo_512_2 <= enable_a when ((address_a >= x"0006000"&"00") and (address_a < x"0007000"&"00")) else '0';
enable_b_lo_512_2 <= enable_b when ((address_b >= x"0006000"&"00") and (address_b < x"0007000"&"00")) else '0';
enable_a_hi_512_2 <= enable_a when ((address_a >= x"0007000"&"00") and (address_a < x"0008000"&"00")) else '0';
enable_b_hi_512_2 <= enable_b when ((address_b >= x"0007000"&"00") and (address_b < x"0008000"&"00")) else '0';
enable_a_lo_1024 <= enable_b when ((address_a >= x"0008000"&"00") and (address_a < x"0009000"&"00")) else '0';
enable_b_lo_1024 <= enable_b when ((address_b >= x"0008000"&"00") and (address_b < x"0009000"&"00")) else '0';
enable_a_hi_1024 <= enable_b when ((address_a >= x"0009000"&"00") and (address_a < x"000A000"&"00")) else '0';
enable_b_hi_1024 <= enable_b when ((address_b >= x"0009000"&"00") and (address_b < x"000A000"&"00")) else '0';
enable_a_lo_1024_2 <= enable_b when ((address_a >= x"000A000"&"00") and (address_a < x"000B000"&"00")) else '0';
enable_b_lo_1024_2 <= enable_b when ((address_b >= x"000A000"&"00") and (address_b < x"000B000"&"00")) else '0';
enable_a_hi_1024_2 <= enable_b when ((address_a >= x"000B000"&"00") and (address_a < x"000C000"&"00")) else '0';
enable_b_hi_1024_2 <= enable_b when ((address_b >= x"000B000"&"00") and (address_b < x"000C000"&"00")) else '0';
enable_a_lo_1024_3 <= enable_b when ((address_a >= x"000C000"&"00") and (address_a < x"000D000"&"00")) else '0';
enable_b_lo_1024_3 <= enable_b when ((address_b >= x"000C000"&"00") and (address_b < x"000D000"&"00")) else '0';
enable_a_hi_1024_3 <= enable_b when ((address_a >= x"000D000"&"00") and (address_a < x"000E000"&"00")) else '0';
enable_b_hi_1024_3 <= enable_b when ((address_b >= x"000D000"&"00") and (address_b < x"000E000"&"00")) else '0';
enable_a_lo_1024_4 <= enable_b when ((address_a >= x"000E000"&"00") and (address_a < x"000F000"&"00")) else '0';
enable_b_lo_1024_4 <= enable_b when ((address_b >= x"000E000"&"00") and (address_b < x"000F000"&"00")) else '0';
enable_a_hi_1024_4 <= enable_b when ((address_a >= x"000F000"&"00") and (address_a < x"0010000"&"00")) else '0';
enable_b_hi_1024_4 <= enable_b when ((address_b >= x"000F000"&"00") and (address_b < x"0010000"&"00")) else '0';
wbe_a_lo <= wbe_a when  enable_a_lo='1' else x"0";
wbe_a_hi <= wbe_a when  enable_a_hi='1' else x"0";
wbe_b_lo <= wbe_b when  enable_b_lo='1' else x"0";
wbe_b_hi <= wbe_b when  enable_b_hi='1' else x"0";
wbe_a_lo_256 <= wbe_a when  enable_a_lo_256='1' else x"0";
wbe_a_hi_256 <= wbe_a when  enable_a_hi_256='1' else x"0";
wbe_b_lo_256 <= wbe_b when  enable_b_lo_256='1' else x"0";
wbe_b_hi_256 <= wbe_b when  enable_b_hi_256='1' else x"0";
wbe_a_lo_512 <= wbe_a when  enable_a_lo_512='1' else x"0";
wbe_a_hi_512 <= wbe_a when  enable_a_hi_512='1' else x"0";
wbe_b_lo_512 <= wbe_b when  enable_b_lo_512='1' else x"0";
wbe_b_hi_512 <= wbe_b when  enable_b_hi_512='1' else x"0";
wbe_a_lo_512_2 <= wbe_a when  enable_a_lo_512_2='1' else x"0";
wbe_a_hi_512_2 <= wbe_a when  enable_a_hi_512_2='1' else x"0";
wbe_b_lo_512_2 <= wbe_b when  enable_b_lo_512_2='1' else x"0";
wbe_b_hi_512_2 <= wbe_b when  enable_b_hi_512_2='1' else x"0";
wbe_a_lo_1024 <= wbe_b when  enable_a_lo_1024 ='1' else x"0";
wbe_a_hi_1024 <= wbe_b when  enable_a_hi_1024 ='1' else x"0";
wbe_b_lo_1024 <= wbe_b when  enable_b_lo_1024 ='1' else x"0";
wbe_b_hi_1024 <= wbe_b when  enable_b_hi_1024 ='1' else x"0";
wbe_a_lo_1024_2 <= wbe_b when  enable_a_lo_1024_2='1' else x"0";
wbe_a_hi_1024_2 <= wbe_b when  enable_a_hi_1024_2='1' else x"0";
wbe_b_lo_1024_2 <= wbe_b when  enable_b_lo_1024_2='1' else x"0";
wbe_b_hi_1024_2 <= wbe_b when  enable_b_hi_1024_2='1' else x"0";
wbe_a_lo_1024_3 <= wbe_b when  enable_a_lo_1024_3='1' else x"0";
wbe_a_hi_1024_3 <= wbe_b when  enable_a_hi_1024_3='1' else x"0";
wbe_b_lo_1024_3 <= wbe_b when  enable_b_lo_1024_3='1' else x"0";
wbe_b_hi_1024_3 <= wbe_b when  enable_b_hi_1024_3='1' else x"0";
wbe_a_lo_1024_4 <= wbe_b when  enable_a_lo_1024_4='1' else x"0";
wbe_a_hi_1024_4 <= wbe_b when  enable_a_hi_1024_4='1' else x"0";
wbe_b_lo_1024_4 <= wbe_b when  enable_b_lo_1024_4='1' else x"0";
wbe_b_hi_1024_4 <= wbe_b when  enable_b_hi_1024_4='1' else x"0";



ram_bit_0_16 : RAMB16_S1_S1
generic map (
INIT_00 => X"ED39BA795990D275FB4A6E96ACC4731DEA4598B0AFB54867F6EE4618C3749803",
INIT_01 => X"8AA0047D8607944AC7DA180001ECA2444042106208408208C20022E9173734B3",
INIT_02 => X"1A7DDD79F9A73E6CCA7DAAF00001000008478020113D98E382FEDF333027C80F",
INIT_03 => X"75D341110C58F31110C58F32A208921F8051500147A0E4AB3493FB3A01EBE240",
INIT_04 => X"86424001531009B100425A97B2AA0001E03501D0A39C8F0078420001106D0C4C",
INIT_05 => X"BCC8CA2EBF03400700402BB20F00239E20341699198600000B08694B16434804",
INIT_06 => X"103FB860B2800161F8432200012DA185F80F24081C3C0707800E600056881308",
INIT_07 => X"B24197ABCDA467F9A73E6CCAFDC3870EEEEC44E2BDFE220094D03022210C011C",
INIT_08 => X"240581B5695EAA80262C080032BF07C7C1FC3F8E94F65B11555EAFFC1C306758",
INIT_09 => X"7E40000BEC004170040DB60017FED1CC0001045002984202003DB931192D60A5",
INIT_0A => X"120071411A74315881A28C141118000C5A85A60444210123820B43B40804674D",
INIT_0B => X"0820008E514045BB514F0106D1D8599581D3A958BC104A89215AC14C48898403",
INIT_0C => X"C261C01C48B1584A0CA3E2687A9A1E2687A9A1E2687A9A1E26870CD061343885",
INIT_0D => X"D274E93A758FA8683AC54B287522E10A74AF4AA59C568752662F5AC218000002",
INIT_0E => X"FF83C002783A0904231C70470C7E0B92800224008AE09FAD4BD48D1FC5D3A4E9",
INIT_0F => X"5BFF078004F075885DFBF7E15C06101C55E921F1F80FAB7FE0F0009E0E903EAD",
INIT_10 => X"F12E0380231F13978FF023FAFDBD9870380230F2D6081F56FFC1E0013C1D207D",
INIT_11 => X"DE7F263C0C8700125C0F8F3C43F1F10BBF7EFC61E01804E1E6C8F8FE807F67FB",
INIT_12 => X"02BE00017C17C1007E5E2E3081C5AC007E6F0E3081C5AC44418D65FE45DEE55B",
INIT_13 => X"61E0042786F103E9F01F9BC3C120C5A703E9F01F978B8C20666703E9F8A0FFED",
INIT_14 => X"FA7E283FFB414F80005F05F10FA7E283F78F6511C048278DCA174FF038FF15B4",
INIT_15 => X"0066A20B61692F293185D8D724E15D3FCC6B7C236FE0691B0700132C1F0EF880",
INIT_16 => X"3A4E93A4E93A4E93A4E93A4E93A4E93A4F942F92E9628540AD2A91442525A000",
INIT_17 => X"A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E9",
INIT_18 => X"4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93",
INIT_19 => X"55F3898E09B56C74DAB15D1CF13501AA495000000000000000003A4E93A4E93A",
INIT_1A => X"082082082082082082082082082082082082082082082082082084E41DC71C71",
INIT_1B => X"E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F82082",
INIT_1C => X"FFFFFFFFFFFFFFF94A5294A5294A5294A5294A52800003E1F0F87C3E1F0F87C3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"3060C183060C187FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"BDEBA0000000000000000000000000000000000000000000003060C183060C18",
INIT_28 => X"168ABA002E82145085155545F7AA975EFFFAABDE00FFAEBDFFF5D2EAAAAAF7AE",
INIT_29 => X"7FFFE10005542145557FD5545FF8000155087FC0155F7D168B55007BFDF45085",
INIT_2A => X"7FFC0010080017555555568AAAFFFFD7545AA8028A00A2802AABAFF8028BEF5D",
INIT_2B => X"FF842AABAA2AE95545FFD168ABAF7AEAAAAAA2FFFDF4500043FE105D2E954BAF",
INIT_2C => X"5007FD7400550415410002E974BA5D5168A00A2D142155005142010FFAE820AA",
INIT_2D => X"FFF780000BA007FE8AAAFF803FFFF5D2A821550000000BA007FD55FF5D7FC014",
INIT_2E => X"000AAFBEAA00007BFDFFF082EBDF455D5142000082E82145FFD17DFEFFFD168B",
INIT_2F => X"DFD75D2AA8A80EA8E2FE3F000000000000000000000000000000000000000000",
INIT_30 => X"68B551475FAF6D1C556F0AA1C24AABEA495FC716F002A975FFE3AA95E00EBAEB",
INIT_31 => X"42A0070071C50BAFEF1FAE0016D56A16D557BC257D415E0216FA3F1E8FC0145B",
INIT_32 => X"8010E004924874825D7FEAA85487FD24AFE3D02DAAAE12BD5545A2803AA00005",
INIT_33 => X"120155EA568E870BAEB8A05A2AEA8B50F55A2F150005A3A438BD04AFAB8F550A",
INIT_34 => X"545E055FFBE81D0BE8EA8A3AA05A2A5504001C74BA42A1571E8028E3DB7816D0",
INIT_35 => X"A5C7E3DFFFE90B45B47ABA497A82FFAFD2A82485FD2415A105C21451ED42A002",
INIT_36 => X"00000000000000000000B55EAAA100AA1D0F6F480B6A555A2A57A002A3D5FDB6",
INIT_37 => X"5EFAAAAB5E1AF3AABFF45592E88A0AFE80A8B0A0000000000000000000000000",
INIT_38 => X"65F520EBE9EF67D7BEA1FD5D556ABEF5D557FEBA55022A3F70C6B405F4D2AE97",
INIT_39 => X"C114728007521170821CE0FDE69411A8DED57CE1055555E5F58EFFC01FE2CACB",
INIT_3A => X"42341D5DEEBEF55080034E0A592A4AD0079C75D6070CC5CBB0280C029ABAA3EB",
INIT_3B => X"7F353AAF6C77F7F20D968BF57812A95E02A2AAB5EB0F280800EFAEE9F5D18F31",
INIT_3C => X"C91565455C141E41887D58AC448B69C30E02116220415A9540AA854140A0A204",
INIT_3D => X"DE6BE93172D7D625B556EEAB157ABEBE1B4D792A4AD1183454180DD3FDCAAAB7",
INIT_3E => X"F0000001FF0000001FF0000001FF0000001FF01EABC4B8014174FF7DA80F52FE",
INIT_3F => X"FF0000001FF0000001FF0000001FF0000001FF0000001FF0000001FF0000001F")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(0),        -- Port A data input
DOA(0)   => data_read_a_lo(0),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(0),        -- Port B data input
DOB(0)   => data_read_b_lo(0),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_1_16 : RAMB16_S1_S1
generic map (
INIT_00 => X"212C001411984004084D000508C53810A03D1450E839B003342114428A000803",
INIT_01 => X"00000019400B100A8196000000CC004400400002000000000000028001340000",
INIT_02 => X"052137AE8031800C0044009000000000061800001CD4019802AD04CCCFC20004",
INIT_03 => X"04514108C60C21008C6042108400000201440020505100000043C30E10E9F000",
INIT_04 => X"02104001011DEFE088805681920000008000004001900800004002108C280008",
INIT_05 => X"040002340105000200000000080001900010000108040000000008411600401C",
INIT_06 => X"1034001042800808201000000001000820020000102000040000000000800180",
INIT_07 => X"64BF81A15EDFDE8031800C00843060C19E030022103600000450020800040004",
INIT_08 => X"00008004691687AA840008000090248CC84E000046000311555521F183060AC5",
INIT_09 => X"0820800D08100171000DB000154440C800400500000852020011200201012021",
INIT_0A => X"02000040001000880A2A04445004000102002041000001008208001440004140",
INIT_0B => X"4820018A1140440078050040511000102000A008183000010002404400000000",
INIT_0C => X"1000C80008000C030030880C2A030A00C28030A80C2A030A00C28018D4061401",
INIT_0D => X"10040802050080200284401C0022880F009E08008205C0020118088018000000",
INIT_0E => X"0F03C00280000000420860C60C0C0B92C0000000004000010042000040102008",
INIT_0F => X"001E078005000108400005E11C0610000000288058000003C0F000A000100000",
INIT_10 => X"F10E0380000000C202300000008D187038000000480800000781E00140002000",
INIT_11 => X"806302380C870010000004400100110800007861E0180000000C400680000001",
INIT_12 => X"023E00000000018000580C308000050000610C30800005000215006800000101",
INIT_13 => X"61E0000000018100B0001843812000014100B00016030C20000141002880026D",
INIT_14 => X"400A20009B404F80000000018400A20044096111C04000000304026000501580",
INIT_15 => X"0046820040082300218450C2800010094000482141E060190700100000002200",
INIT_16 => X"020080200802008020080200802008020080008008600500A82A1100A8000000",
INIT_17 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_18 => X"0080200802008020080200802008020080200802008020080200802008020080",
INIT_19 => X"81328A46BABEFC54A0810C7452B4428A14000000000000000000020080200802",
INIT_1A => X"AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA28A28A28A28A2A8218D2C0C924925",
INIT_1B => X"E974BA5D2E974BA5D2E974BA5D2E974BA5D2E975BADD6EB75BADD6EB75BAAAAA",
INIT_1C => X"FFFFFFFFFFFFFFFD8C6318C6318C6318C6318C63000002E974BA5D2E974BA5D2",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"70E1C3870E1C387FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"5555500000000000000000000000000000000000000000000070E1C3870E1C38",
INIT_28 => X"EBDF455D2EAABEFF7FFE8BFF5D0002155557FFFFFF007FC21EFA2FFD74AAAAD5",
INIT_29 => X"AA95400552AAAABAFFD1574105D7FD75FFAAAA800AAF7AA974BAFFFBE8B45F7A",
INIT_2A => X"0517DF555D2EAAA1055000015500557DF45AAD1400BAA2AE801550051555EFF7",
INIT_2B => X"FFD540155557FD5400F78028BFFFFFBEAB55F780020AAAA80020AA082EAAB550",
INIT_2C => X"AFF842ABEF5D517DF55552A974AAF7AE820AA0851574BAA2D1574AA5D7BFDEBA",
INIT_2D => X"EFAAD1575EF557FFFE10557FFFFFFFFD56AAAAFFFFD7555AAD168B45AAAEAAAB",
INIT_2E => X"0005D7FFDF4500043FE105D2E954BAF7AE80010082A97410557FEABFFAAFBE8B",
INIT_2F => X"51C7A2FBD5490BFD1C056A000000000000000000000000000000000000000000",
INIT_30 => X"974BAF7FFEFB45FFAABDF55492AA8BC2EBDFEAF7F1F840017D4975D2FEF147FC",
INIT_31 => X"080BEF495FC71D54124924385FAAA8AAAE3D145410F7F1D55D71C002DABAEBAA",
INIT_32 => X"002D082082AB8B6DBEDB7DF7F540E2AE85028B40155145F7AF6DBED5450AA1C2",
INIT_33 => X"78E021FF1471FDEAAFFD56F16D5571D2E28E38E0216FA2D1E8E80140F45082B4",
INIT_34 => X"A2DA3FB7DAAD4AAAAF487BC70BFA97F7AF6D417E92482BF84020BA495557E3FF",
INIT_35 => X"55554ADBD7A2FFC7BEFF6FFD7FC7002FD74951D71EDFFABFD16FAAAE92BD5545",
INIT_36 => X"00000000000000000000547AB8F550A8010E00492487482FFFE82A85EBAE2FFC",
INIT_37 => X"1EF005162BEF047FD5545AAFBF7400FBF9424F70000000000000000000000000",
INIT_38 => X"714F8338AAAA1D0AE974AAF7FFFDF55F7AABFF55082CA8B4DF6C1E8F5E540002",
INIT_39 => X"EABEF75550ACBB7582225FF5843404547184164AA5D2EBEEB0A2D555410D3555",
INIT_3A => X"FEAAEB083BC1000FF8409000512AEABFFDF79DCBF755962010BDCBBC21455D7F",
INIT_3B => X"801F8BA0C57740BDAA0688E5405D57D412F7D55F5E50C7F401BAAE8403CF5A3F",
INIT_3C => X"5D16BABAA3EBC3157ABD5FFE55F2AA9FEAFDF7F431A9F7FFE81FF013A8001AFF",
INIT_3D => X"FB863550229BCABEB7DA403FFFDA2FBF7FED2C7F955445079E280A00C56145EF",
INIT_3E => X"0000000000000000000000000000000000000596EBEF55080034E0A592A4AD00",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(1),        -- Port A data input
DOA(0)   => data_read_a_lo(1),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(1),        -- Port B data input
DOB(0)   => data_read_b_lo(1),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_2_16 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10E006600180111284380310006289800480032283E000A34301002001A0817",
INIT_01 => X"0005A00810790848048044A54E404350404000720885800802000906E4910200",
INIT_02 => X"407004208400408044C600C50AA055254010541A110222841200000002402544",
INIT_03 => X"0600011004182401004102408C28414043101000408118000145840440F5C415",
INIT_04 => X"5035855703A2900A000CD3088400F40688C9844409060850925E58A4081A0221",
INIT_05 => X"0200840D1021A15AC50494894850890540D1E12020C6E510818500440A280090",
INIT_06 => X"113044094002801020440090A8011A1224AB9380552102442884882A20004097",
INIT_07 => X"000100880004428400408044860000008C022402102100AA40004404B5075460",
INIT_08 => X"15C23440408C862A2A12382A8A5244145048C06085008010141521F000001240",
INIT_09 => X"400582B9033AA0E7AA4110B0506744810554542450694E710A836188C2C00222",
INIT_0A => X"443518360012C2210B020414109130A28038188096A06B8C120CA440A9C00802",
INIT_0B => X"1345E53300EC68005605002964AF222A5704004D080211121C80024200821780",
INIT_0C => X"181080C1110C882202211488452213C88472213C88472213488441109A442231",
INIT_0D => X"008204440210091341208041000810C00000300220201800A908000038AD0284",
INIT_0E => X"00040002804180300E88D28D206A40000554815500481440300000C44A081100",
INIT_0F => X"000008000500828700000000010000000002380000A00000010000A010050000",
INIT_10 => X"00010000000004CA000214000000020000000000684280000002000140200500",
INIT_11 => X"000000000020000000000442100002840000000800000000010C000026000000",
INIT_12 => X"00000000000805A4800000000000152300000000000015801272000100210020",
INIT_13 => X"000000000101C00000C000000000000940000120000000000009600004050000",
INIT_14 => X"0000130000000000000002018000106000000000000000002380000141000000",
INIT_15 => X"55000190000000000002000280000000011080C0000000000000000000002310",
INIT_16 => X"40902409064190641906419024090244902A9003004800415120D4A190804241",
INIT_17 => X"0900409004090641906419064190240902409024090641906419064190240902",
INIT_18 => X"9044090040900409004190441904419044090040900409004190441904419044",
INIT_19 => X"75960040138D70C030B51C50C7D100A2052F81F81F83F03F03F0419044190441",
INIT_1A => X"0410410410410410410410410410410410410410410410410248602081659659",
INIT_1B => X"5128944A25128944A25128944A25128944A25128944A25128944A25128941041",
INIT_1C => X"FFFFFFFFFFFFFFFE1084210842108421084210843FFF825128944A25128944A2",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"7FD5FF555815607FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"2AA000000000000000000000000000000000000000000000007FD5FF55581560",
INIT_28 => X"FC21EFA2FFD75EFAA8415410AA8415555087BFFF55A2AA800BAFFAE954000800",
INIT_29 => X"84155EFA2AEBDEAAA2FBEAABA5D7FE8B555551421455D0002145552EBFEBA007",
INIT_2A => X"2AEBDF555D2E954BAA2AA974BAFFFFE8B45552EBDF45FFAEAABFFF7FFE8B55F7",
INIT_2B => X"AAAAAAAAAFFD1574105D7FFFF555D2AAAAAA5D2E820BAA2FBEAB5555557DF55A",
INIT_2C => X"50055575EFFF84021555D043DEAA5D04021EF557FC21FFAA8428BFFAAAA954AA",
INIT_2D => X"10085568A00FF80175FFA2D17DFEFF7800215500557DF55AA80001FFAA800015",
INIT_2E => X"0005D00020AAAA80020AA082EAAB5500517DF555D042AA10A284154005D00154",
INIT_2F => X"00AAFFAA9543A080038A2A000000000000000000000000000000000000000000",
INIT_30 => X"0017D5D20B8EAA007FC51C7A2FBD55D2BE800042AFE8E1557D0075D2F45BEAA8",
INIT_31 => X"AA8BC7EBDFEAFEFFD00105FFBC20BDEAAA2FBF8AAA557BE8B6D5D5FFABEF4904",
INIT_32 => X"FFEFB6D555578F7DB6A0BDF7D480E174BFA02A974BAF7F5EFB455D2ABDF55492",
INIT_33 => X"ED1FDE90E3A497492B6AAADAAAE3D155E105571D55D71C002DABA5524820BAB6",
INIT_34 => X"BE8F401D7B6A0001470155C51D0092A071555D5E3AE821D00001FF0871C016DB",
INIT_35 => X"5BE8555400550A38428007FED000E3DA3DFD5E3DFFFBD5A38A021551C5F7AF6D",
INIT_36 => X"00000000000000000000410F45082B4002D082082AB8B6D1C5B7DF7FF78E075C",
INIT_37 => X"5EF005560B55F7AA800AAF7AA954AA00042AAA20000000000000000000000000",
INIT_38 => X"ABEF057D68F5F5A00021EF55042AAAA007FD5555AAFBD7545FBB8020A3F7AE97",
INIT_39 => X"7DF55D7AABFF5428ACA8F45A6C1E8F5EFF84165EFF7802BAB0A2FFEAABA557BE",
INIT_3A => X"CA8AA80800020AAF7FBFFFEF04552ABFFFF841FFE75CA882108202E974AAF7D5",
INIT_3B => X"00151FF0C57401E5F3D1E00A1A884174A8FFAEBFEB0A2D55541051555694F002",
INIT_3C => X"2AA801455D7FE8BFFF680800FFF7AAA155F595542455512A975455D3AA8A0055",
INIT_3D => X"5D79FCAF774AE005BE7895554005D2A8A0B882FFFFE10AAAAAB755A66B6AF56A",
INIT_3E => X"00000000000000000000000000000000000000C3BC1000FF8409000512AEABFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(2),        -- Port A data input
DOA(0)   => data_read_a_lo(2),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(2),        -- Port B data input
DOB(0)   => data_read_b_lo(2),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_3_16 : RAMB16_S1_S1
generic map (
INIT_00 => X"210C00A20020000108430020001600B8156021104940741B3530400E02B92203",
INIT_01 => X"014C9BCA58B1296D24A402C992500B69404040028804A0080A000416A8D90A08",
INIT_02 => X"C12026A484318004404405C9C66E331352180D468B8203980300204442E02B34",
INIT_03 => X"04000748D60D24648D60524C88804D0215011020D15018148040C10A70E1D58C",
INIT_04 => X"18283333240FE41244187308C9104D70944852640901083801750EB0A418C220",
INIT_05 => X"0613142D01912CC2A1B4140528348900C612A104201C689044340ED413A07649",
INIT_06 => X"119000034019881822104C5E68035250A222829710A0A02C18C01A9920842413",
INIT_07 => X"402F00AB0016CA0431800444841020509D038B021230C1990001C644C8273200",
INIT_08 => X"16905000408482088290E8E64010248C4A5AA840C2000110001521F0810A92E7",
INIT_09 => X"0003CE6581BD016342A951AB146C4480530C3B2A8088D3542651670200C1826A",
INIT_0A => X"00735D36209A8A20020894004284B660821030C8990467401218004041020002",
INIT_0B => X"512445B740457154562F957CC08B00093700080D0A4851001D8302D20A0A1530",
INIT_0C => X"00508650008008021021A40861021840869021A408610218C0869810D6043095",
INIT_0D => X"1C8508438450801043A08090380A8834207007022209038080190000999C8F84",
INIT_0E => X"000400200000C0002A48A206204C4205F3304B33004C0041006240140A1C310A",
INIT_0F => X"0000080040000083800400000100000000008400018040000100080000510100",
INIT_10 => X"0001000000000800000244040000020000000100002A0080000200100000A702",
INIT_11 => X"000000000020000000200000080002C000800008000000000022000006808000",
INIT_12 => X"0000000000000A2281000000000040A3810000000000402001400000022002A0",
INIT_13 => X"000000000004200001C0400000000010200001C0400000000010000004490010",
INIT_14 => X"0001070004000000000000060000104C08000000000000001000000903008000",
INIT_15 => X"CC004050CA0C00020220200070040000010401C4000000000000000000100008",
INIT_16 => X"4310E4310A4210A4210A4210A4210A4210A8D0830A68010001B4DA881048061C",
INIT_17 => X"21084290A4210A4210A4210A4210A4210A4210A4210E4310E4310E4310E4310E",
INIT_18 => X"90A421084290A421084390E4310C4390E4310C4390E4310C4290A421084290A4",
INIT_19 => X"015303C0C78C706428A14C586291000A044001FFE000003FFC004290A4210842",
INIT_1A => X"2492492492492492492492492492492492410410410410412821600001249249",
INIT_1B => X"51A8D46A351A8D46A351A8D46A351A8D46A351A9D4EA753A9D4EA753A9D49249",
INIT_1C => X"FFFFFFFFFFFFFFFC00000000000000000000000038F56351A8D46A351A8D46A3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"55AB02055AB0207FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"420000000000000000000000000000000000000000000000007FFFAB57FFFAB5",
INIT_28 => X"A800BAFFAE9554508002AA00AA843DF55FFAA955EFA2D168B55557BEAA000055",
INIT_29 => X"002AB55AAAA955EF005568A00087BE8BFFA2D155410AA8415555087BFFF55A2A",
INIT_2A => X"AAABFF5508003FF555D0002145552ABFEBA007FC21EF007FD75FFAA841541008",
INIT_2B => X"082EBDEAAA2FBEAABA5D7FC0155005168B455D042AB45F7FFD741000042AA10A",
INIT_2C => X"FF7FBEAB55F7AABDEBA5D7FC2010A2D1575FFF7AA975555D2E80145F78415545",
INIT_2D => X"EF5555554AA087BC01FFFFAAAAB55552A954BAFFFFE8B55552EBDE00F7AEAABF",
INIT_2E => X"000082E820BAA2FBEAB5555557DF55A2AEBDF555D2E954BA002EAAABA002A821",
INIT_2F => X"FB7D5D7FEAA3808554203A000000000000000000000000000000000000000000",
INIT_30 => X"1557D1475FAF45BEAA800AAFFAA95578080038A2AA28E3AF55E3A0BA5D7AADB6",
INIT_31 => X"BD55D7BE80004AA1E8E2AB55B6A0925D7085F6AA10087FEABD7AAD57AEBAB68E",
INIT_32 => X"F5D0438140E2FA38B6AEBFF6D1D04AAFFA41040017D5D20B8EAA007FC51C7A2F",
INIT_33 => X"D0A901FFFF801557D1C20B8EAAA2FBE80AA557BE8B6D5D5FFABEF49002FB55FF",
INIT_34 => X"5D20BDE00EBAAA8BC7EBDFEAFEFAB8ABAE925D21C7010EADB525D7FFAE975C75",
INIT_35 => X"F002EADA921420871D74971D24820875C21D5EB8AA8FFF012A954BAFFF5EFB45",
INIT_36 => X"000000000000000000001C24820BAB6FFEFB6D555578F7DB6A0BDF7DEB8E125F",
INIT_37 => X"B55A28408145AAFFFFFFF5D7FEAABA0051400A20000000000000000000000000",
INIT_38 => X"AB55FAD568AA2AFAE975EF555168B55F7AA800BAF7AA955EF00042AAA2A2AEAA",
INIT_39 => X"2AAAA007FD55558A7BD7145FBB8020A35D2ABEF55F7800015F087FEAA00007FE",
INIT_3A => X"968F575D003FF55F7D5420BA5D2ABFEAAF7AE9DFF759A82AEF70800021EF5504",
INIT_3B => X"FFD5145FBAC9755F05040255FFD84175EF55002AAB0A2FFEAABA557BEA3EF057",
INIT_3C => X"82E974AAF7D57DF45552A3FF10AA8429F45A7D5EAF5FFBAEAAA10554155400AA",
INIT_3D => X"FF843FFE77C80825BC052ABFE10550415557085540000005156155FE90A8F5C0",
INIT_3E => X"00000000000000000000000000000000000005500020AAF7FBFFFEF04552ABFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(3),        -- Port A data input
DOA(0)   => data_read_a_lo(3),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(3),        -- Port B data input
DOB(0)   => data_read_b_lo(3),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_4_16 : RAMB16_S1_S1
generic map (
INIT_00 => X"A108400020612C80284210081034849800A00030300004833522C82D04A16002",
INIT_01 => X"2043998A1839284D1CA0650E1E504368403008418984014902030806A0D10200",
INIT_02 => X"C120042200000000044441CE01E80F00A49043118680008002000000026208E4",
INIT_03 => X"040001020019200020011209CC0164C060000000690111040144800042F5C403",
INIT_04 => X"7029AF0F81A00010CCA47700CC513CAC0D0B8E02010740E19754080108988021",
INIT_05 => X"02139405007133C0712244CD20F20105D583000020E9892201D304D42A9835E1",
INIT_06 => X"9190440300078002014405D9EE814C0284A883B6D7038AE079059B7800048092",
INIT_07 => X"000100AA0004408000000004840400008D200102503000782000C00C8025C000",
INIT_08 => X"00728A00408403220811991E02120C044058080004000001101121F220000260",
INIT_09 => X"811001E1185B38AD23C3707AD46440818F3CF80EC423CA7D01D123C80200816A",
INIT_0A => X"45810810A01B40216361056D6150F41200280001900439001FD8A00041400000",
INIT_0B => X"11FC88076266E800D605402962A820211500024808010512C40106D222223B14",
INIT_0C => X"0408804116040B02C02C500B0C02C100B0C02C100B0402C300B0401618058611",
INIT_0D => X"040200050200501301208482200D00D0A0408402C4282200A84800009B878680",
INIT_0E => X"00000020000100024AC88300300060090F0D830F00025400300204D018000804",
INIT_0F => X"8000000040000206A2000800000000000000950002E010000000080000588040",
INIT_10 => X"0000000000000808000554000200000000000100006D0020000000100000BB00",
INIT_11 => X"0000400000000000002000001A0002504001000000000000002280000D800800",
INIT_12 => X"0800000000000E2C802000000000408D801000000000408012440000200110A0",
INIT_13 => X"000000000004680003A0040000000010280003800800000000102800000B0000",
INIT_14 => X"000005C0002000000000000620000158000010000000000010A0000B00000200",
INIT_15 => X"C30146200400104002602600400000000294004000000004000000000010001A",
INIT_16 => X"0080200000008020000000802000000080080000004090014134DA101288C6DB",
INIT_17 => X"0802000000000401806010040180601004018060100000802000000080200000",
INIT_18 => X"8060180601004010040080200802000000000000802008020000000000008020",
INIT_19 => X"C0A28A063807E0500014063450404882846FFE000003FFC00000010040100401",
INIT_1A => X"AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA28A28A28A28A2934C8D0CCD145144",
INIT_1B => X"68341A0D068341A0D068341A0D068341A0D068351A8D46A351A8D46A351AAAAA",
INIT_1C => X"FFFFFFFFFFFFFFFC0000000000000000000000001FE32068341A0D068341A0D0",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"408102040810207FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"800AA00000000000000000000000000000000000000000000040810204081020",
INIT_28 => X"168B55557BEAB4500554200000557FE10FFFBEAA10007FD7410FFAA97555082A",
INIT_29 => X"55574105D2A800AA00043FEBA5D7FEAA00007BE8AAAAA843DF55FFAA955EFA2D",
INIT_2A => X"57BC00AAA2FFEAAAAAA8415555087BFFF55A2AA800BAFFAE9555508002AA0000",
INIT_2B => X"A2AA955EF005568A00087BE8BFFA2D17DE1000517FE10AAAAA8AAA002E975455",
INIT_2C => X"FAA8417410A2D140000F7FBC2010A2D157400AAAE974AAAAAA974BA08002AB55",
INIT_2D => X"EFA2AABDEAA087BEAAAAA2FBD54BA080002145552ABFEAA007FC21EF007FD75F",
INIT_2E => X"00055042AB45F7FFD741000042AA10AAAABFF5508003FF55F7D568A00552EA8B",
INIT_2F => X"5400F7A49057D0824850B8000000000000000000000000000000000000000000",
INIT_30 => X"3AF55F7A0925D7AADB6FB7D5D7FEAB7808554203A145178E00FFFBE8A101475D",
INIT_31 => X"A9557D080038AAA145157428492E8008200043FE925571EFA380871C7028A28E",
INIT_32 => X"AEA8A9200249056D4175C5092AAF5FDA38BE8E1557D1475FAF45BEAA800AAFFA",
INIT_33 => X"AA4954281C0E2FB55B6A0925D7085F6AA10087FEABD7AAD57AEBA08517DE00AA",
INIT_34 => X"007FC51C7007BD55D7BE80004AAFEDB42028EBFBC2028BED152438AAA092492A",
INIT_35 => X"AF7DF6AA00412EAABFFAA803DEBA0875EDA80BEF1C743840040017D5520B8EAA",
INIT_36 => X"0000000000000000000041002FB55FFF5D0438140E2FA38B6AEBFF6DBE84AAEB",
INIT_37 => X"A00FFFFEAA105D5155410FF84021EF0800154B20000000000000000000000000",
INIT_38 => X"DEBA0851574B2AAAEAAB55F78400145AAFFFFFEF5D7FEABFF0051400A25D5568",
INIT_39 => X"68B55F7AA800BAF7AA955EF00042AAA25555410BA082E8201000043FE005D517",
INIT_3A => X"568AA200557DE00AAAAAAA000804001FF005575408AA557FEB2FFAE975EF5551",
INIT_3B => X"D1550AAAA8002010F2AC154B25F2ABFF55F7800015F087FEAA00007FEAB55FAD",
INIT_3C => X"800021EF55042AAAA007FD5555087BD6145FAAC000A2A6FBC00BAAAFBC00BAF7",
INIT_3D => X"F7AEBDFF779A82AA43F7FBE8A00082EA8BFFAA843FEBA08517DE00F3F9574B30",
INIT_3E => X"000000000000000000000000000000000000008003FF55F7D5420BA5D2ABFEAA",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(4),        -- Port A data input
DOA(0)   => data_read_a_lo(4),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(4),        -- Port B data input
DOB(0)   => data_read_b_lo(4),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_5_16 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50DF4A0791B3FCB694379283C81FD996A091832102004A336A20E03C040C002",
INIT_01 => X"805FBDC69830A84D5C6A60000C34C26841280A00084000C8C212892EEAD53235",
INIT_02 => X"3B2026B578918E640A4F01CF8011FF0002080000082CA9998276DF7772C7C80D",
INIT_03 => X"37134108420D700084205702A4008A1D9100002171C0E0051554D93A11F5D140",
INIT_04 => X"8A41A0FC03A56DA000425A819410E3816C086198A388B702A8CA1210844A0C4C",
INIT_05 => X"B1808A062E8BC835F5E84532D708238A282F00A9291224800A2861490343082C",
INIT_06 => X"903FB8483A90581859050424100940825C6184401CDC451B860A6507160C4100",
INIT_07 => X"D26F068BCC96CDF8918E640E96D1A3469D6300E2FFEA27F8E4D23248130E259C",
INIT_08 => X"0BFA82E568442B2A082C0A7E3014250D49DA37A2420619000002AFF48D1222E5",
INIT_09 => X"3F005001E40969289429360416DCD1C46083030604B1CA20C03DF83B0A2C60A5",
INIT_0A => X"14613C71005A10492B888120288F480D58858449026145B3830F449449062B4F",
INIT_0B => X"11AC04934AC648BFD727C031E64170A137D5AA5C3E4B0F8A3C58C34C002290E3",
INIT_0C => X"CA29C6CC50384B6AC6AC86AB31AACA6AB39AAC86AB39AACA6AB3055643559C31",
INIT_0D => X"C673E33CF28F38603855401985228A0614BD30A0A2819852011E5AC2B87F9182",
INIT_0E => X"FF87C002F87A803E460B2516510CA594FF0044FFA4B08BAC4BB2CD0F09CF84E3",
INIT_0F => X"0DFF0F8005F0F5100DFFF5E15D06101C55EB29F1E00BE53FE1F000BE1E802F94",
INIT_10 => X"F12F0380231F17D78FC029FFF58D9A70380230F2FE0017C37FC3E0017C3D005F",
INIT_11 => X"FC7F023C0CA700125C0F8F7E43F1F001BFFE7C69E01804E1E7CCF8FC003FF5F1",
INIT_12 => X"023E00017C1FC1A4BFD82C3081C5BD27BFE30C3081C5BD00C02365D645CEEF5B",
INIT_13 => X"61E0042787F181E9C1EFD8CB8120C5AF41E9C18FD60F0C20666F41E9F009FFFD",
INIT_14 => X"7A7C077FFF404F80005F07F187A7D14BFFC96111C048278DEB074F9930FF9D80",
INIT_15 => X"C064014B8B652E2B3120C81284641D3E8DBF7D636FE860190700132C1F0EFB80",
INIT_16 => X"38CE1384E3384E338CE138CE1384E33C4E3ECE32E128882551349A1CBAA44103",
INIT_17 => X"84E3384E3384E3384E338CE138CE1384E3384E338CE138CE1384E3384E338CE1",
INIT_18 => X"CE138CE138CE138CE1384E3384E3384E3384E338CE138CE138CE138CE1384E33",
INIT_19 => X"F5E5BB4E7F7B9DB7FF3A1B6DB7E8410A8C000000000000000000384E3384E338",
INIT_1A => X"BEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEF9F7CFDFDDCF3CF3D",
INIT_1B => X"BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEFBEF",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000001711C7BBDDEEF77BBDDEEF77",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"FDFFF00000000000000000000000000000000000000000000080000000000000",
INIT_28 => X"FD7410FFAA97410082A800AAAAAE955450055421FFFFFBC0010AAD5574BA557F",
INIT_29 => X"7FD74000055574BA5D7FD7555A2D5575EF55517FF5500557FE10FFFBEAA10007",
INIT_2A => X"0002AABA5D2ABFFFFAA843DF55FFAA955EFA2D168B55557BEAB5500554200000",
INIT_2B => X"5D2A800AA00043FEBA5D7FEAA00007BC00AAAAAEBDF45A28428B45FFD168BFF0",
INIT_2C => X"5080028A00A2FFFDE00F7D57FEBAFF80174BAAAD1555EF555555555005557410",
INIT_2D => X"BA5D2E821FFA2D5554BA557BD75FFAA8415555087BFFF55A2AA800BAFFAE9555",
INIT_2E => X"00000517FE10AAAAA8AAA002E97545557BC00AAA2FFEAAAA082A97545F7D5420",
INIT_2F => X"7010BEDF524AA5571FDFEF000000000000000000000000000000000000000000",
INIT_30 => X"78E00EBFBE8A101475D5400F7A49043D0824850B8A2AE9756D145B401FFFFFFC",
INIT_31 => X"FEAB7D0855420BA1471D74380851524BA5571D757DB6D5525EF555178F6D1451",
INIT_32 => X"8A28B6DEBDF6DBEF1C0A28AAA5524BFFFFA28E3AF55F7A0925D7AADB6FB7D5D7",
INIT_33 => X"5555057D145152428492E8008200043FE925571EFA380871C7028B6AEBDF45B6",
INIT_34 => X"BEAA800AAFFAA9557D080038AAAA2FBF8E10EBD578EAAFF8415482BED1555EF5",
INIT_35 => X"81C209256DFFDF420BA552A821FFB6DF574A85575C55EFBE8E1557D1475FAF45",
INIT_36 => X"0000000000000000000008517DE00AAAEA8A9200249056D4175C50920875FDA3",
INIT_37 => X"5FF5D7BC21EFF7FBD7400F7FBC00BA55557DFF70000000000000000000000000",
INIT_38 => X"01FF5D5568BE7555568A00AAFFEAA105D5155410FF84020AA0800154B2AAAA97",
INIT_39 => X"00145AAFFFFFEF5D7FEABFF0051400A25551554BA0051400BA5551575EFF7D14",
INIT_3A => X"1574B2FFAABFF45FFAAAABFFAAFFFDFFF552EA8AAA55043DFF7AAAEAAB55F784",
INIT_3B => X"8002410FFD5575EF5555421E75555400BA082E8201000043FE005D517DEBA085",
INIT_3C => X"FAE975EF555168B55F7AA800BAF7AA955EF00002AAA2A2FBE8A00A2D16AAAAFF",
INIT_3D => X"0055554088A557FEB25D00021FFFFFFC00BA552A821EFFFFFD74BA5D51575F7F",
INIT_3E => X"000000000000000000000000000000000000000557DE00AAAAAAA000804001FF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(5),        -- Port A data input
DOA(0)   => data_read_a_lo(5),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(5),        -- Port B data input
DOB(0)   => data_read_b_lo(5),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_6_16 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10800B0061A01002840002C03002818000402322520070B313301C4389B2082",
INIT_01 => X"250041CA3839684D18A160000C52426841000000090800090210080008110200",
INIT_02 => X"0020042080010000044654C0000C008010000000001020900200200002620814",
INIT_03 => X"060881021088200021080200E4000A0891000020610111500104C00000F14400",
INIT_04 => X"0880000100000002000052288144004281C050400100280000C8100000080001",
INIT_05 => X"928080840001100A08009000280201000850E022401400002028214043410820",
INIT_06 => X"10100518090012122100C808049310002040000410A0001400000200120840D2",
INIT_07 => X"000100800004400001000000860408108C22000A502010074120044800040001",
INIT_08 => X"50000040D0C4E2088003FD01C01004044058082004000000000121F020408244",
INIT_09 => X"00BF17E9001205A5204911F814444080400100020000D200DFD16400C2A40AA0",
INIT_0A => X"04611C17849000022862A1596C8B5DF04834948900000100220C244840000880",
INIT_0B => X"03AD0413424E4044D665C070C22602291504400D084915020448114080201000",
INIT_0C => X"5E08864011088B22D22C008B0022C408B1022C208B0822C608B1111600458010",
INIT_0D => X"4251A12CD28A300429688001000800000020280204001000A00804309A002182",
INIT_0E => X"0000000280402400420800000000006200FC10002442042429324294014E8CA7",
INIT_0F => X"A40000000500800840000800000000000002280018001480000000A010100052",
INIT_10 => X"00000000000004C2003000010240000000000000680800290000000140202000",
INIT_11 => X"2000C0000000000000000442000001080001000000000000010C000280001804",
INIT_12 => X"08000000000801C300A010000000156000902000000015101200002800000000",
INIT_13 => X"000000000101800038002408000000094000386028040000000940000ED40000",
INIT_14 => X"0003B000002000000000020180002A24005010000000000023000060C7000A40",
INIT_15 => X"3F0280090321000040A410C28108000160008094000810040000000000002300",
INIT_16 => X"284A5284A728CA5284A528CA728CA52C4A5A0A32A300940101349A0408240818",
INIT_17 => X"9CA1294A329CA5284A728CA7284A5284A728CA5284A528CA728CA5284A728CA7",
INIT_18 => X"CA3294A129CA3294A129CA1294A329CA1294A3294A129CA3294A129CA3294A32",
INIT_19 => X"F5F78BCE7F8FF0F4FA955F7CF7F40A80145D55555556AAAAAAAAA94A329CA129",
INIT_1A => X"8E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E39B6CEDECDDF7DF7D",
INIT_1B => X"F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE38E3",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000001A1A33F9FCFE7F3F9FCFE7F3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"555FF00000000000000000000000000000000000000000000080000000000000",
INIT_28 => X"BC0010AAD5574BA557FFDFFF087BFDF45F7AA974AAAAAA97555F784174BAF7D5",
INIT_29 => X"515555508043FE00F7AA97555A2FBD7410AA8428AAAAAAE955450055421FFFFF",
INIT_2A => X"7D1575EFFFAA9555500557FE10FFFBEAA10007FD7410FFAA97400082A800AA08",
INIT_2B => X"0055574BA5D7FD7555A2D5575EF55517FF55A2AA97400552AAAB45082E80155F",
INIT_2C => X"500554200000003DE10FFD5401FFF7AAA8A10082EAAB45A2FFC2000007FD7400",
INIT_2D => X"10AA803FE105D516AABAFF843FFFFAA843DF55FFAA955EFA2D168B55557BEAB5",
INIT_2E => X"000AAAEBDF45A28428B45FFD168BFF00002AABA5D2ABFFFF087BD5545007BFDE",
INIT_2F => X"256DEB84104BAFFD1525FF000000000000000000000000000000000000000000",
INIT_30 => X"9756D145B401FFFFFFC7010BEDF524AA5571FDFEF1C7BFFF55FFA095482B6A49",
INIT_31 => X"4904380824850381C5B5057D1C003DE28F7A49057DAAF5D2428A2842AAAAA2AE",
INIT_32 => X"2AAFB451C2A8017DE3DF525FFFFA49756D145178E00EBFBE8A101475D5400F7A",
INIT_33 => X"2F1C50381471D74380851524BA5571D757DB6D5525EF555178F6DAAA49542841",
INIT_34 => X"AADB6FB7D5D7FEAB7D0855420BA1C0E3FE00E3DB471EFE3AAAAA00082EA8B6DA",
INIT_35 => X"F1C7BD057D1C71FFE10A28038E1049516AAB8FF8428FEFA28E3AF55F7A0925D7",
INIT_36 => X"00000000000000000000B6AEBDF45B68A28B6DEBDF6DBEF1C0A28AAA5524BFFF",
INIT_37 => X"F55F78017400F780001FFAA84000AAFFD1401E70000000000000000000000000",
INIT_38 => X"20BAAA8428AA2AAAA975FF5D7BC21EFF7FBD7400F7FBC00BA55557DFF7557BFD",
INIT_39 => X"EAA105D5155410FF84020AA0800154B2557FC01EF55043FEAAFF80021EFA2D14",
INIT_3A => X"568BE7AA80174AA082ABDF555D2A821EFAAFBC01FFF780155F7555568A00AAFF",
INIT_3B => X"AEA8A10082EA8BEFAAD5554B25551554BA0051400BA5551575EFF7D1401FF5D5",
INIT_3C => X"AAEAAB55F78400145AAFFFFFEF5D7FEABFF0051400A25D2EBFE10AAFFD55EFA2",
INIT_3D => X"552EA8AAA55043DFF7557BC01EF55557DE00AA842AA0000516AABAFF8428BE7A",
INIT_3E => X"0000000000000000000000000000000000000FFAABFF45FFAAAABFFAAFFFDFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(6),        -- Port A data input
DOA(0)   => data_read_a_lo(6),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(6),        -- Port B data input
DOB(0)   => data_read_b_lo(6),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_7_16 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10844B00482258A2842112C02450418800002300500030B313300C418992002",
INIT_01 => X"000009CA3839684D1CA0E0000E51424840000000080000080200080008510204",
INIT_02 => X"0120042086010000044600C00008000004100000000260900200000002402004",
INIT_03 => X"8628A10000082400000002408400080011000000610008000208C00000E14400",
INIT_04 => X"0911800100A000000000524084000040000050001140200100C8100000080102",
INIT_05 => X"0300812401011000000000002000114008008060441000000020024093000000",
INIT_06 => X"9190431C0D4010100000880804010010800000041080081000000200010424B2",
INIT_07 => X"000100AA0004408601000004860000008C02000A103010006928040800062481",
INIT_08 => X"84000048D484C20888000A0002120484C048007004000000000021F000000244",
INIT_09 => X"00A06009881201A520491004106C48A04040002400A15A208001650004001020",
INIT_0A => X"C99E1060201002044809C1040140A001004808810000459033189C0A400118A0",
INIT_0B => X"102000024040484050050041648A0041140C500B08821054C000264120000400",
INIT_0C => X"0404A083260E0832132011880462011880462051881462051881D31018C40620",
INIT_0D => X"0001000080001000813094801A8F80F00A600B52602801A88848011118003700",
INIT_0E => X"000003C007C002808228010410082042C000C000000004001002000400040002",
INIT_0F => X"A4000007800F80C840000800009864038A1200081C0014800000F001F0200052",
INIT_10 => X"00002C0E00E0E4004038000102400002C0E00E0D20100029000001E003E04000",
INIT_11 => X"2000C04031100E0403D0700300080908000100000661801E1900040380001804",
INIT_12 => X"0840878083E8003780A01043203A101780902043203A10082410082880000000",
INIT_13 => X"0601E0187900181035E0240806483248181035E0280410C8198818100DDD0000",
INIT_14 => X"0403774000201021E020FA006040376C00501022131210722060806D47000A40",
INIT_15 => X"00928A0002000110888600C032128201519480D40009902430160403E0E00506",
INIT_16 => X"01000000020080601802000000000405000A0020020081014134928820480010",
INIT_17 => X"0802018040000000006018020080200804010000000000806018020080000004",
INIT_18 => X"0000000001806008020000001006008020080001004008020080201004000020",
INIT_19 => X"0000000000000000000000000000400A004618618618C30C30C3000020180600",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000000B0840000000000000000000",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"1555500000000000000000000000000000000000000000000080000000000000",
INIT_28 => X"A97555F784174BAF7D5555FFF780155EFAAAEA8ABAAAFBFDE0055556AA005D04",
INIT_29 => X"55555EFAAFFFDFEFAAAAAAB455D556AA00FFAE95555087BFDF45F7AA974AAAAA",
INIT_2A => X"02EAAAAA082EA8A00AAAE955450055421FFFFFBC0010AAD5574BA557FFDFFF55",
INIT_2B => X"08043FE00F7AA97555A2FBD7410AA8428AAA557BFDFFF55003DFFFF7FBEAA000",
INIT_2C => X"0082A800AAF7AE975FFA28000010552EBDE00007BEAAAAA2D140000085155555",
INIT_2D => X"45087FEAB455D516AB55557BD55FF00557FE10FFFBEAA10007FD7410FFAA9740",
INIT_2E => X"000A2AA97400552AAAB45082E80155F7D1575EFFFAA955555D51574AAAAFFD55",
INIT_2F => X"AE105D556AA10410E17555000000000000000000000000000000000000000000",
INIT_30 => X"FFF55FFA095482B6A49256DEB84104BAFFD1525FFFF8E175C7A2AAAAA82A2F1F",
INIT_31 => X"F524AA5571FDFEF415B575D7AAF1FFFD7AAAAAFB7D495F6AA10E3AE905551C7B",
INIT_32 => X"003AFEFEBFBEAA001C2EA8A821C2EAAA00A2AE9756D145B401FFFFFFC7010BED",
INIT_33 => X"EDB470101C5B5057D1C003DE28F7A49057DAAF5D2428A2842AAAA497BFAFFF49",
INIT_34 => X"1475D5400F7A490438082485038F7A4905C7A28A070384120BDE100075EAA82B",
INIT_35 => X"D495150492BEF1D2555087BE8B7D555F6AB57417BC05D7145178E00EBFBE8A10",
INIT_36 => X"00000000000000000000AAA495428412AAFB451C2A8017DE3DF525FFFFA49756",
INIT_37 => X"555A2AEA8A10AAD568A00555168A10002E9754D0000000000000000000000000",
INIT_38 => X"8A10AAAE8215D557BFDF55F78017400F780001FFAA84000AAFFD1401E7FFAA97",
INIT_39 => X"C21EFF7FBD7400F7FBC00BA55557DFF7007BD5555AAD57DF55AAAEBDFEF007BE",
INIT_3A => X"428AA2007FE8BFF080028BFFAAFFEAA105D2EAAA005D2AAAA18AAAA975FF5D7B",
INIT_3B => X"043DE0000516AA10F7FBD7408557FC01EF55043FEAAFF80021EFA2D1420BAAA8",
INIT_3C => X"55568A00AAFFEAA105D5155410FF84020AA0800154B2FF8402145A2AA954AA00",
INIT_3D => X"AAFBC01FFF780155F7005140000FFD140145007FE8BEF557BEAB55087FC215D5",
INIT_3E => X"0000000000000000000000000000000000000AA80174AA082ABDF555D2A821EF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(7),        -- Port A data input
DOA(0)   => data_read_a_lo(7),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(7),        -- Port B data input
DOB(0)   => data_read_b_lo(7),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_8_16 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00000648E2840112C00000418000002700500030B3132000400812082",
INIT_01 => X"100008480009004C04A100000252024840000000180800080200010040110204",
INIT_02 => X"0020042000490000004600804008000005100000000024900200000002400004",
INIT_03 => X"0A0C33400008082400000080A4004B0891000020610112000040C00000E5C000",
INIT_04 => X"18800001000000000000512080000040800150400824280110C8100000120200",
INIT_05 => X"908084A10100100200004080280008240810802206940000012C214451610800",
INIT_06 => X"81B000080860109021400008040000202048020414A0021400040200322824C1",
INIT_07 => X"000000080004408049000004860000008402001A50208000630C040800062483",
INIT_08 => X"440000428644212280800A00021004044048002124000000000021F000000244",
INIT_09 => X"00004009001001010008100414644410400102228000D20080114502006409A2",
INIT_0A => X"000051312000042200294429148A4801C80C8C81000045907118040340020832",
INIT_0B => X"4020000240404140004D0544C4AA0001150410090302500011C813428A000400",
INIT_0C => X"46501090008820240240409000240009000240009000240009000120204808A5",
INIT_0D => X"42D1A168D09A301468402480004780F00140080860280004085904309A002196",
INIT_0E => X"00783FC00044340242280000000000020000C0000442106419120004034685A3",
INIT_0F => X"8000F07F800088A80000081EA2F9EC0000064004081010001E0FF00011104040",
INIT_10 => X"0ED0FC7E00000422201080000202658FC7E0000021882020003C1FE000222080",
INIT_11 => X"018059C3F350FE0C00000002A0040500000103961FE780000110010090000800",
INIT_12 => X"FD41FF80000830200021C1CF600012200010D1CF600012121600100810000004",
INIT_13 => X"9E1FE000010A1802100004343ED8000898021000087073D80008980200800002",
INIT_14 => X"0080200000BEB07FE00002086008020000209AEE3F300000246020200000620B",
INIT_15 => X"0088881903210000440610C8000A808040000208901786E4F0FE0C0000000166",
INIT_16 => X"685A1685A769DA368DA368DA769DA36CDA121A11A141800011309284002C0810",
INIT_17 => X"95A5685A1685A5695A368DA368DA769DA368DA368DA7695A1685A1685A5695A1",
INIT_18 => X"5A1695A568DA368DA369DA768DA1685A1695A5685A168DA369DA768DA368DA16",
INIT_19 => X"A4028A0A543EBC57A10A1E75D64108080468618618630C30C30C69DA5685A168",
INIT_1A => X"9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7BF3CCD8DF5B2DB2C",
INIT_1B => X"F87D3E1F4F87D3E1F4F87D3E1F4F87D3E1F4F87C3E1F0F87C3E1F0F87C3E79E7",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000006A6D4F87D3E1F4F87D3E1F4",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"155FF00000000000000000000000000000000000000000000080000000000000",
INIT_28 => X"BFDE0055556AA005D0415555080000000087BEAA10F7803DE00FFAEBFFFF0800",
INIT_29 => X"2AA8AAA557FC0010F780154105D7FC2145005155555F780155EFAAAEA8ABAAAF",
INIT_2A => X"7FFFFF55AA80155FF087BFDF45F7AA974AAAAAA97555F784174BAF7D5555FF55",
INIT_2B => X"AAFFFDFEFAAAAAAB455D556AA00FFAE95555AAFFE8A00552EBFE00F7D17FF45F",
INIT_2C => X"A557FFDFFF5504000AAAAAAA8B55F7D140010552E821EFAAAABDF555555555EF",
INIT_2D => X"55AA8028A00A2D57FF45557BE8A00AAAE955450055421FFFFFBC0010AAD5574B",
INIT_2E => X"000557BFDFFF55003DFFFF7FBEAA00002EAAAAA082EA8A00002AA8A10F784021",
INIT_2F => X"FE10F7AEBAFFF080A175D7000000000000000000000000000000000000000000",
INIT_30 => X"175C7A2AAAAA82A2F1FAE105D556AA10410E17555080E000280071E8A00EB8E3",
INIT_31 => X"4104BAFFD1525FF492EA8AAA5571C2000FF8A17400557FC015514555757DFF8E",
INIT_32 => X"2ABDE10EBDF7AF6DE3FFF8F7DB68A105D71C7BFFF55FFA095482B6A49256DEB8",
INIT_33 => X"AA0BDF6D415B575D7AAF1FFFD7AAAAAFB7D495F6AA10E3AE90555A2FBE8A3849",
INIT_34 => X"FFFFC7010BEDF524AA5571FDFEF550E00082B6A0AFB55F7D1420104124821D7A",
INIT_35 => X"01C2EA8A00F7800017DA2842FA00B6D578F6D557FFDA00A2AE9756D145B401FF",
INIT_36 => X"00000000000000000000497BFAFFF49003AFEFEBFBEAA001C2EA8A821C2EAAA0",
INIT_37 => X"0BA08556AA00AAAABFE00F7AEAABEF082E955450000000000000000000000000",
INIT_38 => X"21555D51575EFFFAA97555A2AEA8A10AAD568A00555168A10002E9754D082E82",
INIT_39 => X"17400F780001FFAA84000AAFFD1401E7082EAAABA5D5140010F7AE974105D7BC",
INIT_3A => X"E8215DA2FFE8ABA082ABFE00AAFBEABFFAAFBEABFFF7AA80145557BFDF55F780",
INIT_3B => X"D540000000402145AA843FFFF007BD5555AAD57DF55AAAEBDFEF007BE8A10AAA",
INIT_3C => X"AAA975FF5D7BC21EFF7FBD7400F7FBC00BA55557DFF75D2E82010F7843DF45FF",
INIT_3D => X"5D2EAAA005D2AAAA185D2AAAA10F780021FFA2803DE10FFD16ABFF5D7BFDE10A",
INIT_3E => X"0000000000000000000000000000000000000007FE8BFF080028BFFAAFFEAA10",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(8),        -- Port A data input
DOA(0)   => data_read_a_lo(8),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(8),        -- Port B data input
DOB(0)   => data_read_b_lo(8),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_9_16 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00018248A2840112C00002C18000002300500030B3132000400812006",
INIT_01 => X"400008000000004C0020000000100248413C0A61590001D90213C10008110204",
INIT_02 => X"01A0042080010000054600C04008000004100000001020900200200002420804",
INIT_03 => X"024003400008012400000010E4004B0891000020610310000144C00000F5C000",
INIT_04 => X"1801800100E000000000510084000040010050020810200000C8900000320200",
INIT_05 => X"918004311104100000000000200008100800002000100000002C234415610820",
INIT_06 => X"81B00008080010100000980804000008800042041080001000100200322C2481",
INIT_07 => X"0000811800044080010000058600000086020002502080006000040800062C80",
INIT_08 => X"0000004001D4618008800A00061004044048002004000000000061F000000244",
INIT_09 => X"000040090802009420409004104444084001022400214A2080014400026401A2",
INIT_0A => X"04000071200000A003CA294140200800C80C8C8100004590111C040040120800",
INIT_0B => X"12210002404848502847040164880021150400080222000200C8034200000000",
INIT_0C => X"4610088010080421021040841021000841021000841021000841010800420820",
INIT_0D => X"42D0A16C529A321068500484000500D10042080040284000084900001A002196",
INIT_0E => X"00000002804000004228010410082002C000C0002400046419120410034285A1",
INIT_0F => X"A00000000500800800000800000000000002290008001080000000A010100042",
INIT_10 => X"00000000000004C2001000000240000000000000680800280000000140202000",
INIT_11 => X"0000C0000000000000000442020001000001000000000000010C800080000804",
INIT_12 => X"08000000000801A7802010000000152780102000000015000600000800000000",
INIT_13 => X"000000000101900011E0240000000009500011E0280000000009500004DD0000",
INIT_14 => X"000137400020000000000201C000136C00101000000000002340002947000240",
INIT_15 => X"0080881901210000000600C280028000419480D4000010040000000000002304",
INIT_16 => X"68DA368DA1685A1685A1685A1685A16C5A121A13A141950051309284A82C0010",
INIT_17 => X"85A1685A1685A1685A368DA368DA368DA368DA368DA368DA368DA368DA368DA3",
INIT_18 => X"5A1685A168DA368DA368DA368DA368DA368DA368DA3685A1685A1685A1685A16",
INIT_19 => X"0157344CCCF48DE68A895C38E2540A8010100000000000000000685A1685A168",
INIT_1A => X"14514514514514514514514514514514514D34D34D34D34D28E1004039248209",
INIT_1B => X"D268341A4D268341A0D069349A0D069349A0D068341A0D068341A0D068345145",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000014D490D069349A0D068341A4",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"EAABA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"03DE00FFAEBFFFF0800155FFAAFBE8B45002A974AAAA803DFFFAA843DF45FFFF",
INIT_29 => X"7BFDE00A2FBD7400F7FBFDFFFA2AEBDE00AAFBEAABA080000000087BEAA10F78",
INIT_2A => X"055401FFF7AEAAA10F780155EFAAAEA8ABAAAFBFDE0055556AA005D041555508",
INIT_2B => X"557FC0010F780154105D7FC2145005155555557BE8BEF007FFDEAAAAD1555EF0",
INIT_2C => X"AF7D5555FFF780154AA5D2AA8A10F7AA974AA082E80010A2AAAAA10552AA8AAA",
INIT_2D => X"BAF7D17FEBAA2AEBDF45002EAAABA087BFDF45F7AA974AAAAAA97555F784174B",
INIT_2E => X"000AAFFE8A00552EBFE00F7D17FF45F7FFFFF55AA80155FF080400145FFFBEAA",
INIT_2F => X"8FC7BE8A3DF7DF7F5E8A92000000000000000000000000000000000000000000",
INIT_30 => X"000280071E8A00EB8E3FE10F7AEBAFFF080A175D7BEF1E8B6D002090482B68E3",
INIT_31 => X"56AA10410E175550871FFE00A2FBD0400FFF5FDFC7B6A0BDE38B6F5E8A92080E",
INIT_32 => X"7BFAE82A2DB555C71C5B451D7FFAAA8A38FF8E175C7A2AAAAA82A2F1FAE105D5",
INIT_33 => X"2AEADA38492EA8AAA5571C2000FF8A17400557FC015514555757D5D71E8BEF14",
INIT_34 => X"B6A49256DEB84104BAFFD1525FFFF84174BA5D20AAA00E3AA904BA142A87010A",
INIT_35 => X"7000400155FFFBEDA82FFD57DEBAAAA0BFF7D0024ADA921C7BFFF55FFA095482",
INIT_36 => X"00000000000000000000A2FBE8A38492ABDE10EBDF7AF6DE3FFF8F7DB68A105D",
INIT_37 => X"BEF080402000F7AAA8B55FFAABDFEFF7D16AA000000000000000000000000000",
INIT_38 => X"FEAAFFD16AA00082E820BA08556AA00AAAABFE00F7AEAABEF082E95545F7D568",
INIT_39 => X"A8A10AAD568A00555168A10002E9754D00517DE00A2FFC2000F7D17FF55FF803",
INIT_3A => X"1575EF555568BEF5D7FE8A10AAFFD55555D7FD5555FFAAA8AAAFFAA97555A2AE",
INIT_3B => X"AE800AA552A97400A2AEBDEAA082EAAABA5D5140010F7AE974105D7BC21555D5",
INIT_3C => X"57BFDF55F78017400F780001FFAA84000AAFFD1401E7FF80174AA5D0028A00AA",
INIT_3D => X"AAFBEABFFF7AA80145080002145F7FBFFE00FFD17FEAAA2803DFEF08043FE005",
INIT_3E => X"0000000000000000000000000000000000000A2FFE8ABA082ABFE00AAFBEABFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(9),        -- Port A data input
DOA(0)   => data_read_a_lo(9),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(9),        -- Port B data input
DOB(0)   => data_read_b_lo(9),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_10_16 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00018248A2840112C00002C18000202300500030B3132000400992006",
INIT_01 => X"254008000000004C002000000010026840000000080000080200010008110204",
INIT_02 => X"0020042000010000004455800008000004100000000000900200000002400004",
INIT_03 => X"020001021089000021081000C400090011000000610001540104C00000F14400",
INIT_04 => X"0811800101A00002000050088554004200C840000000200080C8100000000001",
INIT_05 => X"030080001000100800009400200000000840E020201000000024024001200020",
INIT_06 => X"81B00008080012120004CC080492500280208004148000100000020020042493",
INIT_07 => X"0000000800044080010000048404081085020002502000006000040800062480",
INIT_08 => X"100202400084410808000A00021004044048000004000000000021F020408264",
INIT_09 => X"010040090002008420401004144440004040022484214A2080110108C2C00320",
INIT_0A => X"04004166A48A0001080000000000080080181881000045901118044040020800",
INIT_0B => X"1201000200484910000F0105602622291404020902005002018002400A022000",
INIT_0C => X"0440001011808020120004801120044800120004801120044800110002400884",
INIT_0D => X"008000440210100041308480800F82F00040180260A808008848000018002104",
INIT_0E => X"000000028040000002280104100820020000400020000440100204100A000100",
INIT_0F => X"040000000500800800000000000000000002280008000400000000A010100010",
INIT_10 => X"00000000000004C2001000010000000000000000680800010000000140202000",
INIT_11 => X"200000000000000000000442000001000000000000000000010C000080001000",
INIT_12 => X"00000000000801C0008000000000154000800000000015000410000800000000",
INIT_13 => X"0000000001019800180000080000000958001800000400000009580002800000",
INIT_14 => X"0000A0000000000000000201E0000A0000400000000000002360002080000800",
INIT_15 => X"0080881000000000000600C28102800060000000000800000000000000002306",
INIT_16 => X"401004010040100401004010040100441020D0030008840051309A90BA884010",
INIT_17 => X"0902409024090240900401004010040100401004010040100401004010040100",
INIT_18 => X"1004010040902409024090240902409024090240902409024090240902409024",
INIT_19 => X"F546890A940FE0D3971243555205428290100000000000000000401004010040",
INIT_1A => X"8A28A28A28A28A28A28A28A28A28A28A28A28A28A28A28A29554199854514514",
INIT_1B => X"2B95CAE532994CA6532995CAE572B94CA6532994CA6532994CA6532994CA28A2",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000002718E72B94CA6532994CA657",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"FDE1000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"03DFFFAA843DF45FFFFEAABA007FC2155F7D155545AA80001EFAAFBEAB45557F",
INIT_29 => X"042AB55FFD168B55AA8000010FFFBE8BFFF78402155AAFBE8B45002A974AAAA8",
INIT_2A => X"AD16AABA002ABDE10080000000087BEAA10F7803DE00FFAEBFFFF0800155FF00",
INIT_2B => X"A2FBD7400F7FBFDFFFA2AEBDE00AAFBEAABAA2FFD741055003DFEFF7AA801FFA",
INIT_2C => X"05D0415555007FD74105555555EFF7FBC0145F78028A00A2D142155087BFDE00",
INIT_2D => X"55AAD168ABA002A975FFF7AEBDEBAF780155EFAAAEA8ABAAAFBFDE0055556AA0",
INIT_2E => X"000557BE8BEF007FFDEAAAAD1555EF0055401FFF7AEAAA105D042ABFF5D556AB",
INIT_2F => X"71D7AAFBEFB455D71F8E00000000000000000000000000000000000000000000",
INIT_30 => X"E8B6D002090482B68E38FC7BE8A3DF7DF7F5E8A92007BC217DEBDB55555AA8E0",
INIT_31 => X"EBAFFF080A175D700042AB7DEBDB6DB55BE8E05000EBFFE8BC7E38E07145BEF1",
INIT_32 => X"0A3DFD7F7A4821D7A2D16FA82142EB8E00080E000280071E8A00EB8E3FE10F7A",
INIT_33 => X"ED1421450871FFE00A2FBD0400FFF5FDFC7B6A0BDE38B6F5E8A92B6FBD541049",
INIT_34 => X"A2F1FAE105D556AA10410E175550071D54104951555D7EBF5C5155E3842AA00B",
INIT_35 => X"8410E2ABD749516FB55BED16FA820820955EFE3AEBDEAAFF8E175C7A2AAAAA82",
INIT_36 => X"000000000000000000005D71E8BEF147BFAE82A2DB555C71C5B451D7FFAAA8A3",
INIT_37 => X"1EFA2FFD7545AAAE97555A2FBFDF455D556AA000000000000000000000000000",
INIT_38 => X"8B45AAAA95545F7D568BEF080402000F7AAA8B55FFAABDFEFF7D16AA00087FC0",
INIT_39 => X"6AA00AAAABFE00F7AEAABEF082E9554500042ABFFA2FFFFF45F7AE97400AAFFE",
INIT_3A => X"16AA00FFFBD5400082EBFF45F78400155A2D57FE00552EA8A00082E820BA0855",
INIT_3B => X"D557555A2802AA10FFD54214500517DE00A2FFC2000F7D17FF55FF803FEAAFFD",
INIT_3C => X"FAA97555A2AEA8A10AAD568A00555168A10002E9754D085155410085557555AA",
INIT_3D => X"5D7FD5555FFAAA8AAA002AAAB4508557DF55F7D17FE000804155FFAAAABDEAAF",
INIT_3E => X"0000000000000000000000000000000000000555568BEF5D7FE8A10AAFFD5555",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(10),        -- Port A data input
DOA(0)   => data_read_a_lo(10),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(10),        -- Port B data input
DOB(0)   => data_read_b_lo(10),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_11_16 : RAMB16_S1_S1
generic map (
INIT_00 => X"A101C4B05A0034CA2840712C2D001419000002300500030B31B20084EC992002",
INIT_01 => X"90000986B83028491800E0000C26426040000000080000088200080802512224",
INIT_02 => X"1A2004205E010640024D00800008000004100000040EC090820018003241A00C",
INIT_03 => X"28639100000C5C00000045C08400C8001100000061806A001618C03001E54400",
INIT_04 => X"1A800001000009A0804059A190000040400040008058220008C8100000120D4E",
INIT_05 => X"02000E81080250010000002022000058080400000E1200000020004401000004",
INIT_06 => X"819435143F20101010001008040800B8100102041088011100022200000024B2",
INIT_07 => X"90640D280884453E01064002944180008402001295BA100022E4340800062D82",
INIT_08 => X"400000093204802200280A0012160585C1D808D004000000000323F40C102244",
INIT_09 => X"380040098010001100009204107C5950400000220080C200800900020C006827",
INIT_0A => X"80007100004016EA080801010000080D00200081000045B0511D289940103399",
INIT_0B => X"002000024040410A000D0104408810C115D9C008050042400100D04E88000002",
INIT_0C => X"00655010009264201200C7B421ED0C7B421ED0C7B431ED087B43176843DA1085",
INIT_0D => X"0401020080400A10012494881A4F80F209500BB2602881A488485C1318002000",
INIT_0E => X"6619A540124814800228010410082022C00040002020090020220C9600040802",
INIT_0F => X"ACCC334A802491600C587949B6D0141B4CC600D5761B1599865A500490B86A56",
INIT_10 => X"BAC845542056A61686EC81E3A6CB68AA2C622C9A251C352B330CB4A0092170D8",
INIT_11 => X"BCCAD0B5A81536080CC6B21A21B1FC09CB0F1076D4A200B2AD4068F4101639B5",
INIT_12 => X"4D2CC281E31AA0103AB8D5514066380804B268A2E060901204112566F10AC418",
INIT_13 => X"D551443C47281002540B2C9AAAA8662A1152B202AE3554403028115AA88201A1",
INIT_14 => X"548A20A0492A2724A0621620402A020141F172FB182A32AB6845AB6200251BC9",
INIT_15 => X"00C00A000200074044E6801832728080D00A380B753952C4877E0104DDE4D124",
INIT_16 => X"0080200802008020080200802008020480080022020081010124988800400010",
INIT_17 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_18 => X"0000000000802008020080200802008020080200802008020080200802008020",
INIT_19 => X"55062608804180C0B10A42104201400204000000000000000000000000000000",
INIT_1A => X"00000000000000000000000000000000000820820820820801C4149470000000",
INIT_1B => X"0000000000000000040200000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000007E0F0000000000000100800",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"000AA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0001EFAAFBEAB45557FFDE10082ABDF5508557DF45002ABDFFFF7803DE10AA80",
INIT_29 => X"AEBFF45FFAEBFEAA002A801FFF7FFE8A10A28000000007FC2155F7D155545AA8",
INIT_2A => X"2AABFE10082ABFFEFAAFBE8B45002A974AAAA803DFFFAA843DF45FFFFEAABAA2",
INIT_2B => X"FFD168B55AA8000010FFFBE8BFFF78402155AAD155555A28428BFF002ABDE00A",
INIT_2C => X"F0800155FF00557FF45557FC2010002A80010A2842AAAA007BFFF4500042AB55",
INIT_2D => X"FF5D00154BAF7FBE8BEFFFD540000080000000087BEAA10F7803DE00FFAEBFFF",
INIT_2E => X"000A2FFD741055003DFEFF7AA801FFAAD16AABA002ABDE10A2D168A10A284021",
INIT_2F => X"DFC7F78E3FE28B684070AA000000000000000000000000000000000000000000",
INIT_30 => X"C217DEBDB55555AA8E071D7AAFBEFB455D71F8E00002EBDF6D005B78F7D142AB",
INIT_31 => X"A3DF7DF7F5E8A92BEAEBFF7DEBA0BDEAA1C2A801C7E3FFEFA10B68407038007B",
INIT_32 => X"8A28BFF082ABAE10B6AAB8E280820B8FEFBEF1E8B6D002090482B68E38FC7BE8",
INIT_33 => X"07FF8F7D00042AB7DEBDB6DB55BE8E05000EBFFE8BC7E38E07145B6D15756DA2",
INIT_34 => X"EB8E3FE10F7AEBAFFF080A175D708517DF7D497BC5028142A87000A28A2AA920",
INIT_35 => X"0B6DB6AA28A280001FF5D0A10482FFFFEFBC7E3DF42028080E000280071E8A00",
INIT_36 => X"00000000000000000000B6FBD5410490A3DFD7F7A4821D7A2D16FA82142EB8E0",
INIT_37 => X"FEF007BE8BFF5D2ABDF55F7AABDEAAF784154BA0000000000000000000000000",
INIT_38 => X"DE00FF84154BA087FC01EFA2FFD7545AAAE97555A2FBFDF455D556AA00082EBF",
INIT_39 => X"02000F7AAA8B55FFAABDFEFF7D16AA00FFAEBFFEFAA803DEBA5D2E82155A2FBF",
INIT_3A => X"A95545F7D5555FFAAAAA8BFF002AAAA00FFAAA8AAA080028BFFF7D568BEF0804",
INIT_3B => X"2E95400A2AEA8A00007FEABFF00042ABFFA2FFFFF45F7AE97400AAFFE8B45AAA",
INIT_3C => X"82E820BA08556AA00AAAABFE00F7AEAABEF082E9554508557DFFF007BD54BA5D",
INIT_3D => X"A2D57FE00552EA8A00FFFFE8AAAAA80001FF5D2E82000F7FFFFF45AAFFC20BA0",
INIT_3E => X"0000000000000000000000000000000000000FFFBD5400082EBFF45F78400155",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(11),        -- Port A data input
DOA(0)   => data_read_a_lo(11),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(11),        -- Port B data input
DOB(0)   => data_read_b_lo(11),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_12_16 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50080B01BC002006940202C0DE041196A83183000000023322287E0FC000006",
INIT_01 => X"75400D849830C84C5823E0000C17424840000000080000088200002802153231",
INIT_02 => X"18A026B43ED180040147558040090000061800000C06ED9802768F4472C52005",
INIT_03 => X"2A67E34A528D0524A52850528400C8001100000171C02B550618C91A10E55440",
INIT_04 => X"1BC0000100056C8280825DE98154004300C840800850240080CA921084520A07",
INIT_05 => X"02000F832000500C0000941024000852084060202E100001002000448100000C",
INIT_06 => X"819A1D1C3FE01A1A40045408049A50BA4020C6041090001200006200000000F2",
INIT_07 => X"C26A0719CC96CC6ED18A64019695A854870300FA3968B20068FC06080106249F",
INIT_08 => X"D002024B3E040800008C0A002610240D494A06F3460409000000E3F0AD5282E5",
INIT_09 => X"27A06009200040000400120412445D78400001000410420080218029CC807A27",
INIT_0A => X"18000006848A026F000000000000080000F010C100204593F11A6CDF48003BF8",
INIT_0B => X"000000820040402B28050400400432C9349DF21A31A00ACC0000F04F80020001",
INIT_0C => X"00357804611AE45D05D0833430CD0833420CD0C33420CD0833430668619A1000",
INIT_0D => X"0000000000000A74812DF00E87E80A079F9F90FA0280E87E800C7FF3B8002000",
INIT_0E => X"3B6B0E404D26160682082002000401EA0000C40000800A006002818808000000",
INIT_0F => X"A476D61C809A4DA84272592D6246FC1B17B541F97E1B348EDA93900B2B286C56",
INIT_10 => X"30C669E622DBC325CFD881A962454CFBE5403AB99594362B1DB52720165650D9",
INIT_11 => X"F8D2D39A3745261E4A95A110A3F855000E4B1D32BAB504BB7490FCFF912A3834",
INIT_12 => X"B90E9B018C7530200AB8F8BF41F9A22006B37DC8E1F9A21A70116D4C5080651C",
INIT_13 => X"118780319CCA08AB1001ACDF34B8F1C688AB1002AE3F7B807B6289F368828C4C",
INIT_14 => X"2AF020233376A5ECC016B1A827CDA21160F051DE610A34C50427E6E220323E4A",
INIT_15 => X"0077020000000439FDC05C5806781FAB46095A0B5199B0AC55521524F1864022",
INIT_16 => X"000000000000000000000000000000000026C000002884000130921092804010",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"8020080200000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0051B946088881360A95090CB054420290100000000000000000008020080200",
INIT_1A => X"041041041041041041041041041041041049249249249249200100002D451451",
INIT_1B => X"92C964B2592C964B2592C964B2592C964B2592C86432190C86432190C8641041",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000003800F592C964B2592C964B25",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"7DE1000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"ABDFFFF7803DE10AA80000AAAA843FE0008557DFFF0800020105D557FEAA0055",
INIT_29 => X"D5420000051555FFA2AA8200000557DFFFF7AA80000082ABDF5508557DF45002",
INIT_2A => X"82AA8AAAAAFFC00BA007FC2155F7D155545AA80001EFAAFBEAB45557FFDE10AA",
INIT_2B => X"FFAEBFEAA002A801FFF7FFE8A10A28000000A2D155410F7FFFFEBA08003FE000",
INIT_2C => X"5FFFFEAABA000028A105D2ABFE10A2AABFE1055516ABEF5D517DEAAA2AEBFF45",
INIT_2D => X"55002A820AA08557DFFFF7AA82155AAFBE8B45002A974AAAA803DFFFAA843DF4",
INIT_2E => X"000AAD155555A28428BFF002ABDE00A2AABFE10082ABFFEF0855420000004175",
INIT_2F => X"5010495B7AE921C517DE10000000000000000000000000000000000000000000",
INIT_30 => X"BDF6D005B78F7D142ABDFC7F78E3FE28B684070AABE803AE38145B78FD700000",
INIT_31 => X"BEFB455D71F8E00BED547038145B505FFB6A487000005F7AFD7F7A482038002E",
INIT_32 => X"F1FDE821C003FE001C2EAAAAAB6F5C2082007BC217DEBDB55555AA8E071D7AAF",
INIT_33 => X"D517DEAABEAEBFF7DEBA0BDEAA1C2A801C7E3FFEFA10B68407038B6D550428FF",
INIT_34 => X"B68E38FC7BE8A3DF7DF7F5E8A9200002FA285D20BDE28A2A4B8E10555B68BEF5",
INIT_35 => X"F085F47038140010555142082082005F7DFD7F7A482155BEF1E8B6D002090482",
INIT_36 => X"00000000000000000000B6D15756DA28A28BFF082ABAE10B6AAB8E280820B8FE",
INIT_37 => X"ABA5D7FEAB45080015410007FEAA0055517DE000000000000000000000000000",
INIT_38 => X"AB45F780020BA082EBFFEF007BE8BFF5D2ABDF55F7AABDEAAF784154BAF7802A",
INIT_39 => X"D7545AAAE97555A2FBFDF455D556AA00F7D1554BA5D7BC01FFFF8015410007FE",
INIT_3A => X"4154BAF7D1400BAFFD57FE005D043FE10552EAAAAAFFD140000087FC01EFA2FF",
INIT_3B => X"8428A105D7FEABEF55557DEBAFFAEBFFEFAA803DEBA5D2E82155A2FBFDE00FF8",
INIT_3C => X"7D568BEF080402000F7AAA8B55FFAABDFEFF7D16AA0008003FEBA55003DEBAA2",
INIT_3D => X"FFAAA8AAA080028BFF087BD54AA550402145550000010087FFFF45F78402145F",
INIT_3E => X"0000000000000000000000000000000000000F7D5555FFAAAAA8BFF002AAAA00",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(12),        -- Port A data input
DOA(0)   => data_read_a_lo(12),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(12),        -- Port B data input
DOB(0)   => data_read_b_lo(12),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_13_16 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10154A0441836CA2840512822007C18000E02700500030B31B300040081A042",
INIT_01 => X"00000804A000C04800020000000002404001000008220008A200100802110204",
INIT_02 => X"02200430000104000A4700804008000004100000000420918204D3033240400D",
INIT_03 => X"AA4003400008592400000590C40009141100000C6180C0000000C00001E14000",
INIT_04 => X"0800000102400120088054019000004160004190BAA0270000C8100000600206",
INIT_05 => X"21000012040610050040000227003AA0082400E94C1200000824424005220020",
INIT_06 => X"81963B180C001010580000080400000058000004109C00138000020024142581",
INIT_07 => X"002C8008000441600106400A9600010494020002B8AAA000EF003408000E2580",
INIT_08 => X"000000E48194408000A00A001210040441C80320040210000002ABF004102244",
INIT_09 => X"2A004009640040100400940412D4C4004000022000104200802D983000480120",
INIT_0A => X"8000202020401480000000000000080C90090881000145B0111A14004015080D",
INIT_0B => X"00000002004040AA08050400404040C11444000805200A402090024000008002",
INIT_0C => X"8410000A00280020020040800020040800020000801020000800010020400000",
INIT_0D => X"84A14250A055100050100490000500D00040080040290000084E4000B800610C",
INIT_0E => X"DCD13042BEDA36820228000000000000C000400081A08BC812A2092B02850942",
INIT_0F => X"89B9A260857DB400431969CA985D480949D32804A40AB137341C10B7D6A02EC0",
INIT_10 => X"E6ACA678001CE7D0296C213A460CA4271CA2168AEC1017606E6838216FAD4055",
INIT_11 => X"84AD4961C281B20213073C5FC0058008632D30D522CE80239DCC01AB013A4D20",
INIT_12 => X"2E6B13804A4B01D83461299900F6BD583A519104A0EEBD1A141010B2A4C8E116",
INIT_13 => X"89E5E40913419151EE0E94641828F72B5151EE0D184B321037AF5158BB02D085",
INIT_14 => X"562EC0B42162D68EE0073AE1C562EC13D521921A4170300B2B458B56B01C2280",
INIT_15 => X"00888A120240034000E6DC8285028014B82372011FC1E4F5E0A00929684EAF84",
INIT_16 => X"50942509425094250942509425094254940A1421420082020120908800480030",
INIT_17 => X"0942509425094250942509425094250942509425094250942509425094250942",
INIT_18 => X"9425094250942509425094250942509425094250942509425094250942509425",
INIT_19 => X"F7EFBBEEFF3F7DF7FF3E9F7DF7E2450228000000000000000000509425094250",
INIT_1A => X"BAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBF7DFDFDDD555555",
INIT_1B => X"EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAEBAE",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000000000F7EBF5FAFD7EBF5FAFD7",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"2ABEF00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0020105D557FEAA00557DE10AAD5554BA087FFFF55557BD54AAF7FBC01FFA280",
INIT_29 => X"7BD75EF087FFFFEF557BEAB45552E80155AA802AB45AA843FE0008557DFFF080",
INIT_2A => X"FAE820AA5D5557555082ABDF5508557DF45002ABDFFFF7803DE10AA80000AA08",
INIT_2B => X"0051555FFA2AA8200000557DFFFF7AA80000AAD1420AA087BD7555FFD168AAAF",
INIT_2C => X"5557FFDE10AAAEA8BFFA2FBD7545FFD157555085140010F7AEAABFFAAD542000",
INIT_2D => X"BA557BE8A10A284154BAFFAAAAB45007FC2155F7D155545AA80001EFAAFBEAB4",
INIT_2E => X"000A2D155410F7FFFFEBA08003FE00082AA8AAAAAFFC00BA00002AAAAF7D5574",
INIT_2F => X"0492E3F1C71C7BE8A2ABD7000000000000000000000000000000000000000000",
INIT_30 => X"3AE38145B78FD7000005010495B7AE921C517DE10A2DB50482147FFAF554971D",
INIT_31 => X"E3FE28B684070AA1C71D25D7007FFAFD7497BE8B5555208217DBE8A2AB45BE80",
INIT_32 => X"7FD257DFFD568A82FFA4870BA555F5056D002EBDF6D005B78F7D142ABDFC7F78",
INIT_33 => X"FAAAFBFFBED547038145B505FFB6A487000005F7AFD7F7A482038AADF4709214",
INIT_34 => X"AA8E071D7AAFBEFB455D71F8E00A2A0ADBC7A2FFD257DE3DF52555085142000F",
INIT_35 => X"21C002AA92FFDF574824171EAA10B680124BAFFAAAFB45007BC217DEBDB55555",
INIT_36 => X"00000000000000000000B6D550428FFF1FDE821C003FE001C2EAAAAAB6F5C208",
INIT_37 => X"0105D7BE8B55085142010AAD157545F7AEA8B550000000000000000000000000",
INIT_38 => X"01EFF7AAA8B55F7802AABA5D7FEAB45080015410007FEAA0055517DE00A2FFC0",
INIT_39 => X"E8BFF5D2ABDF55F7AABDEAAF784154BA5D5140145007BE8B55087BEAB555D040",
INIT_3A => X"0020BAA2FFD54105D7FC21EFFFD16AA10FF80174AA557FC21EF082EBFFEF007B",
INIT_3B => X"FBC0155085540000FFAEBFFEFF7D1554BA5D7BC01FFFF8015410007FEAB45F78",
INIT_3C => X"87FC01EFA2FFD7545AAAE97555A2FBFDF455D556AA00A2803FF45AAFFC21EFAA",
INIT_3D => X"552EAAAAAFFD1400005D042AA00F7FBD5410085568A10FF80020AAFFAABFF550",
INIT_3E => X"0000000000000000000000000000000000000F7D1400BAFFD57FE005D043FE10",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(13),        -- Port A data input
DOA(0)   => data_read_a_lo(13),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(13),        -- Port B data input
DOB(0)   => data_read_b_lo(13),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_14_16 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10020A000180000284008280000281800000030000000033022000000580002",
INIT_01 => X"000008020000204D006800000030824840000000084000084200090008510200",
INIT_02 => X"0220043170010A600A4D008040080000041000000028009002000F333240800C",
INIT_03 => X"111813400008002400000000C400090011000000610200001104D83000F14000",
INIT_04 => X"0801800100A000000000540084000040000040000800200000C8100000000748",
INIT_05 => X"0100000000001000000000002000080008000000001000000024024001200020",
INIT_06 => X"819EB84028001010000000080400000000000004108000100000020020040081",
INIT_07 => X"92040608000440100102400A94810206844200021DA2A0002000340800062C80",
INIT_08 => X"000000000084400008800A001214040441481500040000000000A7F408002244",
INIT_09 => X"0A0040090002008420401004104444004000020400214A208001000002400120",
INIT_0A => X"0400002020000000000000000000080C8008088100004590111B480040120000",
INIT_0B => X"1000000200404800000504016000002114000008020000020080024000000000",
INIT_0C => X"0410000010000000000040001000000000000040000000000001000000000000",
INIT_0D => X"04810244825010004010000000000000000000000000000000080000B8002104",
INIT_0E => X"0002C38280001202020800000000001000004000000000401022000002040902",
INIT_0F => X"20000587050001404E8084341CBA3404800828805200008000E0E0A000080002",
INIT_10 => X"4D18178E012010C00224004091C3514072C000444A0400080001C1C140001000",
INIT_11 => X"51709A07424142084458476001003809D0104B01C5710044020C4006010500C5",
INIT_12 => X"C26EE3803180C18006519462A00005001460E4730000050A1011004001060049",
INIT_13 => X"01F9E00660318000000538318740000140000001B4600CE80001400000002B62",
INIT_14 => X"0000000AD89857B0E0684411800000003799EB764D000330C300000000E3554B",
INIT_15 => X"0000021002002C000024008284001A0902000422E3F5960080480A0216A07240",
INIT_16 => X"4090240902409024090240902409024090081021020080015134920800480010",
INIT_17 => X"0902409024090240902409024090240902409024090240902409024090240902",
INIT_18 => X"9024090240902409024090240902409024090240902409024090240902409024",
INIT_19 => X"F5579B4E5C8FF0F7BE9D5F7DF650400200000000000000000000409024090240",
INIT_1A => X"9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7BF7DDDDDFCF3CF3D",
INIT_1B => X"F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE79E7",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000003FFF03F9FCFE7F3F9FCFE7F3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"420BA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"BD54AAF7FBC01FFA2802ABEFA2FBE8B55A2AE80000F7D5555555D2AAAABAAAD1",
INIT_29 => X"AA801FFA28402000AAAE955455500155EF0804155EFAAD5554BA087FFFF55557",
INIT_2A => X"7AEA8B45080417400AA843FE0008557DFFF0800020105D557FEAA00557DE10A2",
INIT_2B => X"087FFFFEF557BEAB45552E80155AA802AB4500516AA00A2AE800BAFFFFC20BAF",
INIT_2C => X"0AA80000AA005568ABAA28402010A2843FEBAFFFBD7410A2D168BFF087BD75EF",
INIT_2D => X"005D7FFDF4555517DFEF00043FEAA082ABDF5508557DF45002ABDFFFF7803DE1",
INIT_2E => X"000AAD1420AA087BD7555FFD168AAAFFAE820AA5D5557555002E80155A280000",
INIT_2F => X"0555412AA8ABAAADB40092000000000000000000000000000000000000000000",
INIT_30 => X"50482147FFAF554971D0492E3F1C71C7BE8A2ABD7A2FFEDB55B6A080038E3DB5",
INIT_31 => X"B7AE921C517DE10A2AE851FFB68402038AAAA955554900105FF0800175D7A2DB",
INIT_32 => X"A0800BAE3F1C0092EBAAADB6D080A12410BE803AE38145B78FD7000005010495",
INIT_33 => X"2D568BC71C71D25D7007FFAFD7497BE8B5555208217DBE8A2AB451C556FA00A2",
INIT_34 => X"142ABDFC7F78E3FE28B684070AA00516DABAA28402038B6803DE82F7F5D5410A",
INIT_35 => X"D002A80155B680000105D7FF8F455D5F78FD7000E3FEAA002EBDF6D005B78F7D",
INIT_36 => X"00000000000000000000AADF47092147FD257DFFD568A82FFA4870BA555F5056",
INIT_37 => X"F55FF84000AAAAFBC0145002AA8AAAAAFFC20000000000000000000000000000",
INIT_38 => X"01EF080417555A2FFC00105D7BE8B55085142010AAD157545F7AEA8B55A2FBFF",
INIT_39 => X"EAB45080015410007FEAA0055517DE00A2AA955FFFF80020BAAAAA9754508000",
INIT_3A => X"AA8B555D557FE00A280020BAAAD140000A2AEBFFEF082A82010F7802AABA5D7F",
INIT_3B => X"803DE00FFD557400AAD56AB455D5140145007BE8B55087BEAB555D04001EFF7A",
INIT_3C => X"82EBFFEF007BE8BFF5D2ABDF55F7AABDEAAF784154BA08557FEAAA284000AAFF",
INIT_3D => X"FF80174AA557FC21EF082A80145F780020105D7BEAB45557BE8B45082EBFEBA0",
INIT_3E => X"0000000000000000000000000000000000000A2FFD54105D7FC21EFFFD16AA10",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(14),        -- Port A data input
DOA(0)   => data_read_a_lo(14),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(14),        -- Port B data input
DOB(0)   => data_read_b_lo(14),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_15_16 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000A000000000284000280000001800020030000000033022000000180002",
INIT_01 => X"8000080000000048000000000000026040000000080000080200000000110200",
INIT_02 => X"0020042004010E60004C0080000800000410000000020090020000300245E005",
INIT_03 => X"0000010000080400000000408400480111000000610008000000C00000E54400",
INIT_04 => X"980000010000000088C2550080000040000040000008A00028C8100000120000",
INIT_05 => X"020004012E025000000001322000000A28008000011000000220004D41000000",
INIT_06 => X"819588000800101000011008040000100001060418800510000A620000000092",
INIT_07 => X"0000000800044004010C20008440810284020002102220002000340800062480",
INIT_08 => X"0000000001140800002C0A001214050540C800400406180000002DF004000244",
INIT_09 => X"1E00400900000000000016041044400440000000000042008001000000000022",
INIT_0A => X"0000000000000220000000000000080C00000081000045901118000040000000",
INIT_0B => X"0000000200404000010500004000000114000009000000000000004200000000",
INIT_0C => X"0000000000000000000040001000040001000000000000000001000020000800",
INIT_0D => X"000000000000001001208000180800000000030200000180800C400030002000",
INIT_0E => X"0000000000002600020800000000001080004000000000000002000000000000",
INIT_0F => X"A400000000000000000008000000000000000000000014800000000000000052",
INIT_10 => X"0000000000000000000000010240000000000000000000290000000000000000",
INIT_11 => X"2001C05838120800000000000000000000010000000000000000000000001804",
INIT_12 => X"081004000000000000A010000000000000902000000000180010002020000000",
INIT_13 => X"6600000000000000000024080000000000000000280400000000000000000000",
INIT_14 => X"0000000000200801000000000000000000501001920000000000000000000A40",
INIT_15 => X"0000020000000000000000003000000000000000000A101C3614000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000080000120980000000010",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000400200000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"28BEF00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"5555555D2AAAABAAAD1420BAFF8000010082A954BA00003DFEF085155400F784",
INIT_29 => X"AE95555A2FBE8BEFA2843DE00AA8015400FF84001EFA2FBE8B55A2AE80000F7D",
INIT_2A => X"2FBEAB45F7D56AABAAAD5554BA087FFFF55557BD54AAF7FBC01FFA2802ABEFF7",
INIT_2B => X"A28402000AAAE955455500155EF0804155EFFFFBE8BFF0800174AA557BFDE10A",
INIT_2C => X"A00557DE10F7D1574AAA2D16AB55FFD568BEF087FE8A1055003FE00A2AA801FF",
INIT_2D => X"00AA802AA00AAAE800BA5D0015545AA843FE0008557DFFF0800020105D557FEA",
INIT_2E => X"00000516AA00A2AE800BAFFFFC20BAF7AEA8B45080417400FFFFC21450800154",
INIT_2F => X"8FD7005150438F78A2DBFF000000000000000000000000000000000000000000",
INIT_30 => X"EDB55B6A080038E3DB50555412AA8ABAAADB40092E38E070280024904AA1C043",
INIT_31 => X"1C71C7BE8A2ABD7E3AA9257DA2FFE8BC7BE8E38E10A28017400E38A051FFA2FF",
INIT_32 => X"00124AA557FFDE10A2FBEDB6DF7D16AABAA2DB50482147FFAF554971D0492E3F",
INIT_33 => X"10038E38A2AE851FFB68402038AAAA955554900105FF0800175D7E3FFEFBD700",
INIT_34 => X"000005010495B7AE921C517DE10FFDF50482A2DB6AB45FFD56DBD7087BEAA384",
INIT_35 => X"0FFF1C017D140410400BE8E28A10AAA085082550A1057DBE803AE38145B78FD7",
INIT_36 => X"000000000000000000001C556FA00A2A0800BAE3F1C0092EBAAADB6D080A1241",
INIT_37 => X"4AA0800020BA550028B550855400AAF7AEBDFEF0000000000000000000000000",
INIT_38 => X"7400AAAE975EFA2FBFFF55FF84000AAAAFBC0145002AA8AAAAAFFC2000AAAA97",
INIT_39 => X"E8B55085142010AAD157545F7AEA8B55AAAE821EFAAFBEAB55F7AAA8A00AA841",
INIT_3A => X"417555AAFFFDF450804020AA557BFFE10A2FFFFFEFF7D568ABAA2FFC00105D7B",
INIT_3B => X"D17DF45007FE8AAA08002AAAAA2AA955FFFF80020BAAAAA975450800001EF080",
INIT_3C => X"7802AABA5D7FEAB45080015410007FEAA0055517DE00FFFBC2000AAFBE8B55F7",
INIT_3D => X"A2AEBFFEF082A82010FFD5421EF5D0000010F7AAA8A10AA8017400552A801EFF",
INIT_3E => X"00000000000000000000000000000000000005D557FE00A280020BAAAD140000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(15),        -- Port A data input
DOA(0)   => data_read_a_lo(15),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(15),        -- Port B data input
DOB(0)   => data_read_b_lo(15),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_16_16 : RAMB16_S1_S1
generic map (
INIT_00 => X"DA22C618B1000482B688B186588884862A400438255FC38381441205BA803003",
INIT_01 => X"7045A80028404C211203A952A90341080B173340412000E1005D628000820484",
INIT_02 => X"428406A4000850848330118D0AAC55001349B108818005460229044001C01784",
INIT_03 => X"092C4020000500020000500986812C405000001A48202050000A214AC0650115",
INIT_04 => X"4804A55440256F504025E003A054F46415A4E62B6FE3307943965A00001A1152",
INIT_05 => X"0000001C40A5B950ADB8EA097057ECE14C86D2B7F85AAD17F4B100000B88148C",
INIT_06 => X"415401DCDCF2C0A8030140BCB0820A200342A1C641C1E8782F508F2B00003584",
INIT_07 => X"002701881A3202080AE00480A2002840BE1480FA004342AA6F12000054004867",
INIT_08 => X"08C54828091002000002B32A8C19064E486A8001510000014140C1E2A14891E0",
INIT_09 => X"015452B103020814004088B64102680B6596594800400413CAC0208944800000",
INIT_0A => X"96AA000484094C000000000000012C9000A0000D0A80000BF8028E87C1B99270",
INIT_0B => X"014808A02004200E540480212000A448C0082024AE50064B44000000000002A2",
INIT_0C => X"0004000D5846256AAEA811150445411150445411150445411150422A088A8200",
INIT_0D => X"00000004010042A204A0C5817D00005034052E40000817D00440004004AD3240",
INIT_0E => X"632B2673FA4587978A2004102800809225545155121740000004900090000000",
INIT_0F => X"00C6564CE7F4EA4B940076D296D003030800462CBD320018CAAAACFE9164C800",
INIT_10 => X"28834ADB1440A114793A4A30A40839AA14910D08DCB2640031955559FD3AC990",
INIT_11 => X"594AB0B1A025371CA0E034E8443C097A800EB090D4AAC91208ED2FA0CE5E09B1",
INIT_12 => X"7B50446083001B94BB38C540EBE61284BB304880E3E4579EDC00992980D58033",
INIT_13 => X"5511121840E7A2CD952ECC12ABC3E6ACB3DFB12ECE315000F61FF1727A85FDBC",
INIT_14 => X"75DEB07F6F2E7084517F126F8395CB2BEFBAB8BA8AF698228CC5E2F08ECA5159",
INIT_15 => X"5580A840A8009F8B108C80A1021B080AFC0DF6422C6077F4A77F20D0C0E21084",
INIT_16 => X"0000000000000000000000000000000000044000102A0001148442A110810359",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"558D11544C690DA64C1C4F68A360400000000000000000000000000000000000",
INIT_1A => X"14D14D14D14D14D14D14D14D14D14D14D14514514514514529E5F87869E79E78",
INIT_1B => X"D1E8F47A3D1E8F47A7D3E9F4FA7D3E9F4FA7D3E9F47A7D1E9F47A7D1E9F4D14D",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000007D3E9F4FA7D3E8F47A3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"C00AA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"03DFEF085155400F78428BEF087FFFFEFF7D168B55AAD17FFFF552EBFE00007F",
INIT_29 => X"2E975EFF7D568BFFFF80175EF0004000BA552A821FFFF8000010082A954BA000",
INIT_2A => X"55540000082EAABFFA2FBE8B55A2AE80000F7D5555555D2AAAABAAAD1420BA5D",
INIT_2B => X"A2FBE8BEFA2843DE00AA8015400FF84001EF0000020AA5D00154005D043FF455",
INIT_2C => X"FA2802ABEF557BEABEF5D0415410087FD74BAAAAEBFFEF557FC00AAF7AE95555",
INIT_2D => X"FFFFAABFEAAFF84001FF002A821FFAAD5554BA087FFFF55557BD54AAF7FBC01F",
INIT_2E => X"000FFFBE8BFF0800174AA557BFDE10A2FBEAB45F7D56AABA082A97545F7D16AB",
INIT_2F => X"FFEF552AB8E38087FC2092000000000000000000000000000000000000000000",
INIT_30 => X"070280024904AA1C0438FD7005150438F78A2DBFF0871F8FC7E3D56AB6DBEDB7",
INIT_31 => X"AA8ABAAADB400924920925EFF7D16ABFFE38E175EF1400000BA412E871FFE38E",
INIT_32 => X"0A1240055003FF6D5551420101C2EAFBD7A2FFEDB55B6A080038E3DB50555412",
INIT_33 => X"57FC00BAE3AA9257DA2FFE8BC7BE8E38E10A28017400E38A051FF0804050BA41",
INIT_34 => X"4971D0492E3F1C71C7BE8A2ABD74975EDBC7550E12410087FD74AAB6AABFFC75",
INIT_35 => X"A08249756DF7D168BC7F7AABAEAAF780051C70824851D7A2DB50482147FFAF55",
INIT_36 => X"00000000000000000000E3FFEFBD70000124AA557FFDE10A2FBEDB6DF7D16AAB",
INIT_37 => X"B55A2D16ABEFFFFBFDFFF552AAAAAA007BC00000000000000000000000000000",
INIT_38 => X"20AA002A955EFAAAA974AA0800020BA550028B550855400AAF7AEBDFEF08516A",
INIT_39 => X"000AAAAFBC0145002AA8AAAAAFFC20000000021EFF7D568BFFA2AA955FF5D040",
INIT_3A => X"E975EF0800174BA002E820105D003DFEF5D51420005D2ABFF45A2FBFFF55FF84",
INIT_3B => X"7BD74AAF7AEBDF455D7BC20BAAAAE821EFAAFBEAB55F7AAA8A00AA8417400AAA",
INIT_3C => X"2FFC00105D7BE8B55085142010AAD157545F7AEA8B5500557DF45552A8200000",
INIT_3D => X"A2FFFFFEFF7D568ABA0804155FFF7D568B55FFAAAAABAFF8415545000015555A",
INIT_3E => X"0000000000000000000000000000000000000AAFFFDF450804020AA557BFFE10",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(16),        -- Port A data input
DOA(0)   => data_read_a_lo(16),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(16),        -- Port B data input
DOB(0)   => data_read_b_lo(16),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_17_16 : RAMB16_S1_S1
generic map (
INIT_00 => X"5284CE4FB7BD2C8994A13392DBD02E14006B82AC7E800D44D3DD2FD5F9B961C0",
INIT_01 => X"2EACD01F7E03FC6793F2199B39FC233C11D93AE6F3BB92B32091DBC339B24542",
INIT_02 => X"E63CCCC00A82C08092A2AFAE667033DB50853379C10BFDC5C6F4044443C817C6",
INIT_03 => X"7FF183635AEF9E3635AEF9E18E237040404446965C0607EE6DB7854AC4DE060C",
INIT_04 => X"D78AC33FB604488B000892EF17BE6D84196482236FE100294152E294350FB697",
INIT_05 => X"081B5F9B409420D0CDB47A05403F6CE0C08A4AB7F840EDB6F48100DFC8081081",
INIT_06 => X"768465354781CBC30316367077B4BDB50646E8D87100A8201ED01C19C020F71A",
INIT_07 => X"4002A110C922480A82D0841147162C48EBB9537A0022DC67987042EE976ABEA7",
INIT_08 => X"DB931BFEF91C00002CC0E019C0C82A4E4820C15A2330E004401891181168C4D1",
INIT_09 => X"09F3A1BC11EFBC66DB65307071477FF1030C397C060B4254064302042F803A69",
INIT_0A => X"3F330802162F3B7EE3F3EC7C7DEF207000F00059D2ED56D7EED2ED3C9A867DC0",
INIT_0B => X"185C44B91BC1740B7605040BE0018CFC7429F326B9E822FFC00074D5A0AB033A",
INIT_0C => X"00367A28FC1B7F7FEFFCFBFF3EFFCFBFF3EFFCFBFF3EFFCFBFF3EFFE7DFF9E00",
INIT_0D => X"0000000008004BA78428C7AD7FC94B533F5B4FFBD2FAD7FCCA786D43FE67C218",
INIT_0E => X"BA494CEBFD4F2667ABB6F68B29760593F33FA0CF170F40006001B1A05C000000",
INIT_0F => X"7F749299D7FAEB237DFE5865B6D2BF23265CBACE542A6FEE92333AFF33E0A9BF",
INIT_10 => X"F6C24B6D18C3C9F8E2881F3F787D776B5DB94A09955054DFDD246675FE7AC153",
INIT_11 => X"BFB349E08FF9A27EDE9FA8AEFD9E7467BFCB195CFEB56A1A70D34D1706FFFA3E",
INIT_12 => X"6FE219CA80725B875EED723FF7FCB2875EDAAFEAF7FD929BFD55BBC71D79F639",
INIT_13 => X"546670D018E7A6E581D7B6AB75FDFCECA6E581D7BB5DDFC6FF0EB7D7E859FDB5",
INIT_14 => X"B978177F6D6AF5ECDB5FB76A5F5FA165B456E0FB308710C49FCFB741598B9C7E",
INIT_15 => X"CFDAAB00AC00A8BBFC8B501CF7A0FED9A540EA1952586CEB54D143ACFF9A3BA9",
INIT_16 => X"000000000000000000000000000000000026E100002F382DBD9ECFE117805F20",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"4372003009EDCC4052E917114F981800C0000000000000000000000000000000",
INIT_1A => X"BA69A69AEBA69AEBA69A69AEBA69AEBA69A69A69A69A69A68698686981D75D74",
INIT_1B => X"6A351A8D46A351A8D068341A0D068341A0D068341A0D46A341A0D46A341A69AE",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000000000046A351A8D46A351A8D4",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"7FEAA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"17FFFF552EBFE00007FC00AA087FFFFFFFFFFFFFEFF7FBEAB450804001EFAAD5",
INIT_29 => X"D168A000004020AA5D7BE8B450051401EF087FD74AA087FFFFEFF7D168B55AAD",
INIT_2A => X"D7FEAB55FF80175EFFF8000010082A954BA00003DFEF085155400F78428BEFAA",
INIT_2B => X"F7D568BFFFF80175EF0004000BA552A821FF5D00020BA552A82000552A821555",
INIT_2C => X"AAAD1420BAFFFFFDF45AAD17FFFFAAFBC01EF5D0015555557BFDEBA5D2E975EF",
INIT_2D => X"BA007FEABEF005555555A2D1554BAA2FBE8B55A2AE80000F7D5555555D2AAAAB",
INIT_2E => X"0000000020AA5D00154005D043FF45555540000082EAABFF00516AA10552E820",
INIT_2F => X"8B550000071EFB6DF7AE92000000000000000000000000000000000000000000",
INIT_30 => X"F8FC7E3D56AB6DBEDB7FFEF552AB8E38087FC2092147FFFFFFFFFBFDFC7EBF5E",
INIT_31 => X"150438F78A2DBFFBED16AA381C0A07082497FEFB6D1451471EF007BD04920871",
INIT_32 => X"2A850105D2A80155417BEFB6DEB8E175FFE38E070280024904AA1C0438FD7005",
INIT_33 => X"D7BFAEBA4920925EFF7D16ABFFE38E175EF1400000BA412E871FF550A0009249",
INIT_34 => X"E3DB50555412AA8ABAAADB40092FFF5FFF6DAADF7FFD7B6F1C71EF55001756D5",
INIT_35 => X"7145B6AA28492487082007FEDBD700515556DA2DF50492A2FFEDB55B6A080038",
INIT_36 => X"000000000000000000000804050BA410A1240055003FF6D5551420101C2EAFBD",
INIT_37 => X"FEFF7FBFFF55A2D16AB550000175EFFFFBEAA000000000000000000000000000",
INIT_38 => X"55EF087FC200008516AB55A2D16ABEFFFFBFDFFF552AAAAAA007BC0000557FFD",
INIT_39 => X"020BA550028B550855400AAF7AEBDFEFF7D568AAA5D2A97410007BFFFFF55515",
INIT_3A => X"A955EF5D2E80010002A954005D2A82155087FFFFEFAAAA975EFAAAA974AA0800",
INIT_3B => X"D1575FF5504175EF5D7FEAAAA0000021EFF7D568BFFA2AA955FF5D04020AA002",
INIT_3C => X"2FBFFF55FF84000AAAAFBC0145002AA8AAAAAFFC2000FFD57DFFFAAFFFDF55FF",
INIT_3D => X"5D51420005D2ABFF45557FE8AAA000415410007BFFF450051555EFA2FBC0000A",
INIT_3E => X"00000000000000000000000000000000000000800174BA002E820105D003DFEF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(17),        -- Port A data input
DOA(0)   => data_read_a_lo(17),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(17),        -- Port B data input
DOB(0)   => data_read_b_lo(17),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_18_16 : RAMB16_S1_S1
generic map (
INIT_00 => X"69844019080000A21A611406840014122A641074155FC28A2024001001801003",
INIT_01 => X"7443D920034004180005E9E3C90360C0041C0181002001602025800008440084",
INIT_02 => X"E2DCCCE61D5C008103F2000781FC0FEDEAC2161B0B8FB0008620044443006010",
INIT_03 => X"884E300802006900802006995C896D605200000856E24A040000640052141103",
INIT_04 => X"480520FC026125AC0025C9122644E3E40EC8E2001001302281841A009038A86A",
INIT_05 => X"432000040089983070019400F01010004C8DB841405A80A100B586200FAC24AE",
INIT_06 => X"09044359DC7040000000002C109B0E0A00A1104641C0803804000707284600E1",
INIT_07 => X"400D10100400481D5EB08501620000007500CE801241021FE78E404860140060",
INIT_08 => X"00880C0106A0528020019307CC082A0A4A6A01ED725021400040D028000A9729",
INIT_09 => X"00117063038000282081402E4106400B6186128040600C10C1C0200950508110",
INIT_0A => X"C0C30C2E21580C874004008080003C32A10A19090C02010E1022944061688000",
INIT_0B => X"0180A8062026000DC425C0301311324AA2373088479105D044A1022000001835",
INIT_0C => X"0D89844703649000000200000000000000000000000000000000000000000010",
INIT_0D => X"0D8306C182701404C1973010802020404084001E00010802046092B5001FB365",
INIT_0E => X"528EB314068AB8B803DB00002900800400FC503F08180050942E4200020C1B06",
INIT_0F => X"40A51D66280D6032C5F96D3C51555D5D7D5AA87285820814A3CCC501C2A60820",
INIT_10 => X"8B35A3FEBF1FEDFD9C2B30E0468AAAD5D48F37E8FC1304102947998A03984C10",
INIT_11 => X"440FE1DD772D37A0A321BC6968F32658BF2D4F2A80BF8FE3F9FE3AC362080529",
INIT_12 => X"5487910D7E5A6D961A28456A1832E5161A100DD5182BC54020EA67A189C6ED36",
INIT_13 => X"AA444CAF91EDD1B725868403BE06323551B725868A100ABD119753B70964122B",
INIT_14 => X"EDC259048ACD868EE3803D65CEDC258A8F80D55E007C3F8EBB56F4C5362C978F",
INIT_15 => X"3F240014BE84370001B6922070440556B15F7FABBC0031BCF2257C41634B14D4",
INIT_16 => X"C1B06C1B06C1B06C1B06C1B06C1B06C1B0491069068000004060300A005A0118",
INIT_17 => X"1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06",
INIT_18 => X"B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C",
INIT_19 => X"B28BBECEB80EE173C2300F7DF16000000000000000000000000041B06C1B06C1",
INIT_1A => X"8A28A28AAAAAAA28A28A28AAAAAAA28A28A28A28A28A28A2910591505C104104",
INIT_1B => X"28944A25128944A25128944A25128944A25128944A2552A954AA5128944AAAA2",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000128944A25128944A251",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"9540000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"BEAB450804001EFAAD57FEAA087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974BA082E",
INIT_29 => X"7FFFFFFFFFBFDF45AAD568B55080028B55002E82000087FFFFFFFFFFFFFEFF7F",
INIT_2A => X"0043DE10AA843DE00087FFFFEFF7D168B55AAD17FFFF552EBFE00007FC00AA08",
INIT_2B => X"0004020AA5D7BE8B450051401EF087FD74AAAAFFFDF45A2D16AB55F7FFFFFFF0",
INIT_2C => X"0F78428BEFAA80000000804154BA55042ABEF5D7FD75FFAAD540145AAD168A00",
INIT_2D => X"00082E95555085168A10557FD7545FF8000010082A954BA00003DFEF08515540",
INIT_2E => X"0005D00020BA552A82000552A821555D7FEAB55FF80175EF5D00020105D2A974",
INIT_2F => X"DFFF5D2A954AA082A92428000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFBFDFC7EBF5E8B550000071EFB6DF7AE921C7FFFFFFFFFFFFFFFF7FBF",
INIT_31 => X"AB8E38087FC2092087FFDFC7E3F1FAF55A2DF6DB7D1C002AB7D002A82028147F",
INIT_32 => X"DF6DB7DE3F5FAFC708003DE28B68E38E280871F8FC7E3D56AB6DBEDB7FFEF552",
INIT_33 => X"ADF4516DBED16AA381C0A07082497FEFB6D1451471EF007BD0492B6F1F8F55AA",
INIT_34 => X"1C0438FD7005150438F78A2DBFFA28407038140410492550A2ABC7497BD25FFA",
INIT_35 => X"F5D0E05000492097428002E9557D1C516FA28417BD5545E38E070280024904AA",
INIT_36 => X"00000000000000000000550A00092492A850105D2A80155417BEFB6DEB8E175F",
INIT_37 => X"FFFFFFFFDFEFF7FBFFFEF552E974AA082A820AA0000000000000000000000000",
INIT_38 => X"ABEF002A800AA557FFDFEFF7FBFFF55A2D16AB550000175EFFFFBEAA00557FFF",
INIT_39 => X"6ABEFFFFBFDFFF552AAAAAA007BC0000087BFDF45AAD568B55AAFBFDFEF55042",
INIT_3A => X"FC2000FFD56AB45A2FFFDFFFAAD16AB4500043DEAAFFAEAAAAA08516AB55A2D1",
INIT_3B => X"2AA8B45087FC01EFA2FFD55EFF7D568AAA5D2A97410007BFFFFF5551555EF087",
INIT_3C => X"AAA974AA0800020BA550028B550855400AAF7AEBDFEFA280154BA55040000055",
INIT_3D => X"087FFFFEFAAAA975EF5D2E974000804154BA082A975EF5D517DEAA007BD5545A",
INIT_3E => X"00000000000000000000000000000000000005D2E80010002A954005D2A82155",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(18),        -- Port A data input
DOA(0)   => data_read_a_lo(18),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(18),        -- Port B data input
DOB(0)   => data_read_b_lo(18),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_19_16 : RAMB16_S1_S1
generic map (
INIT_00 => X"042200000000000041088001001AA00000000000000000000000500802000003",
INIT_01 => X"040048000024000000000404000000000A22000800000800004A200000000001",
INIT_02 => X"200C8840085EB00480060000001C008002489E0F000405EA0004040404000000",
INIT_03 => X"24004000000000000000000900002C4050000000000069500208400002E14100",
INIT_04 => X"4800200C0000000044002000C80020E40000E200000130200188000000800100",
INIT_05 => X"000000000080181000000000701000004C8000000058800000B1000009880480",
INIT_06 => X"80500081081040000000002C100040400000004641C080380400070100000000",
INIT_07 => X"4020109801A4CE005C00048380142810010564C4100114012002402028044808",
INIT_08 => X"0070700000000000000083004C3902420062000020E0000100004082A140102B",
INIT_09 => X"001150200000000000000026400000016186100000000010C04002C000000000",
INIT_0A => X"007C00008082C0002000000000002C3000000004050001030102040000000000",
INIT_0B => X"0000000000000000000000000000010000800011000000000000000000000BC0",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"000000000000000000000000000000042000760000000000000000010004B200",
INIT_0E => X"0D74002280300F0002FB069040000060000C5003000800000000000000000000",
INIT_0F => X"C01AE8004500744C780687DBA828008080A5FC0D385598035D0008A00C015660",
INIT_10 => X"39D8140040201BF861F0E7D693E6170022408116DFE0AB3006BA0011401D02AC",
INIT_11 => X"5412E4997F5249FD005043B8680CC98F00D0F2DD0140100406FE053A98F6ECC7",
INIT_12 => X"7418663001858040E153888000010840E165D0000000285C246A181C03FE4662",
INIT_13 => X"8199830066F0020858385974000001260208583854E2200000660208D6B1423F",
INIT_14 => X"8235AC508FCE8811042040F008235AE04420C040CF00C031C80009B8F224978B",
INIT_15 => X"030004E00000C220010808C10D9A92A74CD7CF4A09051110AD5A3C9200B7F280",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000118",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"07208BBA3F0C7010C660C7441920000000000000000000000000000000000000",
INIT_1A => X"861869A61861861861869A61861861861861861861861861A8208C4C1534D34C",
INIT_1B => X"984C26130984C26130984C26130984C26130984D26930984C26130984C261861",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000984C26130984C26130",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"174BA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFDFEF5D2A974BA082E95400F7FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0004",
INIT_29 => X"FFFFFFFFFFFFFFFFF7FBFDFFF552E974BAA2FFFFE10087FFFFFFFFFFFFFFFFFF",
INIT_2A => X"004001EFAAAEA8ABA087FFFFFFFFFFFFFEFF7FBEAB450804001EFAAD57FEAAF7",
INIT_2B => X"FFFBFDF45AAD568B55080028B55002E82000F7FFFFFFFFFFFFDFEFA2D568B550",
INIT_2C => X"0007FC00AAF7FFFFFFFF7FBE8B55AAD16ABEF5D2ABFF55080402010087FFFFFF",
INIT_2D => X"55A2FFFDFEF5D2EBFE00AAFFFFEBA087FFFFEFF7D168B55AAD17FFFF552EBFE0",
INIT_2E => X"000AAFFFDF45A2D16AB55F7FFFFFFF00043DE10AA843DE00557FFDFEFA2D16AB",
INIT_2F => X"FFEF552A974AA0000104AA000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFF7FBFDFFF5D2A954AA082A92428E3FFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"0071EFB6DF7AE92EBFFFFFFFFFFFFDFEFF7F5FAFC7492A974AAB6F5F8E101C7F",
INIT_32 => X"F1F8FD7AAD16AB450000001FFBEA4A8AAA147FFFFFFFFFBFDFC7EBF5E8B55000",
INIT_33 => X"00000010087FFDFC7E3F1FAF55A2DF6DB7D1C002AB7D002A82028FFFFFFFEFF7",
INIT_34 => X"BEDB7FFEF552AB8E38087FC2092F7FBF8FC7E3F5EAB45B6DF6FBEF5D2AB8F7D0",
INIT_35 => X"84971F8FC7AAD56DB6DBEF5F8FD7412ABFE28B6F5F8E820871F8FC7E3D56AB6D",
INIT_36 => X"00000000000000000000B6F1F8F55AADF6DB7DE3F5FAFC708003DE28B68E38E2",
INIT_37 => X"FFFFFFFFFFFFFFFFFDFEF552E954AA0004000AA0000000000000000000000000",
INIT_38 => X"54AAF7D568A00557FFFFFFFFFFFDFEFF7FBFFFEF552E974AA082A820AAA2FFFF",
INIT_39 => X"FFF55A2D16AB550000175EFFFFBEAA00A2FFFFFFFF7FBFDFFFFFD568B55002A9",
INIT_3A => X"A800AAF7FBFDFEFF7D56AB45AAD56AB450004001EFFF842AAAA557FFDFEFF7FB",
INIT_3B => X"FFFFFFF552AA8BEF080402000087BFDF45AAD568B55AAFBFDFEF55042ABEF002",
INIT_3C => X"8516AB55A2D16ABEFFFFBFDFFF552AAAAAA007BC0000FFFBE8B55AAD168B55F7",
INIT_3D => X"00043DEAAFFAEAAAAA08556AB55A2D57FFFFF7D568B45002ABDEAAFFD16AA000",
INIT_3E => X"0000000000000000000000000000000000000FFD56AB45A2FFFDFFFAAD16AB45",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(19),        -- Port A data input
DOA(0)   => data_read_a_lo(19),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(19),        -- Port B data input
DOB(0)   => data_read_b_lo(19),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_20_16 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000003",
INIT_01 => X"F55FF80000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"E05022020800008400F655001FFCFF80018FA804400000000000004400000001",
INIT_03 => X"00000000000000000000000900002CC07000000000000000000000000000013F",
INIT_04 => X"68002FFE40900010000180000001FFEC0012EE0C001370F40780000000000000",
INIT_05 => X"0840000880FCBBF0100E204DF0F88311DD8005080679800000F3000029980580",
INIT_06 => X"001000030817C8E8840155FDF9001001050023F6C3C3D0F87FA19F7F011000E4",
INIT_07 => X"000000090492260800008000EE00000000000000002101FF2002C00000004018",
INIT_08 => X"2A040001071004000013FF7FCA302C0C0008214800002101554031F800000000",
INIT_09 => X"801F57F200000090000489FEC0000001EFBEF0040008023FDFC0000000004006",
INIT_0A => X"0000000008000000000000000000ADF000000200000008000008028300110230",
INIT_0B => X"0000000000000800080000000000000000000000000000000800800A40000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"000000040900005C848538000020000000800000080000020000800101FFB600",
INIT_0E => X"00800000003A010003000000000000600FFC53FF001800000002004080000000",
INIT_0F => X"0001000000007408040000004000000004E9000008020000200000000E800800",
INIT_10 => X"00200000000313100010002000008000000000129600040000400000001D0010",
INIT_11 => X"81C012060000000000218F7840000100800004000000000066C0000080080000",
INIT_12 => X"800000000017C000100000000001A800080000000001A8040000002840008185",
INIT_13 => X"0000000006F00000100200000000012600001004000000000066000000801040",
INIT_14 => X"0000200410100000000005F00000020080090A0000000085C800002000586000",
INIT_15 => X"FF00400000000000020020020001000040283024E4F2860400008000030ED080",
INIT_16 => X"00000000000000000000000000000004010201001003020200000000000127DB",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"A0700030038200010089120104D2040020000000000000000000000000000000",
INIT_1A => X"2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2C30C30C30C30C306982121A1E79E79",
INIT_1B => X"32190C86432190C86432190C86432190C86432190C86432190C86432190CB2CB",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000432190C86432190C864",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0201000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF552A974AA0004174BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA0804",
INIT_29 => X"7FFFFFFFFFFFFFFFFFFFFFFEF552E954AA000400000F7FFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E954BA007FC00BA087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974BA082E9540000",
INIT_2B => X"FFFFFFFFFF7FBFDFFF552E974BAA2FFFFE10FFFFFFFFFFFFFFFFFFFFFBFDFFF5",
INIT_2C => X"FAAD57FEAA007FFFFFFFFFFFFFEFF7FBFFF550800020BAAAD56AAAAF7FFFFFFF",
INIT_2D => X"EFF7D56AB450000021EFA2D57DE10087FFFFFFFFFFFFFEFF7FBEAB450804001E",
INIT_2E => X"000F7FFFFFFFFFFFFDFEFA2D568B550004001EFAAAEA8ABA5D7FFFFFFFFFFFDF",
INIT_2F => X"FFFF5D2E954AA080005000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFEF552A974AA0000104AAFFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"A954AA082A92428087FFFFFFFFFFFFFFFFFFBFDFEF5D2E974AA000A07000E3FF",
INIT_32 => X"FFFFFEFF7FBFFFFF552E974AA0071C50BA1C7FFFFFFFFFFFFFFFF7FBFDFFF5D2",
INIT_33 => X"EDF6FABAEBFFFFFFFFFFFFDFEFF7F5FAFC7492A974AAB6F5F8E10E3FFFFFFFFF",
INIT_34 => X"EBF5E8B550000071EFB6DF7AE921C7FFFFFFFFFBFDFEFE3F5F8F450004050AAB",
INIT_35 => X"A497FFFFFFF7FBF8FC7EBD168B450804021FFB6D57DE28147FFFFFFFFFBFDFC7",
INIT_36 => X"00000000000000000000FFFFFFFEFF7F1F8FD7AAD16AB450000001FFBEA4A8AA",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2A954AA0800174100000000000000000000000000",
INIT_38 => X"74AA002E95410A2FFFFFFFFFFFFFFFFFFFFFDFEF552E954AA0004000AAFFFFFF",
INIT_39 => X"FDFEFF7FBFFFEF552E974AA082A820AA087FFFFFFFFFFFFFEFF7FBFDFFF5D2A9",
INIT_3A => X"568A00AAFFFFFFFFFFBFDFEFFFFFFDFEF5D2E954AA0051554BA557FFFFFFFFFF",
INIT_3B => X"D16AB450804174AAFFFFFFEBAA2FFFFFFFF7FBFDFFFFFD568B55002A954AAF7D",
INIT_3C => X"57FFDFEFF7FBFFF55A2D16AB550000175EFFFFBEAA005D7FFFFEFF7FBFDFFFAA",
INIT_3D => X"0004001EFFF842AAAA087BFDFEFF7FFEAB45A2D568B550804001EFF7D57DEBA5",
INIT_3E => X"0000000000000000000000000000000000000F7FBFDFEFF7D56AB45AAD56AB45",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(20),        -- Port A data input
DOA(0)   => data_read_a_lo(20),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(20),        -- Port B data input
DOB(0)   => data_read_b_lo(20),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_21_16 : RAMB16_S1_S1
generic map (
INIT_00 => X"4A302428B824900A128C090A5C1800261500213C005FE812D10420054085A202",
INIT_01 => X"001FFE3440B609703B0427F801A40B8115BC4F655300340288A40D30040E4DD8",
INIT_02 => X"E00424256888D8819801000F9FFFFFFFF149FF1FCA448046C60A0D2437C517F9",
INIT_03 => X"20030640003250640003250F06002CC1740002019824E001CD357832440001FF",
INIT_04 => X"EA2C3FFD400006E04401A8837001FFFC004AEF00080B70E08FB5789421007C5C",
INIT_05 => X"00011A0C40F9FFF80920954FF0F00809DF84A0202879800000F3000029980780",
INIT_06 => X"0805984B7A1FC0A0000101FFF0480080002281F7C3C381F87C03DFFF00009004",
INIT_07 => X"B424068086A205481A60A19000908204A855B000A08A61FF20C3D004D331D340",
INIT_08 => X"1BFA0001600802000023F7FFC08D234B40C2028253000040114200000D0226C0",
INIT_09 => X"EF1F5FF054096C6ADBA169FFC202B1C1FFBEF0440021083DFFCE22DC2880E24D",
INIT_0A => X"45FF0C004041D84862A28C54518DBFF00020004C0A6044901112A0908AA0A300",
INIT_0B => X"018C241102068006C620C03882019480E63180855A492712CC01C49C20201BFE",
INIT_0C => X"08A9464116544302C02D92236488D92236488D92236488D922366446C911B210",
INIT_0D => X"08800444021048034004001890000806002804A0822189000900D80621FFBE00",
INIT_0E => X"060580261013813A2CC396506102C4053FFD5BFF00A04A00200602CA52001100",
INIT_0F => X"080C0B004C202621A85C09411500135844C196D3606941018150098404C1A304",
INIT_10 => X"B02901013416181C96C2C9C600890A2028172192C460D1820302A0130809834A",
INIT_11 => X"9C5E803408250180AC268D185DB3F4350B811068C00049A0A4AA68F05C96A001",
INIT_12 => X"002C006560138F032B1804101244C883052208209040CC849063A747512B7678",
INIT_13 => X"41401E240665750440C9488280254530314080C2C601040420352148A00501B1",
INIT_14 => X"500811204D000700114204A70422016149916011008CAA8858850B00C32591C0",
INIT_15 => X"FFC06E60AC0496022300233104663040808E991765205000070121D41D18D098",
INIT_16 => X"40100401004010040100401004010040102090010008000001C0E010020007DF",
INIT_17 => X"0100401004010040100401004010040100401004010040100401004010040100",
INIT_18 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_19 => X"FFEF9FEEFF7FFDF7FF3E3DFDF7E0000000000000000000000000401004010040",
INIT_1A => X"BEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBFFDFDFFFCF3CF3F",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFEFF7FBFDFEFF7FBFDFEFBEF",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000FFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0001000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E954AA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0004",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA0004154BAFFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"52E974BA0804000AAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0004174BAFF",
INIT_2B => X"FFFFFFFFFFFFFFFFEF552E954AA000400000007FFFFFFFFFFFFFFFFFFFFFFEF5",
INIT_2C => X"A082E95400007FFFFFFFFFFFFFFFFFFFFDFEF5D2E974BA002E97400007FFFFFF",
INIT_2D => X"FFFFFBFDFEF5D2A954AA002E974BA087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFBFDFFF5D2E954BA007FC00BA5D7FFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA000002000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080005000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"A974AA0000104AAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974BA0000174AAFFFF",
INIT_32 => X"FFFFFFFFFFFFDFEF552E954BA080A000AAE3FFFFFFFFFFFFFFFFFFFFFFFEF552",
INIT_33 => X"02A95400087FFFFFFFFFFFFFFFFFFBFDFEF5D2E974AA000A07000007FFFFFFFF",
INIT_34 => X"F7FBFDFFF5D2A954AA082A924281C7FFFFFFFFFFFFFFFFFFBFDFEF5D2A974BA0",
INIT_35 => X"A557FFFFFFFFFFFFFFFF7FBFDFFF552E974BA0020924BA1C7FFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000E3FFFFFFFFFFFFFFEFF7FBFFFFF552E974AA0071C50B",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0000020000000000000000000000000000",
INIT_38 => X"74BA0000174BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954AA080017410FFFFFF",
INIT_39 => X"FFFFFFFFFFDFEF552E954AA0004000AAF7FFFFFFFFFFFFFFFFFFFFFFFEF552A9",
INIT_3A => X"E95410087FFFFFFFFFFFFFFFF7FBFDFEF5D2A954BA082E800AAA2FFFFFFFFFFF",
INIT_3B => X"FBFFFFF552E954BA002E97410087FFFFFFFFFFFFFEFF7FBFDFFF5D2A974AA002",
INIT_3C => X"57FFFFFFFFFFFDFEFF7FBFFFEF552E974AA082A820AA557FFFFFFFFFFFFFEFF7",
INIT_3D => X"5D2E954AA0051554BA5D7FFFFFFFFFBFDFEFF7FFFFFEF5D2A974BA0000020AA5",
INIT_3E => X"0000000000000000000000000000000000000AAFFFFFFFFFFBFDFEFFFFFFDFEF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(21),        -- Port A data input
DOA(0)   => data_read_a_lo(21),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(21),        -- Port B data input
DOB(0)   => data_read_b_lo(21),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_22_16 : RAMB16_S1_S1
generic map (
INIT_00 => X"5290F4CDE914905A14A43D33F488243E17122300F55FEB189B343A1140548380",
INIT_01 => X"A54007B259F6A975386262000C344BA9573C6FF57B18A5FB0ABFCD3C2C5F4F0C",
INIT_02 => X"021DFF8C38B3C009D203551040030071869D0040180AA2DC53DB89BEA8204001",
INIT_03 => X"2603475A969D0475A969D0460EAA401005111011BD506954EDB40F5EF41434C0",
INIT_04 => X"922D9002100ED69E443D988B0D5400103E48003D0800011E803B06B5B9125A15",
INIT_05 => X"281B5A0C06000408F4DF9422010D8802022F2124A8022492580040440002021C",
INIT_06 => X"F780C4C052881ADA0E05440205DA50930FA182010004700083E220800440B588",
INIT_07 => X"049D028B93FB561833D8094A02F5EA92FD7247E10305C40040D136E6A023F7FC",
INIT_08 => X"00028241680A0E002A9400803A884B5B5206B7C2E53CA25144009007A64EBD64",
INIT_09 => X"41008810240240C6694008010392354010000560141801002028A83D2A08E06D",
INIT_0A => X"34000000848BCA6902A29C54539C020E11810098D4067EFF9FF284D483E2AB41",
INIT_0B => X"500001840000C80B410014088040F4A944B1AA313C0022AA0011C0DC00028001",
INIT_0C => X"80B14004D158C8CA24A1C2A870AA1C2A870AA1C2A870AA1C2A872550E1543800",
INIT_0D => X"80A14050A01509E050854498B5281A1C34E506A2C6898B52A154DAC6B6000850",
INIT_0E => X"0B03001A483A4146603050080410089180008800143D83888281A2034A850142",
INIT_0F => X"A4160600349075238473F1210006133835E92273612B3482C090068A0E84AC56",
INIT_10 => X"30060181BA1B13959DC08DA902458870201970B29602562B0581200D141D0959",
INIT_11 => X"E042021C040D0152C8058B3840F044708E7E1C20A0106EA166C13AFC14AA3804",
INIT_12 => X"080E004B0C17C1439A9838301DC1A8438EA32C009DC1A8255300650458A1D588",
INIT_13 => X"018010E186F110A908E3A8CB0026C9A610A908E6A60F0807626610E160589C4C",
INIT_14 => X"2A701667334005800B1605F043858125E0D04110408D2485CA034681E43A1E40",
INIT_15 => X"00646002304244A91102C93A2D608D2A258DF8034188200C050171A41108F084",
INIT_16 => X"110441104411044110441104411044110466C440446CA06951D4EA8010009804",
INIT_17 => X"0040100401004411044110441104411044110441104411044110441104411044",
INIT_18 => X"0401004010040100401004010040100401004010040100401004010040100401",
INIT_19 => X"F7DFBFDEFE8FF1F7DEBDDF7DF7D05122890000000003FFFFFFFF900401004010",
INIT_1A => X"9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7BFFDFD7DDDF7DF7D",
INIT_1B => X"F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE79E7",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000003F9FCFE7F3F9FCFE7F3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA000400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0800",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000002000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2A954BA000015400FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080402010FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2A954BA0004154BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A0004174BAFFFFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0800154AAFFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF552A974AA0000174BAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974A",
INIT_2E => X"000007FFFFFFFFFFFFFFFFFFFFFFEF552E974BA0804000AAA2FFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080400010000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E954AA080005000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000402010FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2A954BA000417410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"804154BAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974BA0000174AAFFFFFFFFFFF",
INIT_34 => X"FFFFFFFEF552A974AA0000104AAE3FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0",
INIT_35 => X"AA2FFFFFFFFFFFFFFFFFFFFFFFEF552E954BA000E124BAE3FFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000007FFFFFFFFFFFFFFFFFFFFDFEF552E954BA080A000A",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804000100000000000000000000000000",
INIT_38 => X"54AA000400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2A954AA080017410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"0174BAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A954BA000415400FFFFFFFFFFFFF",
INIT_3B => X"FFFDFEF552E974AA0804174AAF7FFFFFFFFFFFFFFFFFFFFFFFEF552A974BA000",
INIT_3C => X"2FFFFFFFFFFFFFFFFFFFFFDFEF552E954AA0004000AAA2FFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2A954BA082E800AAAAFFFFFFFFFFFFFFFFFFFBFDFEF5D2E954BA002A820BAA",
INIT_3E => X"0000000000000000000000000000000000000087FFFFFFFFFFFFFFFF7FBFDFEF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(22),        -- Port A data input
DOA(0)   => data_read_a_lo(22),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(22),        -- Port B data input
DOB(0)   => data_read_b_lo(22),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_23_16 : RAMB16_S1_S1
generic map (
INIT_00 => X"EF20906D902424807BC8241BC81801B97D38AD3C0800103362A6741C80A12A02",
INIT_01 => X"001FFF8409F089003B4422000D80C80106804A7951C5B9D1C828043EA28838F9",
INIT_02 => X"E01CEE21649C82C40800000F9FFEFF8E72CA7F5FC2E22809925A0D3611C877F8",
INIT_03 => X"24000400402670400402670D48222DC1764446838624000080007460C40001BF",
INIT_04 => X"68403FFC020560E0443E21037C01FFFC0002EE00628BF0E02FAD781014085014",
INIT_05 => X"0112000202FBFFF00920017FF0F0628BFF8488890979800002F702002BB807A0",
INIT_06 => X"EF85788B681FC000000001FFF0010000000001F7CBC385F87C0BFFFF20040001",
INIT_07 => X"F6E200000000C1440E3AE408009120071070FA07A1CB23FFA403F0C4D23BF7C0",
INIT_08 => X"0BF87CA400804000003FF7FFD8880A034AC09662305AB10555421006891A1089",
INIT_09 => X"BE1F5FEA10092C0896A243FFC0008087FFBEF2000000001DFFC612C0C0400100",
INIT_0A => X"41FF0C2060501000600000000001BFFA800808189A657EF81DD0C00079CC8001",
INIT_0B => X"018C24110A860006C620C0312241C482B20400CC52492710CC80060020A81BFE",
INIT_0C => X"0C08866907048320C20C10030400C10030400C10030400C10030400608018210",
INIT_0D => X"040002000041500300100040000500C000801000C02400000952800001FFBF04",
INIT_0E => X"FC850015385380380CDB86106502C5043FFD5FFF00A04BC010A7724B10000800",
INIT_0F => X"89F90A002A70A710A51C01C05904014861433602A1CAF13F2110055614C72FC0",
INIT_10 => X"E02D02001C1E14981B43253EE50C8220180F1082E06397E07E42200AAC298E57",
INIT_11 => X"8421802400A90022B0070FAE18019214A380344920080B21A58B02AC60BACDF0",
INIT_12 => X"0A2A000C480B0704B54028101AC49C84BB4100009AC49C80857A82D20CE8CB22",
INIT_13 => X"01E00C8103416445C12ED0400027C5292445C12D500B0005A62D344CB241D095",
INIT_14 => X"132C907425604680038706A35132C94BDD011010404428886AC91B11311C8280",
INIT_15 => X"FF000470BE0692020328CA0028042054A92771C50FC070110001C1680809591D",
INIT_16 => X"00802008020080200802008020080200800800200200000000000008004807DF",
INIT_17 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_18 => X"8020080200802008020080200802008020080200802008020080200802008020",
INIT_19 => X"0000000000000000000000000000000000000000000000000000008020080200",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080002010FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974AA000400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000400010FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974AA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080000010FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E954AA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954A",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA000015400FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080002010FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974AA000400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000402010FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E954AA080005000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA080407000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA00041741",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080000010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000402010FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2A954AA080002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954AA080017410FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"552A954BA000415400F7FFFFFFFFFFFFFFFFFFFFFFFFF552A954BA080015410F",
INIT_3E => X"0000000000000000000000000000000000000F7FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(23),        -- Port A data input
DOA(0)   => data_read_a_lo(23),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(23),        -- Port B data input
DOB(0)   => data_read_b_lo(23),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_24_16 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100600007FFF000080108004000800020000840041000080808",
INIT_02 => X"FC5CA803400EB8209000000F9FFEFF8E7240FF1FC22409EA04018E50074017F0",
INIT_03 => X"11100400000000400000000D00002CC07400000090C080019001010A000001BF",
INIT_04 => X"68003FFC00040000000000008001FFFC0002EE00000370E007A100000000E468",
INIT_05 => X"0000000000F8BFF00920004DF0F00001DF8000000079800000F3000029980780",
INIT_06 => X"6E461803081FC000000001FFF0000000000001F7C3C380F87C019FFF00000000",
INIT_07 => X"600C2400013649609C8000980040814210254000A00B21FF2003F2A80D500000",
INIT_08 => X"0BF80000000000000003F7FFD88D2B4A02C0940062EC2804001610020408178B",
INIT_09 => X"8E1F5FE010092C0892A041FFC0000001FFBEF0000000001DFFC002C000000000",
INIT_0A => X"41FF0C0000000000600000000001BFFA0000005501AA00000CE2000009400000",
INIT_0B => X"018C0411020600048620C030020502000200000400490510CC00040020201BF4",
INIT_0C => X"0808064106040300C00C10030400C10030400C10030400C10030400608018210",
INIT_0D => X"0000000000004003000000000000001200580000000000000000000001FFBE00",
INIT_0E => X"0086C022005381380FDB96516140C6043FFD5BFF000041000000004110000000",
INIT_0F => X"80010D804400A7240C840C201D0210840043B4804012500021E0088014C04940",
INIT_10 => X"4109038041021C980200D06410C1924030008142E06024A00043C01100298092",
INIT_11 => X"587CC200002100C14428090A1D02348190814C09C010104025AA40041A0D8005",
INIT_12 => X"022E0030300B0E46177004208000D8C61D7004300000D884817B00011306B2D9",
INIT_13 => X"01E003060344710009875C018100013831000985DC000C20003C310006143B70",
INIT_14 => X"4001850EDC004780144806A64400186CBF8961104000C3807884000846EB9500",
INIT_15 => X"FF0006E08C063C0220002201490418082010A57263E0100008000290161E711C",
INIT_16 => X"00000000000000000000000000000000000000000000000000000000000007DF",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"F2D0AEEAF6E7CC1132CDB4441990000000000000000000000000000000000000",
INIT_1A => X"BEFBE79E79E79E79E79EFBEFBEFBEFBEFBEF9EF9EF9EF9EFA69861219575D75F",
INIT_1B => X"783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1EFBEF",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000783C1E0F0783C1E0F0",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0201000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A000400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA000400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000400000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402010000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"00002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080002010FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000400010FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA00040000",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020100000000000000000000000000",
INIT_38 => X"74BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"000010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA000002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974AA000402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000002010F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(24),        -- Port A data input
DOA(0)   => data_read_a_lo(24),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(24),        -- Port B data input
DOB(0)   => data_read_b_lo(24),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_25_16 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100200002000000080100004000000020000800041000080808",
INIT_02 => X"FC400086000000800000000F9FFEFF8E738FFF1FC204010000000111568DD7F8",
INIT_03 => X"00000400000000400000000D00002CC4740000008000000080000000000001BF",
INIT_04 => X"68003FFF64A564AC000000000001FFFE0082EF00010370E007A1000000004000",
INIT_05 => X"0A00040148F8BFF80920804DF0F00101DFC040000079C92484F30499299837C1",
INIT_06 => X"66041803081FC0E0801101FFFD000E41002299F7E3C380F87C019FFF81200096",
INIT_07 => X"000000080480AE00000080000000000000000000A00B21FF2003E00000000000",
INIT_08 => X"1BF80000400A02000003F7FFFA0008000200A0400008A0000014100200081000",
INIT_09 => X"8E1F5FFA53EFBCACB2E369FFE0010001FFBEF80C40630C7DFFEEBAF000800202",
INIT_0A => X"41FF0C0600000000600000000001BFFE00301000000000000CC020000140000C",
INIT_0B => X"01DCCC31222730A49620C030020100000200000400490D10EC00040220201BF4",
INIT_0C => X"0808064106240300C00C10030400C10030400C10030400C10030400608018210",
INIT_0D => X"0883044582114013412080000000000000000000000000000012800001FFBE00",
INIT_0E => X"00040020000180380FC386106140C6043FFD5BFF00A04B80608003CB120C1106",
INIT_0F => X"0000080040000200040400000100000000009480000240000100080000400900",
INIT_10 => X"0001000000000808000000240000020000000100006004800002001000008012",
INIT_11 => X"0001001808220000002004001900000080800008000000000022400000088000",
INIT_12 => X"0010000000000E00110000000000408009000000000040808063004000008200",
INIT_13 => X"6000000000046100000240000000001021000004400000000010210000001010",
INIT_14 => X"4000000404000800000000060400000088000001800000001084000000088000",
INIT_15 => X"FF800C608C041002000002000006100000002100000000180600000000100018",
INIT_16 => X"4110441104411044110441104411044510629041040D180400000010028047DF",
INIT_17 => X"1104411044110441104411044110441104411044110441104411044110441104",
INIT_18 => X"1044110441104411044110441104411044110441104411044110441104411044",
INIT_19 => X"FBA2894A196A8C5A2932EC15DA080800002FFFFFFFFFFFFFFFFFC11044110441",
INIT_1A => X"2492492492492492492410410410410410410492410492412000531215A69A6B",
INIT_1B => X"158AC562B158AC562B158AC562B158AC562B1588C46231188C46231188C49249",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000B158AC562B158AC562B",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080000010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000010FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08000000",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(25),        -- Port A data input
DOA(0)   => data_read_a_lo(25),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(25),        -- Port B data input
DOB(0)   => data_read_b_lo(25),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_26_16 : RAMB16_S1_S1
generic map (
INIT_00 => X"E9264EAB20190CA3BA4997AA9002AE9C001006B0778015CFA17E0811039879C7",
INIT_01 => X"2FFFF9BB1F773C7F9BB07DFFFDD863FC5FFF3FEFFBBF9FFB22FFFBC7B9F30686",
INIT_02 => X"E06CCC62052E708180F6FFBFFFFCFFFFF9C7FF7FC24332E642090000074037F6",
INIT_03 => X"428003739CD9863739CD9869FE2B7DEAF300029E4E300DFE69A6E644E6FF473F",
INIT_04 => X"7C2FEFFFF5BA124F003DD31EAFFFFFEE9FF7EE6F4C0770FFD7DC7CA53997B2B1",
INIT_05 => X"DFFB5421C1F8BBFAFDBFFACDF0FFCC05DDDBFF3690F9EDB7F5F7AFF639BD7DE3",
INIT_06 => X"EFD044ABC817C3E3A74667FDFFB6FF5727CC3BFEF7C3FAF87FF59F7FFBFEF69F",
INIT_07 => X"00003002132462052E708180EF060C18E5BEFB051225CDFF7002C4EEDE77F6E0",
INIT_08 => X"3FFF7D5000EC75088ED3FF7FC8790E46426CE06CB1F8E041051831FA3068D77E",
INIT_09 => X"C05FD7FF9BEFBDCEFBEE59FEF44F6603EFBEFAFCC2E35E7FDFD147CCF3F583FA",
INIT_0A => X"67FF1C7FBFADEB31E35768E8ED6BFDF3EB3EBF9DDBCE7FDC1DF8A760F3EACC02",
INIT_0B => X"5BDDCC3B336F7C548667D47B7737AF3FD62601EDC25B3533DCEB07F262213FFC",
INIT_0C => X"5F9A06E19F4D93A0EA0F78C35E30D78C35E30D78C35E30D78C35E986BC61AE31",
INIT_0D => X"5FD7AFEFDFFAF59B6FF28FE1D80D73D840607307DCFE1D80EF69A004DFFFF7FF",
INIT_0E => X"0004001F8041897B2FFFC6D86D70CE04FFFFF3FF1F5F5475BD7F72E4D75EBFAF",
INIT_0F => X"F60008003F008237B0040A00010003E020023E0201F45EC0010007E01047D17B",
INIT_10 => X"00010001DC0004C81003DE050A700200001DC0006863E8BD8002000FC0208FA2",
INIT_11 => X"2200E400002801E1A00004C21C0206F60081800800007B00010F02007EC09A0E",
INIT_12 => X"0880007E000807C7C1A612001E0015C7C19C22001E0015C59DFE82011A311AA0",
INIT_13 => X"00001BC00101F60409F0670840070809760409F06984800780097604067D0010",
INIT_14 => X"81019F40042100001F800203D81019EC085614000085C80023D81009CF008A74",
INIT_15 => X"FF802FFDFFAFD082003B032FB987E04021D481D4000819060801E0D00001231D",
INIT_16 => X"EBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEFFBFBFBFBBFCFBB0FFDFEFFEF2DFFFFFB",
INIT_17 => X"BFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAF",
INIT_18 => X"FAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFE",
INIT_19 => X"475B15BCF491E166CC8553F86EDB5C88646FFFFFFFFFFFFFFFFFEBFAFEBFAFEB",
INIT_1A => X"861861861861861861861861861861861861869A69A61861AFBD54D5F871C71D",
INIT_1B => X"984C26130984C26130984C26130984C26130984C26130984C26130984C261861",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000984C26130984C26130",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040201",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(26),        -- Port A data input
DOA(0)   => data_read_a_lo(26),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(26),        -- Port B data input
DOB(0)   => data_read_b_lo(26),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_27_16 : RAMB16_S1_S1
generic map (
INIT_00 => X"00080A40000A41248002029000050A088000008242A0004404480002000A1155",
INIT_01 => X"2FFFF1C11F781C129C107DFFFE0860941E81258CA2B71C2220EC1B86E1A00002",
INIT_02 => X"E1000000810000014400FF6FFFF0FFFFF8007F1FC21110005080200000221FF0",
INIT_03 => X"4080026318C18226318C1821302232EAE00002BE001115FE48620040840A863F",
INIT_04 => X"643D4FFC2530000F003D821C0BFFFF8E9EF79E6D440748FED70060842105B0B0",
INIT_05 => X"D6F39020D1F8A3FAFDBFBACDC8FDC405D1DB7F1490E5EDB7D5CBADB2385D79C3",
INIT_06 => X"6FE000A38007C3032646EFF1F0B6FF46A78C39F8E723F2E47FE59C7F9ADA2612",
INIT_07 => X"00002820000000810000014401060C180190310540118DFF1000C0849673F6C0",
INIT_08 => X"3FF779100062B12A8EC3F47FC80208808210880C00082050000110023068D030",
INIT_09 => X"005F07E09BFFBD07FBAC09F8E42922038F7DF8BEC2E39C5F1FD047CEF1B582D8",
INIT_0A => X"63FF5D5F9FADE911E81C09818109E1F16B16B71092CE7ED81CF403601228C402",
INIT_0B => X"1BFDCC39732F3554866AD57C37BEAF1C152201A4C05B7531D56B05B06A213FF8",
INIT_0C => X"5BCA06F18FC59380F00E34430D10C34430D10C34430D10C34430F0861A2186B5",
INIT_0D => X"5B56ADAB5FAAE58B2F628EA0C80FA3F04040510768EA0C80CC61A0044DFFC6EB",
INIT_0E => X"0004001D800188792CE79715710AE4047FFD23FF315D54358D593474955AB6AD",
INIT_0F => X"520008003B000297B0040200010003E020001F0201E44A400100076000579129",
INIT_10 => X"00010001DC00004A10035E0408300200001DC000086BC8948002000EC000AF22",
INIT_11 => X"02002400002801E1A00000C01E0202F60080800800007B00000782006EC0820A",
INIT_12 => X"0080007E000006A7C10602001E0001A7C10C02001E0001C18DE282010A311AA0",
INIT_13 => X"00001BC00000FE0401F04300400708007E0401F04180800780007E04047D0010",
INIT_14 => X"81011F40040100001F800002F81011EC080604000085C80001F810094F008034",
INIT_15 => X"FF800C6DDDAFD082001B03249887E04001D481D4000009020801E0D00001021F",
INIT_16 => X"AB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6BF1EBDABD8E270BF84A25C6ACB777E3",
INIT_17 => X"B6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6AD",
INIT_18 => X"6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADA",
INIT_19 => X"490E2168100481CA860402104A471688747FFFFFFFFFFFFFFFFFAB6ADAB6ADAB",
INIT_1A => X"000000000000000000000000000000000008200000000000200072F210000001",
INIT_1B => X"05028140A05028140A05028140A05028140A0500804020100804020100800000",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000A05028140A05028140A",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040201",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(27),        -- Port A data input
DOA(0)   => data_read_a_lo(27),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(27),        -- Port B data input
DOB(0)   => data_read_b_lo(27),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_28_16 : RAMB16_S1_S1
generic map (
INIT_00 => X"02200AA400180030808802A900002A08001280A08A801044104A1000001818C3",
INIT_01 => X"0AA00011460214428114180000882214413D0A71592A01D92213D28005210202",
INIT_02 => X"0451110A012100884000AA30200000000C100040104112101100008888200000",
INIT_03 => X"448000318C52A20318C52A20148810200111100C211004AA00034204200A2200",
INIT_04 => X"04004001001A90110000121402AA0000003C00000500000040080421080D0080",
INIT_05 => X"4060000C8001000000002E000000050000001610300000010000802202040012",
INIT_06 => X"1000002080001111001222000425A1040026A008000000000000000009328280",
INIT_07 => X"2491008A00491201210088400122448908A20402000408001000040820000000",
INIT_08 => X"20058310402A160026500000028040101004200C840082115554000112244814",
INIT_09 => X"4140000800000060000720000102028000000490160801020002200011100010",
INIT_0A => X"020000081B34211082B694D4D294000020020381040000000200032040004400",
INIT_0B => X"4800210C19808400500010009110091500020B408810000100200020408B0000",
INIT_0C => X"01028000080118020023604858121604858121604858121604858090B0242C00",
INIT_0D => X"010000800920040804020A6058003108402043058C460580653020005A004039",
INIT_0E => X"00000002800008014004104104420A00C000200005000010040A0020CC000200",
INIT_0F => X"520000000500000010000200000000000000280000040A40000000A000001029",
INIT_10 => X"00000000000000C0000002000830000000000000480008148000000140000020",
INIT_11 => X"020024000000000000000440000000020000800000000000000C00000040020A",
INIT_12 => X"00800000000001804006020000000500400C0200000005400A90000000100000",
INIT_13 => X"0000000000018200001003004000000142000010018080000001420000200000",
INIT_14 => X"8000080000010000000000018800008000060400000000000310000008000034",
INIT_15 => X"000002040080000000110006B081400000400000000009020000000000002200",
INIT_16 => X"802008020080200802008020080200802101210810C39A66A90A85420413A820",
INIT_17 => X"0200802008020080200802008020080200802008020080200802008020080200",
INIT_18 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_19 => X"DE21102C110A00246972BD89A40A0C22E1000000000000000000002008020080",
INIT_1A => X"2082082082082082082082082082082082082082082082080D35050758C30C31",
INIT_1B => X"0582C160B0582C160B0582C160B0582C160B0580C06030180C06030180C08208",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000B0582C160B0582C160B",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(28),        -- Port A data input
DOA(0)   => data_read_a_lo(28),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(28),        -- Port B data input
DOB(0)   => data_read_b_lo(28),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_29_16 : RAMB16_S1_S1
generic map (
INIT_00 => X"79964E4BA01DACAB9E659792D00AAE160002829C7FDFEFCEE97C2815039D70C3",
INIT_01 => X"0ABFF9AB0775343F9AB01DF80D5821FC0FFF3FEFD1AF9FF1207FFBC7B9720586",
INIT_02 => X"002CCC60050E700080F6AAA7BFFC007189C7FF2FC00330E602800000074037F6",
INIT_03 => X"468003210868A63210868A68DA017D207200021C4E200CAA6186A40042FF4300",
INIT_04 => X"7C2FE002F0900001003C5316A6ABFFE21F36E02F0D03701F47D41800109FB281",
INIT_05 => X"4979440580F9B808F49F6A4DF00F8D01DC4B97369078249370F482E62BA41462",
INIT_06 => X"B250442BC81001E1870223FC0BF7F11507C423FE33C078F803F19F00E936721D",
INIT_07 => X"00011080012460050E700080EF020408EC8CFA01122149FF700200665A35D260",
INIT_08 => X"2BFD055040A452000443FF00007906464068406C31F84000000831FA1028575A",
INIT_09 => X"805FD017102690AA694551FE30444681E0820AD40201423FC00122C493500172",
INIT_0A => X"0600002AFFBE2330815568A8AD6ABC02A02A0B0CCB463B4C0748A720B1EA4C00",
INIT_0B => X"0850400A11414C005005000B51158936D20601A98A10200308A002E240010BFC",
INIT_0C => X"05928020194918A22A2268C81A32068C81A32068C81A32068C81A99034640C00",
INIT_0D => X"058102C48970541944B20FA1580561D040406305587A158046282000DBFFF13D",
INIT_0E => X"000000028040890327DCD28928324400DFFFF0001F1F0050342D42A086040B02",
INIT_0F => X"F60000000500802010000A000000000000022A0000141EC0000000A01000507B",
INIT_10 => X"00000000000004C0000082010A700000000000006800283D80000001402000A0",
INIT_11 => X"2200E4000000000000000442040004020001800000000000010D000010401A0E",
INIT_12 => X"08800000000801C040A6120000001540409C2200000015441DAC800010100000",
INIT_13 => X"0000000001019600081027084000000956000810298480000009560002200000",
INIT_14 => X"800088000021000000000201D800088000561400000000002358000088000A74",
INIT_15 => X"00802594A282C0000033010FB181E00020400000000819060000000000002305",
INIT_16 => X"C0B02C0B02C0B02C0B02C0B02C0B02C4B12B312912831A27FCFE7FFB175B6FF8",
INIT_17 => X"0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02",
INIT_18 => X"B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C",
INIT_19 => X"BBCF9F96EE7FFDF7FE783FFDFFEA0C00602FFFFFFFFFFFFFFFFFC0B02C0B02C0",
INIT_1A => X"EFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEEBAEBAEBAEBAEBBFFDF9FBEFFFFFFE",
INIT_1B => X"BFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFBEFB",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000FBFDFEFF7FBFDFEFF7F",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(29),        -- Port A data input
DOA(0)   => data_read_a_lo(29),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(29),        -- Port B data input
DOB(0)   => data_read_b_lo(29),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_30_16 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"F7FFBFFEFF9FE1F7FFBFFFFDFFD0000000000000000000000000000000000000",
INIT_1A => X"9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7AFBD75F5FDF7DF7F",
INIT_1B => X"F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE79E7",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000003F9FCFE7F3F9FCFE7F3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(30),        -- Port A data input
DOA(0)   => data_read_a_lo(30),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(30),        -- Port B data input
DOB(0)   => data_read_b_lo(30),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_31_16 : RAMB16_S1_S1
generic map (
INIT_00 => X"129000008004A00804A40000400800020000000C005FEA005800200400050100",
INIT_01 => X"255FF18019700810180065FFFC0040801E80258CA2951C2200EC0906A0804140",
INIT_02 => X"E0000000000000011000550FDFF0FFFFF0007F1FC200000044000000000817F0",
INIT_03 => X"0000024210A30024210A3001002220C06044469200040154482000408400043F",
INIT_04 => X"602D0FFC2420000E003D80080955FF8E1ECA8E2D400340FE870060842100B030",
INIT_05 => X"0213100040F8A3F8FDBF944DC0FDC001D1CB6904A061EDB6D4C30490281831C1",
INIT_06 => X"6FC000830007C202060445F1F0D25E4207A099F0E303F0E07FE19C7F80402412",
INIT_07 => X"0000200000000000000001100004081001103107000185FF0000C0849673F6C0",
INIT_08 => X"1BF27A00000000000883F47FC800080002008000000820440000100220489020",
INIT_09 => X"011F07E013EFBC06FBA009F8E00120038F3CF82C44630C5D1FC002CCE0808248",
INIT_0A => X"61FF0C06C48BC801600000000001A1F00110101092CE7ED81CF0004012288000",
INIT_0B => X"11DCCC31222730048620C4382204A608142002A440492530C401049020221BF8",
INIT_0C => X"0888066187448380E00C10030400C10030400C10030400C10030600608018210",
INIT_0D => X"080204010200418301208480800D02D00040100240A808008840800405FF8640",
INIT_0E => X"0004001D000180780CE386106100C4043FFD03FF101D40008001304018081004",
INIT_0F => X"000008003A000217A0040000010003E02000160201E040000100074000478100",
INIT_10 => X"00010001DC00000810035C0400000200001DC0000063C0800002000E80008F02",
INIT_11 => X"00000000002801E1A00000801C0202F40080000800007B00000302006E808000",
INIT_12 => X"0000007E00000607810000001E000087810000001E000081846282010A211AA0",
INIT_13 => X"00001BC00000740401E0400000070800340401E04000000780003404045D0010",
INIT_14 => X"01011740040000001F8000025010116C080000000085C80000C8100947008000",
INIT_15 => X"FF800C609C06D082000A03200806A040019481D4000000000801E0D00001001D",
INIT_16 => X"010040100401004010040100401004010060C040040C200950402090128057C3",
INIT_17 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_18 => X"0040100401004010040100401004010040100401004010040100401004010040",
INIT_19 => X"00000000000000000000000000001000802FFFFFFFFFFFFFFFFF810040100401",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(31),        -- Port A data input
DOA(0)   => data_read_a_lo(31),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(31),        -- Port B data input
DOB(0)   => data_read_b_lo(31),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_0_15 : RAMB16_S1_S1
generic map (
INIT_00 => X"ED39BA795990D275FB4A6E96ACC4731DEA4598B0AFB54867F6EE4618C3749803",
INIT_01 => X"8AA0047D8607944AC7DA180001ECA2444042106208408208C20022E9173734B3",
INIT_02 => X"1A7DDD79F9A73E6CCA7DAAF00001000008478020113D98E382FEDF333027C80F",
INIT_03 => X"75D341110C58F31110C58F32A208921F8051500147A0E4AB3493FB3A01EBE240",
INIT_04 => X"86424001531009B100425A97B2AA0001E03501D0A39C8F0078420001106D0C4C",
INIT_05 => X"BCC8CA2EBF03400700402BB20F00239E20341699198600000B08694B16434804",
INIT_06 => X"103FB860B2800161F8432200012DA185F80F24081C3C0707800E600056881308",
INIT_07 => X"B24197ABCDA467F9A73E6CCAFDC3870EEEEC44E2BDFE220094D03022210C011C",
INIT_08 => X"240581B5695EAA80262C080032BF07C7C1FC3F8E94F65B11555EAFFC1C306758",
INIT_09 => X"7E40000BEC004170040DB60017FED1CC0001045002984202003DB931192D60A5",
INIT_0A => X"120071411A74315881A28C141118000C5A85A60444210123820B43B40804674D",
INIT_0B => X"0820008E514045BB514F0106D1D8599581D3A958BC104A89215AC14C48898403",
INIT_0C => X"C261C01C48B1584A0CA3E2687A9A1E2687A9A1E2687A9A1E26870CD061343885",
INIT_0D => X"D274E93A758FA8683AC54B287522E10A74AF4AA59C568752662F5AC218000002",
INIT_0E => X"FF83C002783A0904231C70470C7E0B92800224008AE09FAD4BD48D1FC5D3A4E9",
INIT_0F => X"5BFF078004F075885DFBF7E15C06101C55E921F1F80FAB7FE0F0009E0E903EAD",
INIT_10 => X"F12E0380231F13978FF023FAFDBD9870380230F2D6081F56FFC1E0013C1D207D",
INIT_11 => X"DE7F263C0C8700125C0F8F3C43F1F10BBF7EFC61E01804E1E6C8F8FE807F67FB",
INIT_12 => X"02BE00017C17C1007E5E2E3081C5AC007E6F0E3081C5AC44418D65FE45DEE55B",
INIT_13 => X"61E0042786F103E9F01F9BC3C120C5A703E9F01F978B8C20666703E9F8A0FFED",
INIT_14 => X"FA7E283FFB414F80005F05F10FA7E283F78F6511C048278DCA174FF038FF15B4",
INIT_15 => X"0066A20B61692F293185D8D724E15D3FCC6B7C236FE0691B0700132C1F0EF880",
INIT_16 => X"3A4E93A4E93A4E93A4E93A4E93A4E93A4F942F92E9628540AD2A91442525A000",
INIT_17 => X"A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E9",
INIT_18 => X"4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93",
INIT_19 => X"55F3898E09B56C74DAB15D1CF13501AA495000000000000000003A4E93A4E93A",
INIT_1A => X"082082082082082082082082082082082082082082082082082084E41DC71C71",
INIT_1B => X"E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F82082",
INIT_1C => X"FFFFFFFFFFFFFFF94A5294A5294A5294A5294A52800003E1F0F87C3E1F0F87C3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"3060C183060C187FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"BDEBA0000000000000000000000000000000000000000000003060C183060C18",
INIT_28 => X"168ABA002E82145085155545F7AA975EFFFAABDE00FFAEBDFFF5D2EAAAAAF7AE",
INIT_29 => X"7FFFE10005542145557FD5545FF8000155087FC0155F7D168B55007BFDF45085",
INIT_2A => X"7FFC0010080017555555568AAAFFFFD7545AA8028A00A2802AABAFF8028BEF5D",
INIT_2B => X"FF842AABAA2AE95545FFD168ABAF7AEAAAAAA2FFFDF4500043FE105D2E954BAF",
INIT_2C => X"5007FD7400550415410002E974BA5D5168A00A2D142155005142010FFAE820AA",
INIT_2D => X"FFF780000BA007FE8AAAFF803FFFF5D2A821550000000BA007FD55FF5D7FC014",
INIT_2E => X"000AAFBEAA00007BFDFFF082EBDF455D5142000082E82145FFD17DFEFFFD168B",
INIT_2F => X"DFD75D2AA8A80EA8E2FE3F000000000000000000000000000000000000000000",
INIT_30 => X"68B551475FAF6D1C556F0AA1C24AABEA495FC716F002A975FFE3AA95E00EBAEB",
INIT_31 => X"42A0070071C50BAFEF1FAE0016D56A16D557BC257D415E0216FA3F1E8FC0145B",
INIT_32 => X"8010E004924874825D7FEAA85487FD24AFE3D02DAAAE12BD5545A2803AA00005",
INIT_33 => X"120155EA568E870BAEB8A05A2AEA8B50F55A2F150005A3A438BD04AFAB8F550A",
INIT_34 => X"545E055FFBE81D0BE8EA8A3AA05A2A5504001C74BA42A1571E8028E3DB7816D0",
INIT_35 => X"A5C7E3DFFFE90B45B47ABA497A82FFAFD2A82485FD2415A105C21451ED42A002",
INIT_36 => X"00000000000000000000B55EAAA100AA1D0F6F480B6A555A2A57A002A3D5FDB6",
INIT_37 => X"5EFAAAAB5E1AF3AABFF45592E88A0AFE80A8B0A0000000000000000000000000",
INIT_38 => X"65F520EBE9EF67D7BEA1FD5D556ABEF5D557FEBA55022A3F70C6B405F4D2AE97",
INIT_39 => X"C114728007521170821CE0FDE69411A8DED57CE1055555E5F58EFFC01FE2CACB",
INIT_3A => X"42341D5DEEBEF55080034E0A592A4AD0079C75D6070CC5CBB0280C029ABAA3EB",
INIT_3B => X"7F353AAF6C77F7F20D968BF57812A95E02A2AAB5EB0F280800EFAEE9F5D18F31",
INIT_3C => X"C91565455C141E41887D58AC448B69C30E02116220415A9540AA854140A0A204",
INIT_3D => X"DE6BE93172D7D625B556EEAB157ABEBE1B4D792A4AD1183454180DD3FDCAAAB7",
INIT_3E => X"F0000001FF0000001FF0000001FF0000001FF01EABC4B8014174FF7DA80F52FE",
INIT_3F => X"FF0000001FF0000001FF0000001FF0000001FF0000001FF0000001FF0000001F")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(0),        -- Port A data input
DOA(0)   => data_read_a_hi(0),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(0),        -- Port B data input
DOB(0)   => data_read_b_hi(0),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_1_15 : RAMB16_S1_S1
generic map (
INIT_00 => X"212C001411984004084D000508C53810A03D1450E839B003342114428A000803",
INIT_01 => X"00000019400B100A8196000000CC004400400002000000000000028001340000",
INIT_02 => X"052137AE8031800C0044009000000000061800001CD4019802AD04CCCFC20004",
INIT_03 => X"04514108C60C21008C6042108400000201440020505100000043C30E10E9F000",
INIT_04 => X"02104001011DEFE088805681920000008000004001900800004002108C280008",
INIT_05 => X"040002340105000200000000080001900010000108040000000008411600401C",
INIT_06 => X"1034001042800808201000000001000820020000102000040000000000800180",
INIT_07 => X"64BF81A15EDFDE8031800C00843060C19E030022103600000450020800040004",
INIT_08 => X"00008004691687AA840008000090248CC84E000046000311555521F183060AC5",
INIT_09 => X"0820800D08100171000DB000154440C800400500000852020011200201012021",
INIT_0A => X"02000040001000880A2A04445004000102002041000001008208001440004140",
INIT_0B => X"4820018A1140440078050040511000102000A008183000010002404400000000",
INIT_0C => X"1000C80008000C030030880C2A030A00C28030A80C2A030A00C28018D4061401",
INIT_0D => X"10040802050080200284401C0022880F009E08008205C0020118088018000000",
INIT_0E => X"0F03C00280000000420860C60C0C0B92C0000000004000010042000040102008",
INIT_0F => X"001E078005000108400005E11C0610000000288058000003C0F000A000100000",
INIT_10 => X"F10E0380000000C202300000008D187038000000480800000781E00140002000",
INIT_11 => X"806302380C870010000004400100110800007861E0180000000C400680000001",
INIT_12 => X"023E00000000018000580C308000050000610C30800005000215006800000101",
INIT_13 => X"61E0000000018100B0001843812000014100B00016030C20000141002880026D",
INIT_14 => X"400A20009B404F80000000018400A20044096111C04000000304026000501580",
INIT_15 => X"0046820040082300218450C2800010094000482141E060190700100000002200",
INIT_16 => X"020080200802008020080200802008020080008008600500A82A1100A8000000",
INIT_17 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_18 => X"0080200802008020080200802008020080200802008020080200802008020080",
INIT_19 => X"81328A46BABEFC54A0810C7452B4428A14000000000000000000020080200802",
INIT_1A => X"AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA28A28A28A28A2A8218D2C0C924925",
INIT_1B => X"E974BA5D2E974BA5D2E974BA5D2E974BA5D2E975BADD6EB75BADD6EB75BAAAAA",
INIT_1C => X"FFFFFFFFFFFFFFFD8C6318C6318C6318C6318C63000002E974BA5D2E974BA5D2",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"70E1C3870E1C387FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"5555500000000000000000000000000000000000000000000070E1C3870E1C38",
INIT_28 => X"EBDF455D2EAABEFF7FFE8BFF5D0002155557FFFFFF007FC21EFA2FFD74AAAAD5",
INIT_29 => X"AA95400552AAAABAFFD1574105D7FD75FFAAAA800AAF7AA974BAFFFBE8B45F7A",
INIT_2A => X"0517DF555D2EAAA1055000015500557DF45AAD1400BAA2AE801550051555EFF7",
INIT_2B => X"FFD540155557FD5400F78028BFFFFFBEAB55F780020AAAA80020AA082EAAB550",
INIT_2C => X"AFF842ABEF5D517DF55552A974AAF7AE820AA0851574BAA2D1574AA5D7BFDEBA",
INIT_2D => X"EFAAD1575EF557FFFE10557FFFFFFFFD56AAAAFFFFD7555AAD168B45AAAEAAAB",
INIT_2E => X"0005D7FFDF4500043FE105D2E954BAF7AE80010082A97410557FEABFFAAFBE8B",
INIT_2F => X"51C7A2FBD5490BFD1C056A000000000000000000000000000000000000000000",
INIT_30 => X"974BAF7FFEFB45FFAABDF55492AA8BC2EBDFEAF7F1F840017D4975D2FEF147FC",
INIT_31 => X"080BEF495FC71D54124924385FAAA8AAAE3D145410F7F1D55D71C002DABAEBAA",
INIT_32 => X"002D082082AB8B6DBEDB7DF7F540E2AE85028B40155145F7AF6DBED5450AA1C2",
INIT_33 => X"78E021FF1471FDEAAFFD56F16D5571D2E28E38E0216FA2D1E8E80140F45082B4",
INIT_34 => X"A2DA3FB7DAAD4AAAAF487BC70BFA97F7AF6D417E92482BF84020BA495557E3FF",
INIT_35 => X"55554ADBD7A2FFC7BEFF6FFD7FC7002FD74951D71EDFFABFD16FAAAE92BD5545",
INIT_36 => X"00000000000000000000547AB8F550A8010E00492487482FFFE82A85EBAE2FFC",
INIT_37 => X"1EF005162BEF047FD5545AAFBF7400FBF9424F70000000000000000000000000",
INIT_38 => X"714F8338AAAA1D0AE974AAF7FFFDF55F7AABFF55082CA8B4DF6C1E8F5E540002",
INIT_39 => X"EABEF75550ACBB7582225FF5843404547184164AA5D2EBEEB0A2D555410D3555",
INIT_3A => X"FEAAEB083BC1000FF8409000512AEABFFDF79DCBF755962010BDCBBC21455D7F",
INIT_3B => X"801F8BA0C57740BDAA0688E5405D57D412F7D55F5E50C7F401BAAE8403CF5A3F",
INIT_3C => X"5D16BABAA3EBC3157ABD5FFE55F2AA9FEAFDF7F431A9F7FFE81FF013A8001AFF",
INIT_3D => X"FB863550229BCABEB7DA403FFFDA2FBF7FED2C7F955445079E280A00C56145EF",
INIT_3E => X"0000000000000000000000000000000000000596EBEF55080034E0A592A4AD00",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(1),        -- Port A data input
DOA(0)   => data_read_a_hi(1),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(1),        -- Port B data input
DOB(0)   => data_read_b_hi(1),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_2_15 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10E006600180111284380310006289800480032283E000A34301002001A0817",
INIT_01 => X"0005A00810790848048044A54E404350404000720885800802000906E4910200",
INIT_02 => X"407004208400408044C600C50AA055254010541A110222841200000002402544",
INIT_03 => X"0600011004182401004102408C28414043101000408118000145840440F5C415",
INIT_04 => X"5035855703A2900A000CD3088400F40688C9844409060850925E58A4081A0221",
INIT_05 => X"0200840D1021A15AC50494894850890540D1E12020C6E510818500440A280090",
INIT_06 => X"113044094002801020440090A8011A1224AB9380552102442884882A20004097",
INIT_07 => X"000100880004428400408044860000008C022402102100AA40004404B5075460",
INIT_08 => X"15C23440408C862A2A12382A8A5244145048C06085008010141521F000001240",
INIT_09 => X"400582B9033AA0E7AA4110B0506744810554542450694E710A836188C2C00222",
INIT_0A => X"443518360012C2210B020414109130A28038188096A06B8C120CA440A9C00802",
INIT_0B => X"1345E53300EC68005605002964AF222A5704004D080211121C80024200821780",
INIT_0C => X"181080C1110C882202211488452213C88472213C88472213488441109A442231",
INIT_0D => X"008204440210091341208041000810C00000300220201800A908000038AD0284",
INIT_0E => X"00040002804180300E88D28D206A40000554815500481440300000C44A081100",
INIT_0F => X"000008000500828700000000010000000002380000A00000010000A010050000",
INIT_10 => X"00010000000004CA000214000000020000000000684280000002000140200500",
INIT_11 => X"000000000020000000000442100002840000000800000000010C000026000000",
INIT_12 => X"00000000000805A4800000000000152300000000000015801272000100210020",
INIT_13 => X"000000000101C00000C000000000000940000120000000000009600004050000",
INIT_14 => X"0000130000000000000002018000106000000000000000002380000141000000",
INIT_15 => X"55000190000000000002000280000000011080C0000000000000000000002310",
INIT_16 => X"40902409064190641906419024090244902A9003004800415120D4A190804241",
INIT_17 => X"0900409004090641906419064190240902409024090641906419064190240902",
INIT_18 => X"9044090040900409004190441904419044090040900409004190441904419044",
INIT_19 => X"75960040138D70C030B51C50C7D100A2052F81F81F83F03F03F0419044190441",
INIT_1A => X"0410410410410410410410410410410410410410410410410248602081659659",
INIT_1B => X"5128944A25128944A25128944A25128944A25128944A25128944A25128941041",
INIT_1C => X"FFFFFFFFFFFFFFFE1084210842108421084210843FFF825128944A25128944A2",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"7FD5FF555815607FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"2AA000000000000000000000000000000000000000000000007FD5FF55581560",
INIT_28 => X"FC21EFA2FFD75EFAA8415410AA8415555087BFFF55A2AA800BAFFAE954000800",
INIT_29 => X"84155EFA2AEBDEAAA2FBEAABA5D7FE8B555551421455D0002145552EBFEBA007",
INIT_2A => X"2AEBDF555D2E954BAA2AA974BAFFFFE8B45552EBDF45FFAEAABFFF7FFE8B55F7",
INIT_2B => X"AAAAAAAAAFFD1574105D7FFFF555D2AAAAAA5D2E820BAA2FBEAB5555557DF55A",
INIT_2C => X"50055575EFFF84021555D043DEAA5D04021EF557FC21FFAA8428BFFAAAA954AA",
INIT_2D => X"10085568A00FF80175FFA2D17DFEFF7800215500557DF55AA80001FFAA800015",
INIT_2E => X"0005D00020AAAA80020AA082EAAB5500517DF555D042AA10A284154005D00154",
INIT_2F => X"00AAFFAA9543A080038A2A000000000000000000000000000000000000000000",
INIT_30 => X"0017D5D20B8EAA007FC51C7A2FBD55D2BE800042AFE8E1557D0075D2F45BEAA8",
INIT_31 => X"AA8BC7EBDFEAFEFFD00105FFBC20BDEAAA2FBF8AAA557BE8B6D5D5FFABEF4904",
INIT_32 => X"FFEFB6D555578F7DB6A0BDF7D480E174BFA02A974BAF7F5EFB455D2ABDF55492",
INIT_33 => X"ED1FDE90E3A497492B6AAADAAAE3D155E105571D55D71C002DABA5524820BAB6",
INIT_34 => X"BE8F401D7B6A0001470155C51D0092A071555D5E3AE821D00001FF0871C016DB",
INIT_35 => X"5BE8555400550A38428007FED000E3DA3DFD5E3DFFFBD5A38A021551C5F7AF6D",
INIT_36 => X"00000000000000000000410F45082B4002D082082AB8B6D1C5B7DF7FF78E075C",
INIT_37 => X"5EF005560B55F7AA800AAF7AA954AA00042AAA20000000000000000000000000",
INIT_38 => X"ABEF057D68F5F5A00021EF55042AAAA007FD5555AAFBD7545FBB8020A3F7AE97",
INIT_39 => X"7DF55D7AABFF5428ACA8F45A6C1E8F5EFF84165EFF7802BAB0A2FFEAABA557BE",
INIT_3A => X"CA8AA80800020AAF7FBFFFEF04552ABFFFF841FFE75CA882108202E974AAF7D5",
INIT_3B => X"00151FF0C57401E5F3D1E00A1A884174A8FFAEBFEB0A2D55541051555694F002",
INIT_3C => X"2AA801455D7FE8BFFF680800FFF7AAA155F595542455512A975455D3AA8A0055",
INIT_3D => X"5D79FCAF774AE005BE7895554005D2A8A0B882FFFFE10AAAAAB755A66B6AF56A",
INIT_3E => X"00000000000000000000000000000000000000C3BC1000FF8409000512AEABFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(2),        -- Port A data input
DOA(0)   => data_read_a_hi(2),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(2),        -- Port B data input
DOB(0)   => data_read_b_hi(2),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_3_15 : RAMB16_S1_S1
generic map (
INIT_00 => X"210C00A20020000108430020001600B8156021104940741B3530400E02B92203",
INIT_01 => X"014C9BCA58B1296D24A402C992500B69404040028804A0080A000416A8D90A08",
INIT_02 => X"C12026A484318004404405C9C66E331352180D468B8203980300204442E02B34",
INIT_03 => X"04000748D60D24648D60524C88804D0215011020D15018148040C10A70E1D58C",
INIT_04 => X"18283333240FE41244187308C9104D70944852640901083801750EB0A418C220",
INIT_05 => X"0613142D01912CC2A1B4140528348900C612A104201C689044340ED413A07649",
INIT_06 => X"119000034019881822104C5E68035250A222829710A0A02C18C01A9920842413",
INIT_07 => X"402F00AB0016CA0431800444841020509D038B021230C1990001C644C8273200",
INIT_08 => X"16905000408482088290E8E64010248C4A5AA840C2000110001521F0810A92E7",
INIT_09 => X"0003CE6581BD016342A951AB146C4480530C3B2A8088D3542651670200C1826A",
INIT_0A => X"00735D36209A8A20020894004284B660821030C8990467401218004041020002",
INIT_0B => X"512445B740457154562F957CC08B00093700080D0A4851001D8302D20A0A1530",
INIT_0C => X"00508650008008021021A40861021840869021A408610218C0869810D6043095",
INIT_0D => X"1C8508438450801043A08090380A8834207007022209038080190000999C8F84",
INIT_0E => X"000400200000C0002A48A206204C4205F3304B33004C0041006240140A1C310A",
INIT_0F => X"0000080040000083800400000100000000008400018040000100080000510100",
INIT_10 => X"0001000000000800000244040000020000000100002A0080000200100000A702",
INIT_11 => X"000000000020000000200000080002C000800008000000000022000006808000",
INIT_12 => X"0000000000000A2281000000000040A3810000000000402001400000022002A0",
INIT_13 => X"000000000004200001C0400000000010200001C0400000000010000004490010",
INIT_14 => X"0001070004000000000000060000104C08000000000000001000000903008000",
INIT_15 => X"CC004050CA0C00020220200070040000010401C4000000000000000000100008",
INIT_16 => X"4310E4310A4210A4210A4210A4210A4210A8D0830A68010001B4DA881048061C",
INIT_17 => X"21084290A4210A4210A4210A4210A4210A4210A4210E4310E4310E4310E4310E",
INIT_18 => X"90A421084290A421084390E4310C4390E4310C4390E4310C4290A421084290A4",
INIT_19 => X"015303C0C78C706428A14C586291000A044001FFE000003FFC004290A4210842",
INIT_1A => X"2492492492492492492492492492492492410410410410412821600001249249",
INIT_1B => X"51A8D46A351A8D46A351A8D46A351A8D46A351A9D4EA753A9D4EA753A9D49249",
INIT_1C => X"FFFFFFFFFFFFFFFC00000000000000000000000038F56351A8D46A351A8D46A3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"55AB02055AB0207FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"420000000000000000000000000000000000000000000000007FFFAB57FFFAB5",
INIT_28 => X"A800BAFFAE9554508002AA00AA843DF55FFAA955EFA2D168B55557BEAA000055",
INIT_29 => X"002AB55AAAA955EF005568A00087BE8BFFA2D155410AA8415555087BFFF55A2A",
INIT_2A => X"AAABFF5508003FF555D0002145552ABFEBA007FC21EF007FD75FFAA841541008",
INIT_2B => X"082EBDEAAA2FBEAABA5D7FC0155005168B455D042AB45F7FFD741000042AA10A",
INIT_2C => X"FF7FBEAB55F7AABDEBA5D7FC2010A2D1575FFF7AA975555D2E80145F78415545",
INIT_2D => X"EF5555554AA087BC01FFFFAAAAB55552A954BAFFFFE8B55552EBDE00F7AEAABF",
INIT_2E => X"000082E820BAA2FBEAB5555557DF55A2AEBDF555D2E954BA002EAAABA002A821",
INIT_2F => X"FB7D5D7FEAA3808554203A000000000000000000000000000000000000000000",
INIT_30 => X"1557D1475FAF45BEAA800AAFFAA95578080038A2AA28E3AF55E3A0BA5D7AADB6",
INIT_31 => X"BD55D7BE80004AA1E8E2AB55B6A0925D7085F6AA10087FEABD7AAD57AEBAB68E",
INIT_32 => X"F5D0438140E2FA38B6AEBFF6D1D04AAFFA41040017D5D20B8EAA007FC51C7A2F",
INIT_33 => X"D0A901FFFF801557D1C20B8EAAA2FBE80AA557BE8B6D5D5FFABEF49002FB55FF",
INIT_34 => X"5D20BDE00EBAAA8BC7EBDFEAFEFAB8ABAE925D21C7010EADB525D7FFAE975C75",
INIT_35 => X"F002EADA921420871D74971D24820875C21D5EB8AA8FFF012A954BAFFF5EFB45",
INIT_36 => X"000000000000000000001C24820BAB6FFEFB6D555578F7DB6A0BDF7DEB8E125F",
INIT_37 => X"B55A28408145AAFFFFFFF5D7FEAABA0051400A20000000000000000000000000",
INIT_38 => X"AB55FAD568AA2AFAE975EF555168B55F7AA800BAF7AA955EF00042AAA2A2AEAA",
INIT_39 => X"2AAAA007FD55558A7BD7145FBB8020A35D2ABEF55F7800015F087FEAA00007FE",
INIT_3A => X"968F575D003FF55F7D5420BA5D2ABFEAAF7AE9DFF759A82AEF70800021EF5504",
INIT_3B => X"FFD5145FBAC9755F05040255FFD84175EF55002AAB0A2FFEAABA557BEA3EF057",
INIT_3C => X"82E974AAF7D57DF45552A3FF10AA8429F45A7D5EAF5FFBAEAAA10554155400AA",
INIT_3D => X"FF843FFE77C80825BC052ABFE10550415557085540000005156155FE90A8F5C0",
INIT_3E => X"00000000000000000000000000000000000005500020AAF7FBFFFEF04552ABFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(3),        -- Port A data input
DOA(0)   => data_read_a_hi(3),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(3),        -- Port B data input
DOB(0)   => data_read_b_hi(3),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_4_15 : RAMB16_S1_S1
generic map (
INIT_00 => X"A108400020612C80284210081034849800A00030300004833522C82D04A16002",
INIT_01 => X"2043998A1839284D1CA0650E1E504368403008418984014902030806A0D10200",
INIT_02 => X"C120042200000000044441CE01E80F00A49043118680008002000000026208E4",
INIT_03 => X"040001020019200020011209CC0164C060000000690111040144800042F5C403",
INIT_04 => X"7029AF0F81A00010CCA47700CC513CAC0D0B8E02010740E19754080108988021",
INIT_05 => X"02139405007133C0712244CD20F20105D583000020E9892201D304D42A9835E1",
INIT_06 => X"9190440300078002014405D9EE814C0284A883B6D7038AE079059B7800048092",
INIT_07 => X"000100AA0004408000000004840400008D200102503000782000C00C8025C000",
INIT_08 => X"00728A00408403220811991E02120C044058080004000001101121F220000260",
INIT_09 => X"811001E1185B38AD23C3707AD46440818F3CF80EC423CA7D01D123C80200816A",
INIT_0A => X"45810810A01B40216361056D6150F41200280001900439001FD8A00041400000",
INIT_0B => X"11FC88076266E800D605402962A820211500024808010512C40106D222223B14",
INIT_0C => X"0408804116040B02C02C500B0C02C100B0C02C100B0402C300B0401618058611",
INIT_0D => X"040200050200501301208482200D00D0A0408402C4282200A84800009B878680",
INIT_0E => X"00000020000100024AC88300300060090F0D830F00025400300204D018000804",
INIT_0F => X"8000000040000206A2000800000000000000950002E010000000080000588040",
INIT_10 => X"0000000000000808000554000200000000000100006D0020000000100000BB00",
INIT_11 => X"0000400000000000002000001A0002504001000000000000002280000D800800",
INIT_12 => X"0800000000000E2C802000000000408D801000000000408012440000200110A0",
INIT_13 => X"000000000004680003A0040000000010280003800800000000102800000B0000",
INIT_14 => X"000005C0002000000000000620000158000010000000000010A0000B00000200",
INIT_15 => X"C30146200400104002602600400000000294004000000004000000000010001A",
INIT_16 => X"0080200000008020000000802000000080080000004090014134DA101288C6DB",
INIT_17 => X"0802000000000401806010040180601004018060100000802000000080200000",
INIT_18 => X"8060180601004010040080200802000000000000802008020000000000008020",
INIT_19 => X"C0A28A063807E0500014063450404882846FFE000003FFC00000010040100401",
INIT_1A => X"AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA28A28A28A28A2934C8D0CCD145144",
INIT_1B => X"68341A0D068341A0D068341A0D068341A0D068351A8D46A351A8D46A351AAAAA",
INIT_1C => X"FFFFFFFFFFFFFFFC0000000000000000000000001FE32068341A0D068341A0D0",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"408102040810207FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"800AA00000000000000000000000000000000000000000000040810204081020",
INIT_28 => X"168B55557BEAB4500554200000557FE10FFFBEAA10007FD7410FFAA97555082A",
INIT_29 => X"55574105D2A800AA00043FEBA5D7FEAA00007BE8AAAAA843DF55FFAA955EFA2D",
INIT_2A => X"57BC00AAA2FFEAAAAAA8415555087BFFF55A2AA800BAFFAE9555508002AA0000",
INIT_2B => X"A2AA955EF005568A00087BE8BFFA2D17DE1000517FE10AAAAA8AAA002E975455",
INIT_2C => X"FAA8417410A2D140000F7FBC2010A2D157400AAAE974AAAAAA974BA08002AB55",
INIT_2D => X"EFA2AABDEAA087BEAAAAA2FBD54BA080002145552ABFEAA007FC21EF007FD75F",
INIT_2E => X"00055042AB45F7FFD741000042AA10AAAABFF5508003FF55F7D568A00552EA8B",
INIT_2F => X"5400F7A49057D0824850B8000000000000000000000000000000000000000000",
INIT_30 => X"3AF55F7A0925D7AADB6FB7D5D7FEAB7808554203A145178E00FFFBE8A101475D",
INIT_31 => X"A9557D080038AAA145157428492E8008200043FE925571EFA380871C7028A28E",
INIT_32 => X"AEA8A9200249056D4175C5092AAF5FDA38BE8E1557D1475FAF45BEAA800AAFFA",
INIT_33 => X"AA4954281C0E2FB55B6A0925D7085F6AA10087FEABD7AAD57AEBA08517DE00AA",
INIT_34 => X"007FC51C7007BD55D7BE80004AAFEDB42028EBFBC2028BED152438AAA092492A",
INIT_35 => X"AF7DF6AA00412EAABFFAA803DEBA0875EDA80BEF1C743840040017D5520B8EAA",
INIT_36 => X"0000000000000000000041002FB55FFF5D0438140E2FA38B6AEBFF6DBE84AAEB",
INIT_37 => X"A00FFFFEAA105D5155410FF84021EF0800154B20000000000000000000000000",
INIT_38 => X"DEBA0851574B2AAAEAAB55F78400145AAFFFFFEF5D7FEABFF0051400A25D5568",
INIT_39 => X"68B55F7AA800BAF7AA955EF00042AAA25555410BA082E8201000043FE005D517",
INIT_3A => X"568AA200557DE00AAAAAAA000804001FF005575408AA557FEB2FFAE975EF5551",
INIT_3B => X"D1550AAAA8002010F2AC154B25F2ABFF55F7800015F087FEAA00007FEAB55FAD",
INIT_3C => X"800021EF55042AAAA007FD5555087BD6145FAAC000A2A6FBC00BAAAFBC00BAF7",
INIT_3D => X"F7AEBDFF779A82AA43F7FBE8A00082EA8BFFAA843FEBA08517DE00F3F9574B30",
INIT_3E => X"000000000000000000000000000000000000008003FF55F7D5420BA5D2ABFEAA",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(4),        -- Port A data input
DOA(0)   => data_read_a_hi(4),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(4),        -- Port B data input
DOB(0)   => data_read_b_hi(4),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_5_15 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50DF4A0791B3FCB694379283C81FD996A091832102004A336A20E03C040C002",
INIT_01 => X"805FBDC69830A84D5C6A60000C34C26841280A00084000C8C212892EEAD53235",
INIT_02 => X"3B2026B578918E640A4F01CF8011FF0002080000082CA9998276DF7772C7C80D",
INIT_03 => X"37134108420D700084205702A4008A1D9100002171C0E0051554D93A11F5D140",
INIT_04 => X"8A41A0FC03A56DA000425A819410E3816C086198A388B702A8CA1210844A0C4C",
INIT_05 => X"B1808A062E8BC835F5E84532D708238A282F00A9291224800A2861490343082C",
INIT_06 => X"903FB8483A90581859050424100940825C6184401CDC451B860A6507160C4100",
INIT_07 => X"D26F068BCC96CDF8918E640E96D1A3469D6300E2FFEA27F8E4D23248130E259C",
INIT_08 => X"0BFA82E568442B2A082C0A7E3014250D49DA37A2420619000002AFF48D1222E5",
INIT_09 => X"3F005001E40969289429360416DCD1C46083030604B1CA20C03DF83B0A2C60A5",
INIT_0A => X"14613C71005A10492B888120288F480D58858449026145B3830F449449062B4F",
INIT_0B => X"11AC04934AC648BFD727C031E64170A137D5AA5C3E4B0F8A3C58C34C002290E3",
INIT_0C => X"CA29C6CC50384B6AC6AC86AB31AACA6AB39AAC86AB39AACA6AB3055643559C31",
INIT_0D => X"C673E33CF28F38603855401985228A0614BD30A0A2819852011E5AC2B87F9182",
INIT_0E => X"FF87C002F87A803E460B2516510CA594FF0044FFA4B08BAC4BB2CD0F09CF84E3",
INIT_0F => X"0DFF0F8005F0F5100DFFF5E15D06101C55EB29F1E00BE53FE1F000BE1E802F94",
INIT_10 => X"F12F0380231F17D78FC029FFF58D9A70380230F2FE0017C37FC3E0017C3D005F",
INIT_11 => X"FC7F023C0CA700125C0F8F7E43F1F001BFFE7C69E01804E1E7CCF8FC003FF5F1",
INIT_12 => X"023E00017C1FC1A4BFD82C3081C5BD27BFE30C3081C5BD00C02365D645CEEF5B",
INIT_13 => X"61E0042787F181E9C1EFD8CB8120C5AF41E9C18FD60F0C20666F41E9F009FFFD",
INIT_14 => X"7A7C077FFF404F80005F07F187A7D14BFFC96111C048278DEB074F9930FF9D80",
INIT_15 => X"C064014B8B652E2B3120C81284641D3E8DBF7D636FE860190700132C1F0EFB80",
INIT_16 => X"38CE1384E3384E338CE138CE1384E33C4E3ECE32E128882551349A1CBAA44103",
INIT_17 => X"84E3384E3384E3384E338CE138CE1384E3384E338CE138CE1384E3384E338CE1",
INIT_18 => X"CE138CE138CE138CE1384E3384E3384E3384E338CE138CE138CE138CE1384E33",
INIT_19 => X"F5E5BB4E7F7B9DB7FF3A1B6DB7E8410A8C000000000000000000384E3384E338",
INIT_1A => X"BEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEF9F7CFDFDDCF3CF3D",
INIT_1B => X"BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEFBEF",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000001711C7BBDDEEF77BBDDEEF77",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"FDFFF00000000000000000000000000000000000000000000080000000000000",
INIT_28 => X"FD7410FFAA97410082A800AAAAAE955450055421FFFFFBC0010AAD5574BA557F",
INIT_29 => X"7FD74000055574BA5D7FD7555A2D5575EF55517FF5500557FE10FFFBEAA10007",
INIT_2A => X"0002AABA5D2ABFFFFAA843DF55FFAA955EFA2D168B55557BEAB5500554200000",
INIT_2B => X"5D2A800AA00043FEBA5D7FEAA00007BC00AAAAAEBDF45A28428B45FFD168BFF0",
INIT_2C => X"5080028A00A2FFFDE00F7D57FEBAFF80174BAAAD1555EF555555555005557410",
INIT_2D => X"BA5D2E821FFA2D5554BA557BD75FFAA8415555087BFFF55A2AA800BAFFAE9555",
INIT_2E => X"00000517FE10AAAAA8AAA002E97545557BC00AAA2FFEAAAA082A97545F7D5420",
INIT_2F => X"7010BEDF524AA5571FDFEF000000000000000000000000000000000000000000",
INIT_30 => X"78E00EBFBE8A101475D5400F7A49043D0824850B8A2AE9756D145B401FFFFFFC",
INIT_31 => X"FEAB7D0855420BA1471D74380851524BA5571D757DB6D5525EF555178F6D1451",
INIT_32 => X"8A28B6DEBDF6DBEF1C0A28AAA5524BFFFFA28E3AF55F7A0925D7AADB6FB7D5D7",
INIT_33 => X"5555057D145152428492E8008200043FE925571EFA380871C7028B6AEBDF45B6",
INIT_34 => X"BEAA800AAFFAA9557D080038AAAA2FBF8E10EBD578EAAFF8415482BED1555EF5",
INIT_35 => X"81C209256DFFDF420BA552A821FFB6DF574A85575C55EFBE8E1557D1475FAF45",
INIT_36 => X"0000000000000000000008517DE00AAAEA8A9200249056D4175C50920875FDA3",
INIT_37 => X"5FF5D7BC21EFF7FBD7400F7FBC00BA55557DFF70000000000000000000000000",
INIT_38 => X"01FF5D5568BE7555568A00AAFFEAA105D5155410FF84020AA0800154B2AAAA97",
INIT_39 => X"00145AAFFFFFEF5D7FEABFF0051400A25551554BA0051400BA5551575EFF7D14",
INIT_3A => X"1574B2FFAABFF45FFAAAABFFAAFFFDFFF552EA8AAA55043DFF7AAAEAAB55F784",
INIT_3B => X"8002410FFD5575EF5555421E75555400BA082E8201000043FE005D517DEBA085",
INIT_3C => X"FAE975EF555168B55F7AA800BAF7AA955EF00002AAA2A2FBE8A00A2D16AAAAFF",
INIT_3D => X"0055554088A557FEB25D00021FFFFFFC00BA552A821EFFFFFD74BA5D51575F7F",
INIT_3E => X"000000000000000000000000000000000000000557DE00AAAAAAA000804001FF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(5),        -- Port A data input
DOA(0)   => data_read_a_hi(5),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(5),        -- Port B data input
DOB(0)   => data_read_b_hi(5),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_6_15 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10800B0061A01002840002C03002818000402322520070B313301C4389B2082",
INIT_01 => X"250041CA3839684D18A160000C52426841000000090800090210080008110200",
INIT_02 => X"0020042080010000044654C0000C008010000000001020900200200002620814",
INIT_03 => X"060881021088200021080200E4000A0891000020610111500104C00000F14400",
INIT_04 => X"0880000100000002000052288144004281C050400100280000C8100000080001",
INIT_05 => X"928080840001100A08009000280201000850E022401400002028214043410820",
INIT_06 => X"10100518090012122100C808049310002040000410A0001400000200120840D2",
INIT_07 => X"000100800004400001000000860408108C22000A502010074120044800040001",
INIT_08 => X"50000040D0C4E2088003FD01C01004044058082004000000000121F020408244",
INIT_09 => X"00BF17E9001205A5204911F814444080400100020000D200DFD16400C2A40AA0",
INIT_0A => X"04611C17849000022862A1596C8B5DF04834948900000100220C244840000880",
INIT_0B => X"03AD0413424E4044D665C070C22602291504400D084915020448114080201000",
INIT_0C => X"5E08864011088B22D22C008B0022C408B1022C208B0822C608B1111600458010",
INIT_0D => X"4251A12CD28A300429688001000800000020280204001000A00804309A002182",
INIT_0E => X"0000000280402400420800000000006200FC10002442042429324294014E8CA7",
INIT_0F => X"A40000000500800840000800000000000002280018001480000000A010100052",
INIT_10 => X"00000000000004C2003000010240000000000000680800290000000140202000",
INIT_11 => X"2000C0000000000000000442000001080001000000000000010C000280001804",
INIT_12 => X"08000000000801C300A010000000156000902000000015101200002800000000",
INIT_13 => X"000000000101800038002408000000094000386028040000000940000ED40000",
INIT_14 => X"0003B000002000000000020180002A24005010000000000023000060C7000A40",
INIT_15 => X"3F0280090321000040A410C28108000160008094000810040000000000002300",
INIT_16 => X"284A5284A728CA5284A528CA728CA52C4A5A0A32A300940101349A0408240818",
INIT_17 => X"9CA1294A329CA5284A728CA7284A5284A728CA5284A528CA728CA5284A728CA7",
INIT_18 => X"CA3294A129CA3294A129CA1294A329CA1294A3294A129CA3294A129CA3294A32",
INIT_19 => X"F5F78BCE7F8FF0F4FA955F7CF7F40A80145D55555556AAAAAAAAA94A329CA129",
INIT_1A => X"8E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E39B6CEDECDDF7DF7D",
INIT_1B => X"F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE38E3",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000001A1A33F9FCFE7F3F9FCFE7F3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"555FF00000000000000000000000000000000000000000000080000000000000",
INIT_28 => X"BC0010AAD5574BA557FFDFFF087BFDF45F7AA974AAAAAA97555F784174BAF7D5",
INIT_29 => X"515555508043FE00F7AA97555A2FBD7410AA8428AAAAAAE955450055421FFFFF",
INIT_2A => X"7D1575EFFFAA9555500557FE10FFFBEAA10007FD7410FFAA97400082A800AA08",
INIT_2B => X"0055574BA5D7FD7555A2D5575EF55517FF55A2AA97400552AAAB45082E80155F",
INIT_2C => X"500554200000003DE10FFD5401FFF7AAA8A10082EAAB45A2FFC2000007FD7400",
INIT_2D => X"10AA803FE105D516AABAFF843FFFFAA843DF55FFAA955EFA2D168B55557BEAB5",
INIT_2E => X"000AAAEBDF45A28428B45FFD168BFF00002AABA5D2ABFFFF087BD5545007BFDE",
INIT_2F => X"256DEB84104BAFFD1525FF000000000000000000000000000000000000000000",
INIT_30 => X"9756D145B401FFFFFFC7010BEDF524AA5571FDFEF1C7BFFF55FFA095482B6A49",
INIT_31 => X"4904380824850381C5B5057D1C003DE28F7A49057DAAF5D2428A2842AAAAA2AE",
INIT_32 => X"2AAFB451C2A8017DE3DF525FFFFA49756D145178E00EBFBE8A101475D5400F7A",
INIT_33 => X"2F1C50381471D74380851524BA5571D757DB6D5525EF555178F6DAAA49542841",
INIT_34 => X"AADB6FB7D5D7FEAB7D0855420BA1C0E3FE00E3DB471EFE3AAAAA00082EA8B6DA",
INIT_35 => X"F1C7BD057D1C71FFE10A28038E1049516AAB8FF8428FEFA28E3AF55F7A0925D7",
INIT_36 => X"00000000000000000000B6AEBDF45B68A28B6DEBDF6DBEF1C0A28AAA5524BFFF",
INIT_37 => X"F55F78017400F780001FFAA84000AAFFD1401E70000000000000000000000000",
INIT_38 => X"20BAAA8428AA2AAAA975FF5D7BC21EFF7FBD7400F7FBC00BA55557DFF7557BFD",
INIT_39 => X"EAA105D5155410FF84020AA0800154B2557FC01EF55043FEAAFF80021EFA2D14",
INIT_3A => X"568BE7AA80174AA082ABDF555D2A821EFAAFBC01FFF780155F7555568A00AAFF",
INIT_3B => X"AEA8A10082EA8BEFAAD5554B25551554BA0051400BA5551575EFF7D1401FF5D5",
INIT_3C => X"AAEAAB55F78400145AAFFFFFEF5D7FEABFF0051400A25D2EBFE10AAFFD55EFA2",
INIT_3D => X"552EA8AAA55043DFF7557BC01EF55557DE00AA842AA0000516AABAFF8428BE7A",
INIT_3E => X"0000000000000000000000000000000000000FFAABFF45FFAAAABFFAAFFFDFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(6),        -- Port A data input
DOA(0)   => data_read_a_hi(6),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(6),        -- Port B data input
DOB(0)   => data_read_b_hi(6),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_7_15 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10844B00482258A2842112C02450418800002300500030B313300C418992002",
INIT_01 => X"000009CA3839684D1CA0E0000E51424840000000080000080200080008510204",
INIT_02 => X"0120042086010000044600C00008000004100000000260900200000002402004",
INIT_03 => X"8628A10000082400000002408400080011000000610008000208C00000E14400",
INIT_04 => X"0911800100A000000000524084000040000050001140200100C8100000080102",
INIT_05 => X"0300812401011000000000002000114008008060441000000020024093000000",
INIT_06 => X"9190431C0D4010100000880804010010800000041080081000000200010424B2",
INIT_07 => X"000100AA0004408601000004860000008C02000A103010006928040800062481",
INIT_08 => X"84000048D484C20888000A0002120484C048007004000000000021F000000244",
INIT_09 => X"00A06009881201A520491004106C48A04040002400A15A208001650004001020",
INIT_0A => X"C99E1060201002044809C1040140A001004808810000459033189C0A400118A0",
INIT_0B => X"102000024040484050050041648A0041140C500B08821054C000264120000400",
INIT_0C => X"0404A083260E0832132011880462011880462051881462051881D31018C40620",
INIT_0D => X"0001000080001000813094801A8F80F00A600B52602801A88848011118003700",
INIT_0E => X"000003C007C002808228010410082042C000C000000004001002000400040002",
INIT_0F => X"A4000007800F80C840000800009864038A1200081C0014800000F001F0200052",
INIT_10 => X"00002C0E00E0E4004038000102400002C0E00E0D20100029000001E003E04000",
INIT_11 => X"2000C04031100E0403D0700300080908000100000661801E1900040380001804",
INIT_12 => X"0840878083E8003780A01043203A101780902043203A10082410082880000000",
INIT_13 => X"0601E0187900181035E0240806483248181035E0280410C8198818100DDD0000",
INIT_14 => X"0403774000201021E020FA006040376C00501022131210722060806D47000A40",
INIT_15 => X"00928A0002000110888600C032128201519480D40009902430160403E0E00506",
INIT_16 => X"01000000020080601802000000000405000A0020020081014134928820480010",
INIT_17 => X"0802018040000000006018020080200804010000000000806018020080000004",
INIT_18 => X"0000000001806008020000001006008020080001004008020080201004000020",
INIT_19 => X"0000000000000000000000000000400A004618618618C30C30C3000020180600",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000000B0840000000000000000000",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"1555500000000000000000000000000000000000000000000080000000000000",
INIT_28 => X"A97555F784174BAF7D5555FFF780155EFAAAEA8ABAAAFBFDE0055556AA005D04",
INIT_29 => X"55555EFAAFFFDFEFAAAAAAB455D556AA00FFAE95555087BFDF45F7AA974AAAAA",
INIT_2A => X"02EAAAAA082EA8A00AAAE955450055421FFFFFBC0010AAD5574BA557FFDFFF55",
INIT_2B => X"08043FE00F7AA97555A2FBD7410AA8428AAA557BFDFFF55003DFFFF7FBEAA000",
INIT_2C => X"0082A800AAF7AE975FFA28000010552EBDE00007BEAAAAA2D140000085155555",
INIT_2D => X"45087FEAB455D516AB55557BD55FF00557FE10FFFBEAA10007FD7410FFAA9740",
INIT_2E => X"000A2AA97400552AAAB45082E80155F7D1575EFFFAA955555D51574AAAAFFD55",
INIT_2F => X"AE105D556AA10410E17555000000000000000000000000000000000000000000",
INIT_30 => X"FFF55FFA095482B6A49256DEB84104BAFFD1525FFFF8E175C7A2AAAAA82A2F1F",
INIT_31 => X"F524AA5571FDFEF415B575D7AAF1FFFD7AAAAAFB7D495F6AA10E3AE905551C7B",
INIT_32 => X"003AFEFEBFBEAA001C2EA8A821C2EAAA00A2AE9756D145B401FFFFFFC7010BED",
INIT_33 => X"EDB470101C5B5057D1C003DE28F7A49057DAAF5D2428A2842AAAA497BFAFFF49",
INIT_34 => X"1475D5400F7A490438082485038F7A4905C7A28A070384120BDE100075EAA82B",
INIT_35 => X"D495150492BEF1D2555087BE8B7D555F6AB57417BC05D7145178E00EBFBE8A10",
INIT_36 => X"00000000000000000000AAA495428412AAFB451C2A8017DE3DF525FFFFA49756",
INIT_37 => X"555A2AEA8A10AAD568A00555168A10002E9754D0000000000000000000000000",
INIT_38 => X"8A10AAAE8215D557BFDF55F78017400F780001FFAA84000AAFFD1401E7FFAA97",
INIT_39 => X"C21EFF7FBD7400F7FBC00BA55557DFF7007BD5555AAD57DF55AAAEBDFEF007BE",
INIT_3A => X"428AA2007FE8BFF080028BFFAAFFEAA105D2EAAA005D2AAAA18AAAA975FF5D7B",
INIT_3B => X"043DE0000516AA10F7FBD7408557FC01EF55043FEAAFF80021EFA2D1420BAAA8",
INIT_3C => X"55568A00AAFFEAA105D5155410FF84020AA0800154B2FF8402145A2AA954AA00",
INIT_3D => X"AAFBC01FFF780155F7005140000FFD140145007FE8BEF557BEAB55087FC215D5",
INIT_3E => X"0000000000000000000000000000000000000AA80174AA082ABDF555D2A821EF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(7),        -- Port A data input
DOA(0)   => data_read_a_hi(7),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(7),        -- Port B data input
DOB(0)   => data_read_b_hi(7),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_8_15 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00000648E2840112C00000418000002700500030B3132000400812082",
INIT_01 => X"100008480009004C04A100000252024840000000180800080200010040110204",
INIT_02 => X"0020042000490000004600804008000005100000000024900200000002400004",
INIT_03 => X"0A0C33400008082400000080A4004B0891000020610112000040C00000E5C000",
INIT_04 => X"18800001000000000000512080000040800150400824280110C8100000120200",
INIT_05 => X"908084A10100100200004080280008240810802206940000012C214451610800",
INIT_06 => X"81B000080860109021400008040000202048020414A0021400040200322824C1",
INIT_07 => X"000000080004408049000004860000008402001A50208000630C040800062483",
INIT_08 => X"440000428644212280800A00021004044048002124000000000021F000000244",
INIT_09 => X"00004009001001010008100414644410400102228000D20080114502006409A2",
INIT_0A => X"000051312000042200294429148A4801C80C8C81000045907118040340020832",
INIT_0B => X"4020000240404140004D0544C4AA0001150410090302500011C813428A000400",
INIT_0C => X"46501090008820240240409000240009000240009000240009000120204808A5",
INIT_0D => X"42D1A168D09A301468402480004780F00140080860280004085904309A002196",
INIT_0E => X"00783FC00044340242280000000000020000C0000442106419120004034685A3",
INIT_0F => X"8000F07F800088A80000081EA2F9EC0000064004081010001E0FF00011104040",
INIT_10 => X"0ED0FC7E00000422201080000202658FC7E0000021882020003C1FE000222080",
INIT_11 => X"018059C3F350FE0C00000002A0040500000103961FE780000110010090000800",
INIT_12 => X"FD41FF80000830200021C1CF600012200010D1CF600012121600100810000004",
INIT_13 => X"9E1FE000010A1802100004343ED8000898021000087073D80008980200800002",
INIT_14 => X"0080200000BEB07FE00002086008020000209AEE3F300000246020200000620B",
INIT_15 => X"0088881903210000440610C8000A808040000208901786E4F0FE0C0000000166",
INIT_16 => X"685A1685A769DA368DA368DA769DA36CDA121A11A141800011309284002C0810",
INIT_17 => X"95A5685A1685A5695A368DA368DA769DA368DA368DA7695A1685A1685A5695A1",
INIT_18 => X"5A1695A568DA368DA369DA768DA1685A1695A5685A168DA369DA768DA368DA16",
INIT_19 => X"A4028A0A543EBC57A10A1E75D64108080468618618630C30C30C69DA5685A168",
INIT_1A => X"9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7BF3CCD8DF5B2DB2C",
INIT_1B => X"F87D3E1F4F87D3E1F4F87D3E1F4F87D3E1F4F87C3E1F0F87C3E1F0F87C3E79E7",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000006A6D4F87D3E1F4F87D3E1F4",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"155FF00000000000000000000000000000000000000000000080000000000000",
INIT_28 => X"BFDE0055556AA005D0415555080000000087BEAA10F7803DE00FFAEBFFFF0800",
INIT_29 => X"2AA8AAA557FC0010F780154105D7FC2145005155555F780155EFAAAEA8ABAAAF",
INIT_2A => X"7FFFFF55AA80155FF087BFDF45F7AA974AAAAAA97555F784174BAF7D5555FF55",
INIT_2B => X"AAFFFDFEFAAAAAAB455D556AA00FFAE95555AAFFE8A00552EBFE00F7D17FF45F",
INIT_2C => X"A557FFDFFF5504000AAAAAAA8B55F7D140010552E821EFAAAABDF555555555EF",
INIT_2D => X"55AA8028A00A2D57FF45557BE8A00AAAE955450055421FFFFFBC0010AAD5574B",
INIT_2E => X"000557BFDFFF55003DFFFF7FBEAA00002EAAAAA082EA8A00002AA8A10F784021",
INIT_2F => X"FE10F7AEBAFFF080A175D7000000000000000000000000000000000000000000",
INIT_30 => X"175C7A2AAAAA82A2F1FAE105D556AA10410E17555080E000280071E8A00EB8E3",
INIT_31 => X"4104BAFFD1525FF492EA8AAA5571C2000FF8A17400557FC015514555757DFF8E",
INIT_32 => X"2ABDE10EBDF7AF6DE3FFF8F7DB68A105D71C7BFFF55FFA095482B6A49256DEB8",
INIT_33 => X"AA0BDF6D415B575D7AAF1FFFD7AAAAAFB7D495F6AA10E3AE90555A2FBE8A3849",
INIT_34 => X"FFFFC7010BEDF524AA5571FDFEF550E00082B6A0AFB55F7D1420104124821D7A",
INIT_35 => X"01C2EA8A00F7800017DA2842FA00B6D578F6D557FFDA00A2AE9756D145B401FF",
INIT_36 => X"00000000000000000000497BFAFFF49003AFEFEBFBEAA001C2EA8A821C2EAAA0",
INIT_37 => X"0BA08556AA00AAAABFE00F7AEAABEF082E955450000000000000000000000000",
INIT_38 => X"21555D51575EFFFAA97555A2AEA8A10AAD568A00555168A10002E9754D082E82",
INIT_39 => X"17400F780001FFAA84000AAFFD1401E7082EAAABA5D5140010F7AE974105D7BC",
INIT_3A => X"E8215DA2FFE8ABA082ABFE00AAFBEABFFAAFBEABFFF7AA80145557BFDF55F780",
INIT_3B => X"D540000000402145AA843FFFF007BD5555AAD57DF55AAAEBDFEF007BE8A10AAA",
INIT_3C => X"AAA975FF5D7BC21EFF7FBD7400F7FBC00BA55557DFF75D2E82010F7843DF45FF",
INIT_3D => X"5D2EAAA005D2AAAA185D2AAAA10F780021FFA2803DE10FFD16ABFF5D7BFDE10A",
INIT_3E => X"0000000000000000000000000000000000000007FE8BFF080028BFFAAFFEAA10",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(8),        -- Port A data input
DOA(0)   => data_read_a_hi(8),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(8),        -- Port B data input
DOB(0)   => data_read_b_hi(8),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_9_15 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00018248A2840112C00002C18000002300500030B3132000400812006",
INIT_01 => X"400008000000004C0020000000100248413C0A61590001D90213C10008110204",
INIT_02 => X"01A0042080010000054600C04008000004100000001020900200200002420804",
INIT_03 => X"024003400008012400000010E4004B0891000020610310000144C00000F5C000",
INIT_04 => X"1801800100E000000000510084000040010050020810200000C8900000320200",
INIT_05 => X"918004311104100000000000200008100800002000100000002C234415610820",
INIT_06 => X"81B00008080010100000980804000008800042041080001000100200322C2481",
INIT_07 => X"0000811800044080010000058600000086020002502080006000040800062C80",
INIT_08 => X"0000004001D4618008800A00061004044048002004000000000061F000000244",
INIT_09 => X"000040090802009420409004104444084001022400214A2080014400026401A2",
INIT_0A => X"04000071200000A003CA294140200800C80C8C8100004590111C040040120800",
INIT_0B => X"12210002404848502847040164880021150400080222000200C8034200000000",
INIT_0C => X"4610088010080421021040841021000841021000841021000841010800420820",
INIT_0D => X"42D0A16C529A321068500484000500D10042080040284000084900001A002196",
INIT_0E => X"00000002804000004228010410082002C000C0002400046419120410034285A1",
INIT_0F => X"A00000000500800800000800000000000002290008001080000000A010100042",
INIT_10 => X"00000000000004C2001000000240000000000000680800280000000140202000",
INIT_11 => X"0000C0000000000000000442020001000001000000000000010C800080000804",
INIT_12 => X"08000000000801A7802010000000152780102000000015000600000800000000",
INIT_13 => X"000000000101900011E0240000000009500011E0280000000009500004DD0000",
INIT_14 => X"000137400020000000000201C000136C00101000000000002340002947000240",
INIT_15 => X"0080881901210000000600C280028000419480D4000010040000000000002304",
INIT_16 => X"68DA368DA1685A1685A1685A1685A16C5A121A13A141950051309284A82C0010",
INIT_17 => X"85A1685A1685A1685A368DA368DA368DA368DA368DA368DA368DA368DA368DA3",
INIT_18 => X"5A1685A168DA368DA368DA368DA368DA368DA368DA3685A1685A1685A1685A16",
INIT_19 => X"0157344CCCF48DE68A895C38E2540A8010100000000000000000685A1685A168",
INIT_1A => X"14514514514514514514514514514514514D34D34D34D34D28E1004039248209",
INIT_1B => X"D268341A4D268341A0D069349A0D069349A0D068341A0D068341A0D068345145",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000014D490D069349A0D068341A4",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"EAABA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"03DE00FFAEBFFFF0800155FFAAFBE8B45002A974AAAA803DFFFAA843DF45FFFF",
INIT_29 => X"7BFDE00A2FBD7400F7FBFDFFFA2AEBDE00AAFBEAABA080000000087BEAA10F78",
INIT_2A => X"055401FFF7AEAAA10F780155EFAAAEA8ABAAAFBFDE0055556AA005D041555508",
INIT_2B => X"557FC0010F780154105D7FC2145005155555557BE8BEF007FFDEAAAAD1555EF0",
INIT_2C => X"AF7D5555FFF780154AA5D2AA8A10F7AA974AA082E80010A2AAAAA10552AA8AAA",
INIT_2D => X"BAF7D17FEBAA2AEBDF45002EAAABA087BFDF45F7AA974AAAAAA97555F784174B",
INIT_2E => X"000AAFFE8A00552EBFE00F7D17FF45F7FFFFF55AA80155FF080400145FFFBEAA",
INIT_2F => X"8FC7BE8A3DF7DF7F5E8A92000000000000000000000000000000000000000000",
INIT_30 => X"000280071E8A00EB8E3FE10F7AEBAFFF080A175D7BEF1E8B6D002090482B68E3",
INIT_31 => X"56AA10410E175550871FFE00A2FBD0400FFF5FDFC7B6A0BDE38B6F5E8A92080E",
INIT_32 => X"7BFAE82A2DB555C71C5B451D7FFAAA8A38FF8E175C7A2AAAAA82A2F1FAE105D5",
INIT_33 => X"2AEADA38492EA8AAA5571C2000FF8A17400557FC015514555757D5D71E8BEF14",
INIT_34 => X"B6A49256DEB84104BAFFD1525FFFF84174BA5D20AAA00E3AA904BA142A87010A",
INIT_35 => X"7000400155FFFBEDA82FFD57DEBAAAA0BFF7D0024ADA921C7BFFF55FFA095482",
INIT_36 => X"00000000000000000000A2FBE8A38492ABDE10EBDF7AF6DE3FFF8F7DB68A105D",
INIT_37 => X"BEF080402000F7AAA8B55FFAABDFEFF7D16AA000000000000000000000000000",
INIT_38 => X"FEAAFFD16AA00082E820BA08556AA00AAAABFE00F7AEAABEF082E95545F7D568",
INIT_39 => X"A8A10AAD568A00555168A10002E9754D00517DE00A2FFC2000F7D17FF55FF803",
INIT_3A => X"1575EF555568BEF5D7FE8A10AAFFD55555D7FD5555FFAAA8AAAFFAA97555A2AE",
INIT_3B => X"AE800AA552A97400A2AEBDEAA082EAAABA5D5140010F7AE974105D7BC21555D5",
INIT_3C => X"57BFDF55F78017400F780001FFAA84000AAFFD1401E7FF80174AA5D0028A00AA",
INIT_3D => X"AAFBEABFFF7AA80145080002145F7FBFFE00FFD17FEAAA2803DFEF08043FE005",
INIT_3E => X"0000000000000000000000000000000000000A2FFE8ABA082ABFE00AAFBEABFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(9),        -- Port A data input
DOA(0)   => data_read_a_hi(9),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(9),        -- Port B data input
DOB(0)   => data_read_b_hi(9),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_10_15 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00018248A2840112C00002C18000202300500030B3132000400992006",
INIT_01 => X"254008000000004C002000000010026840000000080000080200010008110204",
INIT_02 => X"0020042000010000004455800008000004100000000000900200000002400004",
INIT_03 => X"020001021089000021081000C400090011000000610001540104C00000F14400",
INIT_04 => X"0811800101A00002000050088554004200C840000000200080C8100000000001",
INIT_05 => X"030080001000100800009400200000000840E020201000000024024001200020",
INIT_06 => X"81B00008080012120004CC080492500280208004148000100000020020042493",
INIT_07 => X"0000000800044080010000048404081085020002502000006000040800062480",
INIT_08 => X"100202400084410808000A00021004044048000004000000000021F020408264",
INIT_09 => X"010040090002008420401004144440004040022484214A2080110108C2C00320",
INIT_0A => X"04004166A48A0001080000000000080080181881000045901118044040020800",
INIT_0B => X"1201000200484910000F0105602622291404020902005002018002400A022000",
INIT_0C => X"0440001011808020120004801120044800120004801120044800110002400884",
INIT_0D => X"008000440210100041308480800F82F00040180260A808008848000018002104",
INIT_0E => X"000000028040000002280104100820020000400020000440100204100A000100",
INIT_0F => X"040000000500800800000000000000000002280008000400000000A010100010",
INIT_10 => X"00000000000004C2001000010000000000000000680800010000000140202000",
INIT_11 => X"200000000000000000000442000001000000000000000000010C000080001000",
INIT_12 => X"00000000000801C0008000000000154000800000000015000410000800000000",
INIT_13 => X"0000000001019800180000080000000958001800000400000009580002800000",
INIT_14 => X"0000A0000000000000000201E0000A0000400000000000002360002080000800",
INIT_15 => X"0080881000000000000600C28102800060000000000800000000000000002306",
INIT_16 => X"401004010040100401004010040100441020D0030008840051309A90BA884010",
INIT_17 => X"0902409024090240900401004010040100401004010040100401004010040100",
INIT_18 => X"1004010040902409024090240902409024090240902409024090240902409024",
INIT_19 => X"F546890A940FE0D3971243555205428290100000000000000000401004010040",
INIT_1A => X"8A28A28A28A28A28A28A28A28A28A28A28A28A28A28A28A29554199854514514",
INIT_1B => X"2B95CAE532994CA6532995CAE572B94CA6532994CA6532994CA6532994CA28A2",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000002718E72B94CA6532994CA657",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"FDE1000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"03DFFFAA843DF45FFFFEAABA007FC2155F7D155545AA80001EFAAFBEAB45557F",
INIT_29 => X"042AB55FFD168B55AA8000010FFFBE8BFFF78402155AAFBE8B45002A974AAAA8",
INIT_2A => X"AD16AABA002ABDE10080000000087BEAA10F7803DE00FFAEBFFFF0800155FF00",
INIT_2B => X"A2FBD7400F7FBFDFFFA2AEBDE00AAFBEAABAA2FFD741055003DFEFF7AA801FFA",
INIT_2C => X"05D0415555007FD74105555555EFF7FBC0145F78028A00A2D142155087BFDE00",
INIT_2D => X"55AAD168ABA002A975FFF7AEBDEBAF780155EFAAAEA8ABAAAFBFDE0055556AA0",
INIT_2E => X"000557BE8BEF007FFDEAAAAD1555EF0055401FFF7AEAAA105D042ABFF5D556AB",
INIT_2F => X"71D7AAFBEFB455D71F8E00000000000000000000000000000000000000000000",
INIT_30 => X"E8B6D002090482B68E38FC7BE8A3DF7DF7F5E8A92007BC217DEBDB55555AA8E0",
INIT_31 => X"EBAFFF080A175D700042AB7DEBDB6DB55BE8E05000EBFFE8BC7E38E07145BEF1",
INIT_32 => X"0A3DFD7F7A4821D7A2D16FA82142EB8E00080E000280071E8A00EB8E3FE10F7A",
INIT_33 => X"ED1421450871FFE00A2FBD0400FFF5FDFC7B6A0BDE38B6F5E8A92B6FBD541049",
INIT_34 => X"A2F1FAE105D556AA10410E175550071D54104951555D7EBF5C5155E3842AA00B",
INIT_35 => X"8410E2ABD749516FB55BED16FA820820955EFE3AEBDEAAFF8E175C7A2AAAAA82",
INIT_36 => X"000000000000000000005D71E8BEF147BFAE82A2DB555C71C5B451D7FFAAA8A3",
INIT_37 => X"1EFA2FFD7545AAAE97555A2FBFDF455D556AA000000000000000000000000000",
INIT_38 => X"8B45AAAA95545F7D568BEF080402000F7AAA8B55FFAABDFEFF7D16AA00087FC0",
INIT_39 => X"6AA00AAAABFE00F7AEAABEF082E9554500042ABFFA2FFFFF45F7AE97400AAFFE",
INIT_3A => X"16AA00FFFBD5400082EBFF45F78400155A2D57FE00552EA8A00082E820BA0855",
INIT_3B => X"D557555A2802AA10FFD54214500517DE00A2FFC2000F7D17FF55FF803FEAAFFD",
INIT_3C => X"FAA97555A2AEA8A10AAD568A00555168A10002E9754D085155410085557555AA",
INIT_3D => X"5D7FD5555FFAAA8AAA002AAAB4508557DF55F7D17FE000804155FFAAAABDEAAF",
INIT_3E => X"0000000000000000000000000000000000000555568BEF5D7FE8A10AAFFD5555",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(10),        -- Port A data input
DOA(0)   => data_read_a_hi(10),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(10),        -- Port B data input
DOB(0)   => data_read_b_hi(10),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_11_15 : RAMB16_S1_S1
generic map (
INIT_00 => X"A101C4B05A0034CA2840712C2D001419000002300500030B31B20084EC992002",
INIT_01 => X"90000986B83028491800E0000C26426040000000080000088200080802512224",
INIT_02 => X"1A2004205E010640024D00800008000004100000040EC090820018003241A00C",
INIT_03 => X"28639100000C5C00000045C08400C8001100000061806A001618C03001E54400",
INIT_04 => X"1A800001000009A0804059A190000040400040008058220008C8100000120D4E",
INIT_05 => X"02000E81080250010000002022000058080400000E1200000020004401000004",
INIT_06 => X"819435143F20101010001008040800B8100102041088011100022200000024B2",
INIT_07 => X"90640D280884453E01064002944180008402001295BA100022E4340800062D82",
INIT_08 => X"400000093204802200280A0012160585C1D808D004000000000323F40C102244",
INIT_09 => X"380040098010001100009204107C5950400000220080C200800900020C006827",
INIT_0A => X"80007100004016EA080801010000080D00200081000045B0511D289940103399",
INIT_0B => X"002000024040410A000D0104408810C115D9C008050042400100D04E88000002",
INIT_0C => X"00655010009264201200C7B421ED0C7B421ED0C7B431ED087B43176843DA1085",
INIT_0D => X"0401020080400A10012494881A4F80F209500BB2602881A488485C1318002000",
INIT_0E => X"6619A540124814800228010410082022C00040002020090020220C9600040802",
INIT_0F => X"ACCC334A802491600C587949B6D0141B4CC600D5761B1599865A500490B86A56",
INIT_10 => X"BAC845542056A61686EC81E3A6CB68AA2C622C9A251C352B330CB4A0092170D8",
INIT_11 => X"BCCAD0B5A81536080CC6B21A21B1FC09CB0F1076D4A200B2AD4068F4101639B5",
INIT_12 => X"4D2CC281E31AA0103AB8D5514066380804B268A2E060901204112566F10AC418",
INIT_13 => X"D551443C47281002540B2C9AAAA8662A1152B202AE3554403028115AA88201A1",
INIT_14 => X"548A20A0492A2724A0621620402A020141F172FB182A32AB6845AB6200251BC9",
INIT_15 => X"00C00A000200074044E6801832728080D00A380B753952C4877E0104DDE4D124",
INIT_16 => X"0080200802008020080200802008020480080022020081010124988800400010",
INIT_17 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_18 => X"0000000000802008020080200802008020080200802008020080200802008020",
INIT_19 => X"55062608804180C0B10A42104201400204000000000000000000000000000000",
INIT_1A => X"00000000000000000000000000000000000820820820820801C4149470000000",
INIT_1B => X"0000000000000000040200000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000007E0F0000000000000100800",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"000AA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0001EFAAFBEAB45557FFDE10082ABDF5508557DF45002ABDFFFF7803DE10AA80",
INIT_29 => X"AEBFF45FFAEBFEAA002A801FFF7FFE8A10A28000000007FC2155F7D155545AA8",
INIT_2A => X"2AABFE10082ABFFEFAAFBE8B45002A974AAAA803DFFFAA843DF45FFFFEAABAA2",
INIT_2B => X"FFD168B55AA8000010FFFBE8BFFF78402155AAD155555A28428BFF002ABDE00A",
INIT_2C => X"F0800155FF00557FF45557FC2010002A80010A2842AAAA007BFFF4500042AB55",
INIT_2D => X"FF5D00154BAF7FBE8BEFFFD540000080000000087BEAA10F7803DE00FFAEBFFF",
INIT_2E => X"000A2FFD741055003DFEFF7AA801FFAAD16AABA002ABDE10A2D168A10A284021",
INIT_2F => X"DFC7F78E3FE28B684070AA000000000000000000000000000000000000000000",
INIT_30 => X"C217DEBDB55555AA8E071D7AAFBEFB455D71F8E00002EBDF6D005B78F7D142AB",
INIT_31 => X"A3DF7DF7F5E8A92BEAEBFF7DEBA0BDEAA1C2A801C7E3FFEFA10B68407038007B",
INIT_32 => X"8A28BFF082ABAE10B6AAB8E280820B8FEFBEF1E8B6D002090482B68E38FC7BE8",
INIT_33 => X"07FF8F7D00042AB7DEBDB6DB55BE8E05000EBFFE8BC7E38E07145B6D15756DA2",
INIT_34 => X"EB8E3FE10F7AEBAFFF080A175D708517DF7D497BC5028142A87000A28A2AA920",
INIT_35 => X"0B6DB6AA28A280001FF5D0A10482FFFFEFBC7E3DF42028080E000280071E8A00",
INIT_36 => X"00000000000000000000B6FBD5410490A3DFD7F7A4821D7A2D16FA82142EB8E0",
INIT_37 => X"FEF007BE8BFF5D2ABDF55F7AABDEAAF784154BA0000000000000000000000000",
INIT_38 => X"DE00FF84154BA087FC01EFA2FFD7545AAAE97555A2FBFDF455D556AA00082EBF",
INIT_39 => X"02000F7AAA8B55FFAABDFEFF7D16AA00FFAEBFFEFAA803DEBA5D2E82155A2FBF",
INIT_3A => X"A95545F7D5555FFAAAAA8BFF002AAAA00FFAAA8AAA080028BFFF7D568BEF0804",
INIT_3B => X"2E95400A2AEA8A00007FEABFF00042ABFFA2FFFFF45F7AE97400AAFFE8B45AAA",
INIT_3C => X"82E820BA08556AA00AAAABFE00F7AEAABEF082E9554508557DFFF007BD54BA5D",
INIT_3D => X"A2D57FE00552EA8A00FFFFE8AAAAA80001FF5D2E82000F7FFFFF45AAFFC20BA0",
INIT_3E => X"0000000000000000000000000000000000000FFFBD5400082EBFF45F78400155",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(11),        -- Port A data input
DOA(0)   => data_read_a_hi(11),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(11),        -- Port B data input
DOB(0)   => data_read_b_hi(11),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_12_15 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50080B01BC002006940202C0DE041196A83183000000023322287E0FC000006",
INIT_01 => X"75400D849830C84C5823E0000C17424840000000080000088200002802153231",
INIT_02 => X"18A026B43ED180040147558040090000061800000C06ED9802768F4472C52005",
INIT_03 => X"2A67E34A528D0524A52850528400C8001100000171C02B550618C91A10E55440",
INIT_04 => X"1BC0000100056C8280825DE98154004300C840800850240080CA921084520A07",
INIT_05 => X"02000F832000500C0000941024000852084060202E100001002000448100000C",
INIT_06 => X"819A1D1C3FE01A1A40045408049A50BA4020C6041090001200006200000000F2",
INIT_07 => X"C26A0719CC96CC6ED18A64019695A854870300FA3968B20068FC06080106249F",
INIT_08 => X"D002024B3E040800008C0A002610240D494A06F3460409000000E3F0AD5282E5",
INIT_09 => X"27A06009200040000400120412445D78400001000410420080218029CC807A27",
INIT_0A => X"18000006848A026F000000000000080000F010C100204593F11A6CDF48003BF8",
INIT_0B => X"000000820040402B28050400400432C9349DF21A31A00ACC0000F04F80020001",
INIT_0C => X"00357804611AE45D05D0833430CD0833420CD0C33420CD0833430668619A1000",
INIT_0D => X"0000000000000A74812DF00E87E80A079F9F90FA0280E87E800C7FF3B8002000",
INIT_0E => X"3B6B0E404D26160682082002000401EA0000C40000800A006002818808000000",
INIT_0F => X"A476D61C809A4DA84272592D6246FC1B17B541F97E1B348EDA93900B2B286C56",
INIT_10 => X"30C669E622DBC325CFD881A962454CFBE5403AB99594362B1DB52720165650D9",
INIT_11 => X"F8D2D39A3745261E4A95A110A3F855000E4B1D32BAB504BB7490FCFF912A3834",
INIT_12 => X"B90E9B018C7530200AB8F8BF41F9A22006B37DC8E1F9A21A70116D4C5080651C",
INIT_13 => X"118780319CCA08AB1001ACDF34B8F1C688AB1002AE3F7B807B6289F368828C4C",
INIT_14 => X"2AF020233376A5ECC016B1A827CDA21160F051DE610A34C50427E6E220323E4A",
INIT_15 => X"0077020000000439FDC05C5806781FAB46095A0B5199B0AC55521524F1864022",
INIT_16 => X"000000000000000000000000000000000026C000002884000130921092804010",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"8020080200000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0051B946088881360A95090CB054420290100000000000000000008020080200",
INIT_1A => X"041041041041041041041041041041041049249249249249200100002D451451",
INIT_1B => X"92C964B2592C964B2592C964B2592C964B2592C86432190C86432190C8641041",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000003800F592C964B2592C964B25",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"7DE1000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"ABDFFFF7803DE10AA80000AAAA843FE0008557DFFF0800020105D557FEAA0055",
INIT_29 => X"D5420000051555FFA2AA8200000557DFFFF7AA80000082ABDF5508557DF45002",
INIT_2A => X"82AA8AAAAAFFC00BA007FC2155F7D155545AA80001EFAAFBEAB45557FFDE10AA",
INIT_2B => X"FFAEBFEAA002A801FFF7FFE8A10A28000000A2D155410F7FFFFEBA08003FE000",
INIT_2C => X"5FFFFEAABA000028A105D2ABFE10A2AABFE1055516ABEF5D517DEAAA2AEBFF45",
INIT_2D => X"55002A820AA08557DFFFF7AA82155AAFBE8B45002A974AAAA803DFFFAA843DF4",
INIT_2E => X"000AAD155555A28428BFF002ABDE00A2AABFE10082ABFFEF0855420000004175",
INIT_2F => X"5010495B7AE921C517DE10000000000000000000000000000000000000000000",
INIT_30 => X"BDF6D005B78F7D142ABDFC7F78E3FE28B684070AABE803AE38145B78FD700000",
INIT_31 => X"BEFB455D71F8E00BED547038145B505FFB6A487000005F7AFD7F7A482038002E",
INIT_32 => X"F1FDE821C003FE001C2EAAAAAB6F5C2082007BC217DEBDB55555AA8E071D7AAF",
INIT_33 => X"D517DEAABEAEBFF7DEBA0BDEAA1C2A801C7E3FFEFA10B68407038B6D550428FF",
INIT_34 => X"B68E38FC7BE8A3DF7DF7F5E8A9200002FA285D20BDE28A2A4B8E10555B68BEF5",
INIT_35 => X"F085F47038140010555142082082005F7DFD7F7A482155BEF1E8B6D002090482",
INIT_36 => X"00000000000000000000B6D15756DA28A28BFF082ABAE10B6AAB8E280820B8FE",
INIT_37 => X"ABA5D7FEAB45080015410007FEAA0055517DE000000000000000000000000000",
INIT_38 => X"AB45F780020BA082EBFFEF007BE8BFF5D2ABDF55F7AABDEAAF784154BAF7802A",
INIT_39 => X"D7545AAAE97555A2FBFDF455D556AA00F7D1554BA5D7BC01FFFF8015410007FE",
INIT_3A => X"4154BAF7D1400BAFFD57FE005D043FE10552EAAAAAFFD140000087FC01EFA2FF",
INIT_3B => X"8428A105D7FEABEF55557DEBAFFAEBFFEFAA803DEBA5D2E82155A2FBFDE00FF8",
INIT_3C => X"7D568BEF080402000F7AAA8B55FFAABDFEFF7D16AA0008003FEBA55003DEBAA2",
INIT_3D => X"FFAAA8AAA080028BFF087BD54AA550402145550000010087FFFF45F78402145F",
INIT_3E => X"0000000000000000000000000000000000000F7D5555FFAAAAA8BFF002AAAA00",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(12),        -- Port A data input
DOA(0)   => data_read_a_hi(12),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(12),        -- Port B data input
DOB(0)   => data_read_b_hi(12),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_13_15 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10154A0441836CA2840512822007C18000E02700500030B31B300040081A042",
INIT_01 => X"00000804A000C04800020000000002404001000008220008A200100802110204",
INIT_02 => X"02200430000104000A4700804008000004100000000420918204D3033240400D",
INIT_03 => X"AA4003400008592400000590C40009141100000C6180C0000000C00001E14000",
INIT_04 => X"0800000102400120088054019000004160004190BAA0270000C8100000600206",
INIT_05 => X"21000012040610050040000227003AA0082400E94C1200000824424005220020",
INIT_06 => X"81963B180C001010580000080400000058000004109C00138000020024142581",
INIT_07 => X"002C8008000441600106400A9600010494020002B8AAA000EF003408000E2580",
INIT_08 => X"000000E48194408000A00A001210040441C80320040210000002ABF004102244",
INIT_09 => X"2A004009640040100400940412D4C4004000022000104200802D983000480120",
INIT_0A => X"8000202020401480000000000000080C90090881000145B0111A14004015080D",
INIT_0B => X"00000002004040AA08050400404040C11444000805200A402090024000008002",
INIT_0C => X"8410000A00280020020040800020040800020000801020000800010020400000",
INIT_0D => X"84A14250A055100050100490000500D00040080040290000084E4000B800610C",
INIT_0E => X"DCD13042BEDA36820228000000000000C000400081A08BC812A2092B02850942",
INIT_0F => X"89B9A260857DB400431969CA985D480949D32804A40AB137341C10B7D6A02EC0",
INIT_10 => X"E6ACA678001CE7D0296C213A460CA4271CA2168AEC1017606E6838216FAD4055",
INIT_11 => X"84AD4961C281B20213073C5FC0058008632D30D522CE80239DCC01AB013A4D20",
INIT_12 => X"2E6B13804A4B01D83461299900F6BD583A519104A0EEBD1A141010B2A4C8E116",
INIT_13 => X"89E5E40913419151EE0E94641828F72B5151EE0D184B321037AF5158BB02D085",
INIT_14 => X"562EC0B42162D68EE0073AE1C562EC13D521921A4170300B2B458B56B01C2280",
INIT_15 => X"00888A120240034000E6DC8285028014B82372011FC1E4F5E0A00929684EAF84",
INIT_16 => X"50942509425094250942509425094254940A1421420082020120908800480030",
INIT_17 => X"0942509425094250942509425094250942509425094250942509425094250942",
INIT_18 => X"9425094250942509425094250942509425094250942509425094250942509425",
INIT_19 => X"F7EFBBEEFF3F7DF7FF3E9F7DF7E2450228000000000000000000509425094250",
INIT_1A => X"BAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBF7DFDFDDD555555",
INIT_1B => X"EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAEBAE",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000000000F7EBF5FAFD7EBF5FAFD7",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"2ABEF00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0020105D557FEAA00557DE10AAD5554BA087FFFF55557BD54AAF7FBC01FFA280",
INIT_29 => X"7BD75EF087FFFFEF557BEAB45552E80155AA802AB45AA843FE0008557DFFF080",
INIT_2A => X"FAE820AA5D5557555082ABDF5508557DF45002ABDFFFF7803DE10AA80000AA08",
INIT_2B => X"0051555FFA2AA8200000557DFFFF7AA80000AAD1420AA087BD7555FFD168AAAF",
INIT_2C => X"5557FFDE10AAAEA8BFFA2FBD7545FFD157555085140010F7AEAABFFAAD542000",
INIT_2D => X"BA557BE8A10A284154BAFFAAAAB45007FC2155F7D155545AA80001EFAAFBEAB4",
INIT_2E => X"000A2D155410F7FFFFEBA08003FE00082AA8AAAAAFFC00BA00002AAAAF7D5574",
INIT_2F => X"0492E3F1C71C7BE8A2ABD7000000000000000000000000000000000000000000",
INIT_30 => X"3AE38145B78FD7000005010495B7AE921C517DE10A2DB50482147FFAF554971D",
INIT_31 => X"E3FE28B684070AA1C71D25D7007FFAFD7497BE8B5555208217DBE8A2AB45BE80",
INIT_32 => X"7FD257DFFD568A82FFA4870BA555F5056D002EBDF6D005B78F7D142ABDFC7F78",
INIT_33 => X"FAAAFBFFBED547038145B505FFB6A487000005F7AFD7F7A482038AADF4709214",
INIT_34 => X"AA8E071D7AAFBEFB455D71F8E00A2A0ADBC7A2FFD257DE3DF52555085142000F",
INIT_35 => X"21C002AA92FFDF574824171EAA10B680124BAFFAAAFB45007BC217DEBDB55555",
INIT_36 => X"00000000000000000000B6D550428FFF1FDE821C003FE001C2EAAAAAB6F5C208",
INIT_37 => X"0105D7BE8B55085142010AAD157545F7AEA8B550000000000000000000000000",
INIT_38 => X"01EFF7AAA8B55F7802AABA5D7FEAB45080015410007FEAA0055517DE00A2FFC0",
INIT_39 => X"E8BFF5D2ABDF55F7AABDEAAF784154BA5D5140145007BE8B55087BEAB555D040",
INIT_3A => X"0020BAA2FFD54105D7FC21EFFFD16AA10FF80174AA557FC21EF082EBFFEF007B",
INIT_3B => X"FBC0155085540000FFAEBFFEFF7D1554BA5D7BC01FFFF8015410007FEAB45F78",
INIT_3C => X"87FC01EFA2FFD7545AAAE97555A2FBFDF455D556AA00A2803FF45AAFFC21EFAA",
INIT_3D => X"552EAAAAAFFD1400005D042AA00F7FBD5410085568A10FF80020AAFFAABFF550",
INIT_3E => X"0000000000000000000000000000000000000F7D1400BAFFD57FE005D043FE10",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(13),        -- Port A data input
DOA(0)   => data_read_a_hi(13),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(13),        -- Port B data input
DOB(0)   => data_read_b_hi(13),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_14_15 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10020A000180000284008280000281800000030000000033022000000580002",
INIT_01 => X"000008020000204D006800000030824840000000084000084200090008510200",
INIT_02 => X"0220043170010A600A4D008040080000041000000028009002000F333240800C",
INIT_03 => X"111813400008002400000000C400090011000000610200001104D83000F14000",
INIT_04 => X"0801800100A000000000540084000040000040000800200000C8100000000748",
INIT_05 => X"0100000000001000000000002000080008000000001000000024024001200020",
INIT_06 => X"819EB84028001010000000080400000000000004108000100000020020040081",
INIT_07 => X"92040608000440100102400A94810206844200021DA2A0002000340800062C80",
INIT_08 => X"000000000084400008800A001214040441481500040000000000A7F408002244",
INIT_09 => X"0A0040090002008420401004104444004000020400214A208001000002400120",
INIT_0A => X"0400002020000000000000000000080C8008088100004590111B480040120000",
INIT_0B => X"1000000200404800000504016000002114000008020000020080024000000000",
INIT_0C => X"0410000010000000000040001000000000000040000000000001000000000000",
INIT_0D => X"04810244825010004010000000000000000000000000000000080000B8002104",
INIT_0E => X"0002C38280001202020800000000001000004000000000401022000002040902",
INIT_0F => X"20000587050001404E8084341CBA3404800828805200008000E0E0A000080002",
INIT_10 => X"4D18178E012010C00224004091C3514072C000444A0400080001C1C140001000",
INIT_11 => X"51709A07424142084458476001003809D0104B01C5710044020C4006010500C5",
INIT_12 => X"C26EE3803180C18006519462A00005001460E4730000050A1011004001060049",
INIT_13 => X"01F9E00660318000000538318740000140000001B4600CE80001400000002B62",
INIT_14 => X"0000000AD89857B0E0684411800000003799EB764D000330C300000000E3554B",
INIT_15 => X"0000021002002C000024008284001A0902000422E3F5960080480A0216A07240",
INIT_16 => X"4090240902409024090240902409024090081021020080015134920800480010",
INIT_17 => X"0902409024090240902409024090240902409024090240902409024090240902",
INIT_18 => X"9024090240902409024090240902409024090240902409024090240902409024",
INIT_19 => X"F5579B4E5C8FF0F7BE9D5F7DF650400200000000000000000000409024090240",
INIT_1A => X"9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7BF7DDDDDFCF3CF3D",
INIT_1B => X"F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE79E7",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000003FFF03F9FCFE7F3F9FCFE7F3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"420BA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"BD54AAF7FBC01FFA2802ABEFA2FBE8B55A2AE80000F7D5555555D2AAAABAAAD1",
INIT_29 => X"AA801FFA28402000AAAE955455500155EF0804155EFAAD5554BA087FFFF55557",
INIT_2A => X"7AEA8B45080417400AA843FE0008557DFFF0800020105D557FEAA00557DE10A2",
INIT_2B => X"087FFFFEF557BEAB45552E80155AA802AB4500516AA00A2AE800BAFFFFC20BAF",
INIT_2C => X"0AA80000AA005568ABAA28402010A2843FEBAFFFBD7410A2D168BFF087BD75EF",
INIT_2D => X"005D7FFDF4555517DFEF00043FEAA082ABDF5508557DF45002ABDFFFF7803DE1",
INIT_2E => X"000AAD1420AA087BD7555FFD168AAAFFAE820AA5D5557555002E80155A280000",
INIT_2F => X"0555412AA8ABAAADB40092000000000000000000000000000000000000000000",
INIT_30 => X"50482147FFAF554971D0492E3F1C71C7BE8A2ABD7A2FFEDB55B6A080038E3DB5",
INIT_31 => X"B7AE921C517DE10A2AE851FFB68402038AAAA955554900105FF0800175D7A2DB",
INIT_32 => X"A0800BAE3F1C0092EBAAADB6D080A12410BE803AE38145B78FD7000005010495",
INIT_33 => X"2D568BC71C71D25D7007FFAFD7497BE8B5555208217DBE8A2AB451C556FA00A2",
INIT_34 => X"142ABDFC7F78E3FE28B684070AA00516DABAA28402038B6803DE82F7F5D5410A",
INIT_35 => X"D002A80155B680000105D7FF8F455D5F78FD7000E3FEAA002EBDF6D005B78F7D",
INIT_36 => X"00000000000000000000AADF47092147FD257DFFD568A82FFA4870BA555F5056",
INIT_37 => X"F55FF84000AAAAFBC0145002AA8AAAAAFFC20000000000000000000000000000",
INIT_38 => X"01EF080417555A2FFC00105D7BE8B55085142010AAD157545F7AEA8B55A2FBFF",
INIT_39 => X"EAB45080015410007FEAA0055517DE00A2AA955FFFF80020BAAAAA9754508000",
INIT_3A => X"AA8B555D557FE00A280020BAAAD140000A2AEBFFEF082A82010F7802AABA5D7F",
INIT_3B => X"803DE00FFD557400AAD56AB455D5140145007BE8B55087BEAB555D04001EFF7A",
INIT_3C => X"82EBFFEF007BE8BFF5D2ABDF55F7AABDEAAF784154BA08557FEAAA284000AAFF",
INIT_3D => X"FF80174AA557FC21EF082A80145F780020105D7BEAB45557BE8B45082EBFEBA0",
INIT_3E => X"0000000000000000000000000000000000000A2FFD54105D7FC21EFFFD16AA10",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(14),        -- Port A data input
DOA(0)   => data_read_a_hi(14),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(14),        -- Port B data input
DOB(0)   => data_read_b_hi(14),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_15_15 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000A000000000284000280000001800020030000000033022000000180002",
INIT_01 => X"8000080000000048000000000000026040000000080000080200000000110200",
INIT_02 => X"0020042004010E60004C0080000800000410000000020090020000300245E005",
INIT_03 => X"0000010000080400000000408400480111000000610008000000C00000E54400",
INIT_04 => X"980000010000000088C2550080000040000040000008A00028C8100000120000",
INIT_05 => X"020004012E025000000001322000000A28008000011000000220004D41000000",
INIT_06 => X"819588000800101000011008040000100001060418800510000A620000000092",
INIT_07 => X"0000000800044004010C20008440810284020002102220002000340800062480",
INIT_08 => X"0000000001140800002C0A001214050540C800400406180000002DF004000244",
INIT_09 => X"1E00400900000000000016041044400440000000000042008001000000000022",
INIT_0A => X"0000000000000220000000000000080C00000081000045901118000040000000",
INIT_0B => X"0000000200404000010500004000000114000009000000000000004200000000",
INIT_0C => X"0000000000000000000040001000040001000000000000000001000020000800",
INIT_0D => X"000000000000001001208000180800000000030200000180800C400030002000",
INIT_0E => X"0000000000002600020800000000001080004000000000000002000000000000",
INIT_0F => X"A400000000000000000008000000000000000000000014800000000000000052",
INIT_10 => X"0000000000000000000000010240000000000000000000290000000000000000",
INIT_11 => X"2001C05838120800000000000000000000010000000000000000000000001804",
INIT_12 => X"081004000000000000A010000000000000902000000000180010002020000000",
INIT_13 => X"6600000000000000000024080000000000000000280400000000000000000000",
INIT_14 => X"0000000000200801000000000000000000501001920000000000000000000A40",
INIT_15 => X"0000020000000000000000003000000000000000000A101C3614000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000080000120980000000010",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000400200000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"28BEF00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"5555555D2AAAABAAAD1420BAFF8000010082A954BA00003DFEF085155400F784",
INIT_29 => X"AE95555A2FBE8BEFA2843DE00AA8015400FF84001EFA2FBE8B55A2AE80000F7D",
INIT_2A => X"2FBEAB45F7D56AABAAAD5554BA087FFFF55557BD54AAF7FBC01FFA2802ABEFF7",
INIT_2B => X"A28402000AAAE955455500155EF0804155EFFFFBE8BFF0800174AA557BFDE10A",
INIT_2C => X"A00557DE10F7D1574AAA2D16AB55FFD568BEF087FE8A1055003FE00A2AA801FF",
INIT_2D => X"00AA802AA00AAAE800BA5D0015545AA843FE0008557DFFF0800020105D557FEA",
INIT_2E => X"00000516AA00A2AE800BAFFFFC20BAF7AEA8B45080417400FFFFC21450800154",
INIT_2F => X"8FD7005150438F78A2DBFF000000000000000000000000000000000000000000",
INIT_30 => X"EDB55B6A080038E3DB50555412AA8ABAAADB40092E38E070280024904AA1C043",
INIT_31 => X"1C71C7BE8A2ABD7E3AA9257DA2FFE8BC7BE8E38E10A28017400E38A051FFA2FF",
INIT_32 => X"00124AA557FFDE10A2FBEDB6DF7D16AABAA2DB50482147FFAF554971D0492E3F",
INIT_33 => X"10038E38A2AE851FFB68402038AAAA955554900105FF0800175D7E3FFEFBD700",
INIT_34 => X"000005010495B7AE921C517DE10FFDF50482A2DB6AB45FFD56DBD7087BEAA384",
INIT_35 => X"0FFF1C017D140410400BE8E28A10AAA085082550A1057DBE803AE38145B78FD7",
INIT_36 => X"000000000000000000001C556FA00A2A0800BAE3F1C0092EBAAADB6D080A1241",
INIT_37 => X"4AA0800020BA550028B550855400AAF7AEBDFEF0000000000000000000000000",
INIT_38 => X"7400AAAE975EFA2FBFFF55FF84000AAAAFBC0145002AA8AAAAAFFC2000AAAA97",
INIT_39 => X"E8B55085142010AAD157545F7AEA8B55AAAE821EFAAFBEAB55F7AAA8A00AA841",
INIT_3A => X"417555AAFFFDF450804020AA557BFFE10A2FFFFFEFF7D568ABAA2FFC00105D7B",
INIT_3B => X"D17DF45007FE8AAA08002AAAAA2AA955FFFF80020BAAAAA975450800001EF080",
INIT_3C => X"7802AABA5D7FEAB45080015410007FEAA0055517DE00FFFBC2000AAFBE8B55F7",
INIT_3D => X"A2AEBFFEF082A82010FFD5421EF5D0000010F7AAA8A10AA8017400552A801EFF",
INIT_3E => X"00000000000000000000000000000000000005D557FE00A280020BAAAD140000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(15),        -- Port A data input
DOA(0)   => data_read_a_hi(15),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(15),        -- Port B data input
DOB(0)   => data_read_b_hi(15),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_16_15 : RAMB16_S1_S1
generic map (
INIT_00 => X"DA22C618B1000482B688B186588884862A400438255FC38381441205BA803003",
INIT_01 => X"7045A80028404C211203A952A90341080B173340412000E1005D628000820484",
INIT_02 => X"428406A4000850848330118D0AAC55001349B108818005460229044001C01784",
INIT_03 => X"092C4020000500020000500986812C405000001A48202050000A214AC0650115",
INIT_04 => X"4804A55440256F504025E003A054F46415A4E62B6FE3307943965A00001A1152",
INIT_05 => X"0000001C40A5B950ADB8EA097057ECE14C86D2B7F85AAD17F4B100000B88148C",
INIT_06 => X"415401DCDCF2C0A8030140BCB0820A200342A1C641C1E8782F508F2B00003584",
INIT_07 => X"002701881A3202080AE00480A2002840BE1480FA004342AA6F12000054004867",
INIT_08 => X"08C54828091002000002B32A8C19064E486A8001510000014140C1E2A14891E0",
INIT_09 => X"015452B103020814004088B64102680B6596594800400413CAC0208944800000",
INIT_0A => X"96AA000484094C000000000000012C9000A0000D0A80000BF8028E87C1B99270",
INIT_0B => X"014808A02004200E540480212000A448C0082024AE50064B44000000000002A2",
INIT_0C => X"0004000D5846256AAEA811150445411150445411150445411150422A088A8200",
INIT_0D => X"00000004010042A204A0C5817D00005034052E40000817D00440004004AD3240",
INIT_0E => X"632B2673FA4587978A2004102800809225545155121740000004900090000000",
INIT_0F => X"00C6564CE7F4EA4B940076D296D003030800462CBD320018CAAAACFE9164C800",
INIT_10 => X"28834ADB1440A114793A4A30A40839AA14910D08DCB2640031955559FD3AC990",
INIT_11 => X"594AB0B1A025371CA0E034E8443C097A800EB090D4AAC91208ED2FA0CE5E09B1",
INIT_12 => X"7B50446083001B94BB38C540EBE61284BB304880E3E4579EDC00992980D58033",
INIT_13 => X"5511121840E7A2CD952ECC12ABC3E6ACB3DFB12ECE315000F61FF1727A85FDBC",
INIT_14 => X"75DEB07F6F2E7084517F126F8395CB2BEFBAB8BA8AF698228CC5E2F08ECA5159",
INIT_15 => X"5580A840A8009F8B108C80A1021B080AFC0DF6422C6077F4A77F20D0C0E21084",
INIT_16 => X"0000000000000000000000000000000000044000102A0001148442A110810359",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"558D11544C690DA64C1C4F68A360400000000000000000000000000000000000",
INIT_1A => X"14D14D14D14D14D14D14D14D14D14D14D14514514514514529E5F87869E79E78",
INIT_1B => X"D1E8F47A3D1E8F47A7D3E9F4FA7D3E9F4FA7D3E9F47A7D1E9F47A7D1E9F4D14D",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000007D3E9F4FA7D3E8F47A3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"C00AA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"03DFEF085155400F78428BEF087FFFFEFF7D168B55AAD17FFFF552EBFE00007F",
INIT_29 => X"2E975EFF7D568BFFFF80175EF0004000BA552A821FFFF8000010082A954BA000",
INIT_2A => X"55540000082EAABFFA2FBE8B55A2AE80000F7D5555555D2AAAABAAAD1420BA5D",
INIT_2B => X"A2FBE8BEFA2843DE00AA8015400FF84001EF0000020AA5D00154005D043FF455",
INIT_2C => X"FA2802ABEF557BEABEF5D0415410087FD74BAAAAEBFFEF557FC00AAF7AE95555",
INIT_2D => X"FFFFAABFEAAFF84001FF002A821FFAAD5554BA087FFFF55557BD54AAF7FBC01F",
INIT_2E => X"000FFFBE8BFF0800174AA557BFDE10A2FBEAB45F7D56AABA082A97545F7D16AB",
INIT_2F => X"FFEF552AB8E38087FC2092000000000000000000000000000000000000000000",
INIT_30 => X"070280024904AA1C0438FD7005150438F78A2DBFF0871F8FC7E3D56AB6DBEDB7",
INIT_31 => X"AA8ABAAADB400924920925EFF7D16ABFFE38E175EF1400000BA412E871FFE38E",
INIT_32 => X"0A1240055003FF6D5551420101C2EAFBD7A2FFEDB55B6A080038E3DB50555412",
INIT_33 => X"57FC00BAE3AA9257DA2FFE8BC7BE8E38E10A28017400E38A051FF0804050BA41",
INIT_34 => X"4971D0492E3F1C71C7BE8A2ABD74975EDBC7550E12410087FD74AAB6AABFFC75",
INIT_35 => X"A08249756DF7D168BC7F7AABAEAAF780051C70824851D7A2DB50482147FFAF55",
INIT_36 => X"00000000000000000000E3FFEFBD70000124AA557FFDE10A2FBEDB6DF7D16AAB",
INIT_37 => X"B55A2D16ABEFFFFBFDFFF552AAAAAA007BC00000000000000000000000000000",
INIT_38 => X"20AA002A955EFAAAA974AA0800020BA550028B550855400AAF7AEBDFEF08516A",
INIT_39 => X"000AAAAFBC0145002AA8AAAAAFFC20000000021EFF7D568BFFA2AA955FF5D040",
INIT_3A => X"E975EF0800174BA002E820105D003DFEF5D51420005D2ABFF45A2FBFFF55FF84",
INIT_3B => X"7BD74AAF7AEBDF455D7BC20BAAAAE821EFAAFBEAB55F7AAA8A00AA8417400AAA",
INIT_3C => X"2FFC00105D7BE8B55085142010AAD157545F7AEA8B5500557DF45552A8200000",
INIT_3D => X"A2FFFFFEFF7D568ABA0804155FFF7D568B55FFAAAAABAFF8415545000015555A",
INIT_3E => X"0000000000000000000000000000000000000AAFFFDF450804020AA557BFFE10",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(16),        -- Port A data input
DOA(0)   => data_read_a_hi(16),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(16),        -- Port B data input
DOB(0)   => data_read_b_hi(16),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_17_15 : RAMB16_S1_S1
generic map (
INIT_00 => X"5284CE4FB7BD2C8994A13392DBD02E14006B82AC7E800D44D3DD2FD5F9B961C0",
INIT_01 => X"2EACD01F7E03FC6793F2199B39FC233C11D93AE6F3BB92B32091DBC339B24542",
INIT_02 => X"E63CCCC00A82C08092A2AFAE667033DB50853379C10BFDC5C6F4044443C817C6",
INIT_03 => X"7FF183635AEF9E3635AEF9E18E237040404446965C0607EE6DB7854AC4DE060C",
INIT_04 => X"D78AC33FB604488B000892EF17BE6D84196482236FE100294152E294350FB697",
INIT_05 => X"081B5F9B409420D0CDB47A05403F6CE0C08A4AB7F840EDB6F48100DFC8081081",
INIT_06 => X"768465354781CBC30316367077B4BDB50646E8D87100A8201ED01C19C020F71A",
INIT_07 => X"4002A110C922480A82D0841147162C48EBB9537A0022DC67987042EE976ABEA7",
INIT_08 => X"DB931BFEF91C00002CC0E019C0C82A4E4820C15A2330E004401891181168C4D1",
INIT_09 => X"09F3A1BC11EFBC66DB65307071477FF1030C397C060B4254064302042F803A69",
INIT_0A => X"3F330802162F3B7EE3F3EC7C7DEF207000F00059D2ED56D7EED2ED3C9A867DC0",
INIT_0B => X"185C44B91BC1740B7605040BE0018CFC7429F326B9E822FFC00074D5A0AB033A",
INIT_0C => X"00367A28FC1B7F7FEFFCFBFF3EFFCFBFF3EFFCFBFF3EFFCFBFF3EFFE7DFF9E00",
INIT_0D => X"0000000008004BA78428C7AD7FC94B533F5B4FFBD2FAD7FCCA786D43FE67C218",
INIT_0E => X"BA494CEBFD4F2667ABB6F68B29760593F33FA0CF170F40006001B1A05C000000",
INIT_0F => X"7F749299D7FAEB237DFE5865B6D2BF23265CBACE542A6FEE92333AFF33E0A9BF",
INIT_10 => X"F6C24B6D18C3C9F8E2881F3F787D776B5DB94A09955054DFDD246675FE7AC153",
INIT_11 => X"BFB349E08FF9A27EDE9FA8AEFD9E7467BFCB195CFEB56A1A70D34D1706FFFA3E",
INIT_12 => X"6FE219CA80725B875EED723FF7FCB2875EDAAFEAF7FD929BFD55BBC71D79F639",
INIT_13 => X"546670D018E7A6E581D7B6AB75FDFCECA6E581D7BB5DDFC6FF0EB7D7E859FDB5",
INIT_14 => X"B978177F6D6AF5ECDB5FB76A5F5FA165B456E0FB308710C49FCFB741598B9C7E",
INIT_15 => X"CFDAAB00AC00A8BBFC8B501CF7A0FED9A540EA1952586CEB54D143ACFF9A3BA9",
INIT_16 => X"000000000000000000000000000000000026E100002F382DBD9ECFE117805F20",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"4372003009EDCC4052E917114F981800C0000000000000000000000000000000",
INIT_1A => X"BA69A69AEBA69AEBA69A69AEBA69AEBA69A69A69A69A69A68698686981D75D74",
INIT_1B => X"6A351A8D46A351A8D068341A0D068341A0D068341A0D46A341A0D46A341A69AE",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000000000046A351A8D46A351A8D4",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"7FEAA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"17FFFF552EBFE00007FC00AA087FFFFFFFFFFFFFEFF7FBEAB450804001EFAAD5",
INIT_29 => X"D168A000004020AA5D7BE8B450051401EF087FD74AA087FFFFEFF7D168B55AAD",
INIT_2A => X"D7FEAB55FF80175EFFF8000010082A954BA00003DFEF085155400F78428BEFAA",
INIT_2B => X"F7D568BFFFF80175EF0004000BA552A821FF5D00020BA552A82000552A821555",
INIT_2C => X"AAAD1420BAFFFFFDF45AAD17FFFFAAFBC01EF5D0015555557BFDEBA5D2E975EF",
INIT_2D => X"BA007FEABEF005555555A2D1554BAA2FBE8B55A2AE80000F7D5555555D2AAAAB",
INIT_2E => X"0000000020AA5D00154005D043FF45555540000082EAABFF00516AA10552E820",
INIT_2F => X"8B550000071EFB6DF7AE92000000000000000000000000000000000000000000",
INIT_30 => X"F8FC7E3D56AB6DBEDB7FFEF552AB8E38087FC2092147FFFFFFFFFBFDFC7EBF5E",
INIT_31 => X"150438F78A2DBFFBED16AA381C0A07082497FEFB6D1451471EF007BD04920871",
INIT_32 => X"2A850105D2A80155417BEFB6DEB8E175FFE38E070280024904AA1C0438FD7005",
INIT_33 => X"D7BFAEBA4920925EFF7D16ABFFE38E175EF1400000BA412E871FF550A0009249",
INIT_34 => X"E3DB50555412AA8ABAAADB40092FFF5FFF6DAADF7FFD7B6F1C71EF55001756D5",
INIT_35 => X"7145B6AA28492487082007FEDBD700515556DA2DF50492A2FFEDB55B6A080038",
INIT_36 => X"000000000000000000000804050BA410A1240055003FF6D5551420101C2EAFBD",
INIT_37 => X"FEFF7FBFFF55A2D16AB550000175EFFFFBEAA000000000000000000000000000",
INIT_38 => X"55EF087FC200008516AB55A2D16ABEFFFFBFDFFF552AAAAAA007BC0000557FFD",
INIT_39 => X"020BA550028B550855400AAF7AEBDFEFF7D568AAA5D2A97410007BFFFFF55515",
INIT_3A => X"A955EF5D2E80010002A954005D2A82155087FFFFEFAAAA975EFAAAA974AA0800",
INIT_3B => X"D1575FF5504175EF5D7FEAAAA0000021EFF7D568BFFA2AA955FF5D04020AA002",
INIT_3C => X"2FBFFF55FF84000AAAAFBC0145002AA8AAAAAFFC2000FFD57DFFFAAFFFDF55FF",
INIT_3D => X"5D51420005D2ABFF45557FE8AAA000415410007BFFF450051555EFA2FBC0000A",
INIT_3E => X"00000000000000000000000000000000000000800174BA002E820105D003DFEF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(17),        -- Port A data input
DOA(0)   => data_read_a_hi(17),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(17),        -- Port B data input
DOB(0)   => data_read_b_hi(17),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_18_15 : RAMB16_S1_S1
generic map (
INIT_00 => X"69844019080000A21A611406840014122A641074155FC28A2024001001801003",
INIT_01 => X"7443D920034004180005E9E3C90360C0041C0181002001602025800008440084",
INIT_02 => X"E2DCCCE61D5C008103F2000781FC0FEDEAC2161B0B8FB0008620044443006010",
INIT_03 => X"884E300802006900802006995C896D605200000856E24A040000640052141103",
INIT_04 => X"480520FC026125AC0025C9122644E3E40EC8E2001001302281841A009038A86A",
INIT_05 => X"432000040089983070019400F01010004C8DB841405A80A100B586200FAC24AE",
INIT_06 => X"09044359DC7040000000002C109B0E0A00A1104641C0803804000707284600E1",
INIT_07 => X"400D10100400481D5EB08501620000007500CE801241021FE78E404860140060",
INIT_08 => X"00880C0106A0528020019307CC082A0A4A6A01ED725021400040D028000A9729",
INIT_09 => X"00117063038000282081402E4106400B6186128040600C10C1C0200950508110",
INIT_0A => X"C0C30C2E21580C874004008080003C32A10A19090C02010E1022944061688000",
INIT_0B => X"0180A8062026000DC425C0301311324AA2373088479105D044A1022000001835",
INIT_0C => X"0D89844703649000000200000000000000000000000000000000000000000010",
INIT_0D => X"0D8306C182701404C1973010802020404084001E00010802046092B5001FB365",
INIT_0E => X"528EB314068AB8B803DB00002900800400FC503F08180050942E4200020C1B06",
INIT_0F => X"40A51D66280D6032C5F96D3C51555D5D7D5AA87285820814A3CCC501C2A60820",
INIT_10 => X"8B35A3FEBF1FEDFD9C2B30E0468AAAD5D48F37E8FC1304102947998A03984C10",
INIT_11 => X"440FE1DD772D37A0A321BC6968F32658BF2D4F2A80BF8FE3F9FE3AC362080529",
INIT_12 => X"5487910D7E5A6D961A28456A1832E5161A100DD5182BC54020EA67A189C6ED36",
INIT_13 => X"AA444CAF91EDD1B725868403BE06323551B725868A100ABD119753B70964122B",
INIT_14 => X"EDC259048ACD868EE3803D65CEDC258A8F80D55E007C3F8EBB56F4C5362C978F",
INIT_15 => X"3F240014BE84370001B6922070440556B15F7FABBC0031BCF2257C41634B14D4",
INIT_16 => X"C1B06C1B06C1B06C1B06C1B06C1B06C1B0491069068000004060300A005A0118",
INIT_17 => X"1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06",
INIT_18 => X"B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C",
INIT_19 => X"B28BBECEB80EE173C2300F7DF16000000000000000000000000041B06C1B06C1",
INIT_1A => X"8A28A28AAAAAAA28A28A28AAAAAAA28A28A28A28A28A28A2910591505C104104",
INIT_1B => X"28944A25128944A25128944A25128944A25128944A2552A954AA5128944AAAA2",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000128944A25128944A251",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"9540000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"BEAB450804001EFAAD57FEAA087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974BA082E",
INIT_29 => X"7FFFFFFFFFBFDF45AAD568B55080028B55002E82000087FFFFFFFFFFFFFEFF7F",
INIT_2A => X"0043DE10AA843DE00087FFFFEFF7D168B55AAD17FFFF552EBFE00007FC00AA08",
INIT_2B => X"0004020AA5D7BE8B450051401EF087FD74AAAAFFFDF45A2D16AB55F7FFFFFFF0",
INIT_2C => X"0F78428BEFAA80000000804154BA55042ABEF5D7FD75FFAAD540145AAD168A00",
INIT_2D => X"00082E95555085168A10557FD7545FF8000010082A954BA00003DFEF08515540",
INIT_2E => X"0005D00020BA552A82000552A821555D7FEAB55FF80175EF5D00020105D2A974",
INIT_2F => X"DFFF5D2A954AA082A92428000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFBFDFC7EBF5E8B550000071EFB6DF7AE921C7FFFFFFFFFFFFFFFF7FBF",
INIT_31 => X"AB8E38087FC2092087FFDFC7E3F1FAF55A2DF6DB7D1C002AB7D002A82028147F",
INIT_32 => X"DF6DB7DE3F5FAFC708003DE28B68E38E280871F8FC7E3D56AB6DBEDB7FFEF552",
INIT_33 => X"ADF4516DBED16AA381C0A07082497FEFB6D1451471EF007BD0492B6F1F8F55AA",
INIT_34 => X"1C0438FD7005150438F78A2DBFFA28407038140410492550A2ABC7497BD25FFA",
INIT_35 => X"F5D0E05000492097428002E9557D1C516FA28417BD5545E38E070280024904AA",
INIT_36 => X"00000000000000000000550A00092492A850105D2A80155417BEFB6DEB8E175F",
INIT_37 => X"FFFFFFFFDFEFF7FBFFFEF552E974AA082A820AA0000000000000000000000000",
INIT_38 => X"ABEF002A800AA557FFDFEFF7FBFFF55A2D16AB550000175EFFFFBEAA00557FFF",
INIT_39 => X"6ABEFFFFBFDFFF552AAAAAA007BC0000087BFDF45AAD568B55AAFBFDFEF55042",
INIT_3A => X"FC2000FFD56AB45A2FFFDFFFAAD16AB4500043DEAAFFAEAAAAA08516AB55A2D1",
INIT_3B => X"2AA8B45087FC01EFA2FFD55EFF7D568AAA5D2A97410007BFFFFF5551555EF087",
INIT_3C => X"AAA974AA0800020BA550028B550855400AAF7AEBDFEFA280154BA55040000055",
INIT_3D => X"087FFFFEFAAAA975EF5D2E974000804154BA082A975EF5D517DEAA007BD5545A",
INIT_3E => X"00000000000000000000000000000000000005D2E80010002A954005D2A82155",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(18),        -- Port A data input
DOA(0)   => data_read_a_hi(18),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(18),        -- Port B data input
DOB(0)   => data_read_b_hi(18),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_19_15 : RAMB16_S1_S1
generic map (
INIT_00 => X"042200000000000041088001001AA00000000000000000000000500802000003",
INIT_01 => X"040048000024000000000404000000000A22000800000800004A200000000001",
INIT_02 => X"200C8840085EB00480060000001C008002489E0F000405EA0004040404000000",
INIT_03 => X"24004000000000000000000900002C4050000000000069500208400002E14100",
INIT_04 => X"4800200C0000000044002000C80020E40000E200000130200188000000800100",
INIT_05 => X"000000000080181000000000701000004C8000000058800000B1000009880480",
INIT_06 => X"80500081081040000000002C100040400000004641C080380400070100000000",
INIT_07 => X"4020109801A4CE005C00048380142810010564C4100114012002402028044808",
INIT_08 => X"0070700000000000000083004C3902420062000020E0000100004082A140102B",
INIT_09 => X"001150200000000000000026400000016186100000000010C04002C000000000",
INIT_0A => X"007C00008082C0002000000000002C3000000004050001030102040000000000",
INIT_0B => X"0000000000000000000000000000010000800011000000000000000000000BC0",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"000000000000000000000000000000042000760000000000000000010004B200",
INIT_0E => X"0D74002280300F0002FB069040000060000C5003000800000000000000000000",
INIT_0F => X"C01AE8004500744C780687DBA828008080A5FC0D385598035D0008A00C015660",
INIT_10 => X"39D8140040201BF861F0E7D693E6170022408116DFE0AB3006BA0011401D02AC",
INIT_11 => X"5412E4997F5249FD005043B8680CC98F00D0F2DD0140100406FE053A98F6ECC7",
INIT_12 => X"7418663001858040E153888000010840E165D0000000285C246A181C03FE4662",
INIT_13 => X"8199830066F0020858385974000001260208583854E2200000660208D6B1423F",
INIT_14 => X"8235AC508FCE8811042040F008235AE04420C040CF00C031C80009B8F224978B",
INIT_15 => X"030004E00000C220010808C10D9A92A74CD7CF4A09051110AD5A3C9200B7F280",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000118",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"07208BBA3F0C7010C660C7441920000000000000000000000000000000000000",
INIT_1A => X"861869A61861861861869A61861861861861861861861861A8208C4C1534D34C",
INIT_1B => X"984C26130984C26130984C26130984C26130984D26930984C26130984C261861",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000984C26130984C26130",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"174BA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFDFEF5D2A974BA082E95400F7FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0004",
INIT_29 => X"FFFFFFFFFFFFFFFFF7FBFDFFF552E974BAA2FFFFE10087FFFFFFFFFFFFFFFFFF",
INIT_2A => X"004001EFAAAEA8ABA087FFFFFFFFFFFFFEFF7FBEAB450804001EFAAD57FEAAF7",
INIT_2B => X"FFFBFDF45AAD568B55080028B55002E82000F7FFFFFFFFFFFFDFEFA2D568B550",
INIT_2C => X"0007FC00AAF7FFFFFFFF7FBE8B55AAD16ABEF5D2ABFF55080402010087FFFFFF",
INIT_2D => X"55A2FFFDFEF5D2EBFE00AAFFFFEBA087FFFFEFF7D168B55AAD17FFFF552EBFE0",
INIT_2E => X"000AAFFFDF45A2D16AB55F7FFFFFFF00043DE10AA843DE00557FFDFEFA2D16AB",
INIT_2F => X"FFEF552A974AA0000104AA000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFF7FBFDFFF5D2A954AA082A92428E3FFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"0071EFB6DF7AE92EBFFFFFFFFFFFFDFEFF7F5FAFC7492A974AAB6F5F8E101C7F",
INIT_32 => X"F1F8FD7AAD16AB450000001FFBEA4A8AAA147FFFFFFFFFBFDFC7EBF5E8B55000",
INIT_33 => X"00000010087FFDFC7E3F1FAF55A2DF6DB7D1C002AB7D002A82028FFFFFFFEFF7",
INIT_34 => X"BEDB7FFEF552AB8E38087FC2092F7FBF8FC7E3F5EAB45B6DF6FBEF5D2AB8F7D0",
INIT_35 => X"84971F8FC7AAD56DB6DBEF5F8FD7412ABFE28B6F5F8E820871F8FC7E3D56AB6D",
INIT_36 => X"00000000000000000000B6F1F8F55AADF6DB7DE3F5FAFC708003DE28B68E38E2",
INIT_37 => X"FFFFFFFFFFFFFFFFFDFEF552E954AA0004000AA0000000000000000000000000",
INIT_38 => X"54AAF7D568A00557FFFFFFFFFFFDFEFF7FBFFFEF552E974AA082A820AAA2FFFF",
INIT_39 => X"FFF55A2D16AB550000175EFFFFBEAA00A2FFFFFFFF7FBFDFFFFFD568B55002A9",
INIT_3A => X"A800AAF7FBFDFEFF7D56AB45AAD56AB450004001EFFF842AAAA557FFDFEFF7FB",
INIT_3B => X"FFFFFFF552AA8BEF080402000087BFDF45AAD568B55AAFBFDFEF55042ABEF002",
INIT_3C => X"8516AB55A2D16ABEFFFFBFDFFF552AAAAAA007BC0000FFFBE8B55AAD168B55F7",
INIT_3D => X"00043DEAAFFAEAAAAA08556AB55A2D57FFFFF7D568B45002ABDEAAFFD16AA000",
INIT_3E => X"0000000000000000000000000000000000000FFD56AB45A2FFFDFFFAAD16AB45",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(19),        -- Port A data input
DOA(0)   => data_read_a_hi(19),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(19),        -- Port B data input
DOB(0)   => data_read_b_hi(19),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_20_15 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000003",
INIT_01 => X"F55FF80000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"E05022020800008400F655001FFCFF80018FA804400000000000004400000001",
INIT_03 => X"00000000000000000000000900002CC07000000000000000000000000000013F",
INIT_04 => X"68002FFE40900010000180000001FFEC0012EE0C001370F40780000000000000",
INIT_05 => X"0840000880FCBBF0100E204DF0F88311DD8005080679800000F3000029980580",
INIT_06 => X"001000030817C8E8840155FDF9001001050023F6C3C3D0F87FA19F7F011000E4",
INIT_07 => X"000000090492260800008000EE00000000000000002101FF2002C00000004018",
INIT_08 => X"2A040001071004000013FF7FCA302C0C0008214800002101554031F800000000",
INIT_09 => X"801F57F200000090000489FEC0000001EFBEF0040008023FDFC0000000004006",
INIT_0A => X"0000000008000000000000000000ADF000000200000008000008028300110230",
INIT_0B => X"0000000000000800080000000000000000000000000000000800800A40000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"000000040900005C848538000020000000800000080000020000800101FFB600",
INIT_0E => X"00800000003A010003000000000000600FFC53FF001800000002004080000000",
INIT_0F => X"0001000000007408040000004000000004E9000008020000200000000E800800",
INIT_10 => X"00200000000313100010002000008000000000129600040000400000001D0010",
INIT_11 => X"81C012060000000000218F7840000100800004000000000066C0000080080000",
INIT_12 => X"800000000017C000100000000001A800080000000001A8040000002840008185",
INIT_13 => X"0000000006F00000100200000000012600001004000000000066000000801040",
INIT_14 => X"0000200410100000000005F00000020080090A0000000085C800002000586000",
INIT_15 => X"FF00400000000000020020020001000040283024E4F2860400008000030ED080",
INIT_16 => X"00000000000000000000000000000004010201001003020200000000000127DB",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"A0700030038200010089120104D2040020000000000000000000000000000000",
INIT_1A => X"2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2C30C30C30C30C306982121A1E79E79",
INIT_1B => X"32190C86432190C86432190C86432190C86432190C86432190C86432190CB2CB",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000432190C86432190C864",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0201000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF552A974AA0004174BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA0804",
INIT_29 => X"7FFFFFFFFFFFFFFFFFFFFFFEF552E954AA000400000F7FFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E954BA007FC00BA087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974BA082E9540000",
INIT_2B => X"FFFFFFFFFF7FBFDFFF552E974BAA2FFFFE10FFFFFFFFFFFFFFFFFFFFFBFDFFF5",
INIT_2C => X"FAAD57FEAA007FFFFFFFFFFFFFEFF7FBFFF550800020BAAAD56AAAAF7FFFFFFF",
INIT_2D => X"EFF7D56AB450000021EFA2D57DE10087FFFFFFFFFFFFFEFF7FBEAB450804001E",
INIT_2E => X"000F7FFFFFFFFFFFFDFEFA2D568B550004001EFAAAEA8ABA5D7FFFFFFFFFFFDF",
INIT_2F => X"FFFF5D2E954AA080005000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFEF552A974AA0000104AAFFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"A954AA082A92428087FFFFFFFFFFFFFFFFFFBFDFEF5D2E974AA000A07000E3FF",
INIT_32 => X"FFFFFEFF7FBFFFFF552E974AA0071C50BA1C7FFFFFFFFFFFFFFFF7FBFDFFF5D2",
INIT_33 => X"EDF6FABAEBFFFFFFFFFFFFDFEFF7F5FAFC7492A974AAB6F5F8E10E3FFFFFFFFF",
INIT_34 => X"EBF5E8B550000071EFB6DF7AE921C7FFFFFFFFFBFDFEFE3F5F8F450004050AAB",
INIT_35 => X"A497FFFFFFF7FBF8FC7EBD168B450804021FFB6D57DE28147FFFFFFFFFBFDFC7",
INIT_36 => X"00000000000000000000FFFFFFFEFF7F1F8FD7AAD16AB450000001FFBEA4A8AA",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2A954AA0800174100000000000000000000000000",
INIT_38 => X"74AA002E95410A2FFFFFFFFFFFFFFFFFFFFFDFEF552E954AA0004000AAFFFFFF",
INIT_39 => X"FDFEFF7FBFFFEF552E974AA082A820AA087FFFFFFFFFFFFFEFF7FBFDFFF5D2A9",
INIT_3A => X"568A00AAFFFFFFFFFFBFDFEFFFFFFDFEF5D2E954AA0051554BA557FFFFFFFFFF",
INIT_3B => X"D16AB450804174AAFFFFFFEBAA2FFFFFFFF7FBFDFFFFFD568B55002A954AAF7D",
INIT_3C => X"57FFDFEFF7FBFFF55A2D16AB550000175EFFFFBEAA005D7FFFFEFF7FBFDFFFAA",
INIT_3D => X"0004001EFFF842AAAA087BFDFEFF7FFEAB45A2D568B550804001EFF7D57DEBA5",
INIT_3E => X"0000000000000000000000000000000000000F7FBFDFEFF7D56AB45AAD56AB45",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(20),        -- Port A data input
DOA(0)   => data_read_a_hi(20),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(20),        -- Port B data input
DOB(0)   => data_read_b_hi(20),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_21_15 : RAMB16_S1_S1
generic map (
INIT_00 => X"4A302428B824900A128C090A5C1800261500213C005FE812D10420054085A202",
INIT_01 => X"001FFE3440B609703B0427F801A40B8115BC4F655300340288A40D30040E4DD8",
INIT_02 => X"E00424256888D8819801000F9FFFFFFFF149FF1FCA448046C60A0D2437C517F9",
INIT_03 => X"20030640003250640003250F06002CC1740002019824E001CD357832440001FF",
INIT_04 => X"EA2C3FFD400006E04401A8837001FFFC004AEF00080B70E08FB5789421007C5C",
INIT_05 => X"00011A0C40F9FFF80920954FF0F00809DF84A0202879800000F3000029980780",
INIT_06 => X"0805984B7A1FC0A0000101FFF0480080002281F7C3C381F87C03DFFF00009004",
INIT_07 => X"B424068086A205481A60A19000908204A855B000A08A61FF20C3D004D331D340",
INIT_08 => X"1BFA0001600802000023F7FFC08D234B40C2028253000040114200000D0226C0",
INIT_09 => X"EF1F5FF054096C6ADBA169FFC202B1C1FFBEF0440021083DFFCE22DC2880E24D",
INIT_0A => X"45FF0C004041D84862A28C54518DBFF00020004C0A6044901112A0908AA0A300",
INIT_0B => X"018C241102068006C620C03882019480E63180855A492712CC01C49C20201BFE",
INIT_0C => X"08A9464116544302C02D92236488D92236488D92236488D922366446C911B210",
INIT_0D => X"08800444021048034004001890000806002804A0822189000900D80621FFBE00",
INIT_0E => X"060580261013813A2CC396506102C4053FFD5BFF00A04A00200602CA52001100",
INIT_0F => X"080C0B004C202621A85C09411500135844C196D3606941018150098404C1A304",
INIT_10 => X"B02901013416181C96C2C9C600890A2028172192C460D1820302A0130809834A",
INIT_11 => X"9C5E803408250180AC268D185DB3F4350B811068C00049A0A4AA68F05C96A001",
INIT_12 => X"002C006560138F032B1804101244C883052208209040CC849063A747512B7678",
INIT_13 => X"41401E240665750440C9488280254530314080C2C601040420352148A00501B1",
INIT_14 => X"500811204D000700114204A70422016149916011008CAA8858850B00C32591C0",
INIT_15 => X"FFC06E60AC0496022300233104663040808E991765205000070121D41D18D098",
INIT_16 => X"40100401004010040100401004010040102090010008000001C0E010020007DF",
INIT_17 => X"0100401004010040100401004010040100401004010040100401004010040100",
INIT_18 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_19 => X"FFEF9FEEFF7FFDF7FF3E3DFDF7E0000000000000000000000000401004010040",
INIT_1A => X"BEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBFFDFDFFFCF3CF3F",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFEFF7FBFDFEFF7FBFDFEFBEF",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000FFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0001000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E954AA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0004",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA0004154BAFFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"52E974BA0804000AAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0004174BAFF",
INIT_2B => X"FFFFFFFFFFFFFFFFEF552E954AA000400000007FFFFFFFFFFFFFFFFFFFFFFEF5",
INIT_2C => X"A082E95400007FFFFFFFFFFFFFFFFFFFFDFEF5D2E974BA002E97400007FFFFFF",
INIT_2D => X"FFFFFBFDFEF5D2A954AA002E974BA087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFBFDFFF5D2E954BA007FC00BA5D7FFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA000002000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080005000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"A974AA0000104AAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974BA0000174AAFFFF",
INIT_32 => X"FFFFFFFFFFFFDFEF552E954BA080A000AAE3FFFFFFFFFFFFFFFFFFFFFFFEF552",
INIT_33 => X"02A95400087FFFFFFFFFFFFFFFFFFBFDFEF5D2E974AA000A07000007FFFFFFFF",
INIT_34 => X"F7FBFDFFF5D2A954AA082A924281C7FFFFFFFFFFFFFFFFFFBFDFEF5D2A974BA0",
INIT_35 => X"A557FFFFFFFFFFFFFFFF7FBFDFFF552E974BA0020924BA1C7FFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000E3FFFFFFFFFFFFFFEFF7FBFFFFF552E974AA0071C50B",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0000020000000000000000000000000000",
INIT_38 => X"74BA0000174BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954AA080017410FFFFFF",
INIT_39 => X"FFFFFFFFFFDFEF552E954AA0004000AAF7FFFFFFFFFFFFFFFFFFFFFFFEF552A9",
INIT_3A => X"E95410087FFFFFFFFFFFFFFFF7FBFDFEF5D2A954BA082E800AAA2FFFFFFFFFFF",
INIT_3B => X"FBFFFFF552E954BA002E97410087FFFFFFFFFFFFFEFF7FBFDFFF5D2A974AA002",
INIT_3C => X"57FFFFFFFFFFFDFEFF7FBFFFEF552E974AA082A820AA557FFFFFFFFFFFFFEFF7",
INIT_3D => X"5D2E954AA0051554BA5D7FFFFFFFFFBFDFEFF7FFFFFEF5D2A974BA0000020AA5",
INIT_3E => X"0000000000000000000000000000000000000AAFFFFFFFFFFBFDFEFFFFFFDFEF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(21),        -- Port A data input
DOA(0)   => data_read_a_hi(21),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(21),        -- Port B data input
DOB(0)   => data_read_b_hi(21),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_22_15 : RAMB16_S1_S1
generic map (
INIT_00 => X"5290F4CDE914905A14A43D33F488243E17122300F55FEB189B343A1140548380",
INIT_01 => X"A54007B259F6A975386262000C344BA9573C6FF57B18A5FB0ABFCD3C2C5F4F0C",
INIT_02 => X"021DFF8C38B3C009D203551040030071869D0040180AA2DC53DB89BEA8204001",
INIT_03 => X"2603475A969D0475A969D0460EAA401005111011BD506954EDB40F5EF41434C0",
INIT_04 => X"922D9002100ED69E443D988B0D5400103E48003D0800011E803B06B5B9125A15",
INIT_05 => X"281B5A0C06000408F4DF9422010D8802022F2124A8022492580040440002021C",
INIT_06 => X"F780C4C052881ADA0E05440205DA50930FA182010004700083E220800440B588",
INIT_07 => X"049D028B93FB561833D8094A02F5EA92FD7247E10305C40040D136E6A023F7FC",
INIT_08 => X"00028241680A0E002A9400803A884B5B5206B7C2E53CA25144009007A64EBD64",
INIT_09 => X"41008810240240C6694008010392354010000560141801002028A83D2A08E06D",
INIT_0A => X"34000000848BCA6902A29C54539C020E11810098D4067EFF9FF284D483E2AB41",
INIT_0B => X"500001840000C80B410014088040F4A944B1AA313C0022AA0011C0DC00028001",
INIT_0C => X"80B14004D158C8CA24A1C2A870AA1C2A870AA1C2A870AA1C2A872550E1543800",
INIT_0D => X"80A14050A01509E050854498B5281A1C34E506A2C6898B52A154DAC6B6000850",
INIT_0E => X"0B03001A483A4146603050080410089180008800143D83888281A2034A850142",
INIT_0F => X"A4160600349075238473F1210006133835E92273612B3482C090068A0E84AC56",
INIT_10 => X"30060181BA1B13959DC08DA902458870201970B29602562B0581200D141D0959",
INIT_11 => X"E042021C040D0152C8058B3840F044708E7E1C20A0106EA166C13AFC14AA3804",
INIT_12 => X"080E004B0C17C1439A9838301DC1A8438EA32C009DC1A8255300650458A1D588",
INIT_13 => X"018010E186F110A908E3A8CB0026C9A610A908E6A60F0807626610E160589C4C",
INIT_14 => X"2A701667334005800B1605F043858125E0D04110408D2485CA034681E43A1E40",
INIT_15 => X"00646002304244A91102C93A2D608D2A258DF8034188200C050171A41108F084",
INIT_16 => X"110441104411044110441104411044110466C440446CA06951D4EA8010009804",
INIT_17 => X"0040100401004411044110441104411044110441104411044110441104411044",
INIT_18 => X"0401004010040100401004010040100401004010040100401004010040100401",
INIT_19 => X"F7DFBFDEFE8FF1F7DEBDDF7DF7D05122890000000003FFFFFFFF900401004010",
INIT_1A => X"9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7BFFDFD7DDDF7DF7D",
INIT_1B => X"F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE79E7",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000003F9FCFE7F3F9FCFE7F3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA000400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0800",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000002000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2A954BA000015400FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080402010FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2A954BA0004154BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A0004174BAFFFFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0800154AAFFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF552A974AA0000174BAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974A",
INIT_2E => X"000007FFFFFFFFFFFFFFFFFFFFFFEF552E974BA0804000AAA2FFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080400010000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E954AA080005000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000402010FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2A954BA000417410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"804154BAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974BA0000174AAFFFFFFFFFFF",
INIT_34 => X"FFFFFFFEF552A974AA0000104AAE3FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0",
INIT_35 => X"AA2FFFFFFFFFFFFFFFFFFFFFFFEF552E954BA000E124BAE3FFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000007FFFFFFFFFFFFFFFFFFFFDFEF552E954BA080A000A",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804000100000000000000000000000000",
INIT_38 => X"54AA000400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2A954AA080017410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"0174BAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A954BA000415400FFFFFFFFFFFFF",
INIT_3B => X"FFFDFEF552E974AA0804174AAF7FFFFFFFFFFFFFFFFFFFFFFFEF552A974BA000",
INIT_3C => X"2FFFFFFFFFFFFFFFFFFFFFDFEF552E954AA0004000AAA2FFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2A954BA082E800AAAAFFFFFFFFFFFFFFFFFFFBFDFEF5D2E954BA002A820BAA",
INIT_3E => X"0000000000000000000000000000000000000087FFFFFFFFFFFFFFFF7FBFDFEF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(22),        -- Port A data input
DOA(0)   => data_read_a_hi(22),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(22),        -- Port B data input
DOB(0)   => data_read_b_hi(22),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_23_15 : RAMB16_S1_S1
generic map (
INIT_00 => X"EF20906D902424807BC8241BC81801B97D38AD3C0800103362A6741C80A12A02",
INIT_01 => X"001FFF8409F089003B4422000D80C80106804A7951C5B9D1C828043EA28838F9",
INIT_02 => X"E01CEE21649C82C40800000F9FFEFF8E72CA7F5FC2E22809925A0D3611C877F8",
INIT_03 => X"24000400402670400402670D48222DC1764446838624000080007460C40001BF",
INIT_04 => X"68403FFC020560E0443E21037C01FFFC0002EE00628BF0E02FAD781014085014",
INIT_05 => X"0112000202FBFFF00920017FF0F0628BFF8488890979800002F702002BB807A0",
INIT_06 => X"EF85788B681FC000000001FFF0010000000001F7CBC385F87C0BFFFF20040001",
INIT_07 => X"F6E200000000C1440E3AE408009120071070FA07A1CB23FFA403F0C4D23BF7C0",
INIT_08 => X"0BF87CA400804000003FF7FFD8880A034AC09662305AB10555421006891A1089",
INIT_09 => X"BE1F5FEA10092C0896A243FFC0008087FFBEF2000000001DFFC612C0C0400100",
INIT_0A => X"41FF0C2060501000600000000001BFFA800808189A657EF81DD0C00079CC8001",
INIT_0B => X"018C24110A860006C620C0312241C482B20400CC52492710CC80060020A81BFE",
INIT_0C => X"0C08866907048320C20C10030400C10030400C10030400C10030400608018210",
INIT_0D => X"040002000041500300100040000500C000801000C02400000952800001FFBF04",
INIT_0E => X"FC850015385380380CDB86106502C5043FFD5FFF00A04BC010A7724B10000800",
INIT_0F => X"89F90A002A70A710A51C01C05904014861433602A1CAF13F2110055614C72FC0",
INIT_10 => X"E02D02001C1E14981B43253EE50C8220180F1082E06397E07E42200AAC298E57",
INIT_11 => X"8421802400A90022B0070FAE18019214A380344920080B21A58B02AC60BACDF0",
INIT_12 => X"0A2A000C480B0704B54028101AC49C84BB4100009AC49C80857A82D20CE8CB22",
INIT_13 => X"01E00C8103416445C12ED0400027C5292445C12D500B0005A62D344CB241D095",
INIT_14 => X"132C907425604680038706A35132C94BDD011010404428886AC91B11311C8280",
INIT_15 => X"FF000470BE0692020328CA0028042054A92771C50FC070110001C1680809591D",
INIT_16 => X"00802008020080200802008020080200800800200200000000000008004807DF",
INIT_17 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_18 => X"8020080200802008020080200802008020080200802008020080200802008020",
INIT_19 => X"0000000000000000000000000000000000000000000000000000008020080200",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080002010FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974AA000400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000400010FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974AA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080000010FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E954AA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954A",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA000015400FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080002010FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974AA000400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000402010FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E954AA080005000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA080407000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA00041741",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080000010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000402010FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2A954AA080002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954AA080017410FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"552A954BA000415400F7FFFFFFFFFFFFFFFFFFFFFFFFF552A954BA080015410F",
INIT_3E => X"0000000000000000000000000000000000000F7FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(23),        -- Port A data input
DOA(0)   => data_read_a_hi(23),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(23),        -- Port B data input
DOB(0)   => data_read_b_hi(23),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_24_15 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100600007FFF000080108004000800020000840041000080808",
INIT_02 => X"FC5CA803400EB8209000000F9FFEFF8E7240FF1FC22409EA04018E50074017F0",
INIT_03 => X"11100400000000400000000D00002CC07400000090C080019001010A000001BF",
INIT_04 => X"68003FFC00040000000000008001FFFC0002EE00000370E007A100000000E468",
INIT_05 => X"0000000000F8BFF00920004DF0F00001DF8000000079800000F3000029980780",
INIT_06 => X"6E461803081FC000000001FFF0000000000001F7C3C380F87C019FFF00000000",
INIT_07 => X"600C2400013649609C8000980040814210254000A00B21FF2003F2A80D500000",
INIT_08 => X"0BF80000000000000003F7FFD88D2B4A02C0940062EC2804001610020408178B",
INIT_09 => X"8E1F5FE010092C0892A041FFC0000001FFBEF0000000001DFFC002C000000000",
INIT_0A => X"41FF0C0000000000600000000001BFFA0000005501AA00000CE2000009400000",
INIT_0B => X"018C0411020600048620C030020502000200000400490510CC00040020201BF4",
INIT_0C => X"0808064106040300C00C10030400C10030400C10030400C10030400608018210",
INIT_0D => X"0000000000004003000000000000001200580000000000000000000001FFBE00",
INIT_0E => X"0086C022005381380FDB96516140C6043FFD5BFF000041000000004110000000",
INIT_0F => X"80010D804400A7240C840C201D0210840043B4804012500021E0088014C04940",
INIT_10 => X"4109038041021C980200D06410C1924030008142E06024A00043C01100298092",
INIT_11 => X"587CC200002100C14428090A1D02348190814C09C010104025AA40041A0D8005",
INIT_12 => X"022E0030300B0E46177004208000D8C61D7004300000D884817B00011306B2D9",
INIT_13 => X"01E003060344710009875C018100013831000985DC000C20003C310006143B70",
INIT_14 => X"4001850EDC004780144806A64400186CBF8961104000C3807884000846EB9500",
INIT_15 => X"FF0006E08C063C0220002201490418082010A57263E0100008000290161E711C",
INIT_16 => X"00000000000000000000000000000000000000000000000000000000000007DF",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"F2D0AEEAF6E7CC1132CDB4441990000000000000000000000000000000000000",
INIT_1A => X"BEFBE79E79E79E79E79EFBEFBEFBEFBEFBEF9EF9EF9EF9EFA69861219575D75F",
INIT_1B => X"783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1EFBEF",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000783C1E0F0783C1E0F0",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0201000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A000400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA000400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000400000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402010000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"00002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080002010FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000400010FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA00040000",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020100000000000000000000000000",
INIT_38 => X"74BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"000010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA000002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974AA000402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000002010F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(24),        -- Port A data input
DOA(0)   => data_read_a_hi(24),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(24),        -- Port B data input
DOB(0)   => data_read_b_hi(24),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_25_15 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100200002000000080100004000000020000800041000080808",
INIT_02 => X"FC400086000000800000000F9FFEFF8E738FFF1FC204010000000111568DD7F8",
INIT_03 => X"00000400000000400000000D00002CC4740000008000000080000000000001BF",
INIT_04 => X"68003FFF64A564AC000000000001FFFE0082EF00010370E007A1000000004000",
INIT_05 => X"0A00040148F8BFF80920804DF0F00101DFC040000079C92484F30499299837C1",
INIT_06 => X"66041803081FC0E0801101FFFD000E41002299F7E3C380F87C019FFF81200096",
INIT_07 => X"000000080480AE00000080000000000000000000A00B21FF2003E00000000000",
INIT_08 => X"1BF80000400A02000003F7FFFA0008000200A0400008A0000014100200081000",
INIT_09 => X"8E1F5FFA53EFBCACB2E369FFE0010001FFBEF80C40630C7DFFEEBAF000800202",
INIT_0A => X"41FF0C0600000000600000000001BFFE00301000000000000CC020000140000C",
INIT_0B => X"01DCCC31222730A49620C030020100000200000400490D10EC00040220201BF4",
INIT_0C => X"0808064106240300C00C10030400C10030400C10030400C10030400608018210",
INIT_0D => X"0883044582114013412080000000000000000000000000000012800001FFBE00",
INIT_0E => X"00040020000180380FC386106140C6043FFD5BFF00A04B80608003CB120C1106",
INIT_0F => X"0000080040000200040400000100000000009480000240000100080000400900",
INIT_10 => X"0001000000000808000000240000020000000100006004800002001000008012",
INIT_11 => X"0001001808220000002004001900000080800008000000000022400000088000",
INIT_12 => X"0010000000000E00110000000000408009000000000040808063004000008200",
INIT_13 => X"6000000000046100000240000000001021000004400000000010210000001010",
INIT_14 => X"4000000404000800000000060400000088000001800000001084000000088000",
INIT_15 => X"FF800C608C041002000002000006100000002100000000180600000000100018",
INIT_16 => X"4110441104411044110441104411044510629041040D180400000010028047DF",
INIT_17 => X"1104411044110441104411044110441104411044110441104411044110441104",
INIT_18 => X"1044110441104411044110441104411044110441104411044110441104411044",
INIT_19 => X"FBA2894A196A8C5A2932EC15DA080800002FFFFFFFFFFFFFFFFFC11044110441",
INIT_1A => X"2492492492492492492410410410410410410492410492412000531215A69A6B",
INIT_1B => X"158AC562B158AC562B158AC562B158AC562B1588C46231188C46231188C49249",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000B158AC562B158AC562B",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080000010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000010FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08000000",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(25),        -- Port A data input
DOA(0)   => data_read_a_hi(25),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(25),        -- Port B data input
DOB(0)   => data_read_b_hi(25),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_26_15 : RAMB16_S1_S1
generic map (
INIT_00 => X"E9264EAB20190CA3BA4997AA9002AE9C001006B0778015CFA17E0811039879C7",
INIT_01 => X"2FFFF9BB1F773C7F9BB07DFFFDD863FC5FFF3FEFFBBF9FFB22FFFBC7B9F30686",
INIT_02 => X"E06CCC62052E708180F6FFBFFFFCFFFFF9C7FF7FC24332E642090000074037F6",
INIT_03 => X"428003739CD9863739CD9869FE2B7DEAF300029E4E300DFE69A6E644E6FF473F",
INIT_04 => X"7C2FEFFFF5BA124F003DD31EAFFFFFEE9FF7EE6F4C0770FFD7DC7CA53997B2B1",
INIT_05 => X"DFFB5421C1F8BBFAFDBFFACDF0FFCC05DDDBFF3690F9EDB7F5F7AFF639BD7DE3",
INIT_06 => X"EFD044ABC817C3E3A74667FDFFB6FF5727CC3BFEF7C3FAF87FF59F7FFBFEF69F",
INIT_07 => X"00003002132462052E708180EF060C18E5BEFB051225CDFF7002C4EEDE77F6E0",
INIT_08 => X"3FFF7D5000EC75088ED3FF7FC8790E46426CE06CB1F8E041051831FA3068D77E",
INIT_09 => X"C05FD7FF9BEFBDCEFBEE59FEF44F6603EFBEFAFCC2E35E7FDFD147CCF3F583FA",
INIT_0A => X"67FF1C7FBFADEB31E35768E8ED6BFDF3EB3EBF9DDBCE7FDC1DF8A760F3EACC02",
INIT_0B => X"5BDDCC3B336F7C548667D47B7737AF3FD62601EDC25B3533DCEB07F262213FFC",
INIT_0C => X"5F9A06E19F4D93A0EA0F78C35E30D78C35E30D78C35E30D78C35E986BC61AE31",
INIT_0D => X"5FD7AFEFDFFAF59B6FF28FE1D80D73D840607307DCFE1D80EF69A004DFFFF7FF",
INIT_0E => X"0004001F8041897B2FFFC6D86D70CE04FFFFF3FF1F5F5475BD7F72E4D75EBFAF",
INIT_0F => X"F60008003F008237B0040A00010003E020023E0201F45EC0010007E01047D17B",
INIT_10 => X"00010001DC0004C81003DE050A700200001DC0006863E8BD8002000FC0208FA2",
INIT_11 => X"2200E400002801E1A00004C21C0206F60081800800007B00010F02007EC09A0E",
INIT_12 => X"0880007E000807C7C1A612001E0015C7C19C22001E0015C59DFE82011A311AA0",
INIT_13 => X"00001BC00101F60409F0670840070809760409F06984800780097604067D0010",
INIT_14 => X"81019F40042100001F800203D81019EC085614000085C80023D81009CF008A74",
INIT_15 => X"FF802FFDFFAFD082003B032FB987E04021D481D4000819060801E0D00001231D",
INIT_16 => X"EBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEFFBFBFBFBBFCFBB0FFDFEFFEF2DFFFFFB",
INIT_17 => X"BFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAF",
INIT_18 => X"FAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFE",
INIT_19 => X"475B15BCF491E166CC8553F86EDB5C88646FFFFFFFFFFFFFFFFFEBFAFEBFAFEB",
INIT_1A => X"861861861861861861861861861861861861869A69A61861AFBD54D5F871C71D",
INIT_1B => X"984C26130984C26130984C26130984C26130984C26130984C26130984C261861",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000984C26130984C26130",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040201",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(26),        -- Port A data input
DOA(0)   => data_read_a_hi(26),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(26),        -- Port B data input
DOB(0)   => data_read_b_hi(26),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_27_15 : RAMB16_S1_S1
generic map (
INIT_00 => X"00080A40000A41248002029000050A088000008242A0004404480002000A1155",
INIT_01 => X"2FFFF1C11F781C129C107DFFFE0860941E81258CA2B71C2220EC1B86E1A00002",
INIT_02 => X"E1000000810000014400FF6FFFF0FFFFF8007F1FC21110005080200000221FF0",
INIT_03 => X"4080026318C18226318C1821302232EAE00002BE001115FE48620040840A863F",
INIT_04 => X"643D4FFC2530000F003D821C0BFFFF8E9EF79E6D440748FED70060842105B0B0",
INIT_05 => X"D6F39020D1F8A3FAFDBFBACDC8FDC405D1DB7F1490E5EDB7D5CBADB2385D79C3",
INIT_06 => X"6FE000A38007C3032646EFF1F0B6FF46A78C39F8E723F2E47FE59C7F9ADA2612",
INIT_07 => X"00002820000000810000014401060C180190310540118DFF1000C0849673F6C0",
INIT_08 => X"3FF779100062B12A8EC3F47FC80208808210880C00082050000110023068D030",
INIT_09 => X"005F07E09BFFBD07FBAC09F8E42922038F7DF8BEC2E39C5F1FD047CEF1B582D8",
INIT_0A => X"63FF5D5F9FADE911E81C09818109E1F16B16B71092CE7ED81CF403601228C402",
INIT_0B => X"1BFDCC39732F3554866AD57C37BEAF1C152201A4C05B7531D56B05B06A213FF8",
INIT_0C => X"5BCA06F18FC59380F00E34430D10C34430D10C34430D10C34430F0861A2186B5",
INIT_0D => X"5B56ADAB5FAAE58B2F628EA0C80FA3F04040510768EA0C80CC61A0044DFFC6EB",
INIT_0E => X"0004001D800188792CE79715710AE4047FFD23FF315D54358D593474955AB6AD",
INIT_0F => X"520008003B000297B0040200010003E020001F0201E44A400100076000579129",
INIT_10 => X"00010001DC00004A10035E0408300200001DC000086BC8948002000EC000AF22",
INIT_11 => X"02002400002801E1A00000C01E0202F60080800800007B00000782006EC0820A",
INIT_12 => X"0080007E000006A7C10602001E0001A7C10C02001E0001C18DE282010A311AA0",
INIT_13 => X"00001BC00000FE0401F04300400708007E0401F04180800780007E04047D0010",
INIT_14 => X"81011F40040100001F800002F81011EC080604000085C80001F810094F008034",
INIT_15 => X"FF800C6DDDAFD082001B03249887E04001D481D4000009020801E0D00001021F",
INIT_16 => X"AB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6BF1EBDABD8E270BF84A25C6ACB777E3",
INIT_17 => X"B6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6AD",
INIT_18 => X"6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADA",
INIT_19 => X"490E2168100481CA860402104A471688747FFFFFFFFFFFFFFFFFAB6ADAB6ADAB",
INIT_1A => X"000000000000000000000000000000000008200000000000200072F210000001",
INIT_1B => X"05028140A05028140A05028140A05028140A0500804020100804020100800000",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000A05028140A05028140A",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040201",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(27),        -- Port A data input
DOA(0)   => data_read_a_hi(27),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(27),        -- Port B data input
DOB(0)   => data_read_b_hi(27),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_28_15 : RAMB16_S1_S1
generic map (
INIT_00 => X"02200AA400180030808802A900002A08001280A08A801044104A1000001818C3",
INIT_01 => X"0AA00011460214428114180000882214413D0A71592A01D92213D28005210202",
INIT_02 => X"0451110A012100884000AA30200000000C100040104112101100008888200000",
INIT_03 => X"448000318C52A20318C52A20148810200111100C211004AA00034204200A2200",
INIT_04 => X"04004001001A90110000121402AA0000003C00000500000040080421080D0080",
INIT_05 => X"4060000C8001000000002E000000050000001610300000010000802202040012",
INIT_06 => X"1000002080001111001222000425A1040026A008000000000000000009328280",
INIT_07 => X"2491008A00491201210088400122448908A20402000408001000040820000000",
INIT_08 => X"20058310402A160026500000028040101004200C840082115554000112244814",
INIT_09 => X"4140000800000060000720000102028000000490160801020002200011100010",
INIT_0A => X"020000081B34211082B694D4D294000020020381040000000200032040004400",
INIT_0B => X"4800210C19808400500010009110091500020B408810000100200020408B0000",
INIT_0C => X"01028000080118020023604858121604858121604858121604858090B0242C00",
INIT_0D => X"010000800920040804020A6058003108402043058C460580653020005A004039",
INIT_0E => X"00000002800008014004104104420A00C000200005000010040A0020CC000200",
INIT_0F => X"520000000500000010000200000000000000280000040A40000000A000001029",
INIT_10 => X"00000000000000C0000002000830000000000000480008148000000140000020",
INIT_11 => X"020024000000000000000440000000020000800000000000000C00000040020A",
INIT_12 => X"00800000000001804006020000000500400C0200000005400A90000000100000",
INIT_13 => X"0000000000018200001003004000000142000010018080000001420000200000",
INIT_14 => X"8000080000010000000000018800008000060400000000000310000008000034",
INIT_15 => X"000002040080000000110006B081400000400000000009020000000000002200",
INIT_16 => X"802008020080200802008020080200802101210810C39A66A90A85420413A820",
INIT_17 => X"0200802008020080200802008020080200802008020080200802008020080200",
INIT_18 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_19 => X"DE21102C110A00246972BD89A40A0C22E1000000000000000000002008020080",
INIT_1A => X"2082082082082082082082082082082082082082082082080D35050758C30C31",
INIT_1B => X"0582C160B0582C160B0582C160B0582C160B0580C06030180C06030180C08208",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000B0582C160B0582C160B",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(28),        -- Port A data input
DOA(0)   => data_read_a_hi(28),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(28),        -- Port B data input
DOB(0)   => data_read_b_hi(28),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_29_15 : RAMB16_S1_S1
generic map (
INIT_00 => X"79964E4BA01DACAB9E659792D00AAE160002829C7FDFEFCEE97C2815039D70C3",
INIT_01 => X"0ABFF9AB0775343F9AB01DF80D5821FC0FFF3FEFD1AF9FF1207FFBC7B9720586",
INIT_02 => X"002CCC60050E700080F6AAA7BFFC007189C7FF2FC00330E602800000074037F6",
INIT_03 => X"468003210868A63210868A68DA017D207200021C4E200CAA6186A40042FF4300",
INIT_04 => X"7C2FE002F0900001003C5316A6ABFFE21F36E02F0D03701F47D41800109FB281",
INIT_05 => X"4979440580F9B808F49F6A4DF00F8D01DC4B97369078249370F482E62BA41462",
INIT_06 => X"B250442BC81001E1870223FC0BF7F11507C423FE33C078F803F19F00E936721D",
INIT_07 => X"00011080012460050E700080EF020408EC8CFA01122149FF700200665A35D260",
INIT_08 => X"2BFD055040A452000443FF00007906464068406C31F84000000831FA1028575A",
INIT_09 => X"805FD017102690AA694551FE30444681E0820AD40201423FC00122C493500172",
INIT_0A => X"0600002AFFBE2330815568A8AD6ABC02A02A0B0CCB463B4C0748A720B1EA4C00",
INIT_0B => X"0850400A11414C005005000B51158936D20601A98A10200308A002E240010BFC",
INIT_0C => X"05928020194918A22A2268C81A32068C81A32068C81A32068C81A99034640C00",
INIT_0D => X"058102C48970541944B20FA1580561D040406305587A158046282000DBFFF13D",
INIT_0E => X"000000028040890327DCD28928324400DFFFF0001F1F0050342D42A086040B02",
INIT_0F => X"F60000000500802010000A000000000000022A0000141EC0000000A01000507B",
INIT_10 => X"00000000000004C0000082010A700000000000006800283D80000001402000A0",
INIT_11 => X"2200E4000000000000000442040004020001800000000000010D000010401A0E",
INIT_12 => X"08800000000801C040A6120000001540409C2200000015441DAC800010100000",
INIT_13 => X"0000000001019600081027084000000956000810298480000009560002200000",
INIT_14 => X"800088000021000000000201D800088000561400000000002358000088000A74",
INIT_15 => X"00802594A282C0000033010FB181E00020400000000819060000000000002305",
INIT_16 => X"C0B02C0B02C0B02C0B02C0B02C0B02C4B12B312912831A27FCFE7FFB175B6FF8",
INIT_17 => X"0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02",
INIT_18 => X"B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C",
INIT_19 => X"BBCF9F96EE7FFDF7FE783FFDFFEA0C00602FFFFFFFFFFFFFFFFFC0B02C0B02C0",
INIT_1A => X"EFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEEBAEBAEBAEBAEBBFFDF9FBEFFFFFFE",
INIT_1B => X"BFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFBEFB",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000FBFDFEFF7FBFDFEFF7F",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(29),        -- Port A data input
DOA(0)   => data_read_a_hi(29),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(29),        -- Port B data input
DOB(0)   => data_read_b_hi(29),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_30_15 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"F7FFBFFEFF9FE1F7FFBFFFFDFFD0000000000000000000000000000000000000",
INIT_1A => X"9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7AFBD75F5FDF7DF7F",
INIT_1B => X"F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE79E7",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000003F9FCFE7F3F9FCFE7F3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(30),        -- Port A data input
DOA(0)   => data_read_a_hi(30),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(30),        -- Port B data input
DOB(0)   => data_read_b_hi(30),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_31_15 : RAMB16_S1_S1
generic map (
INIT_00 => X"129000008004A00804A40000400800020000000C005FEA005800200400050100",
INIT_01 => X"255FF18019700810180065FFFC0040801E80258CA2951C2200EC0906A0804140",
INIT_02 => X"E0000000000000011000550FDFF0FFFFF0007F1FC200000044000000000817F0",
INIT_03 => X"0000024210A30024210A3001002220C06044469200040154482000408400043F",
INIT_04 => X"602D0FFC2420000E003D80080955FF8E1ECA8E2D400340FE870060842100B030",
INIT_05 => X"0213100040F8A3F8FDBF944DC0FDC001D1CB6904A061EDB6D4C30490281831C1",
INIT_06 => X"6FC000830007C202060445F1F0D25E4207A099F0E303F0E07FE19C7F80402412",
INIT_07 => X"0000200000000000000001100004081001103107000185FF0000C0849673F6C0",
INIT_08 => X"1BF27A00000000000883F47FC800080002008000000820440000100220489020",
INIT_09 => X"011F07E013EFBC06FBA009F8E00120038F3CF82C44630C5D1FC002CCE0808248",
INIT_0A => X"61FF0C06C48BC801600000000001A1F00110101092CE7ED81CF0004012288000",
INIT_0B => X"11DCCC31222730048620C4382204A608142002A440492530C401049020221BF8",
INIT_0C => X"0888066187448380E00C10030400C10030400C10030400C10030600608018210",
INIT_0D => X"080204010200418301208480800D02D00040100240A808008840800405FF8640",
INIT_0E => X"0004001D000180780CE386106100C4043FFD03FF101D40008001304018081004",
INIT_0F => X"000008003A000217A0040000010003E02000160201E040000100074000478100",
INIT_10 => X"00010001DC00000810035C0400000200001DC0000063C0800002000E80008F02",
INIT_11 => X"00000000002801E1A00000801C0202F40080000800007B00000302006E808000",
INIT_12 => X"0000007E00000607810000001E000087810000001E000081846282010A211AA0",
INIT_13 => X"00001BC00000740401E0400000070800340401E04000000780003404045D0010",
INIT_14 => X"01011740040000001F8000025010116C080000000085C80000C8100947008000",
INIT_15 => X"FF800C609C06D082000A03200806A040019481D4000000000801E0D00001001D",
INIT_16 => X"010040100401004010040100401004010060C040040C200950402090128057C3",
INIT_17 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_18 => X"0040100401004010040100401004010040100401004010040100401004010040",
INIT_19 => X"00000000000000000000000000001000802FFFFFFFFFFFFFFFFF810040100401",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(31),        -- Port A data input
DOA(0)   => data_read_a_hi(31),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(31),        -- Port B data input
DOB(0)   => data_read_b_hi(31),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_0_14 : RAMB16_S1_S1
generic map (
INIT_00 => X"ED39BA795990D275FB4A6E96ACC4731DEA4598B0AFB54867F6EE4618C3749803",
INIT_01 => X"8AA0047D8607944AC7DA180001ECA2444042106208408208C20022E9173734B3",
INIT_02 => X"1A7DDD79F9A73E6CCA7DAAF00001000008478020113D98E382FEDF333027C80F",
INIT_03 => X"75D341110C58F31110C58F32A208921F8051500147A0E4AB3493FB3A01EBE240",
INIT_04 => X"86424001531009B100425A97B2AA0001E03501D0A39C8F0078420001106D0C4C",
INIT_05 => X"BCC8CA2EBF03400700402BB20F00239E20341699198600000B08694B16434804",
INIT_06 => X"103FB860B2800161F8432200012DA185F80F24081C3C0707800E600056881308",
INIT_07 => X"B24197ABCDA467F9A73E6CCAFDC3870EEEEC44E2BDFE220094D03022210C011C",
INIT_08 => X"240581B5695EAA80262C080032BF07C7C1FC3F8E94F65B11555EAFFC1C306758",
INIT_09 => X"7E40000BEC004170040DB60017FED1CC0001045002984202003DB931192D60A5",
INIT_0A => X"120071411A74315881A28C141118000C5A85A60444210123820B43B40804674D",
INIT_0B => X"0820008E514045BB514F0106D1D8599581D3A958BC104A89215AC14C48898403",
INIT_0C => X"C261C01C48B1584A0CA3E2687A9A1E2687A9A1E2687A9A1E26870CD061343885",
INIT_0D => X"D274E93A758FA8683AC54B287522E10A74AF4AA59C568752662F5AC218000002",
INIT_0E => X"FF83C002783A0904231C70470C7E0B92800224008AE09FAD4BD48D1FC5D3A4E9",
INIT_0F => X"5BFF078004F075885DFBF7E15C06101C55E921F1F80FAB7FE0F0009E0E903EAD",
INIT_10 => X"F12E0380231F13978FF023FAFDBD9870380230F2D6081F56FFC1E0013C1D207D",
INIT_11 => X"DE7F263C0C8700125C0F8F3C43F1F10BBF7EFC61E01804E1E6C8F8FE807F67FB",
INIT_12 => X"02BE00017C17C1007E5E2E3081C5AC007E6F0E3081C5AC44418D65FE45DEE55B",
INIT_13 => X"61E0042786F103E9F01F9BC3C120C5A703E9F01F978B8C20666703E9F8A0FFED",
INIT_14 => X"FA7E283FFB414F80005F05F10FA7E283F78F6511C048278DCA174FF038FF15B4",
INIT_15 => X"0066A20B61692F293185D8D724E15D3FCC6B7C236FE0691B0700132C1F0EF880",
INIT_16 => X"3A4E93A4E93A4E93A4E93A4E93A4E93A4F942F92E9628540AD2A91442525A000",
INIT_17 => X"A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E9",
INIT_18 => X"4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93",
INIT_19 => X"55F3898E09B56C74DAB15D1CF13501AA495000000000000000003A4E93A4E93A",
INIT_1A => X"082082082082082082082082082082082082082082082082082084E41DC71C71",
INIT_1B => X"E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F82082",
INIT_1C => X"FFFFFFFFFFFFFFF94A5294A5294A5294A5294A52800003E1F0F87C3E1F0F87C3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"3060C183060C187FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"BDEBA0000000000000000000000000000000000000000000003060C183060C18",
INIT_28 => X"168ABA002E82145085155545F7AA975EFFFAABDE00FFAEBDFFF5D2EAAAAAF7AE",
INIT_29 => X"7FFFE10005542145557FD5545FF8000155087FC0155F7D168B55007BFDF45085",
INIT_2A => X"7FFC0010080017555555568AAAFFFFD7545AA8028A00A2802AABAFF8028BEF5D",
INIT_2B => X"FF842AABAA2AE95545FFD168ABAF7AEAAAAAA2FFFDF4500043FE105D2E954BAF",
INIT_2C => X"5007FD7400550415410002E974BA5D5168A00A2D142155005142010FFAE820AA",
INIT_2D => X"FFF780000BA007FE8AAAFF803FFFF5D2A821550000000BA007FD55FF5D7FC014",
INIT_2E => X"000AAFBEAA00007BFDFFF082EBDF455D5142000082E82145FFD17DFEFFFD168B",
INIT_2F => X"DFD75D2AA8A80EA8E2FE3F000000000000000000000000000000000000000000",
INIT_30 => X"68B551475FAF6D1C556F0AA1C24AABEA495FC716F002A975FFE3AA95E00EBAEB",
INIT_31 => X"42A0070071C50BAFEF1FAE0016D56A16D557BC257D415E0216FA3F1E8FC0145B",
INIT_32 => X"8010E004924874825D7FEAA85487FD24AFE3D02DAAAE12BD5545A2803AA00005",
INIT_33 => X"120155EA568E870BAEB8A05A2AEA8B50F55A2F150005A3A438BD04AFAB8F550A",
INIT_34 => X"545E055FFBE81D0BE8EA8A3AA05A2A5504001C74BA42A1571E8028E3DB7816D0",
INIT_35 => X"A5C7E3DFFFE90B45B47ABA497A82FFAFD2A82485FD2415A105C21451ED42A002",
INIT_36 => X"00000000000000000000B55EAAA100AA1D0F6F480B6A555A2A57A002A3D5FDB6",
INIT_37 => X"5EFAAAAB5E1AF3AABFF45592E88A0AFE80A8B0A0000000000000000000000000",
INIT_38 => X"65F520EBE9EF67D7BEA1FD5D556ABEF5D557FEBA55022A3F70C6B405F4D2AE97",
INIT_39 => X"C114728007521170821CE0FDE69411A8DED57CE1055555E5F58EFFC01FE2CACB",
INIT_3A => X"42341D5DEEBEF55080034E0A592A4AD0079C75D6070CC5CBB0280C029ABAA3EB",
INIT_3B => X"7F353AAF6C77F7F20D968BF57812A95E02A2AAB5EB0F280800EFAEE9F5D18F31",
INIT_3C => X"C91565455C141E41887D58AC448B69C30E02116220415A9540AA854140A0A204",
INIT_3D => X"DE6BE93172D7D625B556EEAB157ABEBE1B4D792A4AD1183454180DD3FDCAAAB7",
INIT_3E => X"F0000001FF0000001FF0000001FF0000001FF01EABC4B8014174FF7DA80F52FE",
INIT_3F => X"FF0000001FF0000001FF0000001FF0000001FF0000001FF0000001FF0000001F")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(0),        -- Port A data input
DOA(0)   => data_read_a_lo_256(0),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(0),        -- Port B data input
DOB(0)   => data_read_b_lo_256(0),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_1_14 : RAMB16_S1_S1
generic map (
INIT_00 => X"212C001411984004084D000508C53810A03D1450E839B003342114428A000803",
INIT_01 => X"00000019400B100A8196000000CC004400400002000000000000028001340000",
INIT_02 => X"052137AE8031800C0044009000000000061800001CD4019802AD04CCCFC20004",
INIT_03 => X"04514108C60C21008C6042108400000201440020505100000043C30E10E9F000",
INIT_04 => X"02104001011DEFE088805681920000008000004001900800004002108C280008",
INIT_05 => X"040002340105000200000000080001900010000108040000000008411600401C",
INIT_06 => X"1034001042800808201000000001000820020000102000040000000000800180",
INIT_07 => X"64BF81A15EDFDE8031800C00843060C19E030022103600000450020800040004",
INIT_08 => X"00008004691687AA840008000090248CC84E000046000311555521F183060AC5",
INIT_09 => X"0820800D08100171000DB000154440C800400500000852020011200201012021",
INIT_0A => X"02000040001000880A2A04445004000102002041000001008208001440004140",
INIT_0B => X"4820018A1140440078050040511000102000A008183000010002404400000000",
INIT_0C => X"1000C80008000C030030880C2A030A00C28030A80C2A030A00C28018D4061401",
INIT_0D => X"10040802050080200284401C0022880F009E08008205C0020118088018000000",
INIT_0E => X"0F03C00280000000420860C60C0C0B92C0000000004000010042000040102008",
INIT_0F => X"001E078005000108400005E11C0610000000288058000003C0F000A000100000",
INIT_10 => X"F10E0380000000C202300000008D187038000000480800000781E00140002000",
INIT_11 => X"806302380C870010000004400100110800007861E0180000000C400680000001",
INIT_12 => X"023E00000000018000580C308000050000610C30800005000215006800000101",
INIT_13 => X"61E0000000018100B0001843812000014100B00016030C20000141002880026D",
INIT_14 => X"400A20009B404F80000000018400A20044096111C04000000304026000501580",
INIT_15 => X"0046820040082300218450C2800010094000482141E060190700100000002200",
INIT_16 => X"020080200802008020080200802008020080008008600500A82A1100A8000000",
INIT_17 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_18 => X"0080200802008020080200802008020080200802008020080200802008020080",
INIT_19 => X"81328A46BABEFC54A0810C7452B4428A14000000000000000000020080200802",
INIT_1A => X"AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA28A28A28A28A2A8218D2C0C924925",
INIT_1B => X"E974BA5D2E974BA5D2E974BA5D2E974BA5D2E975BADD6EB75BADD6EB75BAAAAA",
INIT_1C => X"FFFFFFFFFFFFFFFD8C6318C6318C6318C6318C63000002E974BA5D2E974BA5D2",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"70E1C3870E1C387FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"5555500000000000000000000000000000000000000000000070E1C3870E1C38",
INIT_28 => X"EBDF455D2EAABEFF7FFE8BFF5D0002155557FFFFFF007FC21EFA2FFD74AAAAD5",
INIT_29 => X"AA95400552AAAABAFFD1574105D7FD75FFAAAA800AAF7AA974BAFFFBE8B45F7A",
INIT_2A => X"0517DF555D2EAAA1055000015500557DF45AAD1400BAA2AE801550051555EFF7",
INIT_2B => X"FFD540155557FD5400F78028BFFFFFBEAB55F780020AAAA80020AA082EAAB550",
INIT_2C => X"AFF842ABEF5D517DF55552A974AAF7AE820AA0851574BAA2D1574AA5D7BFDEBA",
INIT_2D => X"EFAAD1575EF557FFFE10557FFFFFFFFD56AAAAFFFFD7555AAD168B45AAAEAAAB",
INIT_2E => X"0005D7FFDF4500043FE105D2E954BAF7AE80010082A97410557FEABFFAAFBE8B",
INIT_2F => X"51C7A2FBD5490BFD1C056A000000000000000000000000000000000000000000",
INIT_30 => X"974BAF7FFEFB45FFAABDF55492AA8BC2EBDFEAF7F1F840017D4975D2FEF147FC",
INIT_31 => X"080BEF495FC71D54124924385FAAA8AAAE3D145410F7F1D55D71C002DABAEBAA",
INIT_32 => X"002D082082AB8B6DBEDB7DF7F540E2AE85028B40155145F7AF6DBED5450AA1C2",
INIT_33 => X"78E021FF1471FDEAAFFD56F16D5571D2E28E38E0216FA2D1E8E80140F45082B4",
INIT_34 => X"A2DA3FB7DAAD4AAAAF487BC70BFA97F7AF6D417E92482BF84020BA495557E3FF",
INIT_35 => X"55554ADBD7A2FFC7BEFF6FFD7FC7002FD74951D71EDFFABFD16FAAAE92BD5545",
INIT_36 => X"00000000000000000000547AB8F550A8010E00492487482FFFE82A85EBAE2FFC",
INIT_37 => X"1EF005162BEF047FD5545AAFBF7400FBF9424F70000000000000000000000000",
INIT_38 => X"714F8338AAAA1D0AE974AAF7FFFDF55F7AABFF55082CA8B4DF6C1E8F5E540002",
INIT_39 => X"EABEF75550ACBB7582225FF5843404547184164AA5D2EBEEB0A2D555410D3555",
INIT_3A => X"FEAAEB083BC1000FF8409000512AEABFFDF79DCBF755962010BDCBBC21455D7F",
INIT_3B => X"801F8BA0C57740BDAA0688E5405D57D412F7D55F5E50C7F401BAAE8403CF5A3F",
INIT_3C => X"5D16BABAA3EBC3157ABD5FFE55F2AA9FEAFDF7F431A9F7FFE81FF013A8001AFF",
INIT_3D => X"FB863550229BCABEB7DA403FFFDA2FBF7FED2C7F955445079E280A00C56145EF",
INIT_3E => X"0000000000000000000000000000000000000596EBEF55080034E0A592A4AD00",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(1),        -- Port A data input
DOA(0)   => data_read_a_lo_256(1),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(1),        -- Port B data input
DOB(0)   => data_read_b_lo_256(1),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_2_14 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10E006600180111284380310006289800480032283E000A34301002001A0817",
INIT_01 => X"0005A00810790848048044A54E404350404000720885800802000906E4910200",
INIT_02 => X"407004208400408044C600C50AA055254010541A110222841200000002402544",
INIT_03 => X"0600011004182401004102408C28414043101000408118000145840440F5C415",
INIT_04 => X"5035855703A2900A000CD3088400F40688C9844409060850925E58A4081A0221",
INIT_05 => X"0200840D1021A15AC50494894850890540D1E12020C6E510818500440A280090",
INIT_06 => X"113044094002801020440090A8011A1224AB9380552102442884882A20004097",
INIT_07 => X"000100880004428400408044860000008C022402102100AA40004404B5075460",
INIT_08 => X"15C23440408C862A2A12382A8A5244145048C06085008010141521F000001240",
INIT_09 => X"400582B9033AA0E7AA4110B0506744810554542450694E710A836188C2C00222",
INIT_0A => X"443518360012C2210B020414109130A28038188096A06B8C120CA440A9C00802",
INIT_0B => X"1345E53300EC68005605002964AF222A5704004D080211121C80024200821780",
INIT_0C => X"181080C1110C882202211488452213C88472213C88472213488441109A442231",
INIT_0D => X"008204440210091341208041000810C00000300220201800A908000038AD0284",
INIT_0E => X"00040002804180300E88D28D206A40000554815500481440300000C44A081100",
INIT_0F => X"000008000500828700000000010000000002380000A00000010000A010050000",
INIT_10 => X"00010000000004CA000214000000020000000000684280000002000140200500",
INIT_11 => X"000000000020000000000442100002840000000800000000010C000026000000",
INIT_12 => X"00000000000805A4800000000000152300000000000015801272000100210020",
INIT_13 => X"000000000101C00000C000000000000940000120000000000009600004050000",
INIT_14 => X"0000130000000000000002018000106000000000000000002380000141000000",
INIT_15 => X"55000190000000000002000280000000011080C0000000000000000000002310",
INIT_16 => X"40902409064190641906419024090244902A9003004800415120D4A190804241",
INIT_17 => X"0900409004090641906419064190240902409024090641906419064190240902",
INIT_18 => X"9044090040900409004190441904419044090040900409004190441904419044",
INIT_19 => X"75960040138D70C030B51C50C7D100A2052F81F81F83F03F03F0419044190441",
INIT_1A => X"0410410410410410410410410410410410410410410410410248602081659659",
INIT_1B => X"5128944A25128944A25128944A25128944A25128944A25128944A25128941041",
INIT_1C => X"FFFFFFFFFFFFFFFE1084210842108421084210843FFF825128944A25128944A2",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"7FD5FF555815607FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"2AA000000000000000000000000000000000000000000000007FD5FF55581560",
INIT_28 => X"FC21EFA2FFD75EFAA8415410AA8415555087BFFF55A2AA800BAFFAE954000800",
INIT_29 => X"84155EFA2AEBDEAAA2FBEAABA5D7FE8B555551421455D0002145552EBFEBA007",
INIT_2A => X"2AEBDF555D2E954BAA2AA974BAFFFFE8B45552EBDF45FFAEAABFFF7FFE8B55F7",
INIT_2B => X"AAAAAAAAAFFD1574105D7FFFF555D2AAAAAA5D2E820BAA2FBEAB5555557DF55A",
INIT_2C => X"50055575EFFF84021555D043DEAA5D04021EF557FC21FFAA8428BFFAAAA954AA",
INIT_2D => X"10085568A00FF80175FFA2D17DFEFF7800215500557DF55AA80001FFAA800015",
INIT_2E => X"0005D00020AAAA80020AA082EAAB5500517DF555D042AA10A284154005D00154",
INIT_2F => X"00AAFFAA9543A080038A2A000000000000000000000000000000000000000000",
INIT_30 => X"0017D5D20B8EAA007FC51C7A2FBD55D2BE800042AFE8E1557D0075D2F45BEAA8",
INIT_31 => X"AA8BC7EBDFEAFEFFD00105FFBC20BDEAAA2FBF8AAA557BE8B6D5D5FFABEF4904",
INIT_32 => X"FFEFB6D555578F7DB6A0BDF7D480E174BFA02A974BAF7F5EFB455D2ABDF55492",
INIT_33 => X"ED1FDE90E3A497492B6AAADAAAE3D155E105571D55D71C002DABA5524820BAB6",
INIT_34 => X"BE8F401D7B6A0001470155C51D0092A071555D5E3AE821D00001FF0871C016DB",
INIT_35 => X"5BE8555400550A38428007FED000E3DA3DFD5E3DFFFBD5A38A021551C5F7AF6D",
INIT_36 => X"00000000000000000000410F45082B4002D082082AB8B6D1C5B7DF7FF78E075C",
INIT_37 => X"5EF005560B55F7AA800AAF7AA954AA00042AAA20000000000000000000000000",
INIT_38 => X"ABEF057D68F5F5A00021EF55042AAAA007FD5555AAFBD7545FBB8020A3F7AE97",
INIT_39 => X"7DF55D7AABFF5428ACA8F45A6C1E8F5EFF84165EFF7802BAB0A2FFEAABA557BE",
INIT_3A => X"CA8AA80800020AAF7FBFFFEF04552ABFFFF841FFE75CA882108202E974AAF7D5",
INIT_3B => X"00151FF0C57401E5F3D1E00A1A884174A8FFAEBFEB0A2D55541051555694F002",
INIT_3C => X"2AA801455D7FE8BFFF680800FFF7AAA155F595542455512A975455D3AA8A0055",
INIT_3D => X"5D79FCAF774AE005BE7895554005D2A8A0B882FFFFE10AAAAAB755A66B6AF56A",
INIT_3E => X"00000000000000000000000000000000000000C3BC1000FF8409000512AEABFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(2),        -- Port A data input
DOA(0)   => data_read_a_lo_256(2),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(2),        -- Port B data input
DOB(0)   => data_read_b_lo_256(2),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_3_14 : RAMB16_S1_S1
generic map (
INIT_00 => X"210C00A20020000108430020001600B8156021104940741B3530400E02B92203",
INIT_01 => X"014C9BCA58B1296D24A402C992500B69404040028804A0080A000416A8D90A08",
INIT_02 => X"C12026A484318004404405C9C66E331352180D468B8203980300204442E02B34",
INIT_03 => X"04000748D60D24648D60524C88804D0215011020D15018148040C10A70E1D58C",
INIT_04 => X"18283333240FE41244187308C9104D70944852640901083801750EB0A418C220",
INIT_05 => X"0613142D01912CC2A1B4140528348900C612A104201C689044340ED413A07649",
INIT_06 => X"119000034019881822104C5E68035250A222829710A0A02C18C01A9920842413",
INIT_07 => X"402F00AB0016CA0431800444841020509D038B021230C1990001C644C8273200",
INIT_08 => X"16905000408482088290E8E64010248C4A5AA840C2000110001521F0810A92E7",
INIT_09 => X"0003CE6581BD016342A951AB146C4480530C3B2A8088D3542651670200C1826A",
INIT_0A => X"00735D36209A8A20020894004284B660821030C8990467401218004041020002",
INIT_0B => X"512445B740457154562F957CC08B00093700080D0A4851001D8302D20A0A1530",
INIT_0C => X"00508650008008021021A40861021840869021A408610218C0869810D6043095",
INIT_0D => X"1C8508438450801043A08090380A8834207007022209038080190000999C8F84",
INIT_0E => X"000400200000C0002A48A206204C4205F3304B33004C0041006240140A1C310A",
INIT_0F => X"0000080040000083800400000100000000008400018040000100080000510100",
INIT_10 => X"0001000000000800000244040000020000000100002A0080000200100000A702",
INIT_11 => X"000000000020000000200000080002C000800008000000000022000006808000",
INIT_12 => X"0000000000000A2281000000000040A3810000000000402001400000022002A0",
INIT_13 => X"000000000004200001C0400000000010200001C0400000000010000004490010",
INIT_14 => X"0001070004000000000000060000104C08000000000000001000000903008000",
INIT_15 => X"CC004050CA0C00020220200070040000010401C4000000000000000000100008",
INIT_16 => X"4310E4310A4210A4210A4210A4210A4210A8D0830A68010001B4DA881048061C",
INIT_17 => X"21084290A4210A4210A4210A4210A4210A4210A4210E4310E4310E4310E4310E",
INIT_18 => X"90A421084290A421084390E4310C4390E4310C4390E4310C4290A421084290A4",
INIT_19 => X"015303C0C78C706428A14C586291000A044001FFE000003FFC004290A4210842",
INIT_1A => X"2492492492492492492492492492492492410410410410412821600001249249",
INIT_1B => X"51A8D46A351A8D46A351A8D46A351A8D46A351A9D4EA753A9D4EA753A9D49249",
INIT_1C => X"FFFFFFFFFFFFFFFC00000000000000000000000038F56351A8D46A351A8D46A3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"55AB02055AB0207FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"420000000000000000000000000000000000000000000000007FFFAB57FFFAB5",
INIT_28 => X"A800BAFFAE9554508002AA00AA843DF55FFAA955EFA2D168B55557BEAA000055",
INIT_29 => X"002AB55AAAA955EF005568A00087BE8BFFA2D155410AA8415555087BFFF55A2A",
INIT_2A => X"AAABFF5508003FF555D0002145552ABFEBA007FC21EF007FD75FFAA841541008",
INIT_2B => X"082EBDEAAA2FBEAABA5D7FC0155005168B455D042AB45F7FFD741000042AA10A",
INIT_2C => X"FF7FBEAB55F7AABDEBA5D7FC2010A2D1575FFF7AA975555D2E80145F78415545",
INIT_2D => X"EF5555554AA087BC01FFFFAAAAB55552A954BAFFFFE8B55552EBDE00F7AEAABF",
INIT_2E => X"000082E820BAA2FBEAB5555557DF55A2AEBDF555D2E954BA002EAAABA002A821",
INIT_2F => X"FB7D5D7FEAA3808554203A000000000000000000000000000000000000000000",
INIT_30 => X"1557D1475FAF45BEAA800AAFFAA95578080038A2AA28E3AF55E3A0BA5D7AADB6",
INIT_31 => X"BD55D7BE80004AA1E8E2AB55B6A0925D7085F6AA10087FEABD7AAD57AEBAB68E",
INIT_32 => X"F5D0438140E2FA38B6AEBFF6D1D04AAFFA41040017D5D20B8EAA007FC51C7A2F",
INIT_33 => X"D0A901FFFF801557D1C20B8EAAA2FBE80AA557BE8B6D5D5FFABEF49002FB55FF",
INIT_34 => X"5D20BDE00EBAAA8BC7EBDFEAFEFAB8ABAE925D21C7010EADB525D7FFAE975C75",
INIT_35 => X"F002EADA921420871D74971D24820875C21D5EB8AA8FFF012A954BAFFF5EFB45",
INIT_36 => X"000000000000000000001C24820BAB6FFEFB6D555578F7DB6A0BDF7DEB8E125F",
INIT_37 => X"B55A28408145AAFFFFFFF5D7FEAABA0051400A20000000000000000000000000",
INIT_38 => X"AB55FAD568AA2AFAE975EF555168B55F7AA800BAF7AA955EF00042AAA2A2AEAA",
INIT_39 => X"2AAAA007FD55558A7BD7145FBB8020A35D2ABEF55F7800015F087FEAA00007FE",
INIT_3A => X"968F575D003FF55F7D5420BA5D2ABFEAAF7AE9DFF759A82AEF70800021EF5504",
INIT_3B => X"FFD5145FBAC9755F05040255FFD84175EF55002AAB0A2FFEAABA557BEA3EF057",
INIT_3C => X"82E974AAF7D57DF45552A3FF10AA8429F45A7D5EAF5FFBAEAAA10554155400AA",
INIT_3D => X"FF843FFE77C80825BC052ABFE10550415557085540000005156155FE90A8F5C0",
INIT_3E => X"00000000000000000000000000000000000005500020AAF7FBFFFEF04552ABFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(3),        -- Port A data input
DOA(0)   => data_read_a_lo_256(3),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(3),        -- Port B data input
DOB(0)   => data_read_b_lo_256(3),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_4_14 : RAMB16_S1_S1
generic map (
INIT_00 => X"A108400020612C80284210081034849800A00030300004833522C82D04A16002",
INIT_01 => X"2043998A1839284D1CA0650E1E504368403008418984014902030806A0D10200",
INIT_02 => X"C120042200000000044441CE01E80F00A49043118680008002000000026208E4",
INIT_03 => X"040001020019200020011209CC0164C060000000690111040144800042F5C403",
INIT_04 => X"7029AF0F81A00010CCA47700CC513CAC0D0B8E02010740E19754080108988021",
INIT_05 => X"02139405007133C0712244CD20F20105D583000020E9892201D304D42A9835E1",
INIT_06 => X"9190440300078002014405D9EE814C0284A883B6D7038AE079059B7800048092",
INIT_07 => X"000100AA0004408000000004840400008D200102503000782000C00C8025C000",
INIT_08 => X"00728A00408403220811991E02120C044058080004000001101121F220000260",
INIT_09 => X"811001E1185B38AD23C3707AD46440818F3CF80EC423CA7D01D123C80200816A",
INIT_0A => X"45810810A01B40216361056D6150F41200280001900439001FD8A00041400000",
INIT_0B => X"11FC88076266E800D605402962A820211500024808010512C40106D222223B14",
INIT_0C => X"0408804116040B02C02C500B0C02C100B0C02C100B0402C300B0401618058611",
INIT_0D => X"040200050200501301208482200D00D0A0408402C4282200A84800009B878680",
INIT_0E => X"00000020000100024AC88300300060090F0D830F00025400300204D018000804",
INIT_0F => X"8000000040000206A2000800000000000000950002E010000000080000588040",
INIT_10 => X"0000000000000808000554000200000000000100006D0020000000100000BB00",
INIT_11 => X"0000400000000000002000001A0002504001000000000000002280000D800800",
INIT_12 => X"0800000000000E2C802000000000408D801000000000408012440000200110A0",
INIT_13 => X"000000000004680003A0040000000010280003800800000000102800000B0000",
INIT_14 => X"000005C0002000000000000620000158000010000000000010A0000B00000200",
INIT_15 => X"C30146200400104002602600400000000294004000000004000000000010001A",
INIT_16 => X"0080200000008020000000802000000080080000004090014134DA101288C6DB",
INIT_17 => X"0802000000000401806010040180601004018060100000802000000080200000",
INIT_18 => X"8060180601004010040080200802000000000000802008020000000000008020",
INIT_19 => X"C0A28A063807E0500014063450404882846FFE000003FFC00000010040100401",
INIT_1A => X"AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA28A28A28A28A2934C8D0CCD145144",
INIT_1B => X"68341A0D068341A0D068341A0D068341A0D068351A8D46A351A8D46A351AAAAA",
INIT_1C => X"FFFFFFFFFFFFFFFC0000000000000000000000001FE32068341A0D068341A0D0",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"408102040810207FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"800AA00000000000000000000000000000000000000000000040810204081020",
INIT_28 => X"168B55557BEAB4500554200000557FE10FFFBEAA10007FD7410FFAA97555082A",
INIT_29 => X"55574105D2A800AA00043FEBA5D7FEAA00007BE8AAAAA843DF55FFAA955EFA2D",
INIT_2A => X"57BC00AAA2FFEAAAAAA8415555087BFFF55A2AA800BAFFAE9555508002AA0000",
INIT_2B => X"A2AA955EF005568A00087BE8BFFA2D17DE1000517FE10AAAAA8AAA002E975455",
INIT_2C => X"FAA8417410A2D140000F7FBC2010A2D157400AAAE974AAAAAA974BA08002AB55",
INIT_2D => X"EFA2AABDEAA087BEAAAAA2FBD54BA080002145552ABFEAA007FC21EF007FD75F",
INIT_2E => X"00055042AB45F7FFD741000042AA10AAAABFF5508003FF55F7D568A00552EA8B",
INIT_2F => X"5400F7A49057D0824850B8000000000000000000000000000000000000000000",
INIT_30 => X"3AF55F7A0925D7AADB6FB7D5D7FEAB7808554203A145178E00FFFBE8A101475D",
INIT_31 => X"A9557D080038AAA145157428492E8008200043FE925571EFA380871C7028A28E",
INIT_32 => X"AEA8A9200249056D4175C5092AAF5FDA38BE8E1557D1475FAF45BEAA800AAFFA",
INIT_33 => X"AA4954281C0E2FB55B6A0925D7085F6AA10087FEABD7AAD57AEBA08517DE00AA",
INIT_34 => X"007FC51C7007BD55D7BE80004AAFEDB42028EBFBC2028BED152438AAA092492A",
INIT_35 => X"AF7DF6AA00412EAABFFAA803DEBA0875EDA80BEF1C743840040017D5520B8EAA",
INIT_36 => X"0000000000000000000041002FB55FFF5D0438140E2FA38B6AEBFF6DBE84AAEB",
INIT_37 => X"A00FFFFEAA105D5155410FF84021EF0800154B20000000000000000000000000",
INIT_38 => X"DEBA0851574B2AAAEAAB55F78400145AAFFFFFEF5D7FEABFF0051400A25D5568",
INIT_39 => X"68B55F7AA800BAF7AA955EF00042AAA25555410BA082E8201000043FE005D517",
INIT_3A => X"568AA200557DE00AAAAAAA000804001FF005575408AA557FEB2FFAE975EF5551",
INIT_3B => X"D1550AAAA8002010F2AC154B25F2ABFF55F7800015F087FEAA00007FEAB55FAD",
INIT_3C => X"800021EF55042AAAA007FD5555087BD6145FAAC000A2A6FBC00BAAAFBC00BAF7",
INIT_3D => X"F7AEBDFF779A82AA43F7FBE8A00082EA8BFFAA843FEBA08517DE00F3F9574B30",
INIT_3E => X"000000000000000000000000000000000000008003FF55F7D5420BA5D2ABFEAA",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(4),        -- Port A data input
DOA(0)   => data_read_a_lo_256(4),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(4),        -- Port B data input
DOB(0)   => data_read_b_lo_256(4),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_5_14 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50DF4A0791B3FCB694379283C81FD996A091832102004A336A20E03C040C002",
INIT_01 => X"805FBDC69830A84D5C6A60000C34C26841280A00084000C8C212892EEAD53235",
INIT_02 => X"3B2026B578918E640A4F01CF8011FF0002080000082CA9998276DF7772C7C80D",
INIT_03 => X"37134108420D700084205702A4008A1D9100002171C0E0051554D93A11F5D140",
INIT_04 => X"8A41A0FC03A56DA000425A819410E3816C086198A388B702A8CA1210844A0C4C",
INIT_05 => X"B1808A062E8BC835F5E84532D708238A282F00A9291224800A2861490343082C",
INIT_06 => X"903FB8483A90581859050424100940825C6184401CDC451B860A6507160C4100",
INIT_07 => X"D26F068BCC96CDF8918E640E96D1A3469D6300E2FFEA27F8E4D23248130E259C",
INIT_08 => X"0BFA82E568442B2A082C0A7E3014250D49DA37A2420619000002AFF48D1222E5",
INIT_09 => X"3F005001E40969289429360416DCD1C46083030604B1CA20C03DF83B0A2C60A5",
INIT_0A => X"14613C71005A10492B888120288F480D58858449026145B3830F449449062B4F",
INIT_0B => X"11AC04934AC648BFD727C031E64170A137D5AA5C3E4B0F8A3C58C34C002290E3",
INIT_0C => X"CA29C6CC50384B6AC6AC86AB31AACA6AB39AAC86AB39AACA6AB3055643559C31",
INIT_0D => X"C673E33CF28F38603855401985228A0614BD30A0A2819852011E5AC2B87F9182",
INIT_0E => X"FF87C002F87A803E460B2516510CA594FF0044FFA4B08BAC4BB2CD0F09CF84E3",
INIT_0F => X"0DFF0F8005F0F5100DFFF5E15D06101C55EB29F1E00BE53FE1F000BE1E802F94",
INIT_10 => X"F12F0380231F17D78FC029FFF58D9A70380230F2FE0017C37FC3E0017C3D005F",
INIT_11 => X"FC7F023C0CA700125C0F8F7E43F1F001BFFE7C69E01804E1E7CCF8FC003FF5F1",
INIT_12 => X"023E00017C1FC1A4BFD82C3081C5BD27BFE30C3081C5BD00C02365D645CEEF5B",
INIT_13 => X"61E0042787F181E9C1EFD8CB8120C5AF41E9C18FD60F0C20666F41E9F009FFFD",
INIT_14 => X"7A7C077FFF404F80005F07F187A7D14BFFC96111C048278DEB074F9930FF9D80",
INIT_15 => X"C064014B8B652E2B3120C81284641D3E8DBF7D636FE860190700132C1F0EFB80",
INIT_16 => X"38CE1384E3384E338CE138CE1384E33C4E3ECE32E128882551349A1CBAA44103",
INIT_17 => X"84E3384E3384E3384E338CE138CE1384E3384E338CE138CE1384E3384E338CE1",
INIT_18 => X"CE138CE138CE138CE1384E3384E3384E3384E338CE138CE138CE138CE1384E33",
INIT_19 => X"F5E5BB4E7F7B9DB7FF3A1B6DB7E8410A8C000000000000000000384E3384E338",
INIT_1A => X"BEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEF9F7CFDFDDCF3CF3D",
INIT_1B => X"BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEFBEF",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000001711C7BBDDEEF77BBDDEEF77",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"FDFFF00000000000000000000000000000000000000000000080000000000000",
INIT_28 => X"FD7410FFAA97410082A800AAAAAE955450055421FFFFFBC0010AAD5574BA557F",
INIT_29 => X"7FD74000055574BA5D7FD7555A2D5575EF55517FF5500557FE10FFFBEAA10007",
INIT_2A => X"0002AABA5D2ABFFFFAA843DF55FFAA955EFA2D168B55557BEAB5500554200000",
INIT_2B => X"5D2A800AA00043FEBA5D7FEAA00007BC00AAAAAEBDF45A28428B45FFD168BFF0",
INIT_2C => X"5080028A00A2FFFDE00F7D57FEBAFF80174BAAAD1555EF555555555005557410",
INIT_2D => X"BA5D2E821FFA2D5554BA557BD75FFAA8415555087BFFF55A2AA800BAFFAE9555",
INIT_2E => X"00000517FE10AAAAA8AAA002E97545557BC00AAA2FFEAAAA082A97545F7D5420",
INIT_2F => X"7010BEDF524AA5571FDFEF000000000000000000000000000000000000000000",
INIT_30 => X"78E00EBFBE8A101475D5400F7A49043D0824850B8A2AE9756D145B401FFFFFFC",
INIT_31 => X"FEAB7D0855420BA1471D74380851524BA5571D757DB6D5525EF555178F6D1451",
INIT_32 => X"8A28B6DEBDF6DBEF1C0A28AAA5524BFFFFA28E3AF55F7A0925D7AADB6FB7D5D7",
INIT_33 => X"5555057D145152428492E8008200043FE925571EFA380871C7028B6AEBDF45B6",
INIT_34 => X"BEAA800AAFFAA9557D080038AAAA2FBF8E10EBD578EAAFF8415482BED1555EF5",
INIT_35 => X"81C209256DFFDF420BA552A821FFB6DF574A85575C55EFBE8E1557D1475FAF45",
INIT_36 => X"0000000000000000000008517DE00AAAEA8A9200249056D4175C50920875FDA3",
INIT_37 => X"5FF5D7BC21EFF7FBD7400F7FBC00BA55557DFF70000000000000000000000000",
INIT_38 => X"01FF5D5568BE7555568A00AAFFEAA105D5155410FF84020AA0800154B2AAAA97",
INIT_39 => X"00145AAFFFFFEF5D7FEABFF0051400A25551554BA0051400BA5551575EFF7D14",
INIT_3A => X"1574B2FFAABFF45FFAAAABFFAAFFFDFFF552EA8AAA55043DFF7AAAEAAB55F784",
INIT_3B => X"8002410FFD5575EF5555421E75555400BA082E8201000043FE005D517DEBA085",
INIT_3C => X"FAE975EF555168B55F7AA800BAF7AA955EF00002AAA2A2FBE8A00A2D16AAAAFF",
INIT_3D => X"0055554088A557FEB25D00021FFFFFFC00BA552A821EFFFFFD74BA5D51575F7F",
INIT_3E => X"000000000000000000000000000000000000000557DE00AAAAAAA000804001FF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(5),        -- Port A data input
DOA(0)   => data_read_a_lo_256(5),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(5),        -- Port B data input
DOB(0)   => data_read_b_lo_256(5),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_6_14 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10800B0061A01002840002C03002818000402322520070B313301C4389B2082",
INIT_01 => X"250041CA3839684D18A160000C52426841000000090800090210080008110200",
INIT_02 => X"0020042080010000044654C0000C008010000000001020900200200002620814",
INIT_03 => X"060881021088200021080200E4000A0891000020610111500104C00000F14400",
INIT_04 => X"0880000100000002000052288144004281C050400100280000C8100000080001",
INIT_05 => X"928080840001100A08009000280201000850E022401400002028214043410820",
INIT_06 => X"10100518090012122100C808049310002040000410A0001400000200120840D2",
INIT_07 => X"000100800004400001000000860408108C22000A502010074120044800040001",
INIT_08 => X"50000040D0C4E2088003FD01C01004044058082004000000000121F020408244",
INIT_09 => X"00BF17E9001205A5204911F814444080400100020000D200DFD16400C2A40AA0",
INIT_0A => X"04611C17849000022862A1596C8B5DF04834948900000100220C244840000880",
INIT_0B => X"03AD0413424E4044D665C070C22602291504400D084915020448114080201000",
INIT_0C => X"5E08864011088B22D22C008B0022C408B1022C208B0822C608B1111600458010",
INIT_0D => X"4251A12CD28A300429688001000800000020280204001000A00804309A002182",
INIT_0E => X"0000000280402400420800000000006200FC10002442042429324294014E8CA7",
INIT_0F => X"A40000000500800840000800000000000002280018001480000000A010100052",
INIT_10 => X"00000000000004C2003000010240000000000000680800290000000140202000",
INIT_11 => X"2000C0000000000000000442000001080001000000000000010C000280001804",
INIT_12 => X"08000000000801C300A010000000156000902000000015101200002800000000",
INIT_13 => X"000000000101800038002408000000094000386028040000000940000ED40000",
INIT_14 => X"0003B000002000000000020180002A24005010000000000023000060C7000A40",
INIT_15 => X"3F0280090321000040A410C28108000160008094000810040000000000002300",
INIT_16 => X"284A5284A728CA5284A528CA728CA52C4A5A0A32A300940101349A0408240818",
INIT_17 => X"9CA1294A329CA5284A728CA7284A5284A728CA5284A528CA728CA5284A728CA7",
INIT_18 => X"CA3294A129CA3294A129CA1294A329CA1294A3294A129CA3294A129CA3294A32",
INIT_19 => X"F5F78BCE7F8FF0F4FA955F7CF7F40A80145D55555556AAAAAAAAA94A329CA129",
INIT_1A => X"8E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E39B6CEDECDDF7DF7D",
INIT_1B => X"F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE38E3",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000001A1A33F9FCFE7F3F9FCFE7F3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"555FF00000000000000000000000000000000000000000000080000000000000",
INIT_28 => X"BC0010AAD5574BA557FFDFFF087BFDF45F7AA974AAAAAA97555F784174BAF7D5",
INIT_29 => X"515555508043FE00F7AA97555A2FBD7410AA8428AAAAAAE955450055421FFFFF",
INIT_2A => X"7D1575EFFFAA9555500557FE10FFFBEAA10007FD7410FFAA97400082A800AA08",
INIT_2B => X"0055574BA5D7FD7555A2D5575EF55517FF55A2AA97400552AAAB45082E80155F",
INIT_2C => X"500554200000003DE10FFD5401FFF7AAA8A10082EAAB45A2FFC2000007FD7400",
INIT_2D => X"10AA803FE105D516AABAFF843FFFFAA843DF55FFAA955EFA2D168B55557BEAB5",
INIT_2E => X"000AAAEBDF45A28428B45FFD168BFF00002AABA5D2ABFFFF087BD5545007BFDE",
INIT_2F => X"256DEB84104BAFFD1525FF000000000000000000000000000000000000000000",
INIT_30 => X"9756D145B401FFFFFFC7010BEDF524AA5571FDFEF1C7BFFF55FFA095482B6A49",
INIT_31 => X"4904380824850381C5B5057D1C003DE28F7A49057DAAF5D2428A2842AAAAA2AE",
INIT_32 => X"2AAFB451C2A8017DE3DF525FFFFA49756D145178E00EBFBE8A101475D5400F7A",
INIT_33 => X"2F1C50381471D74380851524BA5571D757DB6D5525EF555178F6DAAA49542841",
INIT_34 => X"AADB6FB7D5D7FEAB7D0855420BA1C0E3FE00E3DB471EFE3AAAAA00082EA8B6DA",
INIT_35 => X"F1C7BD057D1C71FFE10A28038E1049516AAB8FF8428FEFA28E3AF55F7A0925D7",
INIT_36 => X"00000000000000000000B6AEBDF45B68A28B6DEBDF6DBEF1C0A28AAA5524BFFF",
INIT_37 => X"F55F78017400F780001FFAA84000AAFFD1401E70000000000000000000000000",
INIT_38 => X"20BAAA8428AA2AAAA975FF5D7BC21EFF7FBD7400F7FBC00BA55557DFF7557BFD",
INIT_39 => X"EAA105D5155410FF84020AA0800154B2557FC01EF55043FEAAFF80021EFA2D14",
INIT_3A => X"568BE7AA80174AA082ABDF555D2A821EFAAFBC01FFF780155F7555568A00AAFF",
INIT_3B => X"AEA8A10082EA8BEFAAD5554B25551554BA0051400BA5551575EFF7D1401FF5D5",
INIT_3C => X"AAEAAB55F78400145AAFFFFFEF5D7FEABFF0051400A25D2EBFE10AAFFD55EFA2",
INIT_3D => X"552EA8AAA55043DFF7557BC01EF55557DE00AA842AA0000516AABAFF8428BE7A",
INIT_3E => X"0000000000000000000000000000000000000FFAABFF45FFAAAABFFAAFFFDFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(6),        -- Port A data input
DOA(0)   => data_read_a_lo_256(6),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(6),        -- Port B data input
DOB(0)   => data_read_b_lo_256(6),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_7_14 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10844B00482258A2842112C02450418800002300500030B313300C418992002",
INIT_01 => X"000009CA3839684D1CA0E0000E51424840000000080000080200080008510204",
INIT_02 => X"0120042086010000044600C00008000004100000000260900200000002402004",
INIT_03 => X"8628A10000082400000002408400080011000000610008000208C00000E14400",
INIT_04 => X"0911800100A000000000524084000040000050001140200100C8100000080102",
INIT_05 => X"0300812401011000000000002000114008008060441000000020024093000000",
INIT_06 => X"9190431C0D4010100000880804010010800000041080081000000200010424B2",
INIT_07 => X"000100AA0004408601000004860000008C02000A103010006928040800062481",
INIT_08 => X"84000048D484C20888000A0002120484C048007004000000000021F000000244",
INIT_09 => X"00A06009881201A520491004106C48A04040002400A15A208001650004001020",
INIT_0A => X"C99E1060201002044809C1040140A001004808810000459033189C0A400118A0",
INIT_0B => X"102000024040484050050041648A0041140C500B08821054C000264120000400",
INIT_0C => X"0404A083260E0832132011880462011880462051881462051881D31018C40620",
INIT_0D => X"0001000080001000813094801A8F80F00A600B52602801A88848011118003700",
INIT_0E => X"000003C007C002808228010410082042C000C000000004001002000400040002",
INIT_0F => X"A4000007800F80C840000800009864038A1200081C0014800000F001F0200052",
INIT_10 => X"00002C0E00E0E4004038000102400002C0E00E0D20100029000001E003E04000",
INIT_11 => X"2000C04031100E0403D0700300080908000100000661801E1900040380001804",
INIT_12 => X"0840878083E8003780A01043203A101780902043203A10082410082880000000",
INIT_13 => X"0601E0187900181035E0240806483248181035E0280410C8198818100DDD0000",
INIT_14 => X"0403774000201021E020FA006040376C00501022131210722060806D47000A40",
INIT_15 => X"00928A0002000110888600C032128201519480D40009902430160403E0E00506",
INIT_16 => X"01000000020080601802000000000405000A0020020081014134928820480010",
INIT_17 => X"0802018040000000006018020080200804010000000000806018020080000004",
INIT_18 => X"0000000001806008020000001006008020080001004008020080201004000020",
INIT_19 => X"0000000000000000000000000000400A004618618618C30C30C3000020180600",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000000B0840000000000000000000",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"1555500000000000000000000000000000000000000000000080000000000000",
INIT_28 => X"A97555F784174BAF7D5555FFF780155EFAAAEA8ABAAAFBFDE0055556AA005D04",
INIT_29 => X"55555EFAAFFFDFEFAAAAAAB455D556AA00FFAE95555087BFDF45F7AA974AAAAA",
INIT_2A => X"02EAAAAA082EA8A00AAAE955450055421FFFFFBC0010AAD5574BA557FFDFFF55",
INIT_2B => X"08043FE00F7AA97555A2FBD7410AA8428AAA557BFDFFF55003DFFFF7FBEAA000",
INIT_2C => X"0082A800AAF7AE975FFA28000010552EBDE00007BEAAAAA2D140000085155555",
INIT_2D => X"45087FEAB455D516AB55557BD55FF00557FE10FFFBEAA10007FD7410FFAA9740",
INIT_2E => X"000A2AA97400552AAAB45082E80155F7D1575EFFFAA955555D51574AAAAFFD55",
INIT_2F => X"AE105D556AA10410E17555000000000000000000000000000000000000000000",
INIT_30 => X"FFF55FFA095482B6A49256DEB84104BAFFD1525FFFF8E175C7A2AAAAA82A2F1F",
INIT_31 => X"F524AA5571FDFEF415B575D7AAF1FFFD7AAAAAFB7D495F6AA10E3AE905551C7B",
INIT_32 => X"003AFEFEBFBEAA001C2EA8A821C2EAAA00A2AE9756D145B401FFFFFFC7010BED",
INIT_33 => X"EDB470101C5B5057D1C003DE28F7A49057DAAF5D2428A2842AAAA497BFAFFF49",
INIT_34 => X"1475D5400F7A490438082485038F7A4905C7A28A070384120BDE100075EAA82B",
INIT_35 => X"D495150492BEF1D2555087BE8B7D555F6AB57417BC05D7145178E00EBFBE8A10",
INIT_36 => X"00000000000000000000AAA495428412AAFB451C2A8017DE3DF525FFFFA49756",
INIT_37 => X"555A2AEA8A10AAD568A00555168A10002E9754D0000000000000000000000000",
INIT_38 => X"8A10AAAE8215D557BFDF55F78017400F780001FFAA84000AAFFD1401E7FFAA97",
INIT_39 => X"C21EFF7FBD7400F7FBC00BA55557DFF7007BD5555AAD57DF55AAAEBDFEF007BE",
INIT_3A => X"428AA2007FE8BFF080028BFFAAFFEAA105D2EAAA005D2AAAA18AAAA975FF5D7B",
INIT_3B => X"043DE0000516AA10F7FBD7408557FC01EF55043FEAAFF80021EFA2D1420BAAA8",
INIT_3C => X"55568A00AAFFEAA105D5155410FF84020AA0800154B2FF8402145A2AA954AA00",
INIT_3D => X"AAFBC01FFF780155F7005140000FFD140145007FE8BEF557BEAB55087FC215D5",
INIT_3E => X"0000000000000000000000000000000000000AA80174AA082ABDF555D2A821EF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(7),        -- Port A data input
DOA(0)   => data_read_a_lo_256(7),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(7),        -- Port B data input
DOB(0)   => data_read_b_lo_256(7),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_8_14 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00000648E2840112C00000418000002700500030B3132000400812082",
INIT_01 => X"100008480009004C04A100000252024840000000180800080200010040110204",
INIT_02 => X"0020042000490000004600804008000005100000000024900200000002400004",
INIT_03 => X"0A0C33400008082400000080A4004B0891000020610112000040C00000E5C000",
INIT_04 => X"18800001000000000000512080000040800150400824280110C8100000120200",
INIT_05 => X"908084A10100100200004080280008240810802206940000012C214451610800",
INIT_06 => X"81B000080860109021400008040000202048020414A0021400040200322824C1",
INIT_07 => X"000000080004408049000004860000008402001A50208000630C040800062483",
INIT_08 => X"440000428644212280800A00021004044048002124000000000021F000000244",
INIT_09 => X"00004009001001010008100414644410400102228000D20080114502006409A2",
INIT_0A => X"000051312000042200294429148A4801C80C8C81000045907118040340020832",
INIT_0B => X"4020000240404140004D0544C4AA0001150410090302500011C813428A000400",
INIT_0C => X"46501090008820240240409000240009000240009000240009000120204808A5",
INIT_0D => X"42D1A168D09A301468402480004780F00140080860280004085904309A002196",
INIT_0E => X"00783FC00044340242280000000000020000C0000442106419120004034685A3",
INIT_0F => X"8000F07F800088A80000081EA2F9EC0000064004081010001E0FF00011104040",
INIT_10 => X"0ED0FC7E00000422201080000202658FC7E0000021882020003C1FE000222080",
INIT_11 => X"018059C3F350FE0C00000002A0040500000103961FE780000110010090000800",
INIT_12 => X"FD41FF80000830200021C1CF600012200010D1CF600012121600100810000004",
INIT_13 => X"9E1FE000010A1802100004343ED8000898021000087073D80008980200800002",
INIT_14 => X"0080200000BEB07FE00002086008020000209AEE3F300000246020200000620B",
INIT_15 => X"0088881903210000440610C8000A808040000208901786E4F0FE0C0000000166",
INIT_16 => X"685A1685A769DA368DA368DA769DA36CDA121A11A141800011309284002C0810",
INIT_17 => X"95A5685A1685A5695A368DA368DA769DA368DA368DA7695A1685A1685A5695A1",
INIT_18 => X"5A1695A568DA368DA369DA768DA1685A1695A5685A168DA369DA768DA368DA16",
INIT_19 => X"A4028A0A543EBC57A10A1E75D64108080468618618630C30C30C69DA5685A168",
INIT_1A => X"9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7BF3CCD8DF5B2DB2C",
INIT_1B => X"F87D3E1F4F87D3E1F4F87D3E1F4F87D3E1F4F87C3E1F0F87C3E1F0F87C3E79E7",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000006A6D4F87D3E1F4F87D3E1F4",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"155FF00000000000000000000000000000000000000000000080000000000000",
INIT_28 => X"BFDE0055556AA005D0415555080000000087BEAA10F7803DE00FFAEBFFFF0800",
INIT_29 => X"2AA8AAA557FC0010F780154105D7FC2145005155555F780155EFAAAEA8ABAAAF",
INIT_2A => X"7FFFFF55AA80155FF087BFDF45F7AA974AAAAAA97555F784174BAF7D5555FF55",
INIT_2B => X"AAFFFDFEFAAAAAAB455D556AA00FFAE95555AAFFE8A00552EBFE00F7D17FF45F",
INIT_2C => X"A557FFDFFF5504000AAAAAAA8B55F7D140010552E821EFAAAABDF555555555EF",
INIT_2D => X"55AA8028A00A2D57FF45557BE8A00AAAE955450055421FFFFFBC0010AAD5574B",
INIT_2E => X"000557BFDFFF55003DFFFF7FBEAA00002EAAAAA082EA8A00002AA8A10F784021",
INIT_2F => X"FE10F7AEBAFFF080A175D7000000000000000000000000000000000000000000",
INIT_30 => X"175C7A2AAAAA82A2F1FAE105D556AA10410E17555080E000280071E8A00EB8E3",
INIT_31 => X"4104BAFFD1525FF492EA8AAA5571C2000FF8A17400557FC015514555757DFF8E",
INIT_32 => X"2ABDE10EBDF7AF6DE3FFF8F7DB68A105D71C7BFFF55FFA095482B6A49256DEB8",
INIT_33 => X"AA0BDF6D415B575D7AAF1FFFD7AAAAAFB7D495F6AA10E3AE90555A2FBE8A3849",
INIT_34 => X"FFFFC7010BEDF524AA5571FDFEF550E00082B6A0AFB55F7D1420104124821D7A",
INIT_35 => X"01C2EA8A00F7800017DA2842FA00B6D578F6D557FFDA00A2AE9756D145B401FF",
INIT_36 => X"00000000000000000000497BFAFFF49003AFEFEBFBEAA001C2EA8A821C2EAAA0",
INIT_37 => X"0BA08556AA00AAAABFE00F7AEAABEF082E955450000000000000000000000000",
INIT_38 => X"21555D51575EFFFAA97555A2AEA8A10AAD568A00555168A10002E9754D082E82",
INIT_39 => X"17400F780001FFAA84000AAFFD1401E7082EAAABA5D5140010F7AE974105D7BC",
INIT_3A => X"E8215DA2FFE8ABA082ABFE00AAFBEABFFAAFBEABFFF7AA80145557BFDF55F780",
INIT_3B => X"D540000000402145AA843FFFF007BD5555AAD57DF55AAAEBDFEF007BE8A10AAA",
INIT_3C => X"AAA975FF5D7BC21EFF7FBD7400F7FBC00BA55557DFF75D2E82010F7843DF45FF",
INIT_3D => X"5D2EAAA005D2AAAA185D2AAAA10F780021FFA2803DE10FFD16ABFF5D7BFDE10A",
INIT_3E => X"0000000000000000000000000000000000000007FE8BFF080028BFFAAFFEAA10",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(8),        -- Port A data input
DOA(0)   => data_read_a_lo_256(8),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(8),        -- Port B data input
DOB(0)   => data_read_b_lo_256(8),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_9_14 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00018248A2840112C00002C18000002300500030B3132000400812006",
INIT_01 => X"400008000000004C0020000000100248413C0A61590001D90213C10008110204",
INIT_02 => X"01A0042080010000054600C04008000004100000001020900200200002420804",
INIT_03 => X"024003400008012400000010E4004B0891000020610310000144C00000F5C000",
INIT_04 => X"1801800100E000000000510084000040010050020810200000C8900000320200",
INIT_05 => X"918004311104100000000000200008100800002000100000002C234415610820",
INIT_06 => X"81B00008080010100000980804000008800042041080001000100200322C2481",
INIT_07 => X"0000811800044080010000058600000086020002502080006000040800062C80",
INIT_08 => X"0000004001D4618008800A00061004044048002004000000000061F000000244",
INIT_09 => X"000040090802009420409004104444084001022400214A2080014400026401A2",
INIT_0A => X"04000071200000A003CA294140200800C80C8C8100004590111C040040120800",
INIT_0B => X"12210002404848502847040164880021150400080222000200C8034200000000",
INIT_0C => X"4610088010080421021040841021000841021000841021000841010800420820",
INIT_0D => X"42D0A16C529A321068500484000500D10042080040284000084900001A002196",
INIT_0E => X"00000002804000004228010410082002C000C0002400046419120410034285A1",
INIT_0F => X"A00000000500800800000800000000000002290008001080000000A010100042",
INIT_10 => X"00000000000004C2001000000240000000000000680800280000000140202000",
INIT_11 => X"0000C0000000000000000442020001000001000000000000010C800080000804",
INIT_12 => X"08000000000801A7802010000000152780102000000015000600000800000000",
INIT_13 => X"000000000101900011E0240000000009500011E0280000000009500004DD0000",
INIT_14 => X"000137400020000000000201C000136C00101000000000002340002947000240",
INIT_15 => X"0080881901210000000600C280028000419480D4000010040000000000002304",
INIT_16 => X"68DA368DA1685A1685A1685A1685A16C5A121A13A141950051309284A82C0010",
INIT_17 => X"85A1685A1685A1685A368DA368DA368DA368DA368DA368DA368DA368DA368DA3",
INIT_18 => X"5A1685A168DA368DA368DA368DA368DA368DA368DA3685A1685A1685A1685A16",
INIT_19 => X"0157344CCCF48DE68A895C38E2540A8010100000000000000000685A1685A168",
INIT_1A => X"14514514514514514514514514514514514D34D34D34D34D28E1004039248209",
INIT_1B => X"D268341A4D268341A0D069349A0D069349A0D068341A0D068341A0D068345145",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000014D490D069349A0D068341A4",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"EAABA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"03DE00FFAEBFFFF0800155FFAAFBE8B45002A974AAAA803DFFFAA843DF45FFFF",
INIT_29 => X"7BFDE00A2FBD7400F7FBFDFFFA2AEBDE00AAFBEAABA080000000087BEAA10F78",
INIT_2A => X"055401FFF7AEAAA10F780155EFAAAEA8ABAAAFBFDE0055556AA005D041555508",
INIT_2B => X"557FC0010F780154105D7FC2145005155555557BE8BEF007FFDEAAAAD1555EF0",
INIT_2C => X"AF7D5555FFF780154AA5D2AA8A10F7AA974AA082E80010A2AAAAA10552AA8AAA",
INIT_2D => X"BAF7D17FEBAA2AEBDF45002EAAABA087BFDF45F7AA974AAAAAA97555F784174B",
INIT_2E => X"000AAFFE8A00552EBFE00F7D17FF45F7FFFFF55AA80155FF080400145FFFBEAA",
INIT_2F => X"8FC7BE8A3DF7DF7F5E8A92000000000000000000000000000000000000000000",
INIT_30 => X"000280071E8A00EB8E3FE10F7AEBAFFF080A175D7BEF1E8B6D002090482B68E3",
INIT_31 => X"56AA10410E175550871FFE00A2FBD0400FFF5FDFC7B6A0BDE38B6F5E8A92080E",
INIT_32 => X"7BFAE82A2DB555C71C5B451D7FFAAA8A38FF8E175C7A2AAAAA82A2F1FAE105D5",
INIT_33 => X"2AEADA38492EA8AAA5571C2000FF8A17400557FC015514555757D5D71E8BEF14",
INIT_34 => X"B6A49256DEB84104BAFFD1525FFFF84174BA5D20AAA00E3AA904BA142A87010A",
INIT_35 => X"7000400155FFFBEDA82FFD57DEBAAAA0BFF7D0024ADA921C7BFFF55FFA095482",
INIT_36 => X"00000000000000000000A2FBE8A38492ABDE10EBDF7AF6DE3FFF8F7DB68A105D",
INIT_37 => X"BEF080402000F7AAA8B55FFAABDFEFF7D16AA000000000000000000000000000",
INIT_38 => X"FEAAFFD16AA00082E820BA08556AA00AAAABFE00F7AEAABEF082E95545F7D568",
INIT_39 => X"A8A10AAD568A00555168A10002E9754D00517DE00A2FFC2000F7D17FF55FF803",
INIT_3A => X"1575EF555568BEF5D7FE8A10AAFFD55555D7FD5555FFAAA8AAAFFAA97555A2AE",
INIT_3B => X"AE800AA552A97400A2AEBDEAA082EAAABA5D5140010F7AE974105D7BC21555D5",
INIT_3C => X"57BFDF55F78017400F780001FFAA84000AAFFD1401E7FF80174AA5D0028A00AA",
INIT_3D => X"AAFBEABFFF7AA80145080002145F7FBFFE00FFD17FEAAA2803DFEF08043FE005",
INIT_3E => X"0000000000000000000000000000000000000A2FFE8ABA082ABFE00AAFBEABFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(9),        -- Port A data input
DOA(0)   => data_read_a_lo_256(9),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(9),        -- Port B data input
DOB(0)   => data_read_b_lo_256(9),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_10_14 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00018248A2840112C00002C18000202300500030B3132000400992006",
INIT_01 => X"254008000000004C002000000010026840000000080000080200010008110204",
INIT_02 => X"0020042000010000004455800008000004100000000000900200000002400004",
INIT_03 => X"020001021089000021081000C400090011000000610001540104C00000F14400",
INIT_04 => X"0811800101A00002000050088554004200C840000000200080C8100000000001",
INIT_05 => X"030080001000100800009400200000000840E020201000000024024001200020",
INIT_06 => X"81B00008080012120004CC080492500280208004148000100000020020042493",
INIT_07 => X"0000000800044080010000048404081085020002502000006000040800062480",
INIT_08 => X"100202400084410808000A00021004044048000004000000000021F020408264",
INIT_09 => X"010040090002008420401004144440004040022484214A2080110108C2C00320",
INIT_0A => X"04004166A48A0001080000000000080080181881000045901118044040020800",
INIT_0B => X"1201000200484910000F0105602622291404020902005002018002400A022000",
INIT_0C => X"0440001011808020120004801120044800120004801120044800110002400884",
INIT_0D => X"008000440210100041308480800F82F00040180260A808008848000018002104",
INIT_0E => X"000000028040000002280104100820020000400020000440100204100A000100",
INIT_0F => X"040000000500800800000000000000000002280008000400000000A010100010",
INIT_10 => X"00000000000004C2001000010000000000000000680800010000000140202000",
INIT_11 => X"200000000000000000000442000001000000000000000000010C000080001000",
INIT_12 => X"00000000000801C0008000000000154000800000000015000410000800000000",
INIT_13 => X"0000000001019800180000080000000958001800000400000009580002800000",
INIT_14 => X"0000A0000000000000000201E0000A0000400000000000002360002080000800",
INIT_15 => X"0080881000000000000600C28102800060000000000800000000000000002306",
INIT_16 => X"401004010040100401004010040100441020D0030008840051309A90BA884010",
INIT_17 => X"0902409024090240900401004010040100401004010040100401004010040100",
INIT_18 => X"1004010040902409024090240902409024090240902409024090240902409024",
INIT_19 => X"F546890A940FE0D3971243555205428290100000000000000000401004010040",
INIT_1A => X"8A28A28A28A28A28A28A28A28A28A28A28A28A28A28A28A29554199854514514",
INIT_1B => X"2B95CAE532994CA6532995CAE572B94CA6532994CA6532994CA6532994CA28A2",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000002718E72B94CA6532994CA657",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"FDE1000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"03DFFFAA843DF45FFFFEAABA007FC2155F7D155545AA80001EFAAFBEAB45557F",
INIT_29 => X"042AB55FFD168B55AA8000010FFFBE8BFFF78402155AAFBE8B45002A974AAAA8",
INIT_2A => X"AD16AABA002ABDE10080000000087BEAA10F7803DE00FFAEBFFFF0800155FF00",
INIT_2B => X"A2FBD7400F7FBFDFFFA2AEBDE00AAFBEAABAA2FFD741055003DFEFF7AA801FFA",
INIT_2C => X"05D0415555007FD74105555555EFF7FBC0145F78028A00A2D142155087BFDE00",
INIT_2D => X"55AAD168ABA002A975FFF7AEBDEBAF780155EFAAAEA8ABAAAFBFDE0055556AA0",
INIT_2E => X"000557BE8BEF007FFDEAAAAD1555EF0055401FFF7AEAAA105D042ABFF5D556AB",
INIT_2F => X"71D7AAFBEFB455D71F8E00000000000000000000000000000000000000000000",
INIT_30 => X"E8B6D002090482B68E38FC7BE8A3DF7DF7F5E8A92007BC217DEBDB55555AA8E0",
INIT_31 => X"EBAFFF080A175D700042AB7DEBDB6DB55BE8E05000EBFFE8BC7E38E07145BEF1",
INIT_32 => X"0A3DFD7F7A4821D7A2D16FA82142EB8E00080E000280071E8A00EB8E3FE10F7A",
INIT_33 => X"ED1421450871FFE00A2FBD0400FFF5FDFC7B6A0BDE38B6F5E8A92B6FBD541049",
INIT_34 => X"A2F1FAE105D556AA10410E175550071D54104951555D7EBF5C5155E3842AA00B",
INIT_35 => X"8410E2ABD749516FB55BED16FA820820955EFE3AEBDEAAFF8E175C7A2AAAAA82",
INIT_36 => X"000000000000000000005D71E8BEF147BFAE82A2DB555C71C5B451D7FFAAA8A3",
INIT_37 => X"1EFA2FFD7545AAAE97555A2FBFDF455D556AA000000000000000000000000000",
INIT_38 => X"8B45AAAA95545F7D568BEF080402000F7AAA8B55FFAABDFEFF7D16AA00087FC0",
INIT_39 => X"6AA00AAAABFE00F7AEAABEF082E9554500042ABFFA2FFFFF45F7AE97400AAFFE",
INIT_3A => X"16AA00FFFBD5400082EBFF45F78400155A2D57FE00552EA8A00082E820BA0855",
INIT_3B => X"D557555A2802AA10FFD54214500517DE00A2FFC2000F7D17FF55FF803FEAAFFD",
INIT_3C => X"FAA97555A2AEA8A10AAD568A00555168A10002E9754D085155410085557555AA",
INIT_3D => X"5D7FD5555FFAAA8AAA002AAAB4508557DF55F7D17FE000804155FFAAAABDEAAF",
INIT_3E => X"0000000000000000000000000000000000000555568BEF5D7FE8A10AAFFD5555",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(10),        -- Port A data input
DOA(0)   => data_read_a_lo_256(10),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(10),        -- Port B data input
DOB(0)   => data_read_b_lo_256(10),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_11_14 : RAMB16_S1_S1
generic map (
INIT_00 => X"A101C4B05A0034CA2840712C2D001419000002300500030B31B20084EC992002",
INIT_01 => X"90000986B83028491800E0000C26426040000000080000088200080802512224",
INIT_02 => X"1A2004205E010640024D00800008000004100000040EC090820018003241A00C",
INIT_03 => X"28639100000C5C00000045C08400C8001100000061806A001618C03001E54400",
INIT_04 => X"1A800001000009A0804059A190000040400040008058220008C8100000120D4E",
INIT_05 => X"02000E81080250010000002022000058080400000E1200000020004401000004",
INIT_06 => X"819435143F20101010001008040800B8100102041088011100022200000024B2",
INIT_07 => X"90640D280884453E01064002944180008402001295BA100022E4340800062D82",
INIT_08 => X"400000093204802200280A0012160585C1D808D004000000000323F40C102244",
INIT_09 => X"380040098010001100009204107C5950400000220080C200800900020C006827",
INIT_0A => X"80007100004016EA080801010000080D00200081000045B0511D289940103399",
INIT_0B => X"002000024040410A000D0104408810C115D9C008050042400100D04E88000002",
INIT_0C => X"00655010009264201200C7B421ED0C7B421ED0C7B431ED087B43176843DA1085",
INIT_0D => X"0401020080400A10012494881A4F80F209500BB2602881A488485C1318002000",
INIT_0E => X"6619A540124814800228010410082022C00040002020090020220C9600040802",
INIT_0F => X"ACCC334A802491600C587949B6D0141B4CC600D5761B1599865A500490B86A56",
INIT_10 => X"BAC845542056A61686EC81E3A6CB68AA2C622C9A251C352B330CB4A0092170D8",
INIT_11 => X"BCCAD0B5A81536080CC6B21A21B1FC09CB0F1076D4A200B2AD4068F4101639B5",
INIT_12 => X"4D2CC281E31AA0103AB8D5514066380804B268A2E060901204112566F10AC418",
INIT_13 => X"D551443C47281002540B2C9AAAA8662A1152B202AE3554403028115AA88201A1",
INIT_14 => X"548A20A0492A2724A0621620402A020141F172FB182A32AB6845AB6200251BC9",
INIT_15 => X"00C00A000200074044E6801832728080D00A380B753952C4877E0104DDE4D124",
INIT_16 => X"0080200802008020080200802008020480080022020081010124988800400010",
INIT_17 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_18 => X"0000000000802008020080200802008020080200802008020080200802008020",
INIT_19 => X"55062608804180C0B10A42104201400204000000000000000000000000000000",
INIT_1A => X"00000000000000000000000000000000000820820820820801C4149470000000",
INIT_1B => X"0000000000000000040200000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000007E0F0000000000000100800",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"000AA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0001EFAAFBEAB45557FFDE10082ABDF5508557DF45002ABDFFFF7803DE10AA80",
INIT_29 => X"AEBFF45FFAEBFEAA002A801FFF7FFE8A10A28000000007FC2155F7D155545AA8",
INIT_2A => X"2AABFE10082ABFFEFAAFBE8B45002A974AAAA803DFFFAA843DF45FFFFEAABAA2",
INIT_2B => X"FFD168B55AA8000010FFFBE8BFFF78402155AAD155555A28428BFF002ABDE00A",
INIT_2C => X"F0800155FF00557FF45557FC2010002A80010A2842AAAA007BFFF4500042AB55",
INIT_2D => X"FF5D00154BAF7FBE8BEFFFD540000080000000087BEAA10F7803DE00FFAEBFFF",
INIT_2E => X"000A2FFD741055003DFEFF7AA801FFAAD16AABA002ABDE10A2D168A10A284021",
INIT_2F => X"DFC7F78E3FE28B684070AA000000000000000000000000000000000000000000",
INIT_30 => X"C217DEBDB55555AA8E071D7AAFBEFB455D71F8E00002EBDF6D005B78F7D142AB",
INIT_31 => X"A3DF7DF7F5E8A92BEAEBFF7DEBA0BDEAA1C2A801C7E3FFEFA10B68407038007B",
INIT_32 => X"8A28BFF082ABAE10B6AAB8E280820B8FEFBEF1E8B6D002090482B68E38FC7BE8",
INIT_33 => X"07FF8F7D00042AB7DEBDB6DB55BE8E05000EBFFE8BC7E38E07145B6D15756DA2",
INIT_34 => X"EB8E3FE10F7AEBAFFF080A175D708517DF7D497BC5028142A87000A28A2AA920",
INIT_35 => X"0B6DB6AA28A280001FF5D0A10482FFFFEFBC7E3DF42028080E000280071E8A00",
INIT_36 => X"00000000000000000000B6FBD5410490A3DFD7F7A4821D7A2D16FA82142EB8E0",
INIT_37 => X"FEF007BE8BFF5D2ABDF55F7AABDEAAF784154BA0000000000000000000000000",
INIT_38 => X"DE00FF84154BA087FC01EFA2FFD7545AAAE97555A2FBFDF455D556AA00082EBF",
INIT_39 => X"02000F7AAA8B55FFAABDFEFF7D16AA00FFAEBFFEFAA803DEBA5D2E82155A2FBF",
INIT_3A => X"A95545F7D5555FFAAAAA8BFF002AAAA00FFAAA8AAA080028BFFF7D568BEF0804",
INIT_3B => X"2E95400A2AEA8A00007FEABFF00042ABFFA2FFFFF45F7AE97400AAFFE8B45AAA",
INIT_3C => X"82E820BA08556AA00AAAABFE00F7AEAABEF082E9554508557DFFF007BD54BA5D",
INIT_3D => X"A2D57FE00552EA8A00FFFFE8AAAAA80001FF5D2E82000F7FFFFF45AAFFC20BA0",
INIT_3E => X"0000000000000000000000000000000000000FFFBD5400082EBFF45F78400155",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(11),        -- Port A data input
DOA(0)   => data_read_a_lo_256(11),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(11),        -- Port B data input
DOB(0)   => data_read_b_lo_256(11),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_12_14 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50080B01BC002006940202C0DE041196A83183000000023322287E0FC000006",
INIT_01 => X"75400D849830C84C5823E0000C17424840000000080000088200002802153231",
INIT_02 => X"18A026B43ED180040147558040090000061800000C06ED9802768F4472C52005",
INIT_03 => X"2A67E34A528D0524A52850528400C8001100000171C02B550618C91A10E55440",
INIT_04 => X"1BC0000100056C8280825DE98154004300C840800850240080CA921084520A07",
INIT_05 => X"02000F832000500C0000941024000852084060202E100001002000448100000C",
INIT_06 => X"819A1D1C3FE01A1A40045408049A50BA4020C6041090001200006200000000F2",
INIT_07 => X"C26A0719CC96CC6ED18A64019695A854870300FA3968B20068FC06080106249F",
INIT_08 => X"D002024B3E040800008C0A002610240D494A06F3460409000000E3F0AD5282E5",
INIT_09 => X"27A06009200040000400120412445D78400001000410420080218029CC807A27",
INIT_0A => X"18000006848A026F000000000000080000F010C100204593F11A6CDF48003BF8",
INIT_0B => X"000000820040402B28050400400432C9349DF21A31A00ACC0000F04F80020001",
INIT_0C => X"00357804611AE45D05D0833430CD0833420CD0C33420CD0833430668619A1000",
INIT_0D => X"0000000000000A74812DF00E87E80A079F9F90FA0280E87E800C7FF3B8002000",
INIT_0E => X"3B6B0E404D26160682082002000401EA0000C40000800A006002818808000000",
INIT_0F => X"A476D61C809A4DA84272592D6246FC1B17B541F97E1B348EDA93900B2B286C56",
INIT_10 => X"30C669E622DBC325CFD881A962454CFBE5403AB99594362B1DB52720165650D9",
INIT_11 => X"F8D2D39A3745261E4A95A110A3F855000E4B1D32BAB504BB7490FCFF912A3834",
INIT_12 => X"B90E9B018C7530200AB8F8BF41F9A22006B37DC8E1F9A21A70116D4C5080651C",
INIT_13 => X"118780319CCA08AB1001ACDF34B8F1C688AB1002AE3F7B807B6289F368828C4C",
INIT_14 => X"2AF020233376A5ECC016B1A827CDA21160F051DE610A34C50427E6E220323E4A",
INIT_15 => X"0077020000000439FDC05C5806781FAB46095A0B5199B0AC55521524F1864022",
INIT_16 => X"000000000000000000000000000000000026C000002884000130921092804010",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"8020080200000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0051B946088881360A95090CB054420290100000000000000000008020080200",
INIT_1A => X"041041041041041041041041041041041049249249249249200100002D451451",
INIT_1B => X"92C964B2592C964B2592C964B2592C964B2592C86432190C86432190C8641041",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000003800F592C964B2592C964B25",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"7DE1000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"ABDFFFF7803DE10AA80000AAAA843FE0008557DFFF0800020105D557FEAA0055",
INIT_29 => X"D5420000051555FFA2AA8200000557DFFFF7AA80000082ABDF5508557DF45002",
INIT_2A => X"82AA8AAAAAFFC00BA007FC2155F7D155545AA80001EFAAFBEAB45557FFDE10AA",
INIT_2B => X"FFAEBFEAA002A801FFF7FFE8A10A28000000A2D155410F7FFFFEBA08003FE000",
INIT_2C => X"5FFFFEAABA000028A105D2ABFE10A2AABFE1055516ABEF5D517DEAAA2AEBFF45",
INIT_2D => X"55002A820AA08557DFFFF7AA82155AAFBE8B45002A974AAAA803DFFFAA843DF4",
INIT_2E => X"000AAD155555A28428BFF002ABDE00A2AABFE10082ABFFEF0855420000004175",
INIT_2F => X"5010495B7AE921C517DE10000000000000000000000000000000000000000000",
INIT_30 => X"BDF6D005B78F7D142ABDFC7F78E3FE28B684070AABE803AE38145B78FD700000",
INIT_31 => X"BEFB455D71F8E00BED547038145B505FFB6A487000005F7AFD7F7A482038002E",
INIT_32 => X"F1FDE821C003FE001C2EAAAAAB6F5C2082007BC217DEBDB55555AA8E071D7AAF",
INIT_33 => X"D517DEAABEAEBFF7DEBA0BDEAA1C2A801C7E3FFEFA10B68407038B6D550428FF",
INIT_34 => X"B68E38FC7BE8A3DF7DF7F5E8A9200002FA285D20BDE28A2A4B8E10555B68BEF5",
INIT_35 => X"F085F47038140010555142082082005F7DFD7F7A482155BEF1E8B6D002090482",
INIT_36 => X"00000000000000000000B6D15756DA28A28BFF082ABAE10B6AAB8E280820B8FE",
INIT_37 => X"ABA5D7FEAB45080015410007FEAA0055517DE000000000000000000000000000",
INIT_38 => X"AB45F780020BA082EBFFEF007BE8BFF5D2ABDF55F7AABDEAAF784154BAF7802A",
INIT_39 => X"D7545AAAE97555A2FBFDF455D556AA00F7D1554BA5D7BC01FFFF8015410007FE",
INIT_3A => X"4154BAF7D1400BAFFD57FE005D043FE10552EAAAAAFFD140000087FC01EFA2FF",
INIT_3B => X"8428A105D7FEABEF55557DEBAFFAEBFFEFAA803DEBA5D2E82155A2FBFDE00FF8",
INIT_3C => X"7D568BEF080402000F7AAA8B55FFAABDFEFF7D16AA0008003FEBA55003DEBAA2",
INIT_3D => X"FFAAA8AAA080028BFF087BD54AA550402145550000010087FFFF45F78402145F",
INIT_3E => X"0000000000000000000000000000000000000F7D5555FFAAAAA8BFF002AAAA00",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(12),        -- Port A data input
DOA(0)   => data_read_a_lo_256(12),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(12),        -- Port B data input
DOB(0)   => data_read_b_lo_256(12),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_13_14 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10154A0441836CA2840512822007C18000E02700500030B31B300040081A042",
INIT_01 => X"00000804A000C04800020000000002404001000008220008A200100802110204",
INIT_02 => X"02200430000104000A4700804008000004100000000420918204D3033240400D",
INIT_03 => X"AA4003400008592400000590C40009141100000C6180C0000000C00001E14000",
INIT_04 => X"0800000102400120088054019000004160004190BAA0270000C8100000600206",
INIT_05 => X"21000012040610050040000227003AA0082400E94C1200000824424005220020",
INIT_06 => X"81963B180C001010580000080400000058000004109C00138000020024142581",
INIT_07 => X"002C8008000441600106400A9600010494020002B8AAA000EF003408000E2580",
INIT_08 => X"000000E48194408000A00A001210040441C80320040210000002ABF004102244",
INIT_09 => X"2A004009640040100400940412D4C4004000022000104200802D983000480120",
INIT_0A => X"8000202020401480000000000000080C90090881000145B0111A14004015080D",
INIT_0B => X"00000002004040AA08050400404040C11444000805200A402090024000008002",
INIT_0C => X"8410000A00280020020040800020040800020000801020000800010020400000",
INIT_0D => X"84A14250A055100050100490000500D00040080040290000084E4000B800610C",
INIT_0E => X"DCD13042BEDA36820228000000000000C000400081A08BC812A2092B02850942",
INIT_0F => X"89B9A260857DB400431969CA985D480949D32804A40AB137341C10B7D6A02EC0",
INIT_10 => X"E6ACA678001CE7D0296C213A460CA4271CA2168AEC1017606E6838216FAD4055",
INIT_11 => X"84AD4961C281B20213073C5FC0058008632D30D522CE80239DCC01AB013A4D20",
INIT_12 => X"2E6B13804A4B01D83461299900F6BD583A519104A0EEBD1A141010B2A4C8E116",
INIT_13 => X"89E5E40913419151EE0E94641828F72B5151EE0D184B321037AF5158BB02D085",
INIT_14 => X"562EC0B42162D68EE0073AE1C562EC13D521921A4170300B2B458B56B01C2280",
INIT_15 => X"00888A120240034000E6DC8285028014B82372011FC1E4F5E0A00929684EAF84",
INIT_16 => X"50942509425094250942509425094254940A1421420082020120908800480030",
INIT_17 => X"0942509425094250942509425094250942509425094250942509425094250942",
INIT_18 => X"9425094250942509425094250942509425094250942509425094250942509425",
INIT_19 => X"F7EFBBEEFF3F7DF7FF3E9F7DF7E2450228000000000000000000509425094250",
INIT_1A => X"BAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBF7DFDFDDD555555",
INIT_1B => X"EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAEBAE",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000000000F7EBF5FAFD7EBF5FAFD7",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"2ABEF00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0020105D557FEAA00557DE10AAD5554BA087FFFF55557BD54AAF7FBC01FFA280",
INIT_29 => X"7BD75EF087FFFFEF557BEAB45552E80155AA802AB45AA843FE0008557DFFF080",
INIT_2A => X"FAE820AA5D5557555082ABDF5508557DF45002ABDFFFF7803DE10AA80000AA08",
INIT_2B => X"0051555FFA2AA8200000557DFFFF7AA80000AAD1420AA087BD7555FFD168AAAF",
INIT_2C => X"5557FFDE10AAAEA8BFFA2FBD7545FFD157555085140010F7AEAABFFAAD542000",
INIT_2D => X"BA557BE8A10A284154BAFFAAAAB45007FC2155F7D155545AA80001EFAAFBEAB4",
INIT_2E => X"000A2D155410F7FFFFEBA08003FE00082AA8AAAAAFFC00BA00002AAAAF7D5574",
INIT_2F => X"0492E3F1C71C7BE8A2ABD7000000000000000000000000000000000000000000",
INIT_30 => X"3AE38145B78FD7000005010495B7AE921C517DE10A2DB50482147FFAF554971D",
INIT_31 => X"E3FE28B684070AA1C71D25D7007FFAFD7497BE8B5555208217DBE8A2AB45BE80",
INIT_32 => X"7FD257DFFD568A82FFA4870BA555F5056D002EBDF6D005B78F7D142ABDFC7F78",
INIT_33 => X"FAAAFBFFBED547038145B505FFB6A487000005F7AFD7F7A482038AADF4709214",
INIT_34 => X"AA8E071D7AAFBEFB455D71F8E00A2A0ADBC7A2FFD257DE3DF52555085142000F",
INIT_35 => X"21C002AA92FFDF574824171EAA10B680124BAFFAAAFB45007BC217DEBDB55555",
INIT_36 => X"00000000000000000000B6D550428FFF1FDE821C003FE001C2EAAAAAB6F5C208",
INIT_37 => X"0105D7BE8B55085142010AAD157545F7AEA8B550000000000000000000000000",
INIT_38 => X"01EFF7AAA8B55F7802AABA5D7FEAB45080015410007FEAA0055517DE00A2FFC0",
INIT_39 => X"E8BFF5D2ABDF55F7AABDEAAF784154BA5D5140145007BE8B55087BEAB555D040",
INIT_3A => X"0020BAA2FFD54105D7FC21EFFFD16AA10FF80174AA557FC21EF082EBFFEF007B",
INIT_3B => X"FBC0155085540000FFAEBFFEFF7D1554BA5D7BC01FFFF8015410007FEAB45F78",
INIT_3C => X"87FC01EFA2FFD7545AAAE97555A2FBFDF455D556AA00A2803FF45AAFFC21EFAA",
INIT_3D => X"552EAAAAAFFD1400005D042AA00F7FBD5410085568A10FF80020AAFFAABFF550",
INIT_3E => X"0000000000000000000000000000000000000F7D1400BAFFD57FE005D043FE10",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(13),        -- Port A data input
DOA(0)   => data_read_a_lo_256(13),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(13),        -- Port B data input
DOB(0)   => data_read_b_lo_256(13),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_14_14 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10020A000180000284008280000281800000030000000033022000000580002",
INIT_01 => X"000008020000204D006800000030824840000000084000084200090008510200",
INIT_02 => X"0220043170010A600A4D008040080000041000000028009002000F333240800C",
INIT_03 => X"111813400008002400000000C400090011000000610200001104D83000F14000",
INIT_04 => X"0801800100A000000000540084000040000040000800200000C8100000000748",
INIT_05 => X"0100000000001000000000002000080008000000001000000024024001200020",
INIT_06 => X"819EB84028001010000000080400000000000004108000100000020020040081",
INIT_07 => X"92040608000440100102400A94810206844200021DA2A0002000340800062C80",
INIT_08 => X"000000000084400008800A001214040441481500040000000000A7F408002244",
INIT_09 => X"0A0040090002008420401004104444004000020400214A208001000002400120",
INIT_0A => X"0400002020000000000000000000080C8008088100004590111B480040120000",
INIT_0B => X"1000000200404800000504016000002114000008020000020080024000000000",
INIT_0C => X"0410000010000000000040001000000000000040000000000001000000000000",
INIT_0D => X"04810244825010004010000000000000000000000000000000080000B8002104",
INIT_0E => X"0002C38280001202020800000000001000004000000000401022000002040902",
INIT_0F => X"20000587050001404E8084341CBA3404800828805200008000E0E0A000080002",
INIT_10 => X"4D18178E012010C00224004091C3514072C000444A0400080001C1C140001000",
INIT_11 => X"51709A07424142084458476001003809D0104B01C5710044020C4006010500C5",
INIT_12 => X"C26EE3803180C18006519462A00005001460E4730000050A1011004001060049",
INIT_13 => X"01F9E00660318000000538318740000140000001B4600CE80001400000002B62",
INIT_14 => X"0000000AD89857B0E0684411800000003799EB764D000330C300000000E3554B",
INIT_15 => X"0000021002002C000024008284001A0902000422E3F5960080480A0216A07240",
INIT_16 => X"4090240902409024090240902409024090081021020080015134920800480010",
INIT_17 => X"0902409024090240902409024090240902409024090240902409024090240902",
INIT_18 => X"9024090240902409024090240902409024090240902409024090240902409024",
INIT_19 => X"F5579B4E5C8FF0F7BE9D5F7DF650400200000000000000000000409024090240",
INIT_1A => X"9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7BF7DDDDDFCF3CF3D",
INIT_1B => X"F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE79E7",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000003FFF03F9FCFE7F3F9FCFE7F3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"420BA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"BD54AAF7FBC01FFA2802ABEFA2FBE8B55A2AE80000F7D5555555D2AAAABAAAD1",
INIT_29 => X"AA801FFA28402000AAAE955455500155EF0804155EFAAD5554BA087FFFF55557",
INIT_2A => X"7AEA8B45080417400AA843FE0008557DFFF0800020105D557FEAA00557DE10A2",
INIT_2B => X"087FFFFEF557BEAB45552E80155AA802AB4500516AA00A2AE800BAFFFFC20BAF",
INIT_2C => X"0AA80000AA005568ABAA28402010A2843FEBAFFFBD7410A2D168BFF087BD75EF",
INIT_2D => X"005D7FFDF4555517DFEF00043FEAA082ABDF5508557DF45002ABDFFFF7803DE1",
INIT_2E => X"000AAD1420AA087BD7555FFD168AAAFFAE820AA5D5557555002E80155A280000",
INIT_2F => X"0555412AA8ABAAADB40092000000000000000000000000000000000000000000",
INIT_30 => X"50482147FFAF554971D0492E3F1C71C7BE8A2ABD7A2FFEDB55B6A080038E3DB5",
INIT_31 => X"B7AE921C517DE10A2AE851FFB68402038AAAA955554900105FF0800175D7A2DB",
INIT_32 => X"A0800BAE3F1C0092EBAAADB6D080A12410BE803AE38145B78FD7000005010495",
INIT_33 => X"2D568BC71C71D25D7007FFAFD7497BE8B5555208217DBE8A2AB451C556FA00A2",
INIT_34 => X"142ABDFC7F78E3FE28B684070AA00516DABAA28402038B6803DE82F7F5D5410A",
INIT_35 => X"D002A80155B680000105D7FF8F455D5F78FD7000E3FEAA002EBDF6D005B78F7D",
INIT_36 => X"00000000000000000000AADF47092147FD257DFFD568A82FFA4870BA555F5056",
INIT_37 => X"F55FF84000AAAAFBC0145002AA8AAAAAFFC20000000000000000000000000000",
INIT_38 => X"01EF080417555A2FFC00105D7BE8B55085142010AAD157545F7AEA8B55A2FBFF",
INIT_39 => X"EAB45080015410007FEAA0055517DE00A2AA955FFFF80020BAAAAA9754508000",
INIT_3A => X"AA8B555D557FE00A280020BAAAD140000A2AEBFFEF082A82010F7802AABA5D7F",
INIT_3B => X"803DE00FFD557400AAD56AB455D5140145007BE8B55087BEAB555D04001EFF7A",
INIT_3C => X"82EBFFEF007BE8BFF5D2ABDF55F7AABDEAAF784154BA08557FEAAA284000AAFF",
INIT_3D => X"FF80174AA557FC21EF082A80145F780020105D7BEAB45557BE8B45082EBFEBA0",
INIT_3E => X"0000000000000000000000000000000000000A2FFD54105D7FC21EFFFD16AA10",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(14),        -- Port A data input
DOA(0)   => data_read_a_lo_256(14),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(14),        -- Port B data input
DOB(0)   => data_read_b_lo_256(14),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_15_14 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000A000000000284000280000001800020030000000033022000000180002",
INIT_01 => X"8000080000000048000000000000026040000000080000080200000000110200",
INIT_02 => X"0020042004010E60004C0080000800000410000000020090020000300245E005",
INIT_03 => X"0000010000080400000000408400480111000000610008000000C00000E54400",
INIT_04 => X"980000010000000088C2550080000040000040000008A00028C8100000120000",
INIT_05 => X"020004012E025000000001322000000A28008000011000000220004D41000000",
INIT_06 => X"819588000800101000011008040000100001060418800510000A620000000092",
INIT_07 => X"0000000800044004010C20008440810284020002102220002000340800062480",
INIT_08 => X"0000000001140800002C0A001214050540C800400406180000002DF004000244",
INIT_09 => X"1E00400900000000000016041044400440000000000042008001000000000022",
INIT_0A => X"0000000000000220000000000000080C00000081000045901118000040000000",
INIT_0B => X"0000000200404000010500004000000114000009000000000000004200000000",
INIT_0C => X"0000000000000000000040001000040001000000000000000001000020000800",
INIT_0D => X"000000000000001001208000180800000000030200000180800C400030002000",
INIT_0E => X"0000000000002600020800000000001080004000000000000002000000000000",
INIT_0F => X"A400000000000000000008000000000000000000000014800000000000000052",
INIT_10 => X"0000000000000000000000010240000000000000000000290000000000000000",
INIT_11 => X"2001C05838120800000000000000000000010000000000000000000000001804",
INIT_12 => X"081004000000000000A010000000000000902000000000180010002020000000",
INIT_13 => X"6600000000000000000024080000000000000000280400000000000000000000",
INIT_14 => X"0000000000200801000000000000000000501001920000000000000000000A40",
INIT_15 => X"0000020000000000000000003000000000000000000A101C3614000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000080000120980000000010",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000400200000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"28BEF00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"5555555D2AAAABAAAD1420BAFF8000010082A954BA00003DFEF085155400F784",
INIT_29 => X"AE95555A2FBE8BEFA2843DE00AA8015400FF84001EFA2FBE8B55A2AE80000F7D",
INIT_2A => X"2FBEAB45F7D56AABAAAD5554BA087FFFF55557BD54AAF7FBC01FFA2802ABEFF7",
INIT_2B => X"A28402000AAAE955455500155EF0804155EFFFFBE8BFF0800174AA557BFDE10A",
INIT_2C => X"A00557DE10F7D1574AAA2D16AB55FFD568BEF087FE8A1055003FE00A2AA801FF",
INIT_2D => X"00AA802AA00AAAE800BA5D0015545AA843FE0008557DFFF0800020105D557FEA",
INIT_2E => X"00000516AA00A2AE800BAFFFFC20BAF7AEA8B45080417400FFFFC21450800154",
INIT_2F => X"8FD7005150438F78A2DBFF000000000000000000000000000000000000000000",
INIT_30 => X"EDB55B6A080038E3DB50555412AA8ABAAADB40092E38E070280024904AA1C043",
INIT_31 => X"1C71C7BE8A2ABD7E3AA9257DA2FFE8BC7BE8E38E10A28017400E38A051FFA2FF",
INIT_32 => X"00124AA557FFDE10A2FBEDB6DF7D16AABAA2DB50482147FFAF554971D0492E3F",
INIT_33 => X"10038E38A2AE851FFB68402038AAAA955554900105FF0800175D7E3FFEFBD700",
INIT_34 => X"000005010495B7AE921C517DE10FFDF50482A2DB6AB45FFD56DBD7087BEAA384",
INIT_35 => X"0FFF1C017D140410400BE8E28A10AAA085082550A1057DBE803AE38145B78FD7",
INIT_36 => X"000000000000000000001C556FA00A2A0800BAE3F1C0092EBAAADB6D080A1241",
INIT_37 => X"4AA0800020BA550028B550855400AAF7AEBDFEF0000000000000000000000000",
INIT_38 => X"7400AAAE975EFA2FBFFF55FF84000AAAAFBC0145002AA8AAAAAFFC2000AAAA97",
INIT_39 => X"E8B55085142010AAD157545F7AEA8B55AAAE821EFAAFBEAB55F7AAA8A00AA841",
INIT_3A => X"417555AAFFFDF450804020AA557BFFE10A2FFFFFEFF7D568ABAA2FFC00105D7B",
INIT_3B => X"D17DF45007FE8AAA08002AAAAA2AA955FFFF80020BAAAAA975450800001EF080",
INIT_3C => X"7802AABA5D7FEAB45080015410007FEAA0055517DE00FFFBC2000AAFBE8B55F7",
INIT_3D => X"A2AEBFFEF082A82010FFD5421EF5D0000010F7AAA8A10AA8017400552A801EFF",
INIT_3E => X"00000000000000000000000000000000000005D557FE00A280020BAAAD140000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(15),        -- Port A data input
DOA(0)   => data_read_a_lo_256(15),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(15),        -- Port B data input
DOB(0)   => data_read_b_lo_256(15),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_16_14 : RAMB16_S1_S1
generic map (
INIT_00 => X"DA22C618B1000482B688B186588884862A400438255FC38381441205BA803003",
INIT_01 => X"7045A80028404C211203A952A90341080B173340412000E1005D628000820484",
INIT_02 => X"428406A4000850848330118D0AAC55001349B108818005460229044001C01784",
INIT_03 => X"092C4020000500020000500986812C405000001A48202050000A214AC0650115",
INIT_04 => X"4804A55440256F504025E003A054F46415A4E62B6FE3307943965A00001A1152",
INIT_05 => X"0000001C40A5B950ADB8EA097057ECE14C86D2B7F85AAD17F4B100000B88148C",
INIT_06 => X"415401DCDCF2C0A8030140BCB0820A200342A1C641C1E8782F508F2B00003584",
INIT_07 => X"002701881A3202080AE00480A2002840BE1480FA004342AA6F12000054004867",
INIT_08 => X"08C54828091002000002B32A8C19064E486A8001510000014140C1E2A14891E0",
INIT_09 => X"015452B103020814004088B64102680B6596594800400413CAC0208944800000",
INIT_0A => X"96AA000484094C000000000000012C9000A0000D0A80000BF8028E87C1B99270",
INIT_0B => X"014808A02004200E540480212000A448C0082024AE50064B44000000000002A2",
INIT_0C => X"0004000D5846256AAEA811150445411150445411150445411150422A088A8200",
INIT_0D => X"00000004010042A204A0C5817D00005034052E40000817D00440004004AD3240",
INIT_0E => X"632B2673FA4587978A2004102800809225545155121740000004900090000000",
INIT_0F => X"00C6564CE7F4EA4B940076D296D003030800462CBD320018CAAAACFE9164C800",
INIT_10 => X"28834ADB1440A114793A4A30A40839AA14910D08DCB2640031955559FD3AC990",
INIT_11 => X"594AB0B1A025371CA0E034E8443C097A800EB090D4AAC91208ED2FA0CE5E09B1",
INIT_12 => X"7B50446083001B94BB38C540EBE61284BB304880E3E4579EDC00992980D58033",
INIT_13 => X"5511121840E7A2CD952ECC12ABC3E6ACB3DFB12ECE315000F61FF1727A85FDBC",
INIT_14 => X"75DEB07F6F2E7084517F126F8395CB2BEFBAB8BA8AF698228CC5E2F08ECA5159",
INIT_15 => X"5580A840A8009F8B108C80A1021B080AFC0DF6422C6077F4A77F20D0C0E21084",
INIT_16 => X"0000000000000000000000000000000000044000102A0001148442A110810359",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"558D11544C690DA64C1C4F68A360400000000000000000000000000000000000",
INIT_1A => X"14D14D14D14D14D14D14D14D14D14D14D14514514514514529E5F87869E79E78",
INIT_1B => X"D1E8F47A3D1E8F47A7D3E9F4FA7D3E9F4FA7D3E9F47A7D1E9F47A7D1E9F4D14D",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000007D3E9F4FA7D3E8F47A3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"C00AA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"03DFEF085155400F78428BEF087FFFFEFF7D168B55AAD17FFFF552EBFE00007F",
INIT_29 => X"2E975EFF7D568BFFFF80175EF0004000BA552A821FFFF8000010082A954BA000",
INIT_2A => X"55540000082EAABFFA2FBE8B55A2AE80000F7D5555555D2AAAABAAAD1420BA5D",
INIT_2B => X"A2FBE8BEFA2843DE00AA8015400FF84001EF0000020AA5D00154005D043FF455",
INIT_2C => X"FA2802ABEF557BEABEF5D0415410087FD74BAAAAEBFFEF557FC00AAF7AE95555",
INIT_2D => X"FFFFAABFEAAFF84001FF002A821FFAAD5554BA087FFFF55557BD54AAF7FBC01F",
INIT_2E => X"000FFFBE8BFF0800174AA557BFDE10A2FBEAB45F7D56AABA082A97545F7D16AB",
INIT_2F => X"FFEF552AB8E38087FC2092000000000000000000000000000000000000000000",
INIT_30 => X"070280024904AA1C0438FD7005150438F78A2DBFF0871F8FC7E3D56AB6DBEDB7",
INIT_31 => X"AA8ABAAADB400924920925EFF7D16ABFFE38E175EF1400000BA412E871FFE38E",
INIT_32 => X"0A1240055003FF6D5551420101C2EAFBD7A2FFEDB55B6A080038E3DB50555412",
INIT_33 => X"57FC00BAE3AA9257DA2FFE8BC7BE8E38E10A28017400E38A051FF0804050BA41",
INIT_34 => X"4971D0492E3F1C71C7BE8A2ABD74975EDBC7550E12410087FD74AAB6AABFFC75",
INIT_35 => X"A08249756DF7D168BC7F7AABAEAAF780051C70824851D7A2DB50482147FFAF55",
INIT_36 => X"00000000000000000000E3FFEFBD70000124AA557FFDE10A2FBEDB6DF7D16AAB",
INIT_37 => X"B55A2D16ABEFFFFBFDFFF552AAAAAA007BC00000000000000000000000000000",
INIT_38 => X"20AA002A955EFAAAA974AA0800020BA550028B550855400AAF7AEBDFEF08516A",
INIT_39 => X"000AAAAFBC0145002AA8AAAAAFFC20000000021EFF7D568BFFA2AA955FF5D040",
INIT_3A => X"E975EF0800174BA002E820105D003DFEF5D51420005D2ABFF45A2FBFFF55FF84",
INIT_3B => X"7BD74AAF7AEBDF455D7BC20BAAAAE821EFAAFBEAB55F7AAA8A00AA8417400AAA",
INIT_3C => X"2FFC00105D7BE8B55085142010AAD157545F7AEA8B5500557DF45552A8200000",
INIT_3D => X"A2FFFFFEFF7D568ABA0804155FFF7D568B55FFAAAAABAFF8415545000015555A",
INIT_3E => X"0000000000000000000000000000000000000AAFFFDF450804020AA557BFFE10",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(16),        -- Port A data input
DOA(0)   => data_read_a_lo_256(16),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(16),        -- Port B data input
DOB(0)   => data_read_b_lo_256(16),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_17_14 : RAMB16_S1_S1
generic map (
INIT_00 => X"5284CE4FB7BD2C8994A13392DBD02E14006B82AC7E800D44D3DD2FD5F9B961C0",
INIT_01 => X"2EACD01F7E03FC6793F2199B39FC233C11D93AE6F3BB92B32091DBC339B24542",
INIT_02 => X"E63CCCC00A82C08092A2AFAE667033DB50853379C10BFDC5C6F4044443C817C6",
INIT_03 => X"7FF183635AEF9E3635AEF9E18E237040404446965C0607EE6DB7854AC4DE060C",
INIT_04 => X"D78AC33FB604488B000892EF17BE6D84196482236FE100294152E294350FB697",
INIT_05 => X"081B5F9B409420D0CDB47A05403F6CE0C08A4AB7F840EDB6F48100DFC8081081",
INIT_06 => X"768465354781CBC30316367077B4BDB50646E8D87100A8201ED01C19C020F71A",
INIT_07 => X"4002A110C922480A82D0841147162C48EBB9537A0022DC67987042EE976ABEA7",
INIT_08 => X"DB931BFEF91C00002CC0E019C0C82A4E4820C15A2330E004401891181168C4D1",
INIT_09 => X"09F3A1BC11EFBC66DB65307071477FF1030C397C060B4254064302042F803A69",
INIT_0A => X"3F330802162F3B7EE3F3EC7C7DEF207000F00059D2ED56D7EED2ED3C9A867DC0",
INIT_0B => X"185C44B91BC1740B7605040BE0018CFC7429F326B9E822FFC00074D5A0AB033A",
INIT_0C => X"00367A28FC1B7F7FEFFCFBFF3EFFCFBFF3EFFCFBFF3EFFCFBFF3EFFE7DFF9E00",
INIT_0D => X"0000000008004BA78428C7AD7FC94B533F5B4FFBD2FAD7FCCA786D43FE67C218",
INIT_0E => X"BA494CEBFD4F2667ABB6F68B29760593F33FA0CF170F40006001B1A05C000000",
INIT_0F => X"7F749299D7FAEB237DFE5865B6D2BF23265CBACE542A6FEE92333AFF33E0A9BF",
INIT_10 => X"F6C24B6D18C3C9F8E2881F3F787D776B5DB94A09955054DFDD246675FE7AC153",
INIT_11 => X"BFB349E08FF9A27EDE9FA8AEFD9E7467BFCB195CFEB56A1A70D34D1706FFFA3E",
INIT_12 => X"6FE219CA80725B875EED723FF7FCB2875EDAAFEAF7FD929BFD55BBC71D79F639",
INIT_13 => X"546670D018E7A6E581D7B6AB75FDFCECA6E581D7BB5DDFC6FF0EB7D7E859FDB5",
INIT_14 => X"B978177F6D6AF5ECDB5FB76A5F5FA165B456E0FB308710C49FCFB741598B9C7E",
INIT_15 => X"CFDAAB00AC00A8BBFC8B501CF7A0FED9A540EA1952586CEB54D143ACFF9A3BA9",
INIT_16 => X"000000000000000000000000000000000026E100002F382DBD9ECFE117805F20",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"4372003009EDCC4052E917114F981800C0000000000000000000000000000000",
INIT_1A => X"BA69A69AEBA69AEBA69A69AEBA69AEBA69A69A69A69A69A68698686981D75D74",
INIT_1B => X"6A351A8D46A351A8D068341A0D068341A0D068341A0D46A341A0D46A341A69AE",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000000000046A351A8D46A351A8D4",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"7FEAA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"17FFFF552EBFE00007FC00AA087FFFFFFFFFFFFFEFF7FBEAB450804001EFAAD5",
INIT_29 => X"D168A000004020AA5D7BE8B450051401EF087FD74AA087FFFFEFF7D168B55AAD",
INIT_2A => X"D7FEAB55FF80175EFFF8000010082A954BA00003DFEF085155400F78428BEFAA",
INIT_2B => X"F7D568BFFFF80175EF0004000BA552A821FF5D00020BA552A82000552A821555",
INIT_2C => X"AAAD1420BAFFFFFDF45AAD17FFFFAAFBC01EF5D0015555557BFDEBA5D2E975EF",
INIT_2D => X"BA007FEABEF005555555A2D1554BAA2FBE8B55A2AE80000F7D5555555D2AAAAB",
INIT_2E => X"0000000020AA5D00154005D043FF45555540000082EAABFF00516AA10552E820",
INIT_2F => X"8B550000071EFB6DF7AE92000000000000000000000000000000000000000000",
INIT_30 => X"F8FC7E3D56AB6DBEDB7FFEF552AB8E38087FC2092147FFFFFFFFFBFDFC7EBF5E",
INIT_31 => X"150438F78A2DBFFBED16AA381C0A07082497FEFB6D1451471EF007BD04920871",
INIT_32 => X"2A850105D2A80155417BEFB6DEB8E175FFE38E070280024904AA1C0438FD7005",
INIT_33 => X"D7BFAEBA4920925EFF7D16ABFFE38E175EF1400000BA412E871FF550A0009249",
INIT_34 => X"E3DB50555412AA8ABAAADB40092FFF5FFF6DAADF7FFD7B6F1C71EF55001756D5",
INIT_35 => X"7145B6AA28492487082007FEDBD700515556DA2DF50492A2FFEDB55B6A080038",
INIT_36 => X"000000000000000000000804050BA410A1240055003FF6D5551420101C2EAFBD",
INIT_37 => X"FEFF7FBFFF55A2D16AB550000175EFFFFBEAA000000000000000000000000000",
INIT_38 => X"55EF087FC200008516AB55A2D16ABEFFFFBFDFFF552AAAAAA007BC0000557FFD",
INIT_39 => X"020BA550028B550855400AAF7AEBDFEFF7D568AAA5D2A97410007BFFFFF55515",
INIT_3A => X"A955EF5D2E80010002A954005D2A82155087FFFFEFAAAA975EFAAAA974AA0800",
INIT_3B => X"D1575FF5504175EF5D7FEAAAA0000021EFF7D568BFFA2AA955FF5D04020AA002",
INIT_3C => X"2FBFFF55FF84000AAAAFBC0145002AA8AAAAAFFC2000FFD57DFFFAAFFFDF55FF",
INIT_3D => X"5D51420005D2ABFF45557FE8AAA000415410007BFFF450051555EFA2FBC0000A",
INIT_3E => X"00000000000000000000000000000000000000800174BA002E820105D003DFEF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(17),        -- Port A data input
DOA(0)   => data_read_a_lo_256(17),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(17),        -- Port B data input
DOB(0)   => data_read_b_lo_256(17),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_18_14 : RAMB16_S1_S1
generic map (
INIT_00 => X"69844019080000A21A611406840014122A641074155FC28A2024001001801003",
INIT_01 => X"7443D920034004180005E9E3C90360C0041C0181002001602025800008440084",
INIT_02 => X"E2DCCCE61D5C008103F2000781FC0FEDEAC2161B0B8FB0008620044443006010",
INIT_03 => X"884E300802006900802006995C896D605200000856E24A040000640052141103",
INIT_04 => X"480520FC026125AC0025C9122644E3E40EC8E2001001302281841A009038A86A",
INIT_05 => X"432000040089983070019400F01010004C8DB841405A80A100B586200FAC24AE",
INIT_06 => X"09044359DC7040000000002C109B0E0A00A1104641C0803804000707284600E1",
INIT_07 => X"400D10100400481D5EB08501620000007500CE801241021FE78E404860140060",
INIT_08 => X"00880C0106A0528020019307CC082A0A4A6A01ED725021400040D028000A9729",
INIT_09 => X"00117063038000282081402E4106400B6186128040600C10C1C0200950508110",
INIT_0A => X"C0C30C2E21580C874004008080003C32A10A19090C02010E1022944061688000",
INIT_0B => X"0180A8062026000DC425C0301311324AA2373088479105D044A1022000001835",
INIT_0C => X"0D89844703649000000200000000000000000000000000000000000000000010",
INIT_0D => X"0D8306C182701404C1973010802020404084001E00010802046092B5001FB365",
INIT_0E => X"528EB314068AB8B803DB00002900800400FC503F08180050942E4200020C1B06",
INIT_0F => X"40A51D66280D6032C5F96D3C51555D5D7D5AA87285820814A3CCC501C2A60820",
INIT_10 => X"8B35A3FEBF1FEDFD9C2B30E0468AAAD5D48F37E8FC1304102947998A03984C10",
INIT_11 => X"440FE1DD772D37A0A321BC6968F32658BF2D4F2A80BF8FE3F9FE3AC362080529",
INIT_12 => X"5487910D7E5A6D961A28456A1832E5161A100DD5182BC54020EA67A189C6ED36",
INIT_13 => X"AA444CAF91EDD1B725868403BE06323551B725868A100ABD119753B70964122B",
INIT_14 => X"EDC259048ACD868EE3803D65CEDC258A8F80D55E007C3F8EBB56F4C5362C978F",
INIT_15 => X"3F240014BE84370001B6922070440556B15F7FABBC0031BCF2257C41634B14D4",
INIT_16 => X"C1B06C1B06C1B06C1B06C1B06C1B06C1B0491069068000004060300A005A0118",
INIT_17 => X"1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06",
INIT_18 => X"B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C",
INIT_19 => X"B28BBECEB80EE173C2300F7DF16000000000000000000000000041B06C1B06C1",
INIT_1A => X"8A28A28AAAAAAA28A28A28AAAAAAA28A28A28A28A28A28A2910591505C104104",
INIT_1B => X"28944A25128944A25128944A25128944A25128944A2552A954AA5128944AAAA2",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000128944A25128944A251",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"9540000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"BEAB450804001EFAAD57FEAA087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974BA082E",
INIT_29 => X"7FFFFFFFFFBFDF45AAD568B55080028B55002E82000087FFFFFFFFFFFFFEFF7F",
INIT_2A => X"0043DE10AA843DE00087FFFFEFF7D168B55AAD17FFFF552EBFE00007FC00AA08",
INIT_2B => X"0004020AA5D7BE8B450051401EF087FD74AAAAFFFDF45A2D16AB55F7FFFFFFF0",
INIT_2C => X"0F78428BEFAA80000000804154BA55042ABEF5D7FD75FFAAD540145AAD168A00",
INIT_2D => X"00082E95555085168A10557FD7545FF8000010082A954BA00003DFEF08515540",
INIT_2E => X"0005D00020BA552A82000552A821555D7FEAB55FF80175EF5D00020105D2A974",
INIT_2F => X"DFFF5D2A954AA082A92428000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFBFDFC7EBF5E8B550000071EFB6DF7AE921C7FFFFFFFFFFFFFFFF7FBF",
INIT_31 => X"AB8E38087FC2092087FFDFC7E3F1FAF55A2DF6DB7D1C002AB7D002A82028147F",
INIT_32 => X"DF6DB7DE3F5FAFC708003DE28B68E38E280871F8FC7E3D56AB6DBEDB7FFEF552",
INIT_33 => X"ADF4516DBED16AA381C0A07082497FEFB6D1451471EF007BD0492B6F1F8F55AA",
INIT_34 => X"1C0438FD7005150438F78A2DBFFA28407038140410492550A2ABC7497BD25FFA",
INIT_35 => X"F5D0E05000492097428002E9557D1C516FA28417BD5545E38E070280024904AA",
INIT_36 => X"00000000000000000000550A00092492A850105D2A80155417BEFB6DEB8E175F",
INIT_37 => X"FFFFFFFFDFEFF7FBFFFEF552E974AA082A820AA0000000000000000000000000",
INIT_38 => X"ABEF002A800AA557FFDFEFF7FBFFF55A2D16AB550000175EFFFFBEAA00557FFF",
INIT_39 => X"6ABEFFFFBFDFFF552AAAAAA007BC0000087BFDF45AAD568B55AAFBFDFEF55042",
INIT_3A => X"FC2000FFD56AB45A2FFFDFFFAAD16AB4500043DEAAFFAEAAAAA08516AB55A2D1",
INIT_3B => X"2AA8B45087FC01EFA2FFD55EFF7D568AAA5D2A97410007BFFFFF5551555EF087",
INIT_3C => X"AAA974AA0800020BA550028B550855400AAF7AEBDFEFA280154BA55040000055",
INIT_3D => X"087FFFFEFAAAA975EF5D2E974000804154BA082A975EF5D517DEAA007BD5545A",
INIT_3E => X"00000000000000000000000000000000000005D2E80010002A954005D2A82155",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(18),        -- Port A data input
DOA(0)   => data_read_a_lo_256(18),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(18),        -- Port B data input
DOB(0)   => data_read_b_lo_256(18),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_19_14 : RAMB16_S1_S1
generic map (
INIT_00 => X"042200000000000041088001001AA00000000000000000000000500802000003",
INIT_01 => X"040048000024000000000404000000000A22000800000800004A200000000001",
INIT_02 => X"200C8840085EB00480060000001C008002489E0F000405EA0004040404000000",
INIT_03 => X"24004000000000000000000900002C4050000000000069500208400002E14100",
INIT_04 => X"4800200C0000000044002000C80020E40000E200000130200188000000800100",
INIT_05 => X"000000000080181000000000701000004C8000000058800000B1000009880480",
INIT_06 => X"80500081081040000000002C100040400000004641C080380400070100000000",
INIT_07 => X"4020109801A4CE005C00048380142810010564C4100114012002402028044808",
INIT_08 => X"0070700000000000000083004C3902420062000020E0000100004082A140102B",
INIT_09 => X"001150200000000000000026400000016186100000000010C04002C000000000",
INIT_0A => X"007C00008082C0002000000000002C3000000004050001030102040000000000",
INIT_0B => X"0000000000000000000000000000010000800011000000000000000000000BC0",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"000000000000000000000000000000042000760000000000000000010004B200",
INIT_0E => X"0D74002280300F0002FB069040000060000C5003000800000000000000000000",
INIT_0F => X"C01AE8004500744C780687DBA828008080A5FC0D385598035D0008A00C015660",
INIT_10 => X"39D8140040201BF861F0E7D693E6170022408116DFE0AB3006BA0011401D02AC",
INIT_11 => X"5412E4997F5249FD005043B8680CC98F00D0F2DD0140100406FE053A98F6ECC7",
INIT_12 => X"7418663001858040E153888000010840E165D0000000285C246A181C03FE4662",
INIT_13 => X"8199830066F0020858385974000001260208583854E2200000660208D6B1423F",
INIT_14 => X"8235AC508FCE8811042040F008235AE04420C040CF00C031C80009B8F224978B",
INIT_15 => X"030004E00000C220010808C10D9A92A74CD7CF4A09051110AD5A3C9200B7F280",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000118",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"07208BBA3F0C7010C660C7441920000000000000000000000000000000000000",
INIT_1A => X"861869A61861861861869A61861861861861861861861861A8208C4C1534D34C",
INIT_1B => X"984C26130984C26130984C26130984C26130984D26930984C26130984C261861",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000984C26130984C26130",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"174BA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFDFEF5D2A974BA082E95400F7FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0004",
INIT_29 => X"FFFFFFFFFFFFFFFFF7FBFDFFF552E974BAA2FFFFE10087FFFFFFFFFFFFFFFFFF",
INIT_2A => X"004001EFAAAEA8ABA087FFFFFFFFFFFFFEFF7FBEAB450804001EFAAD57FEAAF7",
INIT_2B => X"FFFBFDF45AAD568B55080028B55002E82000F7FFFFFFFFFFFFDFEFA2D568B550",
INIT_2C => X"0007FC00AAF7FFFFFFFF7FBE8B55AAD16ABEF5D2ABFF55080402010087FFFFFF",
INIT_2D => X"55A2FFFDFEF5D2EBFE00AAFFFFEBA087FFFFEFF7D168B55AAD17FFFF552EBFE0",
INIT_2E => X"000AAFFFDF45A2D16AB55F7FFFFFFF00043DE10AA843DE00557FFDFEFA2D16AB",
INIT_2F => X"FFEF552A974AA0000104AA000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFF7FBFDFFF5D2A954AA082A92428E3FFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"0071EFB6DF7AE92EBFFFFFFFFFFFFDFEFF7F5FAFC7492A974AAB6F5F8E101C7F",
INIT_32 => X"F1F8FD7AAD16AB450000001FFBEA4A8AAA147FFFFFFFFFBFDFC7EBF5E8B55000",
INIT_33 => X"00000010087FFDFC7E3F1FAF55A2DF6DB7D1C002AB7D002A82028FFFFFFFEFF7",
INIT_34 => X"BEDB7FFEF552AB8E38087FC2092F7FBF8FC7E3F5EAB45B6DF6FBEF5D2AB8F7D0",
INIT_35 => X"84971F8FC7AAD56DB6DBEF5F8FD7412ABFE28B6F5F8E820871F8FC7E3D56AB6D",
INIT_36 => X"00000000000000000000B6F1F8F55AADF6DB7DE3F5FAFC708003DE28B68E38E2",
INIT_37 => X"FFFFFFFFFFFFFFFFFDFEF552E954AA0004000AA0000000000000000000000000",
INIT_38 => X"54AAF7D568A00557FFFFFFFFFFFDFEFF7FBFFFEF552E974AA082A820AAA2FFFF",
INIT_39 => X"FFF55A2D16AB550000175EFFFFBEAA00A2FFFFFFFF7FBFDFFFFFD568B55002A9",
INIT_3A => X"A800AAF7FBFDFEFF7D56AB45AAD56AB450004001EFFF842AAAA557FFDFEFF7FB",
INIT_3B => X"FFFFFFF552AA8BEF080402000087BFDF45AAD568B55AAFBFDFEF55042ABEF002",
INIT_3C => X"8516AB55A2D16ABEFFFFBFDFFF552AAAAAA007BC0000FFFBE8B55AAD168B55F7",
INIT_3D => X"00043DEAAFFAEAAAAA08556AB55A2D57FFFFF7D568B45002ABDEAAFFD16AA000",
INIT_3E => X"0000000000000000000000000000000000000FFD56AB45A2FFFDFFFAAD16AB45",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(19),        -- Port A data input
DOA(0)   => data_read_a_lo_256(19),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(19),        -- Port B data input
DOB(0)   => data_read_b_lo_256(19),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_20_14 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000003",
INIT_01 => X"F55FF80000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"E05022020800008400F655001FFCFF80018FA804400000000000004400000001",
INIT_03 => X"00000000000000000000000900002CC07000000000000000000000000000013F",
INIT_04 => X"68002FFE40900010000180000001FFEC0012EE0C001370F40780000000000000",
INIT_05 => X"0840000880FCBBF0100E204DF0F88311DD8005080679800000F3000029980580",
INIT_06 => X"001000030817C8E8840155FDF9001001050023F6C3C3D0F87FA19F7F011000E4",
INIT_07 => X"000000090492260800008000EE00000000000000002101FF2002C00000004018",
INIT_08 => X"2A040001071004000013FF7FCA302C0C0008214800002101554031F800000000",
INIT_09 => X"801F57F200000090000489FEC0000001EFBEF0040008023FDFC0000000004006",
INIT_0A => X"0000000008000000000000000000ADF000000200000008000008028300110230",
INIT_0B => X"0000000000000800080000000000000000000000000000000800800A40000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"000000040900005C848538000020000000800000080000020000800101FFB600",
INIT_0E => X"00800000003A010003000000000000600FFC53FF001800000002004080000000",
INIT_0F => X"0001000000007408040000004000000004E9000008020000200000000E800800",
INIT_10 => X"00200000000313100010002000008000000000129600040000400000001D0010",
INIT_11 => X"81C012060000000000218F7840000100800004000000000066C0000080080000",
INIT_12 => X"800000000017C000100000000001A800080000000001A8040000002840008185",
INIT_13 => X"0000000006F00000100200000000012600001004000000000066000000801040",
INIT_14 => X"0000200410100000000005F00000020080090A0000000085C800002000586000",
INIT_15 => X"FF00400000000000020020020001000040283024E4F2860400008000030ED080",
INIT_16 => X"00000000000000000000000000000004010201001003020200000000000127DB",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"A0700030038200010089120104D2040020000000000000000000000000000000",
INIT_1A => X"2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2C30C30C30C30C306982121A1E79E79",
INIT_1B => X"32190C86432190C86432190C86432190C86432190C86432190C86432190CB2CB",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000432190C86432190C864",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0201000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF552A974AA0004174BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA0804",
INIT_29 => X"7FFFFFFFFFFFFFFFFFFFFFFEF552E954AA000400000F7FFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E954BA007FC00BA087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974BA082E9540000",
INIT_2B => X"FFFFFFFFFF7FBFDFFF552E974BAA2FFFFE10FFFFFFFFFFFFFFFFFFFFFBFDFFF5",
INIT_2C => X"FAAD57FEAA007FFFFFFFFFFFFFEFF7FBFFF550800020BAAAD56AAAAF7FFFFFFF",
INIT_2D => X"EFF7D56AB450000021EFA2D57DE10087FFFFFFFFFFFFFEFF7FBEAB450804001E",
INIT_2E => X"000F7FFFFFFFFFFFFDFEFA2D568B550004001EFAAAEA8ABA5D7FFFFFFFFFFFDF",
INIT_2F => X"FFFF5D2E954AA080005000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFEF552A974AA0000104AAFFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"A954AA082A92428087FFFFFFFFFFFFFFFFFFBFDFEF5D2E974AA000A07000E3FF",
INIT_32 => X"FFFFFEFF7FBFFFFF552E974AA0071C50BA1C7FFFFFFFFFFFFFFFF7FBFDFFF5D2",
INIT_33 => X"EDF6FABAEBFFFFFFFFFFFFDFEFF7F5FAFC7492A974AAB6F5F8E10E3FFFFFFFFF",
INIT_34 => X"EBF5E8B550000071EFB6DF7AE921C7FFFFFFFFFBFDFEFE3F5F8F450004050AAB",
INIT_35 => X"A497FFFFFFF7FBF8FC7EBD168B450804021FFB6D57DE28147FFFFFFFFFBFDFC7",
INIT_36 => X"00000000000000000000FFFFFFFEFF7F1F8FD7AAD16AB450000001FFBEA4A8AA",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2A954AA0800174100000000000000000000000000",
INIT_38 => X"74AA002E95410A2FFFFFFFFFFFFFFFFFFFFFDFEF552E954AA0004000AAFFFFFF",
INIT_39 => X"FDFEFF7FBFFFEF552E974AA082A820AA087FFFFFFFFFFFFFEFF7FBFDFFF5D2A9",
INIT_3A => X"568A00AAFFFFFFFFFFBFDFEFFFFFFDFEF5D2E954AA0051554BA557FFFFFFFFFF",
INIT_3B => X"D16AB450804174AAFFFFFFEBAA2FFFFFFFF7FBFDFFFFFD568B55002A954AAF7D",
INIT_3C => X"57FFDFEFF7FBFFF55A2D16AB550000175EFFFFBEAA005D7FFFFEFF7FBFDFFFAA",
INIT_3D => X"0004001EFFF842AAAA087BFDFEFF7FFEAB45A2D568B550804001EFF7D57DEBA5",
INIT_3E => X"0000000000000000000000000000000000000F7FBFDFEFF7D56AB45AAD56AB45",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(20),        -- Port A data input
DOA(0)   => data_read_a_lo_256(20),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(20),        -- Port B data input
DOB(0)   => data_read_b_lo_256(20),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_21_14 : RAMB16_S1_S1
generic map (
INIT_00 => X"4A302428B824900A128C090A5C1800261500213C005FE812D10420054085A202",
INIT_01 => X"001FFE3440B609703B0427F801A40B8115BC4F655300340288A40D30040E4DD8",
INIT_02 => X"E00424256888D8819801000F9FFFFFFFF149FF1FCA448046C60A0D2437C517F9",
INIT_03 => X"20030640003250640003250F06002CC1740002019824E001CD357832440001FF",
INIT_04 => X"EA2C3FFD400006E04401A8837001FFFC004AEF00080B70E08FB5789421007C5C",
INIT_05 => X"00011A0C40F9FFF80920954FF0F00809DF84A0202879800000F3000029980780",
INIT_06 => X"0805984B7A1FC0A0000101FFF0480080002281F7C3C381F87C03DFFF00009004",
INIT_07 => X"B424068086A205481A60A19000908204A855B000A08A61FF20C3D004D331D340",
INIT_08 => X"1BFA0001600802000023F7FFC08D234B40C2028253000040114200000D0226C0",
INIT_09 => X"EF1F5FF054096C6ADBA169FFC202B1C1FFBEF0440021083DFFCE22DC2880E24D",
INIT_0A => X"45FF0C004041D84862A28C54518DBFF00020004C0A6044901112A0908AA0A300",
INIT_0B => X"018C241102068006C620C03882019480E63180855A492712CC01C49C20201BFE",
INIT_0C => X"08A9464116544302C02D92236488D92236488D92236488D922366446C911B210",
INIT_0D => X"08800444021048034004001890000806002804A0822189000900D80621FFBE00",
INIT_0E => X"060580261013813A2CC396506102C4053FFD5BFF00A04A00200602CA52001100",
INIT_0F => X"080C0B004C202621A85C09411500135844C196D3606941018150098404C1A304",
INIT_10 => X"B02901013416181C96C2C9C600890A2028172192C460D1820302A0130809834A",
INIT_11 => X"9C5E803408250180AC268D185DB3F4350B811068C00049A0A4AA68F05C96A001",
INIT_12 => X"002C006560138F032B1804101244C883052208209040CC849063A747512B7678",
INIT_13 => X"41401E240665750440C9488280254530314080C2C601040420352148A00501B1",
INIT_14 => X"500811204D000700114204A70422016149916011008CAA8858850B00C32591C0",
INIT_15 => X"FFC06E60AC0496022300233104663040808E991765205000070121D41D18D098",
INIT_16 => X"40100401004010040100401004010040102090010008000001C0E010020007DF",
INIT_17 => X"0100401004010040100401004010040100401004010040100401004010040100",
INIT_18 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_19 => X"FFEF9FEEFF7FFDF7FF3E3DFDF7E0000000000000000000000000401004010040",
INIT_1A => X"BEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBFFDFDFFFCF3CF3F",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFEFF7FBFDFEFF7FBFDFEFBEF",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000FFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0001000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E954AA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0004",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA0004154BAFFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"52E974BA0804000AAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0004174BAFF",
INIT_2B => X"FFFFFFFFFFFFFFFFEF552E954AA000400000007FFFFFFFFFFFFFFFFFFFFFFEF5",
INIT_2C => X"A082E95400007FFFFFFFFFFFFFFFFFFFFDFEF5D2E974BA002E97400007FFFFFF",
INIT_2D => X"FFFFFBFDFEF5D2A954AA002E974BA087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFBFDFFF5D2E954BA007FC00BA5D7FFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA000002000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080005000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"A974AA0000104AAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974BA0000174AAFFFF",
INIT_32 => X"FFFFFFFFFFFFDFEF552E954BA080A000AAE3FFFFFFFFFFFFFFFFFFFFFFFEF552",
INIT_33 => X"02A95400087FFFFFFFFFFFFFFFFFFBFDFEF5D2E974AA000A07000007FFFFFFFF",
INIT_34 => X"F7FBFDFFF5D2A954AA082A924281C7FFFFFFFFFFFFFFFFFFBFDFEF5D2A974BA0",
INIT_35 => X"A557FFFFFFFFFFFFFFFF7FBFDFFF552E974BA0020924BA1C7FFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000E3FFFFFFFFFFFFFFEFF7FBFFFFF552E974AA0071C50B",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0000020000000000000000000000000000",
INIT_38 => X"74BA0000174BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954AA080017410FFFFFF",
INIT_39 => X"FFFFFFFFFFDFEF552E954AA0004000AAF7FFFFFFFFFFFFFFFFFFFFFFFEF552A9",
INIT_3A => X"E95410087FFFFFFFFFFFFFFFF7FBFDFEF5D2A954BA082E800AAA2FFFFFFFFFFF",
INIT_3B => X"FBFFFFF552E954BA002E97410087FFFFFFFFFFFFFEFF7FBFDFFF5D2A974AA002",
INIT_3C => X"57FFFFFFFFFFFDFEFF7FBFFFEF552E974AA082A820AA557FFFFFFFFFFFFFEFF7",
INIT_3D => X"5D2E954AA0051554BA5D7FFFFFFFFFBFDFEFF7FFFFFEF5D2A974BA0000020AA5",
INIT_3E => X"0000000000000000000000000000000000000AAFFFFFFFFFFBFDFEFFFFFFDFEF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(21),        -- Port A data input
DOA(0)   => data_read_a_lo_256(21),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(21),        -- Port B data input
DOB(0)   => data_read_b_lo_256(21),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_22_14 : RAMB16_S1_S1
generic map (
INIT_00 => X"5290F4CDE914905A14A43D33F488243E17122300F55FEB189B343A1140548380",
INIT_01 => X"A54007B259F6A975386262000C344BA9573C6FF57B18A5FB0ABFCD3C2C5F4F0C",
INIT_02 => X"021DFF8C38B3C009D203551040030071869D0040180AA2DC53DB89BEA8204001",
INIT_03 => X"2603475A969D0475A969D0460EAA401005111011BD506954EDB40F5EF41434C0",
INIT_04 => X"922D9002100ED69E443D988B0D5400103E48003D0800011E803B06B5B9125A15",
INIT_05 => X"281B5A0C06000408F4DF9422010D8802022F2124A8022492580040440002021C",
INIT_06 => X"F780C4C052881ADA0E05440205DA50930FA182010004700083E220800440B588",
INIT_07 => X"049D028B93FB561833D8094A02F5EA92FD7247E10305C40040D136E6A023F7FC",
INIT_08 => X"00028241680A0E002A9400803A884B5B5206B7C2E53CA25144009007A64EBD64",
INIT_09 => X"41008810240240C6694008010392354010000560141801002028A83D2A08E06D",
INIT_0A => X"34000000848BCA6902A29C54539C020E11810098D4067EFF9FF284D483E2AB41",
INIT_0B => X"500001840000C80B410014088040F4A944B1AA313C0022AA0011C0DC00028001",
INIT_0C => X"80B14004D158C8CA24A1C2A870AA1C2A870AA1C2A870AA1C2A872550E1543800",
INIT_0D => X"80A14050A01509E050854498B5281A1C34E506A2C6898B52A154DAC6B6000850",
INIT_0E => X"0B03001A483A4146603050080410089180008800143D83888281A2034A850142",
INIT_0F => X"A4160600349075238473F1210006133835E92273612B3482C090068A0E84AC56",
INIT_10 => X"30060181BA1B13959DC08DA902458870201970B29602562B0581200D141D0959",
INIT_11 => X"E042021C040D0152C8058B3840F044708E7E1C20A0106EA166C13AFC14AA3804",
INIT_12 => X"080E004B0C17C1439A9838301DC1A8438EA32C009DC1A8255300650458A1D588",
INIT_13 => X"018010E186F110A908E3A8CB0026C9A610A908E6A60F0807626610E160589C4C",
INIT_14 => X"2A701667334005800B1605F043858125E0D04110408D2485CA034681E43A1E40",
INIT_15 => X"00646002304244A91102C93A2D608D2A258DF8034188200C050171A41108F084",
INIT_16 => X"110441104411044110441104411044110466C440446CA06951D4EA8010009804",
INIT_17 => X"0040100401004411044110441104411044110441104411044110441104411044",
INIT_18 => X"0401004010040100401004010040100401004010040100401004010040100401",
INIT_19 => X"F7DFBFDEFE8FF1F7DEBDDF7DF7D05122890000000003FFFFFFFF900401004010",
INIT_1A => X"9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7BFFDFD7DDDF7DF7D",
INIT_1B => X"F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE79E7",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000003F9FCFE7F3F9FCFE7F3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA000400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0800",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000002000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2A954BA000015400FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080402010FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2A954BA0004154BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A0004174BAFFFFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0800154AAFFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF552A974AA0000174BAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974A",
INIT_2E => X"000007FFFFFFFFFFFFFFFFFFFFFFEF552E974BA0804000AAA2FFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080400010000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E954AA080005000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000402010FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2A954BA000417410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"804154BAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974BA0000174AAFFFFFFFFFFF",
INIT_34 => X"FFFFFFFEF552A974AA0000104AAE3FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0",
INIT_35 => X"AA2FFFFFFFFFFFFFFFFFFFFFFFEF552E954BA000E124BAE3FFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000007FFFFFFFFFFFFFFFFFFFFDFEF552E954BA080A000A",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804000100000000000000000000000000",
INIT_38 => X"54AA000400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2A954AA080017410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"0174BAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A954BA000415400FFFFFFFFFFFFF",
INIT_3B => X"FFFDFEF552E974AA0804174AAF7FFFFFFFFFFFFFFFFFFFFFFFEF552A974BA000",
INIT_3C => X"2FFFFFFFFFFFFFFFFFFFFFDFEF552E954AA0004000AAA2FFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2A954BA082E800AAAAFFFFFFFFFFFFFFFFFFFBFDFEF5D2E954BA002A820BAA",
INIT_3E => X"0000000000000000000000000000000000000087FFFFFFFFFFFFFFFF7FBFDFEF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(22),        -- Port A data input
DOA(0)   => data_read_a_lo_256(22),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(22),        -- Port B data input
DOB(0)   => data_read_b_lo_256(22),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_23_14 : RAMB16_S1_S1
generic map (
INIT_00 => X"EF20906D902424807BC8241BC81801B97D38AD3C0800103362A6741C80A12A02",
INIT_01 => X"001FFF8409F089003B4422000D80C80106804A7951C5B9D1C828043EA28838F9",
INIT_02 => X"E01CEE21649C82C40800000F9FFEFF8E72CA7F5FC2E22809925A0D3611C877F8",
INIT_03 => X"24000400402670400402670D48222DC1764446838624000080007460C40001BF",
INIT_04 => X"68403FFC020560E0443E21037C01FFFC0002EE00628BF0E02FAD781014085014",
INIT_05 => X"0112000202FBFFF00920017FF0F0628BFF8488890979800002F702002BB807A0",
INIT_06 => X"EF85788B681FC000000001FFF0010000000001F7CBC385F87C0BFFFF20040001",
INIT_07 => X"F6E200000000C1440E3AE408009120071070FA07A1CB23FFA403F0C4D23BF7C0",
INIT_08 => X"0BF87CA400804000003FF7FFD8880A034AC09662305AB10555421006891A1089",
INIT_09 => X"BE1F5FEA10092C0896A243FFC0008087FFBEF2000000001DFFC612C0C0400100",
INIT_0A => X"41FF0C2060501000600000000001BFFA800808189A657EF81DD0C00079CC8001",
INIT_0B => X"018C24110A860006C620C0312241C482B20400CC52492710CC80060020A81BFE",
INIT_0C => X"0C08866907048320C20C10030400C10030400C10030400C10030400608018210",
INIT_0D => X"040002000041500300100040000500C000801000C02400000952800001FFBF04",
INIT_0E => X"FC850015385380380CDB86106502C5043FFD5FFF00A04BC010A7724B10000800",
INIT_0F => X"89F90A002A70A710A51C01C05904014861433602A1CAF13F2110055614C72FC0",
INIT_10 => X"E02D02001C1E14981B43253EE50C8220180F1082E06397E07E42200AAC298E57",
INIT_11 => X"8421802400A90022B0070FAE18019214A380344920080B21A58B02AC60BACDF0",
INIT_12 => X"0A2A000C480B0704B54028101AC49C84BB4100009AC49C80857A82D20CE8CB22",
INIT_13 => X"01E00C8103416445C12ED0400027C5292445C12D500B0005A62D344CB241D095",
INIT_14 => X"132C907425604680038706A35132C94BDD011010404428886AC91B11311C8280",
INIT_15 => X"FF000470BE0692020328CA0028042054A92771C50FC070110001C1680809591D",
INIT_16 => X"00802008020080200802008020080200800800200200000000000008004807DF",
INIT_17 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_18 => X"8020080200802008020080200802008020080200802008020080200802008020",
INIT_19 => X"0000000000000000000000000000000000000000000000000000008020080200",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080002010FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974AA000400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000400010FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974AA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080000010FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E954AA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954A",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA000015400FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080002010FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974AA000400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000402010FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E954AA080005000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA080407000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA00041741",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080000010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000402010FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2A954AA080002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954AA080017410FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"552A954BA000415400F7FFFFFFFFFFFFFFFFFFFFFFFFF552A954BA080015410F",
INIT_3E => X"0000000000000000000000000000000000000F7FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(23),        -- Port A data input
DOA(0)   => data_read_a_lo_256(23),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(23),        -- Port B data input
DOB(0)   => data_read_b_lo_256(23),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_24_14 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100600007FFF000080108004000800020000840041000080808",
INIT_02 => X"FC5CA803400EB8209000000F9FFEFF8E7240FF1FC22409EA04018E50074017F0",
INIT_03 => X"11100400000000400000000D00002CC07400000090C080019001010A000001BF",
INIT_04 => X"68003FFC00040000000000008001FFFC0002EE00000370E007A100000000E468",
INIT_05 => X"0000000000F8BFF00920004DF0F00001DF8000000079800000F3000029980780",
INIT_06 => X"6E461803081FC000000001FFF0000000000001F7C3C380F87C019FFF00000000",
INIT_07 => X"600C2400013649609C8000980040814210254000A00B21FF2003F2A80D500000",
INIT_08 => X"0BF80000000000000003F7FFD88D2B4A02C0940062EC2804001610020408178B",
INIT_09 => X"8E1F5FE010092C0892A041FFC0000001FFBEF0000000001DFFC002C000000000",
INIT_0A => X"41FF0C0000000000600000000001BFFA0000005501AA00000CE2000009400000",
INIT_0B => X"018C0411020600048620C030020502000200000400490510CC00040020201BF4",
INIT_0C => X"0808064106040300C00C10030400C10030400C10030400C10030400608018210",
INIT_0D => X"0000000000004003000000000000001200580000000000000000000001FFBE00",
INIT_0E => X"0086C022005381380FDB96516140C6043FFD5BFF000041000000004110000000",
INIT_0F => X"80010D804400A7240C840C201D0210840043B4804012500021E0088014C04940",
INIT_10 => X"4109038041021C980200D06410C1924030008142E06024A00043C01100298092",
INIT_11 => X"587CC200002100C14428090A1D02348190814C09C010104025AA40041A0D8005",
INIT_12 => X"022E0030300B0E46177004208000D8C61D7004300000D884817B00011306B2D9",
INIT_13 => X"01E003060344710009875C018100013831000985DC000C20003C310006143B70",
INIT_14 => X"4001850EDC004780144806A64400186CBF8961104000C3807884000846EB9500",
INIT_15 => X"FF0006E08C063C0220002201490418082010A57263E0100008000290161E711C",
INIT_16 => X"00000000000000000000000000000000000000000000000000000000000007DF",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"F2D0AEEAF6E7CC1132CDB4441990000000000000000000000000000000000000",
INIT_1A => X"BEFBE79E79E79E79E79EFBEFBEFBEFBEFBEF9EF9EF9EF9EFA69861219575D75F",
INIT_1B => X"783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1EFBEF",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000783C1E0F0783C1E0F0",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0201000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A000400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA000400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000400000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402010000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"00002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080002010FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000400010FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA00040000",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020100000000000000000000000000",
INIT_38 => X"74BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"000010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA000002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974AA000402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000002010F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(24),        -- Port A data input
DOA(0)   => data_read_a_lo_256(24),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(24),        -- Port B data input
DOB(0)   => data_read_b_lo_256(24),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_25_14 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100200002000000080100004000000020000800041000080808",
INIT_02 => X"FC400086000000800000000F9FFEFF8E738FFF1FC204010000000111568DD7F8",
INIT_03 => X"00000400000000400000000D00002CC4740000008000000080000000000001BF",
INIT_04 => X"68003FFF64A564AC000000000001FFFE0082EF00010370E007A1000000004000",
INIT_05 => X"0A00040148F8BFF80920804DF0F00101DFC040000079C92484F30499299837C1",
INIT_06 => X"66041803081FC0E0801101FFFD000E41002299F7E3C380F87C019FFF81200096",
INIT_07 => X"000000080480AE00000080000000000000000000A00B21FF2003E00000000000",
INIT_08 => X"1BF80000400A02000003F7FFFA0008000200A0400008A0000014100200081000",
INIT_09 => X"8E1F5FFA53EFBCACB2E369FFE0010001FFBEF80C40630C7DFFEEBAF000800202",
INIT_0A => X"41FF0C0600000000600000000001BFFE00301000000000000CC020000140000C",
INIT_0B => X"01DCCC31222730A49620C030020100000200000400490D10EC00040220201BF4",
INIT_0C => X"0808064106240300C00C10030400C10030400C10030400C10030400608018210",
INIT_0D => X"0883044582114013412080000000000000000000000000000012800001FFBE00",
INIT_0E => X"00040020000180380FC386106140C6043FFD5BFF00A04B80608003CB120C1106",
INIT_0F => X"0000080040000200040400000100000000009480000240000100080000400900",
INIT_10 => X"0001000000000808000000240000020000000100006004800002001000008012",
INIT_11 => X"0001001808220000002004001900000080800008000000000022400000088000",
INIT_12 => X"0010000000000E00110000000000408009000000000040808063004000008200",
INIT_13 => X"6000000000046100000240000000001021000004400000000010210000001010",
INIT_14 => X"4000000404000800000000060400000088000001800000001084000000088000",
INIT_15 => X"FF800C608C041002000002000006100000002100000000180600000000100018",
INIT_16 => X"4110441104411044110441104411044510629041040D180400000010028047DF",
INIT_17 => X"1104411044110441104411044110441104411044110441104411044110441104",
INIT_18 => X"1044110441104411044110441104411044110441104411044110441104411044",
INIT_19 => X"FBA2894A196A8C5A2932EC15DA080800002FFFFFFFFFFFFFFFFFC11044110441",
INIT_1A => X"2492492492492492492410410410410410410492410492412000531215A69A6B",
INIT_1B => X"158AC562B158AC562B158AC562B158AC562B1588C46231188C46231188C49249",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000B158AC562B158AC562B",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080000010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000010FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08000000",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(25),        -- Port A data input
DOA(0)   => data_read_a_lo_256(25),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(25),        -- Port B data input
DOB(0)   => data_read_b_lo_256(25),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_26_14 : RAMB16_S1_S1
generic map (
INIT_00 => X"E9264EAB20190CA3BA4997AA9002AE9C001006B0778015CFA17E0811039879C7",
INIT_01 => X"2FFFF9BB1F773C7F9BB07DFFFDD863FC5FFF3FEFFBBF9FFB22FFFBC7B9F30686",
INIT_02 => X"E06CCC62052E708180F6FFBFFFFCFFFFF9C7FF7FC24332E642090000074037F6",
INIT_03 => X"428003739CD9863739CD9869FE2B7DEAF300029E4E300DFE69A6E644E6FF473F",
INIT_04 => X"7C2FEFFFF5BA124F003DD31EAFFFFFEE9FF7EE6F4C0770FFD7DC7CA53997B2B1",
INIT_05 => X"DFFB5421C1F8BBFAFDBFFACDF0FFCC05DDDBFF3690F9EDB7F5F7AFF639BD7DE3",
INIT_06 => X"EFD044ABC817C3E3A74667FDFFB6FF5727CC3BFEF7C3FAF87FF59F7FFBFEF69F",
INIT_07 => X"00003002132462052E708180EF060C18E5BEFB051225CDFF7002C4EEDE77F6E0",
INIT_08 => X"3FFF7D5000EC75088ED3FF7FC8790E46426CE06CB1F8E041051831FA3068D77E",
INIT_09 => X"C05FD7FF9BEFBDCEFBEE59FEF44F6603EFBEFAFCC2E35E7FDFD147CCF3F583FA",
INIT_0A => X"67FF1C7FBFADEB31E35768E8ED6BFDF3EB3EBF9DDBCE7FDC1DF8A760F3EACC02",
INIT_0B => X"5BDDCC3B336F7C548667D47B7737AF3FD62601EDC25B3533DCEB07F262213FFC",
INIT_0C => X"5F9A06E19F4D93A0EA0F78C35E30D78C35E30D78C35E30D78C35E986BC61AE31",
INIT_0D => X"5FD7AFEFDFFAF59B6FF28FE1D80D73D840607307DCFE1D80EF69A004DFFFF7FF",
INIT_0E => X"0004001F8041897B2FFFC6D86D70CE04FFFFF3FF1F5F5475BD7F72E4D75EBFAF",
INIT_0F => X"F60008003F008237B0040A00010003E020023E0201F45EC0010007E01047D17B",
INIT_10 => X"00010001DC0004C81003DE050A700200001DC0006863E8BD8002000FC0208FA2",
INIT_11 => X"2200E400002801E1A00004C21C0206F60081800800007B00010F02007EC09A0E",
INIT_12 => X"0880007E000807C7C1A612001E0015C7C19C22001E0015C59DFE82011A311AA0",
INIT_13 => X"00001BC00101F60409F0670840070809760409F06984800780097604067D0010",
INIT_14 => X"81019F40042100001F800203D81019EC085614000085C80023D81009CF008A74",
INIT_15 => X"FF802FFDFFAFD082003B032FB987E04021D481D4000819060801E0D00001231D",
INIT_16 => X"EBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEFFBFBFBFBBFCFBB0FFDFEFFEF2DFFFFFB",
INIT_17 => X"BFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAF",
INIT_18 => X"FAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFE",
INIT_19 => X"475B15BCF491E166CC8553F86EDB5C88646FFFFFFFFFFFFFFFFFEBFAFEBFAFEB",
INIT_1A => X"861861861861861861861861861861861861869A69A61861AFBD54D5F871C71D",
INIT_1B => X"984C26130984C26130984C26130984C26130984C26130984C26130984C261861",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000984C26130984C26130",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040201",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(26),        -- Port A data input
DOA(0)   => data_read_a_lo_256(26),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(26),        -- Port B data input
DOB(0)   => data_read_b_lo_256(26),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_27_14 : RAMB16_S1_S1
generic map (
INIT_00 => X"00080A40000A41248002029000050A088000008242A0004404480002000A1155",
INIT_01 => X"2FFFF1C11F781C129C107DFFFE0860941E81258CA2B71C2220EC1B86E1A00002",
INIT_02 => X"E1000000810000014400FF6FFFF0FFFFF8007F1FC21110005080200000221FF0",
INIT_03 => X"4080026318C18226318C1821302232EAE00002BE001115FE48620040840A863F",
INIT_04 => X"643D4FFC2530000F003D821C0BFFFF8E9EF79E6D440748FED70060842105B0B0",
INIT_05 => X"D6F39020D1F8A3FAFDBFBACDC8FDC405D1DB7F1490E5EDB7D5CBADB2385D79C3",
INIT_06 => X"6FE000A38007C3032646EFF1F0B6FF46A78C39F8E723F2E47FE59C7F9ADA2612",
INIT_07 => X"00002820000000810000014401060C180190310540118DFF1000C0849673F6C0",
INIT_08 => X"3FF779100062B12A8EC3F47FC80208808210880C00082050000110023068D030",
INIT_09 => X"005F07E09BFFBD07FBAC09F8E42922038F7DF8BEC2E39C5F1FD047CEF1B582D8",
INIT_0A => X"63FF5D5F9FADE911E81C09818109E1F16B16B71092CE7ED81CF403601228C402",
INIT_0B => X"1BFDCC39732F3554866AD57C37BEAF1C152201A4C05B7531D56B05B06A213FF8",
INIT_0C => X"5BCA06F18FC59380F00E34430D10C34430D10C34430D10C34430F0861A2186B5",
INIT_0D => X"5B56ADAB5FAAE58B2F628EA0C80FA3F04040510768EA0C80CC61A0044DFFC6EB",
INIT_0E => X"0004001D800188792CE79715710AE4047FFD23FF315D54358D593474955AB6AD",
INIT_0F => X"520008003B000297B0040200010003E020001F0201E44A400100076000579129",
INIT_10 => X"00010001DC00004A10035E0408300200001DC000086BC8948002000EC000AF22",
INIT_11 => X"02002400002801E1A00000C01E0202F60080800800007B00000782006EC0820A",
INIT_12 => X"0080007E000006A7C10602001E0001A7C10C02001E0001C18DE282010A311AA0",
INIT_13 => X"00001BC00000FE0401F04300400708007E0401F04180800780007E04047D0010",
INIT_14 => X"81011F40040100001F800002F81011EC080604000085C80001F810094F008034",
INIT_15 => X"FF800C6DDDAFD082001B03249887E04001D481D4000009020801E0D00001021F",
INIT_16 => X"AB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6BF1EBDABD8E270BF84A25C6ACB777E3",
INIT_17 => X"B6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6AD",
INIT_18 => X"6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADA",
INIT_19 => X"490E2168100481CA860402104A471688747FFFFFFFFFFFFFFFFFAB6ADAB6ADAB",
INIT_1A => X"000000000000000000000000000000000008200000000000200072F210000001",
INIT_1B => X"05028140A05028140A05028140A05028140A0500804020100804020100800000",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000A05028140A05028140A",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040201",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(27),        -- Port A data input
DOA(0)   => data_read_a_lo_256(27),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(27),        -- Port B data input
DOB(0)   => data_read_b_lo_256(27),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_28_14 : RAMB16_S1_S1
generic map (
INIT_00 => X"02200AA400180030808802A900002A08001280A08A801044104A1000001818C3",
INIT_01 => X"0AA00011460214428114180000882214413D0A71592A01D92213D28005210202",
INIT_02 => X"0451110A012100884000AA30200000000C100040104112101100008888200000",
INIT_03 => X"448000318C52A20318C52A20148810200111100C211004AA00034204200A2200",
INIT_04 => X"04004001001A90110000121402AA0000003C00000500000040080421080D0080",
INIT_05 => X"4060000C8001000000002E000000050000001610300000010000802202040012",
INIT_06 => X"1000002080001111001222000425A1040026A008000000000000000009328280",
INIT_07 => X"2491008A00491201210088400122448908A20402000408001000040820000000",
INIT_08 => X"20058310402A160026500000028040101004200C840082115554000112244814",
INIT_09 => X"4140000800000060000720000102028000000490160801020002200011100010",
INIT_0A => X"020000081B34211082B694D4D294000020020381040000000200032040004400",
INIT_0B => X"4800210C19808400500010009110091500020B408810000100200020408B0000",
INIT_0C => X"01028000080118020023604858121604858121604858121604858090B0242C00",
INIT_0D => X"010000800920040804020A6058003108402043058C460580653020005A004039",
INIT_0E => X"00000002800008014004104104420A00C000200005000010040A0020CC000200",
INIT_0F => X"520000000500000010000200000000000000280000040A40000000A000001029",
INIT_10 => X"00000000000000C0000002000830000000000000480008148000000140000020",
INIT_11 => X"020024000000000000000440000000020000800000000000000C00000040020A",
INIT_12 => X"00800000000001804006020000000500400C0200000005400A90000000100000",
INIT_13 => X"0000000000018200001003004000000142000010018080000001420000200000",
INIT_14 => X"8000080000010000000000018800008000060400000000000310000008000034",
INIT_15 => X"000002040080000000110006B081400000400000000009020000000000002200",
INIT_16 => X"802008020080200802008020080200802101210810C39A66A90A85420413A820",
INIT_17 => X"0200802008020080200802008020080200802008020080200802008020080200",
INIT_18 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_19 => X"DE21102C110A00246972BD89A40A0C22E1000000000000000000002008020080",
INIT_1A => X"2082082082082082082082082082082082082082082082080D35050758C30C31",
INIT_1B => X"0582C160B0582C160B0582C160B0582C160B0580C06030180C06030180C08208",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000B0582C160B0582C160B",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(28),        -- Port A data input
DOA(0)   => data_read_a_lo_256(28),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(28),        -- Port B data input
DOB(0)   => data_read_b_lo_256(28),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_29_14 : RAMB16_S1_S1
generic map (
INIT_00 => X"79964E4BA01DACAB9E659792D00AAE160002829C7FDFEFCEE97C2815039D70C3",
INIT_01 => X"0ABFF9AB0775343F9AB01DF80D5821FC0FFF3FEFD1AF9FF1207FFBC7B9720586",
INIT_02 => X"002CCC60050E700080F6AAA7BFFC007189C7FF2FC00330E602800000074037F6",
INIT_03 => X"468003210868A63210868A68DA017D207200021C4E200CAA6186A40042FF4300",
INIT_04 => X"7C2FE002F0900001003C5316A6ABFFE21F36E02F0D03701F47D41800109FB281",
INIT_05 => X"4979440580F9B808F49F6A4DF00F8D01DC4B97369078249370F482E62BA41462",
INIT_06 => X"B250442BC81001E1870223FC0BF7F11507C423FE33C078F803F19F00E936721D",
INIT_07 => X"00011080012460050E700080EF020408EC8CFA01122149FF700200665A35D260",
INIT_08 => X"2BFD055040A452000443FF00007906464068406C31F84000000831FA1028575A",
INIT_09 => X"805FD017102690AA694551FE30444681E0820AD40201423FC00122C493500172",
INIT_0A => X"0600002AFFBE2330815568A8AD6ABC02A02A0B0CCB463B4C0748A720B1EA4C00",
INIT_0B => X"0850400A11414C005005000B51158936D20601A98A10200308A002E240010BFC",
INIT_0C => X"05928020194918A22A2268C81A32068C81A32068C81A32068C81A99034640C00",
INIT_0D => X"058102C48970541944B20FA1580561D040406305587A158046282000DBFFF13D",
INIT_0E => X"000000028040890327DCD28928324400DFFFF0001F1F0050342D42A086040B02",
INIT_0F => X"F60000000500802010000A000000000000022A0000141EC0000000A01000507B",
INIT_10 => X"00000000000004C0000082010A700000000000006800283D80000001402000A0",
INIT_11 => X"2200E4000000000000000442040004020001800000000000010D000010401A0E",
INIT_12 => X"08800000000801C040A6120000001540409C2200000015441DAC800010100000",
INIT_13 => X"0000000001019600081027084000000956000810298480000009560002200000",
INIT_14 => X"800088000021000000000201D800088000561400000000002358000088000A74",
INIT_15 => X"00802594A282C0000033010FB181E00020400000000819060000000000002305",
INIT_16 => X"C0B02C0B02C0B02C0B02C0B02C0B02C4B12B312912831A27FCFE7FFB175B6FF8",
INIT_17 => X"0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02",
INIT_18 => X"B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C",
INIT_19 => X"BBCF9F96EE7FFDF7FE783FFDFFEA0C00602FFFFFFFFFFFFFFFFFC0B02C0B02C0",
INIT_1A => X"EFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEEBAEBAEBAEBAEBBFFDF9FBEFFFFFFE",
INIT_1B => X"BFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFBEFB",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000FBFDFEFF7FBFDFEFF7F",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(29),        -- Port A data input
DOA(0)   => data_read_a_lo_256(29),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(29),        -- Port B data input
DOB(0)   => data_read_b_lo_256(29),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_30_14 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"F7FFBFFEFF9FE1F7FFBFFFFDFFD0000000000000000000000000000000000000",
INIT_1A => X"9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7AFBD75F5FDF7DF7F",
INIT_1B => X"F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE79E7",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000003F9FCFE7F3F9FCFE7F3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(30),        -- Port A data input
DOA(0)   => data_read_a_lo_256(30),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(30),        -- Port B data input
DOB(0)   => data_read_b_lo_256(30),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_31_14 : RAMB16_S1_S1
generic map (
INIT_00 => X"129000008004A00804A40000400800020000000C005FEA005800200400050100",
INIT_01 => X"255FF18019700810180065FFFC0040801E80258CA2951C2200EC0906A0804140",
INIT_02 => X"E0000000000000011000550FDFF0FFFFF0007F1FC200000044000000000817F0",
INIT_03 => X"0000024210A30024210A3001002220C06044469200040154482000408400043F",
INIT_04 => X"602D0FFC2420000E003D80080955FF8E1ECA8E2D400340FE870060842100B030",
INIT_05 => X"0213100040F8A3F8FDBF944DC0FDC001D1CB6904A061EDB6D4C30490281831C1",
INIT_06 => X"6FC000830007C202060445F1F0D25E4207A099F0E303F0E07FE19C7F80402412",
INIT_07 => X"0000200000000000000001100004081001103107000185FF0000C0849673F6C0",
INIT_08 => X"1BF27A00000000000883F47FC800080002008000000820440000100220489020",
INIT_09 => X"011F07E013EFBC06FBA009F8E00120038F3CF82C44630C5D1FC002CCE0808248",
INIT_0A => X"61FF0C06C48BC801600000000001A1F00110101092CE7ED81CF0004012288000",
INIT_0B => X"11DCCC31222730048620C4382204A608142002A440492530C401049020221BF8",
INIT_0C => X"0888066187448380E00C10030400C10030400C10030400C10030600608018210",
INIT_0D => X"080204010200418301208480800D02D00040100240A808008840800405FF8640",
INIT_0E => X"0004001D000180780CE386106100C4043FFD03FF101D40008001304018081004",
INIT_0F => X"000008003A000217A0040000010003E02000160201E040000100074000478100",
INIT_10 => X"00010001DC00000810035C0400000200001DC0000063C0800002000E80008F02",
INIT_11 => X"00000000002801E1A00000801C0202F40080000800007B00000302006E808000",
INIT_12 => X"0000007E00000607810000001E000087810000001E000081846282010A211AA0",
INIT_13 => X"00001BC00000740401E0400000070800340401E04000000780003404045D0010",
INIT_14 => X"01011740040000001F8000025010116C080000000085C80000C8100947008000",
INIT_15 => X"FF800C609C06D082000A03200806A040019481D4000000000801E0D00001001D",
INIT_16 => X"010040100401004010040100401004010060C040040C200950402090128057C3",
INIT_17 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_18 => X"0040100401004010040100401004010040100401004010040100401004010040",
INIT_19 => X"00000000000000000000000000001000802FFFFFFFFFFFFFFFFF810040100401",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(31),        -- Port A data input
DOA(0)   => data_read_a_lo_256(31),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(31),        -- Port B data input
DOB(0)   => data_read_b_lo_256(31),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_0_13 : RAMB16_S1_S1
generic map (
INIT_00 => X"ED39BA795990D275FB4A6E96ACC4731DEA4598B0AFB54867F6EE4618C3749803",
INIT_01 => X"8AA0047D8607944AC7DA180001ECA2444042106208408208C20022E9173734B3",
INIT_02 => X"1A7DDD79F9A73E6CCA7DAAF00001000008478020113D98E382FEDF333027C80F",
INIT_03 => X"75D341110C58F31110C58F32A208921F8051500147A0E4AB3493FB3A01EBE240",
INIT_04 => X"86424001531009B100425A97B2AA0001E03501D0A39C8F0078420001106D0C4C",
INIT_05 => X"BCC8CA2EBF03400700402BB20F00239E20341699198600000B08694B16434804",
INIT_06 => X"103FB860B2800161F8432200012DA185F80F24081C3C0707800E600056881308",
INIT_07 => X"B24197ABCDA467F9A73E6CCAFDC3870EEEEC44E2BDFE220094D03022210C011C",
INIT_08 => X"240581B5695EAA80262C080032BF07C7C1FC3F8E94F65B11555EAFFC1C306758",
INIT_09 => X"7E40000BEC004170040DB60017FED1CC0001045002984202003DB931192D60A5",
INIT_0A => X"120071411A74315881A28C141118000C5A85A60444210123820B43B40804674D",
INIT_0B => X"0820008E514045BB514F0106D1D8599581D3A958BC104A89215AC14C48898403",
INIT_0C => X"C261C01C48B1584A0CA3E2687A9A1E2687A9A1E2687A9A1E26870CD061343885",
INIT_0D => X"D274E93A758FA8683AC54B287522E10A74AF4AA59C568752662F5AC218000002",
INIT_0E => X"FF83C002783A0904231C70470C7E0B92800224008AE09FAD4BD48D1FC5D3A4E9",
INIT_0F => X"5BFF078004F075885DFBF7E15C06101C55E921F1F80FAB7FE0F0009E0E903EAD",
INIT_10 => X"F12E0380231F13978FF023FAFDBD9870380230F2D6081F56FFC1E0013C1D207D",
INIT_11 => X"DE7F263C0C8700125C0F8F3C43F1F10BBF7EFC61E01804E1E6C8F8FE807F67FB",
INIT_12 => X"02BE00017C17C1007E5E2E3081C5AC007E6F0E3081C5AC44418D65FE45DEE55B",
INIT_13 => X"61E0042786F103E9F01F9BC3C120C5A703E9F01F978B8C20666703E9F8A0FFED",
INIT_14 => X"FA7E283FFB414F80005F05F10FA7E283F78F6511C048278DCA174FF038FF15B4",
INIT_15 => X"0066A20B61692F293185D8D724E15D3FCC6B7C236FE0691B0700132C1F0EF880",
INIT_16 => X"3A4E93A4E93A4E93A4E93A4E93A4E93A4F942F92E9628540AD2A91442525A000",
INIT_17 => X"A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E9",
INIT_18 => X"4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93",
INIT_19 => X"55F3898E09B56C74DAB15D1CF13501AA495000000000000000003A4E93A4E93A",
INIT_1A => X"082082082082082082082082082082082082082082082082082084E41DC71C71",
INIT_1B => X"E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F82082",
INIT_1C => X"FFFFFFFFFFFFFFF94A5294A5294A5294A5294A52800003E1F0F87C3E1F0F87C3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"3060C183060C187FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"BDEBA0000000000000000000000000000000000000000000003060C183060C18",
INIT_28 => X"168ABA002E82145085155545F7AA975EFFFAABDE00FFAEBDFFF5D2EAAAAAF7AE",
INIT_29 => X"7FFFE10005542145557FD5545FF8000155087FC0155F7D168B55007BFDF45085",
INIT_2A => X"7FFC0010080017555555568AAAFFFFD7545AA8028A00A2802AABAFF8028BEF5D",
INIT_2B => X"FF842AABAA2AE95545FFD168ABAF7AEAAAAAA2FFFDF4500043FE105D2E954BAF",
INIT_2C => X"5007FD7400550415410002E974BA5D5168A00A2D142155005142010FFAE820AA",
INIT_2D => X"FFF780000BA007FE8AAAFF803FFFF5D2A821550000000BA007FD55FF5D7FC014",
INIT_2E => X"000AAFBEAA00007BFDFFF082EBDF455D5142000082E82145FFD17DFEFFFD168B",
INIT_2F => X"DFD75D2AA8A80EA8E2FE3F000000000000000000000000000000000000000000",
INIT_30 => X"68B551475FAF6D1C556F0AA1C24AABEA495FC716F002A975FFE3AA95E00EBAEB",
INIT_31 => X"42A0070071C50BAFEF1FAE0016D56A16D557BC257D415E0216FA3F1E8FC0145B",
INIT_32 => X"8010E004924874825D7FEAA85487FD24AFE3D02DAAAE12BD5545A2803AA00005",
INIT_33 => X"120155EA568E870BAEB8A05A2AEA8B50F55A2F150005A3A438BD04AFAB8F550A",
INIT_34 => X"545E055FFBE81D0BE8EA8A3AA05A2A5504001C74BA42A1571E8028E3DB7816D0",
INIT_35 => X"A5C7E3DFFFE90B45B47ABA497A82FFAFD2A82485FD2415A105C21451ED42A002",
INIT_36 => X"00000000000000000000B55EAAA100AA1D0F6F480B6A555A2A57A002A3D5FDB6",
INIT_37 => X"5EFAAAAB5E1AF3AABFF45592E88A0AFE80A8B0A0000000000000000000000000",
INIT_38 => X"65F520EBE9EF67D7BEA1FD5D556ABEF5D557FEBA55022A3F70C6B405F4D2AE97",
INIT_39 => X"C114728007521170821CE0FDE69411A8DED57CE1055555E5F58EFFC01FE2CACB",
INIT_3A => X"42341D5DEEBEF55080034E0A592A4AD0079C75D6070CC5CBB0280C029ABAA3EB",
INIT_3B => X"7F353AAF6C77F7F20D968BF57812A95E02A2AAB5EB0F280800EFAEE9F5D18F31",
INIT_3C => X"C91565455C141E41887D58AC448B69C30E02116220415A9540AA854140A0A204",
INIT_3D => X"DE6BE93172D7D625B556EEAB157ABEBE1B4D792A4AD1183454180DD3FDCAAAB7",
INIT_3E => X"F0000001FF0000001FF0000001FF0000001FF01EABC4B8014174FF7DA80F52FE",
INIT_3F => X"FF0000001FF0000001FF0000001FF0000001FF0000001FF0000001FF0000001F")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(0),        -- Port A data input
DOA(0)   => data_read_a_hi_256(0),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(0),        -- Port B data input
DOB(0)   => data_read_b_hi_256(0),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_1_13 : RAMB16_S1_S1
generic map (
INIT_00 => X"212C001411984004084D000508C53810A03D1450E839B003342114428A000803",
INIT_01 => X"00000019400B100A8196000000CC004400400002000000000000028001340000",
INIT_02 => X"052137AE8031800C0044009000000000061800001CD4019802AD04CCCFC20004",
INIT_03 => X"04514108C60C21008C6042108400000201440020505100000043C30E10E9F000",
INIT_04 => X"02104001011DEFE088805681920000008000004001900800004002108C280008",
INIT_05 => X"040002340105000200000000080001900010000108040000000008411600401C",
INIT_06 => X"1034001042800808201000000001000820020000102000040000000000800180",
INIT_07 => X"64BF81A15EDFDE8031800C00843060C19E030022103600000450020800040004",
INIT_08 => X"00008004691687AA840008000090248CC84E000046000311555521F183060AC5",
INIT_09 => X"0820800D08100171000DB000154440C800400500000852020011200201012021",
INIT_0A => X"02000040001000880A2A04445004000102002041000001008208001440004140",
INIT_0B => X"4820018A1140440078050040511000102000A008183000010002404400000000",
INIT_0C => X"1000C80008000C030030880C2A030A00C28030A80C2A030A00C28018D4061401",
INIT_0D => X"10040802050080200284401C0022880F009E08008205C0020118088018000000",
INIT_0E => X"0F03C00280000000420860C60C0C0B92C0000000004000010042000040102008",
INIT_0F => X"001E078005000108400005E11C0610000000288058000003C0F000A000100000",
INIT_10 => X"F10E0380000000C202300000008D187038000000480800000781E00140002000",
INIT_11 => X"806302380C870010000004400100110800007861E0180000000C400680000001",
INIT_12 => X"023E00000000018000580C308000050000610C30800005000215006800000101",
INIT_13 => X"61E0000000018100B0001843812000014100B00016030C20000141002880026D",
INIT_14 => X"400A20009B404F80000000018400A20044096111C04000000304026000501580",
INIT_15 => X"0046820040082300218450C2800010094000482141E060190700100000002200",
INIT_16 => X"020080200802008020080200802008020080008008600500A82A1100A8000000",
INIT_17 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_18 => X"0080200802008020080200802008020080200802008020080200802008020080",
INIT_19 => X"81328A46BABEFC54A0810C7452B4428A14000000000000000000020080200802",
INIT_1A => X"AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA28A28A28A28A2A8218D2C0C924925",
INIT_1B => X"E974BA5D2E974BA5D2E974BA5D2E974BA5D2E975BADD6EB75BADD6EB75BAAAAA",
INIT_1C => X"FFFFFFFFFFFFFFFD8C6318C6318C6318C6318C63000002E974BA5D2E974BA5D2",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"70E1C3870E1C387FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"5555500000000000000000000000000000000000000000000070E1C3870E1C38",
INIT_28 => X"EBDF455D2EAABEFF7FFE8BFF5D0002155557FFFFFF007FC21EFA2FFD74AAAAD5",
INIT_29 => X"AA95400552AAAABAFFD1574105D7FD75FFAAAA800AAF7AA974BAFFFBE8B45F7A",
INIT_2A => X"0517DF555D2EAAA1055000015500557DF45AAD1400BAA2AE801550051555EFF7",
INIT_2B => X"FFD540155557FD5400F78028BFFFFFBEAB55F780020AAAA80020AA082EAAB550",
INIT_2C => X"AFF842ABEF5D517DF55552A974AAF7AE820AA0851574BAA2D1574AA5D7BFDEBA",
INIT_2D => X"EFAAD1575EF557FFFE10557FFFFFFFFD56AAAAFFFFD7555AAD168B45AAAEAAAB",
INIT_2E => X"0005D7FFDF4500043FE105D2E954BAF7AE80010082A97410557FEABFFAAFBE8B",
INIT_2F => X"51C7A2FBD5490BFD1C056A000000000000000000000000000000000000000000",
INIT_30 => X"974BAF7FFEFB45FFAABDF55492AA8BC2EBDFEAF7F1F840017D4975D2FEF147FC",
INIT_31 => X"080BEF495FC71D54124924385FAAA8AAAE3D145410F7F1D55D71C002DABAEBAA",
INIT_32 => X"002D082082AB8B6DBEDB7DF7F540E2AE85028B40155145F7AF6DBED5450AA1C2",
INIT_33 => X"78E021FF1471FDEAAFFD56F16D5571D2E28E38E0216FA2D1E8E80140F45082B4",
INIT_34 => X"A2DA3FB7DAAD4AAAAF487BC70BFA97F7AF6D417E92482BF84020BA495557E3FF",
INIT_35 => X"55554ADBD7A2FFC7BEFF6FFD7FC7002FD74951D71EDFFABFD16FAAAE92BD5545",
INIT_36 => X"00000000000000000000547AB8F550A8010E00492487482FFFE82A85EBAE2FFC",
INIT_37 => X"1EF005162BEF047FD5545AAFBF7400FBF9424F70000000000000000000000000",
INIT_38 => X"714F8338AAAA1D0AE974AAF7FFFDF55F7AABFF55082CA8B4DF6C1E8F5E540002",
INIT_39 => X"EABEF75550ACBB7582225FF5843404547184164AA5D2EBEEB0A2D555410D3555",
INIT_3A => X"FEAAEB083BC1000FF8409000512AEABFFDF79DCBF755962010BDCBBC21455D7F",
INIT_3B => X"801F8BA0C57740BDAA0688E5405D57D412F7D55F5E50C7F401BAAE8403CF5A3F",
INIT_3C => X"5D16BABAA3EBC3157ABD5FFE55F2AA9FEAFDF7F431A9F7FFE81FF013A8001AFF",
INIT_3D => X"FB863550229BCABEB7DA403FFFDA2FBF7FED2C7F955445079E280A00C56145EF",
INIT_3E => X"0000000000000000000000000000000000000596EBEF55080034E0A592A4AD00",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(1),        -- Port A data input
DOA(0)   => data_read_a_hi_256(1),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(1),        -- Port B data input
DOB(0)   => data_read_b_hi_256(1),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_2_13 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10E006600180111284380310006289800480032283E000A34301002001A0817",
INIT_01 => X"0005A00810790848048044A54E404350404000720885800802000906E4910200",
INIT_02 => X"407004208400408044C600C50AA055254010541A110222841200000002402544",
INIT_03 => X"0600011004182401004102408C28414043101000408118000145840440F5C415",
INIT_04 => X"5035855703A2900A000CD3088400F40688C9844409060850925E58A4081A0221",
INIT_05 => X"0200840D1021A15AC50494894850890540D1E12020C6E510818500440A280090",
INIT_06 => X"113044094002801020440090A8011A1224AB9380552102442884882A20004097",
INIT_07 => X"000100880004428400408044860000008C022402102100AA40004404B5075460",
INIT_08 => X"15C23440408C862A2A12382A8A5244145048C06085008010141521F000001240",
INIT_09 => X"400582B9033AA0E7AA4110B0506744810554542450694E710A836188C2C00222",
INIT_0A => X"443518360012C2210B020414109130A28038188096A06B8C120CA440A9C00802",
INIT_0B => X"1345E53300EC68005605002964AF222A5704004D080211121C80024200821780",
INIT_0C => X"181080C1110C882202211488452213C88472213C88472213488441109A442231",
INIT_0D => X"008204440210091341208041000810C00000300220201800A908000038AD0284",
INIT_0E => X"00040002804180300E88D28D206A40000554815500481440300000C44A081100",
INIT_0F => X"000008000500828700000000010000000002380000A00000010000A010050000",
INIT_10 => X"00010000000004CA000214000000020000000000684280000002000140200500",
INIT_11 => X"000000000020000000000442100002840000000800000000010C000026000000",
INIT_12 => X"00000000000805A4800000000000152300000000000015801272000100210020",
INIT_13 => X"000000000101C00000C000000000000940000120000000000009600004050000",
INIT_14 => X"0000130000000000000002018000106000000000000000002380000141000000",
INIT_15 => X"55000190000000000002000280000000011080C0000000000000000000002310",
INIT_16 => X"40902409064190641906419024090244902A9003004800415120D4A190804241",
INIT_17 => X"0900409004090641906419064190240902409024090641906419064190240902",
INIT_18 => X"9044090040900409004190441904419044090040900409004190441904419044",
INIT_19 => X"75960040138D70C030B51C50C7D100A2052F81F81F83F03F03F0419044190441",
INIT_1A => X"0410410410410410410410410410410410410410410410410248602081659659",
INIT_1B => X"5128944A25128944A25128944A25128944A25128944A25128944A25128941041",
INIT_1C => X"FFFFFFFFFFFFFFFE1084210842108421084210843FFF825128944A25128944A2",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"7FD5FF555815607FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"2AA000000000000000000000000000000000000000000000007FD5FF55581560",
INIT_28 => X"FC21EFA2FFD75EFAA8415410AA8415555087BFFF55A2AA800BAFFAE954000800",
INIT_29 => X"84155EFA2AEBDEAAA2FBEAABA5D7FE8B555551421455D0002145552EBFEBA007",
INIT_2A => X"2AEBDF555D2E954BAA2AA974BAFFFFE8B45552EBDF45FFAEAABFFF7FFE8B55F7",
INIT_2B => X"AAAAAAAAAFFD1574105D7FFFF555D2AAAAAA5D2E820BAA2FBEAB5555557DF55A",
INIT_2C => X"50055575EFFF84021555D043DEAA5D04021EF557FC21FFAA8428BFFAAAA954AA",
INIT_2D => X"10085568A00FF80175FFA2D17DFEFF7800215500557DF55AA80001FFAA800015",
INIT_2E => X"0005D00020AAAA80020AA082EAAB5500517DF555D042AA10A284154005D00154",
INIT_2F => X"00AAFFAA9543A080038A2A000000000000000000000000000000000000000000",
INIT_30 => X"0017D5D20B8EAA007FC51C7A2FBD55D2BE800042AFE8E1557D0075D2F45BEAA8",
INIT_31 => X"AA8BC7EBDFEAFEFFD00105FFBC20BDEAAA2FBF8AAA557BE8B6D5D5FFABEF4904",
INIT_32 => X"FFEFB6D555578F7DB6A0BDF7D480E174BFA02A974BAF7F5EFB455D2ABDF55492",
INIT_33 => X"ED1FDE90E3A497492B6AAADAAAE3D155E105571D55D71C002DABA5524820BAB6",
INIT_34 => X"BE8F401D7B6A0001470155C51D0092A071555D5E3AE821D00001FF0871C016DB",
INIT_35 => X"5BE8555400550A38428007FED000E3DA3DFD5E3DFFFBD5A38A021551C5F7AF6D",
INIT_36 => X"00000000000000000000410F45082B4002D082082AB8B6D1C5B7DF7FF78E075C",
INIT_37 => X"5EF005560B55F7AA800AAF7AA954AA00042AAA20000000000000000000000000",
INIT_38 => X"ABEF057D68F5F5A00021EF55042AAAA007FD5555AAFBD7545FBB8020A3F7AE97",
INIT_39 => X"7DF55D7AABFF5428ACA8F45A6C1E8F5EFF84165EFF7802BAB0A2FFEAABA557BE",
INIT_3A => X"CA8AA80800020AAF7FBFFFEF04552ABFFFF841FFE75CA882108202E974AAF7D5",
INIT_3B => X"00151FF0C57401E5F3D1E00A1A884174A8FFAEBFEB0A2D55541051555694F002",
INIT_3C => X"2AA801455D7FE8BFFF680800FFF7AAA155F595542455512A975455D3AA8A0055",
INIT_3D => X"5D79FCAF774AE005BE7895554005D2A8A0B882FFFFE10AAAAAB755A66B6AF56A",
INIT_3E => X"00000000000000000000000000000000000000C3BC1000FF8409000512AEABFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(2),        -- Port A data input
DOA(0)   => data_read_a_hi_256(2),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(2),        -- Port B data input
DOB(0)   => data_read_b_hi_256(2),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_3_13 : RAMB16_S1_S1
generic map (
INIT_00 => X"210C00A20020000108430020001600B8156021104940741B3530400E02B92203",
INIT_01 => X"014C9BCA58B1296D24A402C992500B69404040028804A0080A000416A8D90A08",
INIT_02 => X"C12026A484318004404405C9C66E331352180D468B8203980300204442E02B34",
INIT_03 => X"04000748D60D24648D60524C88804D0215011020D15018148040C10A70E1D58C",
INIT_04 => X"18283333240FE41244187308C9104D70944852640901083801750EB0A418C220",
INIT_05 => X"0613142D01912CC2A1B4140528348900C612A104201C689044340ED413A07649",
INIT_06 => X"119000034019881822104C5E68035250A222829710A0A02C18C01A9920842413",
INIT_07 => X"402F00AB0016CA0431800444841020509D038B021230C1990001C644C8273200",
INIT_08 => X"16905000408482088290E8E64010248C4A5AA840C2000110001521F0810A92E7",
INIT_09 => X"0003CE6581BD016342A951AB146C4480530C3B2A8088D3542651670200C1826A",
INIT_0A => X"00735D36209A8A20020894004284B660821030C8990467401218004041020002",
INIT_0B => X"512445B740457154562F957CC08B00093700080D0A4851001D8302D20A0A1530",
INIT_0C => X"00508650008008021021A40861021840869021A408610218C0869810D6043095",
INIT_0D => X"1C8508438450801043A08090380A8834207007022209038080190000999C8F84",
INIT_0E => X"000400200000C0002A48A206204C4205F3304B33004C0041006240140A1C310A",
INIT_0F => X"0000080040000083800400000100000000008400018040000100080000510100",
INIT_10 => X"0001000000000800000244040000020000000100002A0080000200100000A702",
INIT_11 => X"000000000020000000200000080002C000800008000000000022000006808000",
INIT_12 => X"0000000000000A2281000000000040A3810000000000402001400000022002A0",
INIT_13 => X"000000000004200001C0400000000010200001C0400000000010000004490010",
INIT_14 => X"0001070004000000000000060000104C08000000000000001000000903008000",
INIT_15 => X"CC004050CA0C00020220200070040000010401C4000000000000000000100008",
INIT_16 => X"4310E4310A4210A4210A4210A4210A4210A8D0830A68010001B4DA881048061C",
INIT_17 => X"21084290A4210A4210A4210A4210A4210A4210A4210E4310E4310E4310E4310E",
INIT_18 => X"90A421084290A421084390E4310C4390E4310C4390E4310C4290A421084290A4",
INIT_19 => X"015303C0C78C706428A14C586291000A044001FFE000003FFC004290A4210842",
INIT_1A => X"2492492492492492492492492492492492410410410410412821600001249249",
INIT_1B => X"51A8D46A351A8D46A351A8D46A351A8D46A351A9D4EA753A9D4EA753A9D49249",
INIT_1C => X"FFFFFFFFFFFFFFFC00000000000000000000000038F56351A8D46A351A8D46A3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"55AB02055AB0207FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"420000000000000000000000000000000000000000000000007FFFAB57FFFAB5",
INIT_28 => X"A800BAFFAE9554508002AA00AA843DF55FFAA955EFA2D168B55557BEAA000055",
INIT_29 => X"002AB55AAAA955EF005568A00087BE8BFFA2D155410AA8415555087BFFF55A2A",
INIT_2A => X"AAABFF5508003FF555D0002145552ABFEBA007FC21EF007FD75FFAA841541008",
INIT_2B => X"082EBDEAAA2FBEAABA5D7FC0155005168B455D042AB45F7FFD741000042AA10A",
INIT_2C => X"FF7FBEAB55F7AABDEBA5D7FC2010A2D1575FFF7AA975555D2E80145F78415545",
INIT_2D => X"EF5555554AA087BC01FFFFAAAAB55552A954BAFFFFE8B55552EBDE00F7AEAABF",
INIT_2E => X"000082E820BAA2FBEAB5555557DF55A2AEBDF555D2E954BA002EAAABA002A821",
INIT_2F => X"FB7D5D7FEAA3808554203A000000000000000000000000000000000000000000",
INIT_30 => X"1557D1475FAF45BEAA800AAFFAA95578080038A2AA28E3AF55E3A0BA5D7AADB6",
INIT_31 => X"BD55D7BE80004AA1E8E2AB55B6A0925D7085F6AA10087FEABD7AAD57AEBAB68E",
INIT_32 => X"F5D0438140E2FA38B6AEBFF6D1D04AAFFA41040017D5D20B8EAA007FC51C7A2F",
INIT_33 => X"D0A901FFFF801557D1C20B8EAAA2FBE80AA557BE8B6D5D5FFABEF49002FB55FF",
INIT_34 => X"5D20BDE00EBAAA8BC7EBDFEAFEFAB8ABAE925D21C7010EADB525D7FFAE975C75",
INIT_35 => X"F002EADA921420871D74971D24820875C21D5EB8AA8FFF012A954BAFFF5EFB45",
INIT_36 => X"000000000000000000001C24820BAB6FFEFB6D555578F7DB6A0BDF7DEB8E125F",
INIT_37 => X"B55A28408145AAFFFFFFF5D7FEAABA0051400A20000000000000000000000000",
INIT_38 => X"AB55FAD568AA2AFAE975EF555168B55F7AA800BAF7AA955EF00042AAA2A2AEAA",
INIT_39 => X"2AAAA007FD55558A7BD7145FBB8020A35D2ABEF55F7800015F087FEAA00007FE",
INIT_3A => X"968F575D003FF55F7D5420BA5D2ABFEAAF7AE9DFF759A82AEF70800021EF5504",
INIT_3B => X"FFD5145FBAC9755F05040255FFD84175EF55002AAB0A2FFEAABA557BEA3EF057",
INIT_3C => X"82E974AAF7D57DF45552A3FF10AA8429F45A7D5EAF5FFBAEAAA10554155400AA",
INIT_3D => X"FF843FFE77C80825BC052ABFE10550415557085540000005156155FE90A8F5C0",
INIT_3E => X"00000000000000000000000000000000000005500020AAF7FBFFFEF04552ABFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(3),        -- Port A data input
DOA(0)   => data_read_a_hi_256(3),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(3),        -- Port B data input
DOB(0)   => data_read_b_hi_256(3),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_4_13 : RAMB16_S1_S1
generic map (
INIT_00 => X"A108400020612C80284210081034849800A00030300004833522C82D04A16002",
INIT_01 => X"2043998A1839284D1CA0650E1E504368403008418984014902030806A0D10200",
INIT_02 => X"C120042200000000044441CE01E80F00A49043118680008002000000026208E4",
INIT_03 => X"040001020019200020011209CC0164C060000000690111040144800042F5C403",
INIT_04 => X"7029AF0F81A00010CCA47700CC513CAC0D0B8E02010740E19754080108988021",
INIT_05 => X"02139405007133C0712244CD20F20105D583000020E9892201D304D42A9835E1",
INIT_06 => X"9190440300078002014405D9EE814C0284A883B6D7038AE079059B7800048092",
INIT_07 => X"000100AA0004408000000004840400008D200102503000782000C00C8025C000",
INIT_08 => X"00728A00408403220811991E02120C044058080004000001101121F220000260",
INIT_09 => X"811001E1185B38AD23C3707AD46440818F3CF80EC423CA7D01D123C80200816A",
INIT_0A => X"45810810A01B40216361056D6150F41200280001900439001FD8A00041400000",
INIT_0B => X"11FC88076266E800D605402962A820211500024808010512C40106D222223B14",
INIT_0C => X"0408804116040B02C02C500B0C02C100B0C02C100B0402C300B0401618058611",
INIT_0D => X"040200050200501301208482200D00D0A0408402C4282200A84800009B878680",
INIT_0E => X"00000020000100024AC88300300060090F0D830F00025400300204D018000804",
INIT_0F => X"8000000040000206A2000800000000000000950002E010000000080000588040",
INIT_10 => X"0000000000000808000554000200000000000100006D0020000000100000BB00",
INIT_11 => X"0000400000000000002000001A0002504001000000000000002280000D800800",
INIT_12 => X"0800000000000E2C802000000000408D801000000000408012440000200110A0",
INIT_13 => X"000000000004680003A0040000000010280003800800000000102800000B0000",
INIT_14 => X"000005C0002000000000000620000158000010000000000010A0000B00000200",
INIT_15 => X"C30146200400104002602600400000000294004000000004000000000010001A",
INIT_16 => X"0080200000008020000000802000000080080000004090014134DA101288C6DB",
INIT_17 => X"0802000000000401806010040180601004018060100000802000000080200000",
INIT_18 => X"8060180601004010040080200802000000000000802008020000000000008020",
INIT_19 => X"C0A28A063807E0500014063450404882846FFE000003FFC00000010040100401",
INIT_1A => X"AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA28A28A28A28A2934C8D0CCD145144",
INIT_1B => X"68341A0D068341A0D068341A0D068341A0D068351A8D46A351A8D46A351AAAAA",
INIT_1C => X"FFFFFFFFFFFFFFFC0000000000000000000000001FE32068341A0D068341A0D0",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"408102040810207FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"800AA00000000000000000000000000000000000000000000040810204081020",
INIT_28 => X"168B55557BEAB4500554200000557FE10FFFBEAA10007FD7410FFAA97555082A",
INIT_29 => X"55574105D2A800AA00043FEBA5D7FEAA00007BE8AAAAA843DF55FFAA955EFA2D",
INIT_2A => X"57BC00AAA2FFEAAAAAA8415555087BFFF55A2AA800BAFFAE9555508002AA0000",
INIT_2B => X"A2AA955EF005568A00087BE8BFFA2D17DE1000517FE10AAAAA8AAA002E975455",
INIT_2C => X"FAA8417410A2D140000F7FBC2010A2D157400AAAE974AAAAAA974BA08002AB55",
INIT_2D => X"EFA2AABDEAA087BEAAAAA2FBD54BA080002145552ABFEAA007FC21EF007FD75F",
INIT_2E => X"00055042AB45F7FFD741000042AA10AAAABFF5508003FF55F7D568A00552EA8B",
INIT_2F => X"5400F7A49057D0824850B8000000000000000000000000000000000000000000",
INIT_30 => X"3AF55F7A0925D7AADB6FB7D5D7FEAB7808554203A145178E00FFFBE8A101475D",
INIT_31 => X"A9557D080038AAA145157428492E8008200043FE925571EFA380871C7028A28E",
INIT_32 => X"AEA8A9200249056D4175C5092AAF5FDA38BE8E1557D1475FAF45BEAA800AAFFA",
INIT_33 => X"AA4954281C0E2FB55B6A0925D7085F6AA10087FEABD7AAD57AEBA08517DE00AA",
INIT_34 => X"007FC51C7007BD55D7BE80004AAFEDB42028EBFBC2028BED152438AAA092492A",
INIT_35 => X"AF7DF6AA00412EAABFFAA803DEBA0875EDA80BEF1C743840040017D5520B8EAA",
INIT_36 => X"0000000000000000000041002FB55FFF5D0438140E2FA38B6AEBFF6DBE84AAEB",
INIT_37 => X"A00FFFFEAA105D5155410FF84021EF0800154B20000000000000000000000000",
INIT_38 => X"DEBA0851574B2AAAEAAB55F78400145AAFFFFFEF5D7FEABFF0051400A25D5568",
INIT_39 => X"68B55F7AA800BAF7AA955EF00042AAA25555410BA082E8201000043FE005D517",
INIT_3A => X"568AA200557DE00AAAAAAA000804001FF005575408AA557FEB2FFAE975EF5551",
INIT_3B => X"D1550AAAA8002010F2AC154B25F2ABFF55F7800015F087FEAA00007FEAB55FAD",
INIT_3C => X"800021EF55042AAAA007FD5555087BD6145FAAC000A2A6FBC00BAAAFBC00BAF7",
INIT_3D => X"F7AEBDFF779A82AA43F7FBE8A00082EA8BFFAA843FEBA08517DE00F3F9574B30",
INIT_3E => X"000000000000000000000000000000000000008003FF55F7D5420BA5D2ABFEAA",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(4),        -- Port A data input
DOA(0)   => data_read_a_hi_256(4),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(4),        -- Port B data input
DOB(0)   => data_read_b_hi_256(4),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_5_13 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50DF4A0791B3FCB694379283C81FD996A091832102004A336A20E03C040C002",
INIT_01 => X"805FBDC69830A84D5C6A60000C34C26841280A00084000C8C212892EEAD53235",
INIT_02 => X"3B2026B578918E640A4F01CF8011FF0002080000082CA9998276DF7772C7C80D",
INIT_03 => X"37134108420D700084205702A4008A1D9100002171C0E0051554D93A11F5D140",
INIT_04 => X"8A41A0FC03A56DA000425A819410E3816C086198A388B702A8CA1210844A0C4C",
INIT_05 => X"B1808A062E8BC835F5E84532D708238A282F00A9291224800A2861490343082C",
INIT_06 => X"903FB8483A90581859050424100940825C6184401CDC451B860A6507160C4100",
INIT_07 => X"D26F068BCC96CDF8918E640E96D1A3469D6300E2FFEA27F8E4D23248130E259C",
INIT_08 => X"0BFA82E568442B2A082C0A7E3014250D49DA37A2420619000002AFF48D1222E5",
INIT_09 => X"3F005001E40969289429360416DCD1C46083030604B1CA20C03DF83B0A2C60A5",
INIT_0A => X"14613C71005A10492B888120288F480D58858449026145B3830F449449062B4F",
INIT_0B => X"11AC04934AC648BFD727C031E64170A137D5AA5C3E4B0F8A3C58C34C002290E3",
INIT_0C => X"CA29C6CC50384B6AC6AC86AB31AACA6AB39AAC86AB39AACA6AB3055643559C31",
INIT_0D => X"C673E33CF28F38603855401985228A0614BD30A0A2819852011E5AC2B87F9182",
INIT_0E => X"FF87C002F87A803E460B2516510CA594FF0044FFA4B08BAC4BB2CD0F09CF84E3",
INIT_0F => X"0DFF0F8005F0F5100DFFF5E15D06101C55EB29F1E00BE53FE1F000BE1E802F94",
INIT_10 => X"F12F0380231F17D78FC029FFF58D9A70380230F2FE0017C37FC3E0017C3D005F",
INIT_11 => X"FC7F023C0CA700125C0F8F7E43F1F001BFFE7C69E01804E1E7CCF8FC003FF5F1",
INIT_12 => X"023E00017C1FC1A4BFD82C3081C5BD27BFE30C3081C5BD00C02365D645CEEF5B",
INIT_13 => X"61E0042787F181E9C1EFD8CB8120C5AF41E9C18FD60F0C20666F41E9F009FFFD",
INIT_14 => X"7A7C077FFF404F80005F07F187A7D14BFFC96111C048278DEB074F9930FF9D80",
INIT_15 => X"C064014B8B652E2B3120C81284641D3E8DBF7D636FE860190700132C1F0EFB80",
INIT_16 => X"38CE1384E3384E338CE138CE1384E33C4E3ECE32E128882551349A1CBAA44103",
INIT_17 => X"84E3384E3384E3384E338CE138CE1384E3384E338CE138CE1384E3384E338CE1",
INIT_18 => X"CE138CE138CE138CE1384E3384E3384E3384E338CE138CE138CE138CE1384E33",
INIT_19 => X"F5E5BB4E7F7B9DB7FF3A1B6DB7E8410A8C000000000000000000384E3384E338",
INIT_1A => X"BEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEF9F7CFDFDDCF3CF3D",
INIT_1B => X"BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEFBEF",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000001711C7BBDDEEF77BBDDEEF77",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"FDFFF00000000000000000000000000000000000000000000080000000000000",
INIT_28 => X"FD7410FFAA97410082A800AAAAAE955450055421FFFFFBC0010AAD5574BA557F",
INIT_29 => X"7FD74000055574BA5D7FD7555A2D5575EF55517FF5500557FE10FFFBEAA10007",
INIT_2A => X"0002AABA5D2ABFFFFAA843DF55FFAA955EFA2D168B55557BEAB5500554200000",
INIT_2B => X"5D2A800AA00043FEBA5D7FEAA00007BC00AAAAAEBDF45A28428B45FFD168BFF0",
INIT_2C => X"5080028A00A2FFFDE00F7D57FEBAFF80174BAAAD1555EF555555555005557410",
INIT_2D => X"BA5D2E821FFA2D5554BA557BD75FFAA8415555087BFFF55A2AA800BAFFAE9555",
INIT_2E => X"00000517FE10AAAAA8AAA002E97545557BC00AAA2FFEAAAA082A97545F7D5420",
INIT_2F => X"7010BEDF524AA5571FDFEF000000000000000000000000000000000000000000",
INIT_30 => X"78E00EBFBE8A101475D5400F7A49043D0824850B8A2AE9756D145B401FFFFFFC",
INIT_31 => X"FEAB7D0855420BA1471D74380851524BA5571D757DB6D5525EF555178F6D1451",
INIT_32 => X"8A28B6DEBDF6DBEF1C0A28AAA5524BFFFFA28E3AF55F7A0925D7AADB6FB7D5D7",
INIT_33 => X"5555057D145152428492E8008200043FE925571EFA380871C7028B6AEBDF45B6",
INIT_34 => X"BEAA800AAFFAA9557D080038AAAA2FBF8E10EBD578EAAFF8415482BED1555EF5",
INIT_35 => X"81C209256DFFDF420BA552A821FFB6DF574A85575C55EFBE8E1557D1475FAF45",
INIT_36 => X"0000000000000000000008517DE00AAAEA8A9200249056D4175C50920875FDA3",
INIT_37 => X"5FF5D7BC21EFF7FBD7400F7FBC00BA55557DFF70000000000000000000000000",
INIT_38 => X"01FF5D5568BE7555568A00AAFFEAA105D5155410FF84020AA0800154B2AAAA97",
INIT_39 => X"00145AAFFFFFEF5D7FEABFF0051400A25551554BA0051400BA5551575EFF7D14",
INIT_3A => X"1574B2FFAABFF45FFAAAABFFAAFFFDFFF552EA8AAA55043DFF7AAAEAAB55F784",
INIT_3B => X"8002410FFD5575EF5555421E75555400BA082E8201000043FE005D517DEBA085",
INIT_3C => X"FAE975EF555168B55F7AA800BAF7AA955EF00002AAA2A2FBE8A00A2D16AAAAFF",
INIT_3D => X"0055554088A557FEB25D00021FFFFFFC00BA552A821EFFFFFD74BA5D51575F7F",
INIT_3E => X"000000000000000000000000000000000000000557DE00AAAAAAA000804001FF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(5),        -- Port A data input
DOA(0)   => data_read_a_hi_256(5),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(5),        -- Port B data input
DOB(0)   => data_read_b_hi_256(5),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_6_13 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10800B0061A01002840002C03002818000402322520070B313301C4389B2082",
INIT_01 => X"250041CA3839684D18A160000C52426841000000090800090210080008110200",
INIT_02 => X"0020042080010000044654C0000C008010000000001020900200200002620814",
INIT_03 => X"060881021088200021080200E4000A0891000020610111500104C00000F14400",
INIT_04 => X"0880000100000002000052288144004281C050400100280000C8100000080001",
INIT_05 => X"928080840001100A08009000280201000850E022401400002028214043410820",
INIT_06 => X"10100518090012122100C808049310002040000410A0001400000200120840D2",
INIT_07 => X"000100800004400001000000860408108C22000A502010074120044800040001",
INIT_08 => X"50000040D0C4E2088003FD01C01004044058082004000000000121F020408244",
INIT_09 => X"00BF17E9001205A5204911F814444080400100020000D200DFD16400C2A40AA0",
INIT_0A => X"04611C17849000022862A1596C8B5DF04834948900000100220C244840000880",
INIT_0B => X"03AD0413424E4044D665C070C22602291504400D084915020448114080201000",
INIT_0C => X"5E08864011088B22D22C008B0022C408B1022C208B0822C608B1111600458010",
INIT_0D => X"4251A12CD28A300429688001000800000020280204001000A00804309A002182",
INIT_0E => X"0000000280402400420800000000006200FC10002442042429324294014E8CA7",
INIT_0F => X"A40000000500800840000800000000000002280018001480000000A010100052",
INIT_10 => X"00000000000004C2003000010240000000000000680800290000000140202000",
INIT_11 => X"2000C0000000000000000442000001080001000000000000010C000280001804",
INIT_12 => X"08000000000801C300A010000000156000902000000015101200002800000000",
INIT_13 => X"000000000101800038002408000000094000386028040000000940000ED40000",
INIT_14 => X"0003B000002000000000020180002A24005010000000000023000060C7000A40",
INIT_15 => X"3F0280090321000040A410C28108000160008094000810040000000000002300",
INIT_16 => X"284A5284A728CA5284A528CA728CA52C4A5A0A32A300940101349A0408240818",
INIT_17 => X"9CA1294A329CA5284A728CA7284A5284A728CA5284A528CA728CA5284A728CA7",
INIT_18 => X"CA3294A129CA3294A129CA1294A329CA1294A3294A129CA3294A129CA3294A32",
INIT_19 => X"F5F78BCE7F8FF0F4FA955F7CF7F40A80145D55555556AAAAAAAAA94A329CA129",
INIT_1A => X"8E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E39B6CEDECDDF7DF7D",
INIT_1B => X"F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE38E3",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000001A1A33F9FCFE7F3F9FCFE7F3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"555FF00000000000000000000000000000000000000000000080000000000000",
INIT_28 => X"BC0010AAD5574BA557FFDFFF087BFDF45F7AA974AAAAAA97555F784174BAF7D5",
INIT_29 => X"515555508043FE00F7AA97555A2FBD7410AA8428AAAAAAE955450055421FFFFF",
INIT_2A => X"7D1575EFFFAA9555500557FE10FFFBEAA10007FD7410FFAA97400082A800AA08",
INIT_2B => X"0055574BA5D7FD7555A2D5575EF55517FF55A2AA97400552AAAB45082E80155F",
INIT_2C => X"500554200000003DE10FFD5401FFF7AAA8A10082EAAB45A2FFC2000007FD7400",
INIT_2D => X"10AA803FE105D516AABAFF843FFFFAA843DF55FFAA955EFA2D168B55557BEAB5",
INIT_2E => X"000AAAEBDF45A28428B45FFD168BFF00002AABA5D2ABFFFF087BD5545007BFDE",
INIT_2F => X"256DEB84104BAFFD1525FF000000000000000000000000000000000000000000",
INIT_30 => X"9756D145B401FFFFFFC7010BEDF524AA5571FDFEF1C7BFFF55FFA095482B6A49",
INIT_31 => X"4904380824850381C5B5057D1C003DE28F7A49057DAAF5D2428A2842AAAAA2AE",
INIT_32 => X"2AAFB451C2A8017DE3DF525FFFFA49756D145178E00EBFBE8A101475D5400F7A",
INIT_33 => X"2F1C50381471D74380851524BA5571D757DB6D5525EF555178F6DAAA49542841",
INIT_34 => X"AADB6FB7D5D7FEAB7D0855420BA1C0E3FE00E3DB471EFE3AAAAA00082EA8B6DA",
INIT_35 => X"F1C7BD057D1C71FFE10A28038E1049516AAB8FF8428FEFA28E3AF55F7A0925D7",
INIT_36 => X"00000000000000000000B6AEBDF45B68A28B6DEBDF6DBEF1C0A28AAA5524BFFF",
INIT_37 => X"F55F78017400F780001FFAA84000AAFFD1401E70000000000000000000000000",
INIT_38 => X"20BAAA8428AA2AAAA975FF5D7BC21EFF7FBD7400F7FBC00BA55557DFF7557BFD",
INIT_39 => X"EAA105D5155410FF84020AA0800154B2557FC01EF55043FEAAFF80021EFA2D14",
INIT_3A => X"568BE7AA80174AA082ABDF555D2A821EFAAFBC01FFF780155F7555568A00AAFF",
INIT_3B => X"AEA8A10082EA8BEFAAD5554B25551554BA0051400BA5551575EFF7D1401FF5D5",
INIT_3C => X"AAEAAB55F78400145AAFFFFFEF5D7FEABFF0051400A25D2EBFE10AAFFD55EFA2",
INIT_3D => X"552EA8AAA55043DFF7557BC01EF55557DE00AA842AA0000516AABAFF8428BE7A",
INIT_3E => X"0000000000000000000000000000000000000FFAABFF45FFAAAABFFAAFFFDFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(6),        -- Port A data input
DOA(0)   => data_read_a_hi_256(6),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(6),        -- Port B data input
DOB(0)   => data_read_b_hi_256(6),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_7_13 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10844B00482258A2842112C02450418800002300500030B313300C418992002",
INIT_01 => X"000009CA3839684D1CA0E0000E51424840000000080000080200080008510204",
INIT_02 => X"0120042086010000044600C00008000004100000000260900200000002402004",
INIT_03 => X"8628A10000082400000002408400080011000000610008000208C00000E14400",
INIT_04 => X"0911800100A000000000524084000040000050001140200100C8100000080102",
INIT_05 => X"0300812401011000000000002000114008008060441000000020024093000000",
INIT_06 => X"9190431C0D4010100000880804010010800000041080081000000200010424B2",
INIT_07 => X"000100AA0004408601000004860000008C02000A103010006928040800062481",
INIT_08 => X"84000048D484C20888000A0002120484C048007004000000000021F000000244",
INIT_09 => X"00A06009881201A520491004106C48A04040002400A15A208001650004001020",
INIT_0A => X"C99E1060201002044809C1040140A001004808810000459033189C0A400118A0",
INIT_0B => X"102000024040484050050041648A0041140C500B08821054C000264120000400",
INIT_0C => X"0404A083260E0832132011880462011880462051881462051881D31018C40620",
INIT_0D => X"0001000080001000813094801A8F80F00A600B52602801A88848011118003700",
INIT_0E => X"000003C007C002808228010410082042C000C000000004001002000400040002",
INIT_0F => X"A4000007800F80C840000800009864038A1200081C0014800000F001F0200052",
INIT_10 => X"00002C0E00E0E4004038000102400002C0E00E0D20100029000001E003E04000",
INIT_11 => X"2000C04031100E0403D0700300080908000100000661801E1900040380001804",
INIT_12 => X"0840878083E8003780A01043203A101780902043203A10082410082880000000",
INIT_13 => X"0601E0187900181035E0240806483248181035E0280410C8198818100DDD0000",
INIT_14 => X"0403774000201021E020FA006040376C00501022131210722060806D47000A40",
INIT_15 => X"00928A0002000110888600C032128201519480D40009902430160403E0E00506",
INIT_16 => X"01000000020080601802000000000405000A0020020081014134928820480010",
INIT_17 => X"0802018040000000006018020080200804010000000000806018020080000004",
INIT_18 => X"0000000001806008020000001006008020080001004008020080201004000020",
INIT_19 => X"0000000000000000000000000000400A004618618618C30C30C3000020180600",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000000B0840000000000000000000",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"1555500000000000000000000000000000000000000000000080000000000000",
INIT_28 => X"A97555F784174BAF7D5555FFF780155EFAAAEA8ABAAAFBFDE0055556AA005D04",
INIT_29 => X"55555EFAAFFFDFEFAAAAAAB455D556AA00FFAE95555087BFDF45F7AA974AAAAA",
INIT_2A => X"02EAAAAA082EA8A00AAAE955450055421FFFFFBC0010AAD5574BA557FFDFFF55",
INIT_2B => X"08043FE00F7AA97555A2FBD7410AA8428AAA557BFDFFF55003DFFFF7FBEAA000",
INIT_2C => X"0082A800AAF7AE975FFA28000010552EBDE00007BEAAAAA2D140000085155555",
INIT_2D => X"45087FEAB455D516AB55557BD55FF00557FE10FFFBEAA10007FD7410FFAA9740",
INIT_2E => X"000A2AA97400552AAAB45082E80155F7D1575EFFFAA955555D51574AAAAFFD55",
INIT_2F => X"AE105D556AA10410E17555000000000000000000000000000000000000000000",
INIT_30 => X"FFF55FFA095482B6A49256DEB84104BAFFD1525FFFF8E175C7A2AAAAA82A2F1F",
INIT_31 => X"F524AA5571FDFEF415B575D7AAF1FFFD7AAAAAFB7D495F6AA10E3AE905551C7B",
INIT_32 => X"003AFEFEBFBEAA001C2EA8A821C2EAAA00A2AE9756D145B401FFFFFFC7010BED",
INIT_33 => X"EDB470101C5B5057D1C003DE28F7A49057DAAF5D2428A2842AAAA497BFAFFF49",
INIT_34 => X"1475D5400F7A490438082485038F7A4905C7A28A070384120BDE100075EAA82B",
INIT_35 => X"D495150492BEF1D2555087BE8B7D555F6AB57417BC05D7145178E00EBFBE8A10",
INIT_36 => X"00000000000000000000AAA495428412AAFB451C2A8017DE3DF525FFFFA49756",
INIT_37 => X"555A2AEA8A10AAD568A00555168A10002E9754D0000000000000000000000000",
INIT_38 => X"8A10AAAE8215D557BFDF55F78017400F780001FFAA84000AAFFD1401E7FFAA97",
INIT_39 => X"C21EFF7FBD7400F7FBC00BA55557DFF7007BD5555AAD57DF55AAAEBDFEF007BE",
INIT_3A => X"428AA2007FE8BFF080028BFFAAFFEAA105D2EAAA005D2AAAA18AAAA975FF5D7B",
INIT_3B => X"043DE0000516AA10F7FBD7408557FC01EF55043FEAAFF80021EFA2D1420BAAA8",
INIT_3C => X"55568A00AAFFEAA105D5155410FF84020AA0800154B2FF8402145A2AA954AA00",
INIT_3D => X"AAFBC01FFF780155F7005140000FFD140145007FE8BEF557BEAB55087FC215D5",
INIT_3E => X"0000000000000000000000000000000000000AA80174AA082ABDF555D2A821EF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(7),        -- Port A data input
DOA(0)   => data_read_a_hi_256(7),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(7),        -- Port B data input
DOB(0)   => data_read_b_hi_256(7),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_8_13 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00000648E2840112C00000418000002700500030B3132000400812082",
INIT_01 => X"100008480009004C04A100000252024840000000180800080200010040110204",
INIT_02 => X"0020042000490000004600804008000005100000000024900200000002400004",
INIT_03 => X"0A0C33400008082400000080A4004B0891000020610112000040C00000E5C000",
INIT_04 => X"18800001000000000000512080000040800150400824280110C8100000120200",
INIT_05 => X"908084A10100100200004080280008240810802206940000012C214451610800",
INIT_06 => X"81B000080860109021400008040000202048020414A0021400040200322824C1",
INIT_07 => X"000000080004408049000004860000008402001A50208000630C040800062483",
INIT_08 => X"440000428644212280800A00021004044048002124000000000021F000000244",
INIT_09 => X"00004009001001010008100414644410400102228000D20080114502006409A2",
INIT_0A => X"000051312000042200294429148A4801C80C8C81000045907118040340020832",
INIT_0B => X"4020000240404140004D0544C4AA0001150410090302500011C813428A000400",
INIT_0C => X"46501090008820240240409000240009000240009000240009000120204808A5",
INIT_0D => X"42D1A168D09A301468402480004780F00140080860280004085904309A002196",
INIT_0E => X"00783FC00044340242280000000000020000C0000442106419120004034685A3",
INIT_0F => X"8000F07F800088A80000081EA2F9EC0000064004081010001E0FF00011104040",
INIT_10 => X"0ED0FC7E00000422201080000202658FC7E0000021882020003C1FE000222080",
INIT_11 => X"018059C3F350FE0C00000002A0040500000103961FE780000110010090000800",
INIT_12 => X"FD41FF80000830200021C1CF600012200010D1CF600012121600100810000004",
INIT_13 => X"9E1FE000010A1802100004343ED8000898021000087073D80008980200800002",
INIT_14 => X"0080200000BEB07FE00002086008020000209AEE3F300000246020200000620B",
INIT_15 => X"0088881903210000440610C8000A808040000208901786E4F0FE0C0000000166",
INIT_16 => X"685A1685A769DA368DA368DA769DA36CDA121A11A141800011309284002C0810",
INIT_17 => X"95A5685A1685A5695A368DA368DA769DA368DA368DA7695A1685A1685A5695A1",
INIT_18 => X"5A1695A568DA368DA369DA768DA1685A1695A5685A168DA369DA768DA368DA16",
INIT_19 => X"A4028A0A543EBC57A10A1E75D64108080468618618630C30C30C69DA5685A168",
INIT_1A => X"9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7BF3CCD8DF5B2DB2C",
INIT_1B => X"F87D3E1F4F87D3E1F4F87D3E1F4F87D3E1F4F87C3E1F0F87C3E1F0F87C3E79E7",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000006A6D4F87D3E1F4F87D3E1F4",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"155FF00000000000000000000000000000000000000000000080000000000000",
INIT_28 => X"BFDE0055556AA005D0415555080000000087BEAA10F7803DE00FFAEBFFFF0800",
INIT_29 => X"2AA8AAA557FC0010F780154105D7FC2145005155555F780155EFAAAEA8ABAAAF",
INIT_2A => X"7FFFFF55AA80155FF087BFDF45F7AA974AAAAAA97555F784174BAF7D5555FF55",
INIT_2B => X"AAFFFDFEFAAAAAAB455D556AA00FFAE95555AAFFE8A00552EBFE00F7D17FF45F",
INIT_2C => X"A557FFDFFF5504000AAAAAAA8B55F7D140010552E821EFAAAABDF555555555EF",
INIT_2D => X"55AA8028A00A2D57FF45557BE8A00AAAE955450055421FFFFFBC0010AAD5574B",
INIT_2E => X"000557BFDFFF55003DFFFF7FBEAA00002EAAAAA082EA8A00002AA8A10F784021",
INIT_2F => X"FE10F7AEBAFFF080A175D7000000000000000000000000000000000000000000",
INIT_30 => X"175C7A2AAAAA82A2F1FAE105D556AA10410E17555080E000280071E8A00EB8E3",
INIT_31 => X"4104BAFFD1525FF492EA8AAA5571C2000FF8A17400557FC015514555757DFF8E",
INIT_32 => X"2ABDE10EBDF7AF6DE3FFF8F7DB68A105D71C7BFFF55FFA095482B6A49256DEB8",
INIT_33 => X"AA0BDF6D415B575D7AAF1FFFD7AAAAAFB7D495F6AA10E3AE90555A2FBE8A3849",
INIT_34 => X"FFFFC7010BEDF524AA5571FDFEF550E00082B6A0AFB55F7D1420104124821D7A",
INIT_35 => X"01C2EA8A00F7800017DA2842FA00B6D578F6D557FFDA00A2AE9756D145B401FF",
INIT_36 => X"00000000000000000000497BFAFFF49003AFEFEBFBEAA001C2EA8A821C2EAAA0",
INIT_37 => X"0BA08556AA00AAAABFE00F7AEAABEF082E955450000000000000000000000000",
INIT_38 => X"21555D51575EFFFAA97555A2AEA8A10AAD568A00555168A10002E9754D082E82",
INIT_39 => X"17400F780001FFAA84000AAFFD1401E7082EAAABA5D5140010F7AE974105D7BC",
INIT_3A => X"E8215DA2FFE8ABA082ABFE00AAFBEABFFAAFBEABFFF7AA80145557BFDF55F780",
INIT_3B => X"D540000000402145AA843FFFF007BD5555AAD57DF55AAAEBDFEF007BE8A10AAA",
INIT_3C => X"AAA975FF5D7BC21EFF7FBD7400F7FBC00BA55557DFF75D2E82010F7843DF45FF",
INIT_3D => X"5D2EAAA005D2AAAA185D2AAAA10F780021FFA2803DE10FFD16ABFF5D7BFDE10A",
INIT_3E => X"0000000000000000000000000000000000000007FE8BFF080028BFFAAFFEAA10",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(8),        -- Port A data input
DOA(0)   => data_read_a_hi_256(8),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(8),        -- Port B data input
DOB(0)   => data_read_b_hi_256(8),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_9_13 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00018248A2840112C00002C18000002300500030B3132000400812006",
INIT_01 => X"400008000000004C0020000000100248413C0A61590001D90213C10008110204",
INIT_02 => X"01A0042080010000054600C04008000004100000001020900200200002420804",
INIT_03 => X"024003400008012400000010E4004B0891000020610310000144C00000F5C000",
INIT_04 => X"1801800100E000000000510084000040010050020810200000C8900000320200",
INIT_05 => X"918004311104100000000000200008100800002000100000002C234415610820",
INIT_06 => X"81B00008080010100000980804000008800042041080001000100200322C2481",
INIT_07 => X"0000811800044080010000058600000086020002502080006000040800062C80",
INIT_08 => X"0000004001D4618008800A00061004044048002004000000000061F000000244",
INIT_09 => X"000040090802009420409004104444084001022400214A2080014400026401A2",
INIT_0A => X"04000071200000A003CA294140200800C80C8C8100004590111C040040120800",
INIT_0B => X"12210002404848502847040164880021150400080222000200C8034200000000",
INIT_0C => X"4610088010080421021040841021000841021000841021000841010800420820",
INIT_0D => X"42D0A16C529A321068500484000500D10042080040284000084900001A002196",
INIT_0E => X"00000002804000004228010410082002C000C0002400046419120410034285A1",
INIT_0F => X"A00000000500800800000800000000000002290008001080000000A010100042",
INIT_10 => X"00000000000004C2001000000240000000000000680800280000000140202000",
INIT_11 => X"0000C0000000000000000442020001000001000000000000010C800080000804",
INIT_12 => X"08000000000801A7802010000000152780102000000015000600000800000000",
INIT_13 => X"000000000101900011E0240000000009500011E0280000000009500004DD0000",
INIT_14 => X"000137400020000000000201C000136C00101000000000002340002947000240",
INIT_15 => X"0080881901210000000600C280028000419480D4000010040000000000002304",
INIT_16 => X"68DA368DA1685A1685A1685A1685A16C5A121A13A141950051309284A82C0010",
INIT_17 => X"85A1685A1685A1685A368DA368DA368DA368DA368DA368DA368DA368DA368DA3",
INIT_18 => X"5A1685A168DA368DA368DA368DA368DA368DA368DA3685A1685A1685A1685A16",
INIT_19 => X"0157344CCCF48DE68A895C38E2540A8010100000000000000000685A1685A168",
INIT_1A => X"14514514514514514514514514514514514D34D34D34D34D28E1004039248209",
INIT_1B => X"D268341A4D268341A0D069349A0D069349A0D068341A0D068341A0D068345145",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000014D490D069349A0D068341A4",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"EAABA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"03DE00FFAEBFFFF0800155FFAAFBE8B45002A974AAAA803DFFFAA843DF45FFFF",
INIT_29 => X"7BFDE00A2FBD7400F7FBFDFFFA2AEBDE00AAFBEAABA080000000087BEAA10F78",
INIT_2A => X"055401FFF7AEAAA10F780155EFAAAEA8ABAAAFBFDE0055556AA005D041555508",
INIT_2B => X"557FC0010F780154105D7FC2145005155555557BE8BEF007FFDEAAAAD1555EF0",
INIT_2C => X"AF7D5555FFF780154AA5D2AA8A10F7AA974AA082E80010A2AAAAA10552AA8AAA",
INIT_2D => X"BAF7D17FEBAA2AEBDF45002EAAABA087BFDF45F7AA974AAAAAA97555F784174B",
INIT_2E => X"000AAFFE8A00552EBFE00F7D17FF45F7FFFFF55AA80155FF080400145FFFBEAA",
INIT_2F => X"8FC7BE8A3DF7DF7F5E8A92000000000000000000000000000000000000000000",
INIT_30 => X"000280071E8A00EB8E3FE10F7AEBAFFF080A175D7BEF1E8B6D002090482B68E3",
INIT_31 => X"56AA10410E175550871FFE00A2FBD0400FFF5FDFC7B6A0BDE38B6F5E8A92080E",
INIT_32 => X"7BFAE82A2DB555C71C5B451D7FFAAA8A38FF8E175C7A2AAAAA82A2F1FAE105D5",
INIT_33 => X"2AEADA38492EA8AAA5571C2000FF8A17400557FC015514555757D5D71E8BEF14",
INIT_34 => X"B6A49256DEB84104BAFFD1525FFFF84174BA5D20AAA00E3AA904BA142A87010A",
INIT_35 => X"7000400155FFFBEDA82FFD57DEBAAAA0BFF7D0024ADA921C7BFFF55FFA095482",
INIT_36 => X"00000000000000000000A2FBE8A38492ABDE10EBDF7AF6DE3FFF8F7DB68A105D",
INIT_37 => X"BEF080402000F7AAA8B55FFAABDFEFF7D16AA000000000000000000000000000",
INIT_38 => X"FEAAFFD16AA00082E820BA08556AA00AAAABFE00F7AEAABEF082E95545F7D568",
INIT_39 => X"A8A10AAD568A00555168A10002E9754D00517DE00A2FFC2000F7D17FF55FF803",
INIT_3A => X"1575EF555568BEF5D7FE8A10AAFFD55555D7FD5555FFAAA8AAAFFAA97555A2AE",
INIT_3B => X"AE800AA552A97400A2AEBDEAA082EAAABA5D5140010F7AE974105D7BC21555D5",
INIT_3C => X"57BFDF55F78017400F780001FFAA84000AAFFD1401E7FF80174AA5D0028A00AA",
INIT_3D => X"AAFBEABFFF7AA80145080002145F7FBFFE00FFD17FEAAA2803DFEF08043FE005",
INIT_3E => X"0000000000000000000000000000000000000A2FFE8ABA082ABFE00AAFBEABFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(9),        -- Port A data input
DOA(0)   => data_read_a_hi_256(9),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(9),        -- Port B data input
DOB(0)   => data_read_b_hi_256(9),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_10_13 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00018248A2840112C00002C18000202300500030B3132000400992006",
INIT_01 => X"254008000000004C002000000010026840000000080000080200010008110204",
INIT_02 => X"0020042000010000004455800008000004100000000000900200000002400004",
INIT_03 => X"020001021089000021081000C400090011000000610001540104C00000F14400",
INIT_04 => X"0811800101A00002000050088554004200C840000000200080C8100000000001",
INIT_05 => X"030080001000100800009400200000000840E020201000000024024001200020",
INIT_06 => X"81B00008080012120004CC080492500280208004148000100000020020042493",
INIT_07 => X"0000000800044080010000048404081085020002502000006000040800062480",
INIT_08 => X"100202400084410808000A00021004044048000004000000000021F020408264",
INIT_09 => X"010040090002008420401004144440004040022484214A2080110108C2C00320",
INIT_0A => X"04004166A48A0001080000000000080080181881000045901118044040020800",
INIT_0B => X"1201000200484910000F0105602622291404020902005002018002400A022000",
INIT_0C => X"0440001011808020120004801120044800120004801120044800110002400884",
INIT_0D => X"008000440210100041308480800F82F00040180260A808008848000018002104",
INIT_0E => X"000000028040000002280104100820020000400020000440100204100A000100",
INIT_0F => X"040000000500800800000000000000000002280008000400000000A010100010",
INIT_10 => X"00000000000004C2001000010000000000000000680800010000000140202000",
INIT_11 => X"200000000000000000000442000001000000000000000000010C000080001000",
INIT_12 => X"00000000000801C0008000000000154000800000000015000410000800000000",
INIT_13 => X"0000000001019800180000080000000958001800000400000009580002800000",
INIT_14 => X"0000A0000000000000000201E0000A0000400000000000002360002080000800",
INIT_15 => X"0080881000000000000600C28102800060000000000800000000000000002306",
INIT_16 => X"401004010040100401004010040100441020D0030008840051309A90BA884010",
INIT_17 => X"0902409024090240900401004010040100401004010040100401004010040100",
INIT_18 => X"1004010040902409024090240902409024090240902409024090240902409024",
INIT_19 => X"F546890A940FE0D3971243555205428290100000000000000000401004010040",
INIT_1A => X"8A28A28A28A28A28A28A28A28A28A28A28A28A28A28A28A29554199854514514",
INIT_1B => X"2B95CAE532994CA6532995CAE572B94CA6532994CA6532994CA6532994CA28A2",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000002718E72B94CA6532994CA657",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"FDE1000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"03DFFFAA843DF45FFFFEAABA007FC2155F7D155545AA80001EFAAFBEAB45557F",
INIT_29 => X"042AB55FFD168B55AA8000010FFFBE8BFFF78402155AAFBE8B45002A974AAAA8",
INIT_2A => X"AD16AABA002ABDE10080000000087BEAA10F7803DE00FFAEBFFFF0800155FF00",
INIT_2B => X"A2FBD7400F7FBFDFFFA2AEBDE00AAFBEAABAA2FFD741055003DFEFF7AA801FFA",
INIT_2C => X"05D0415555007FD74105555555EFF7FBC0145F78028A00A2D142155087BFDE00",
INIT_2D => X"55AAD168ABA002A975FFF7AEBDEBAF780155EFAAAEA8ABAAAFBFDE0055556AA0",
INIT_2E => X"000557BE8BEF007FFDEAAAAD1555EF0055401FFF7AEAAA105D042ABFF5D556AB",
INIT_2F => X"71D7AAFBEFB455D71F8E00000000000000000000000000000000000000000000",
INIT_30 => X"E8B6D002090482B68E38FC7BE8A3DF7DF7F5E8A92007BC217DEBDB55555AA8E0",
INIT_31 => X"EBAFFF080A175D700042AB7DEBDB6DB55BE8E05000EBFFE8BC7E38E07145BEF1",
INIT_32 => X"0A3DFD7F7A4821D7A2D16FA82142EB8E00080E000280071E8A00EB8E3FE10F7A",
INIT_33 => X"ED1421450871FFE00A2FBD0400FFF5FDFC7B6A0BDE38B6F5E8A92B6FBD541049",
INIT_34 => X"A2F1FAE105D556AA10410E175550071D54104951555D7EBF5C5155E3842AA00B",
INIT_35 => X"8410E2ABD749516FB55BED16FA820820955EFE3AEBDEAAFF8E175C7A2AAAAA82",
INIT_36 => X"000000000000000000005D71E8BEF147BFAE82A2DB555C71C5B451D7FFAAA8A3",
INIT_37 => X"1EFA2FFD7545AAAE97555A2FBFDF455D556AA000000000000000000000000000",
INIT_38 => X"8B45AAAA95545F7D568BEF080402000F7AAA8B55FFAABDFEFF7D16AA00087FC0",
INIT_39 => X"6AA00AAAABFE00F7AEAABEF082E9554500042ABFFA2FFFFF45F7AE97400AAFFE",
INIT_3A => X"16AA00FFFBD5400082EBFF45F78400155A2D57FE00552EA8A00082E820BA0855",
INIT_3B => X"D557555A2802AA10FFD54214500517DE00A2FFC2000F7D17FF55FF803FEAAFFD",
INIT_3C => X"FAA97555A2AEA8A10AAD568A00555168A10002E9754D085155410085557555AA",
INIT_3D => X"5D7FD5555FFAAA8AAA002AAAB4508557DF55F7D17FE000804155FFAAAABDEAAF",
INIT_3E => X"0000000000000000000000000000000000000555568BEF5D7FE8A10AAFFD5555",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(10),        -- Port A data input
DOA(0)   => data_read_a_hi_256(10),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(10),        -- Port B data input
DOB(0)   => data_read_b_hi_256(10),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_11_13 : RAMB16_S1_S1
generic map (
INIT_00 => X"A101C4B05A0034CA2840712C2D001419000002300500030B31B20084EC992002",
INIT_01 => X"90000986B83028491800E0000C26426040000000080000088200080802512224",
INIT_02 => X"1A2004205E010640024D00800008000004100000040EC090820018003241A00C",
INIT_03 => X"28639100000C5C00000045C08400C8001100000061806A001618C03001E54400",
INIT_04 => X"1A800001000009A0804059A190000040400040008058220008C8100000120D4E",
INIT_05 => X"02000E81080250010000002022000058080400000E1200000020004401000004",
INIT_06 => X"819435143F20101010001008040800B8100102041088011100022200000024B2",
INIT_07 => X"90640D280884453E01064002944180008402001295BA100022E4340800062D82",
INIT_08 => X"400000093204802200280A0012160585C1D808D004000000000323F40C102244",
INIT_09 => X"380040098010001100009204107C5950400000220080C200800900020C006827",
INIT_0A => X"80007100004016EA080801010000080D00200081000045B0511D289940103399",
INIT_0B => X"002000024040410A000D0104408810C115D9C008050042400100D04E88000002",
INIT_0C => X"00655010009264201200C7B421ED0C7B421ED0C7B431ED087B43176843DA1085",
INIT_0D => X"0401020080400A10012494881A4F80F209500BB2602881A488485C1318002000",
INIT_0E => X"6619A540124814800228010410082022C00040002020090020220C9600040802",
INIT_0F => X"ACCC334A802491600C587949B6D0141B4CC600D5761B1599865A500490B86A56",
INIT_10 => X"BAC845542056A61686EC81E3A6CB68AA2C622C9A251C352B330CB4A0092170D8",
INIT_11 => X"BCCAD0B5A81536080CC6B21A21B1FC09CB0F1076D4A200B2AD4068F4101639B5",
INIT_12 => X"4D2CC281E31AA0103AB8D5514066380804B268A2E060901204112566F10AC418",
INIT_13 => X"D551443C47281002540B2C9AAAA8662A1152B202AE3554403028115AA88201A1",
INIT_14 => X"548A20A0492A2724A0621620402A020141F172FB182A32AB6845AB6200251BC9",
INIT_15 => X"00C00A000200074044E6801832728080D00A380B753952C4877E0104DDE4D124",
INIT_16 => X"0080200802008020080200802008020480080022020081010124988800400010",
INIT_17 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_18 => X"0000000000802008020080200802008020080200802008020080200802008020",
INIT_19 => X"55062608804180C0B10A42104201400204000000000000000000000000000000",
INIT_1A => X"00000000000000000000000000000000000820820820820801C4149470000000",
INIT_1B => X"0000000000000000040200000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000007E0F0000000000000100800",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"000AA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0001EFAAFBEAB45557FFDE10082ABDF5508557DF45002ABDFFFF7803DE10AA80",
INIT_29 => X"AEBFF45FFAEBFEAA002A801FFF7FFE8A10A28000000007FC2155F7D155545AA8",
INIT_2A => X"2AABFE10082ABFFEFAAFBE8B45002A974AAAA803DFFFAA843DF45FFFFEAABAA2",
INIT_2B => X"FFD168B55AA8000010FFFBE8BFFF78402155AAD155555A28428BFF002ABDE00A",
INIT_2C => X"F0800155FF00557FF45557FC2010002A80010A2842AAAA007BFFF4500042AB55",
INIT_2D => X"FF5D00154BAF7FBE8BEFFFD540000080000000087BEAA10F7803DE00FFAEBFFF",
INIT_2E => X"000A2FFD741055003DFEFF7AA801FFAAD16AABA002ABDE10A2D168A10A284021",
INIT_2F => X"DFC7F78E3FE28B684070AA000000000000000000000000000000000000000000",
INIT_30 => X"C217DEBDB55555AA8E071D7AAFBEFB455D71F8E00002EBDF6D005B78F7D142AB",
INIT_31 => X"A3DF7DF7F5E8A92BEAEBFF7DEBA0BDEAA1C2A801C7E3FFEFA10B68407038007B",
INIT_32 => X"8A28BFF082ABAE10B6AAB8E280820B8FEFBEF1E8B6D002090482B68E38FC7BE8",
INIT_33 => X"07FF8F7D00042AB7DEBDB6DB55BE8E05000EBFFE8BC7E38E07145B6D15756DA2",
INIT_34 => X"EB8E3FE10F7AEBAFFF080A175D708517DF7D497BC5028142A87000A28A2AA920",
INIT_35 => X"0B6DB6AA28A280001FF5D0A10482FFFFEFBC7E3DF42028080E000280071E8A00",
INIT_36 => X"00000000000000000000B6FBD5410490A3DFD7F7A4821D7A2D16FA82142EB8E0",
INIT_37 => X"FEF007BE8BFF5D2ABDF55F7AABDEAAF784154BA0000000000000000000000000",
INIT_38 => X"DE00FF84154BA087FC01EFA2FFD7545AAAE97555A2FBFDF455D556AA00082EBF",
INIT_39 => X"02000F7AAA8B55FFAABDFEFF7D16AA00FFAEBFFEFAA803DEBA5D2E82155A2FBF",
INIT_3A => X"A95545F7D5555FFAAAAA8BFF002AAAA00FFAAA8AAA080028BFFF7D568BEF0804",
INIT_3B => X"2E95400A2AEA8A00007FEABFF00042ABFFA2FFFFF45F7AE97400AAFFE8B45AAA",
INIT_3C => X"82E820BA08556AA00AAAABFE00F7AEAABEF082E9554508557DFFF007BD54BA5D",
INIT_3D => X"A2D57FE00552EA8A00FFFFE8AAAAA80001FF5D2E82000F7FFFFF45AAFFC20BA0",
INIT_3E => X"0000000000000000000000000000000000000FFFBD5400082EBFF45F78400155",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(11),        -- Port A data input
DOA(0)   => data_read_a_hi_256(11),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(11),        -- Port B data input
DOB(0)   => data_read_b_hi_256(11),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_12_13 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50080B01BC002006940202C0DE041196A83183000000023322287E0FC000006",
INIT_01 => X"75400D849830C84C5823E0000C17424840000000080000088200002802153231",
INIT_02 => X"18A026B43ED180040147558040090000061800000C06ED9802768F4472C52005",
INIT_03 => X"2A67E34A528D0524A52850528400C8001100000171C02B550618C91A10E55440",
INIT_04 => X"1BC0000100056C8280825DE98154004300C840800850240080CA921084520A07",
INIT_05 => X"02000F832000500C0000941024000852084060202E100001002000448100000C",
INIT_06 => X"819A1D1C3FE01A1A40045408049A50BA4020C6041090001200006200000000F2",
INIT_07 => X"C26A0719CC96CC6ED18A64019695A854870300FA3968B20068FC06080106249F",
INIT_08 => X"D002024B3E040800008C0A002610240D494A06F3460409000000E3F0AD5282E5",
INIT_09 => X"27A06009200040000400120412445D78400001000410420080218029CC807A27",
INIT_0A => X"18000006848A026F000000000000080000F010C100204593F11A6CDF48003BF8",
INIT_0B => X"000000820040402B28050400400432C9349DF21A31A00ACC0000F04F80020001",
INIT_0C => X"00357804611AE45D05D0833430CD0833420CD0C33420CD0833430668619A1000",
INIT_0D => X"0000000000000A74812DF00E87E80A079F9F90FA0280E87E800C7FF3B8002000",
INIT_0E => X"3B6B0E404D26160682082002000401EA0000C40000800A006002818808000000",
INIT_0F => X"A476D61C809A4DA84272592D6246FC1B17B541F97E1B348EDA93900B2B286C56",
INIT_10 => X"30C669E622DBC325CFD881A962454CFBE5403AB99594362B1DB52720165650D9",
INIT_11 => X"F8D2D39A3745261E4A95A110A3F855000E4B1D32BAB504BB7490FCFF912A3834",
INIT_12 => X"B90E9B018C7530200AB8F8BF41F9A22006B37DC8E1F9A21A70116D4C5080651C",
INIT_13 => X"118780319CCA08AB1001ACDF34B8F1C688AB1002AE3F7B807B6289F368828C4C",
INIT_14 => X"2AF020233376A5ECC016B1A827CDA21160F051DE610A34C50427E6E220323E4A",
INIT_15 => X"0077020000000439FDC05C5806781FAB46095A0B5199B0AC55521524F1864022",
INIT_16 => X"000000000000000000000000000000000026C000002884000130921092804010",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"8020080200000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0051B946088881360A95090CB054420290100000000000000000008020080200",
INIT_1A => X"041041041041041041041041041041041049249249249249200100002D451451",
INIT_1B => X"92C964B2592C964B2592C964B2592C964B2592C86432190C86432190C8641041",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000003800F592C964B2592C964B25",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"7DE1000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"ABDFFFF7803DE10AA80000AAAA843FE0008557DFFF0800020105D557FEAA0055",
INIT_29 => X"D5420000051555FFA2AA8200000557DFFFF7AA80000082ABDF5508557DF45002",
INIT_2A => X"82AA8AAAAAFFC00BA007FC2155F7D155545AA80001EFAAFBEAB45557FFDE10AA",
INIT_2B => X"FFAEBFEAA002A801FFF7FFE8A10A28000000A2D155410F7FFFFEBA08003FE000",
INIT_2C => X"5FFFFEAABA000028A105D2ABFE10A2AABFE1055516ABEF5D517DEAAA2AEBFF45",
INIT_2D => X"55002A820AA08557DFFFF7AA82155AAFBE8B45002A974AAAA803DFFFAA843DF4",
INIT_2E => X"000AAD155555A28428BFF002ABDE00A2AABFE10082ABFFEF0855420000004175",
INIT_2F => X"5010495B7AE921C517DE10000000000000000000000000000000000000000000",
INIT_30 => X"BDF6D005B78F7D142ABDFC7F78E3FE28B684070AABE803AE38145B78FD700000",
INIT_31 => X"BEFB455D71F8E00BED547038145B505FFB6A487000005F7AFD7F7A482038002E",
INIT_32 => X"F1FDE821C003FE001C2EAAAAAB6F5C2082007BC217DEBDB55555AA8E071D7AAF",
INIT_33 => X"D517DEAABEAEBFF7DEBA0BDEAA1C2A801C7E3FFEFA10B68407038B6D550428FF",
INIT_34 => X"B68E38FC7BE8A3DF7DF7F5E8A9200002FA285D20BDE28A2A4B8E10555B68BEF5",
INIT_35 => X"F085F47038140010555142082082005F7DFD7F7A482155BEF1E8B6D002090482",
INIT_36 => X"00000000000000000000B6D15756DA28A28BFF082ABAE10B6AAB8E280820B8FE",
INIT_37 => X"ABA5D7FEAB45080015410007FEAA0055517DE000000000000000000000000000",
INIT_38 => X"AB45F780020BA082EBFFEF007BE8BFF5D2ABDF55F7AABDEAAF784154BAF7802A",
INIT_39 => X"D7545AAAE97555A2FBFDF455D556AA00F7D1554BA5D7BC01FFFF8015410007FE",
INIT_3A => X"4154BAF7D1400BAFFD57FE005D043FE10552EAAAAAFFD140000087FC01EFA2FF",
INIT_3B => X"8428A105D7FEABEF55557DEBAFFAEBFFEFAA803DEBA5D2E82155A2FBFDE00FF8",
INIT_3C => X"7D568BEF080402000F7AAA8B55FFAABDFEFF7D16AA0008003FEBA55003DEBAA2",
INIT_3D => X"FFAAA8AAA080028BFF087BD54AA550402145550000010087FFFF45F78402145F",
INIT_3E => X"0000000000000000000000000000000000000F7D5555FFAAAAA8BFF002AAAA00",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(12),        -- Port A data input
DOA(0)   => data_read_a_hi_256(12),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(12),        -- Port B data input
DOB(0)   => data_read_b_hi_256(12),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_13_13 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10154A0441836CA2840512822007C18000E02700500030B31B300040081A042",
INIT_01 => X"00000804A000C04800020000000002404001000008220008A200100802110204",
INIT_02 => X"02200430000104000A4700804008000004100000000420918204D3033240400D",
INIT_03 => X"AA4003400008592400000590C40009141100000C6180C0000000C00001E14000",
INIT_04 => X"0800000102400120088054019000004160004190BAA0270000C8100000600206",
INIT_05 => X"21000012040610050040000227003AA0082400E94C1200000824424005220020",
INIT_06 => X"81963B180C001010580000080400000058000004109C00138000020024142581",
INIT_07 => X"002C8008000441600106400A9600010494020002B8AAA000EF003408000E2580",
INIT_08 => X"000000E48194408000A00A001210040441C80320040210000002ABF004102244",
INIT_09 => X"2A004009640040100400940412D4C4004000022000104200802D983000480120",
INIT_0A => X"8000202020401480000000000000080C90090881000145B0111A14004015080D",
INIT_0B => X"00000002004040AA08050400404040C11444000805200A402090024000008002",
INIT_0C => X"8410000A00280020020040800020040800020000801020000800010020400000",
INIT_0D => X"84A14250A055100050100490000500D00040080040290000084E4000B800610C",
INIT_0E => X"DCD13042BEDA36820228000000000000C000400081A08BC812A2092B02850942",
INIT_0F => X"89B9A260857DB400431969CA985D480949D32804A40AB137341C10B7D6A02EC0",
INIT_10 => X"E6ACA678001CE7D0296C213A460CA4271CA2168AEC1017606E6838216FAD4055",
INIT_11 => X"84AD4961C281B20213073C5FC0058008632D30D522CE80239DCC01AB013A4D20",
INIT_12 => X"2E6B13804A4B01D83461299900F6BD583A519104A0EEBD1A141010B2A4C8E116",
INIT_13 => X"89E5E40913419151EE0E94641828F72B5151EE0D184B321037AF5158BB02D085",
INIT_14 => X"562EC0B42162D68EE0073AE1C562EC13D521921A4170300B2B458B56B01C2280",
INIT_15 => X"00888A120240034000E6DC8285028014B82372011FC1E4F5E0A00929684EAF84",
INIT_16 => X"50942509425094250942509425094254940A1421420082020120908800480030",
INIT_17 => X"0942509425094250942509425094250942509425094250942509425094250942",
INIT_18 => X"9425094250942509425094250942509425094250942509425094250942509425",
INIT_19 => X"F7EFBBEEFF3F7DF7FF3E9F7DF7E2450228000000000000000000509425094250",
INIT_1A => X"BAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBF7DFDFDDD555555",
INIT_1B => X"EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAEBAE",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000000000F7EBF5FAFD7EBF5FAFD7",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"2ABEF00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0020105D557FEAA00557DE10AAD5554BA087FFFF55557BD54AAF7FBC01FFA280",
INIT_29 => X"7BD75EF087FFFFEF557BEAB45552E80155AA802AB45AA843FE0008557DFFF080",
INIT_2A => X"FAE820AA5D5557555082ABDF5508557DF45002ABDFFFF7803DE10AA80000AA08",
INIT_2B => X"0051555FFA2AA8200000557DFFFF7AA80000AAD1420AA087BD7555FFD168AAAF",
INIT_2C => X"5557FFDE10AAAEA8BFFA2FBD7545FFD157555085140010F7AEAABFFAAD542000",
INIT_2D => X"BA557BE8A10A284154BAFFAAAAB45007FC2155F7D155545AA80001EFAAFBEAB4",
INIT_2E => X"000A2D155410F7FFFFEBA08003FE00082AA8AAAAAFFC00BA00002AAAAF7D5574",
INIT_2F => X"0492E3F1C71C7BE8A2ABD7000000000000000000000000000000000000000000",
INIT_30 => X"3AE38145B78FD7000005010495B7AE921C517DE10A2DB50482147FFAF554971D",
INIT_31 => X"E3FE28B684070AA1C71D25D7007FFAFD7497BE8B5555208217DBE8A2AB45BE80",
INIT_32 => X"7FD257DFFD568A82FFA4870BA555F5056D002EBDF6D005B78F7D142ABDFC7F78",
INIT_33 => X"FAAAFBFFBED547038145B505FFB6A487000005F7AFD7F7A482038AADF4709214",
INIT_34 => X"AA8E071D7AAFBEFB455D71F8E00A2A0ADBC7A2FFD257DE3DF52555085142000F",
INIT_35 => X"21C002AA92FFDF574824171EAA10B680124BAFFAAAFB45007BC217DEBDB55555",
INIT_36 => X"00000000000000000000B6D550428FFF1FDE821C003FE001C2EAAAAAB6F5C208",
INIT_37 => X"0105D7BE8B55085142010AAD157545F7AEA8B550000000000000000000000000",
INIT_38 => X"01EFF7AAA8B55F7802AABA5D7FEAB45080015410007FEAA0055517DE00A2FFC0",
INIT_39 => X"E8BFF5D2ABDF55F7AABDEAAF784154BA5D5140145007BE8B55087BEAB555D040",
INIT_3A => X"0020BAA2FFD54105D7FC21EFFFD16AA10FF80174AA557FC21EF082EBFFEF007B",
INIT_3B => X"FBC0155085540000FFAEBFFEFF7D1554BA5D7BC01FFFF8015410007FEAB45F78",
INIT_3C => X"87FC01EFA2FFD7545AAAE97555A2FBFDF455D556AA00A2803FF45AAFFC21EFAA",
INIT_3D => X"552EAAAAAFFD1400005D042AA00F7FBD5410085568A10FF80020AAFFAABFF550",
INIT_3E => X"0000000000000000000000000000000000000F7D1400BAFFD57FE005D043FE10",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(13),        -- Port A data input
DOA(0)   => data_read_a_hi_256(13),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(13),        -- Port B data input
DOB(0)   => data_read_b_hi_256(13),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_14_13 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10020A000180000284008280000281800000030000000033022000000580002",
INIT_01 => X"000008020000204D006800000030824840000000084000084200090008510200",
INIT_02 => X"0220043170010A600A4D008040080000041000000028009002000F333240800C",
INIT_03 => X"111813400008002400000000C400090011000000610200001104D83000F14000",
INIT_04 => X"0801800100A000000000540084000040000040000800200000C8100000000748",
INIT_05 => X"0100000000001000000000002000080008000000001000000024024001200020",
INIT_06 => X"819EB84028001010000000080400000000000004108000100000020020040081",
INIT_07 => X"92040608000440100102400A94810206844200021DA2A0002000340800062C80",
INIT_08 => X"000000000084400008800A001214040441481500040000000000A7F408002244",
INIT_09 => X"0A0040090002008420401004104444004000020400214A208001000002400120",
INIT_0A => X"0400002020000000000000000000080C8008088100004590111B480040120000",
INIT_0B => X"1000000200404800000504016000002114000008020000020080024000000000",
INIT_0C => X"0410000010000000000040001000000000000040000000000001000000000000",
INIT_0D => X"04810244825010004010000000000000000000000000000000080000B8002104",
INIT_0E => X"0002C38280001202020800000000001000004000000000401022000002040902",
INIT_0F => X"20000587050001404E8084341CBA3404800828805200008000E0E0A000080002",
INIT_10 => X"4D18178E012010C00224004091C3514072C000444A0400080001C1C140001000",
INIT_11 => X"51709A07424142084458476001003809D0104B01C5710044020C4006010500C5",
INIT_12 => X"C26EE3803180C18006519462A00005001460E4730000050A1011004001060049",
INIT_13 => X"01F9E00660318000000538318740000140000001B4600CE80001400000002B62",
INIT_14 => X"0000000AD89857B0E0684411800000003799EB764D000330C300000000E3554B",
INIT_15 => X"0000021002002C000024008284001A0902000422E3F5960080480A0216A07240",
INIT_16 => X"4090240902409024090240902409024090081021020080015134920800480010",
INIT_17 => X"0902409024090240902409024090240902409024090240902409024090240902",
INIT_18 => X"9024090240902409024090240902409024090240902409024090240902409024",
INIT_19 => X"F5579B4E5C8FF0F7BE9D5F7DF650400200000000000000000000409024090240",
INIT_1A => X"9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7BF7DDDDDFCF3CF3D",
INIT_1B => X"F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE79E7",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000003FFF03F9FCFE7F3F9FCFE7F3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"420BA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"BD54AAF7FBC01FFA2802ABEFA2FBE8B55A2AE80000F7D5555555D2AAAABAAAD1",
INIT_29 => X"AA801FFA28402000AAAE955455500155EF0804155EFAAD5554BA087FFFF55557",
INIT_2A => X"7AEA8B45080417400AA843FE0008557DFFF0800020105D557FEAA00557DE10A2",
INIT_2B => X"087FFFFEF557BEAB45552E80155AA802AB4500516AA00A2AE800BAFFFFC20BAF",
INIT_2C => X"0AA80000AA005568ABAA28402010A2843FEBAFFFBD7410A2D168BFF087BD75EF",
INIT_2D => X"005D7FFDF4555517DFEF00043FEAA082ABDF5508557DF45002ABDFFFF7803DE1",
INIT_2E => X"000AAD1420AA087BD7555FFD168AAAFFAE820AA5D5557555002E80155A280000",
INIT_2F => X"0555412AA8ABAAADB40092000000000000000000000000000000000000000000",
INIT_30 => X"50482147FFAF554971D0492E3F1C71C7BE8A2ABD7A2FFEDB55B6A080038E3DB5",
INIT_31 => X"B7AE921C517DE10A2AE851FFB68402038AAAA955554900105FF0800175D7A2DB",
INIT_32 => X"A0800BAE3F1C0092EBAAADB6D080A12410BE803AE38145B78FD7000005010495",
INIT_33 => X"2D568BC71C71D25D7007FFAFD7497BE8B5555208217DBE8A2AB451C556FA00A2",
INIT_34 => X"142ABDFC7F78E3FE28B684070AA00516DABAA28402038B6803DE82F7F5D5410A",
INIT_35 => X"D002A80155B680000105D7FF8F455D5F78FD7000E3FEAA002EBDF6D005B78F7D",
INIT_36 => X"00000000000000000000AADF47092147FD257DFFD568A82FFA4870BA555F5056",
INIT_37 => X"F55FF84000AAAAFBC0145002AA8AAAAAFFC20000000000000000000000000000",
INIT_38 => X"01EF080417555A2FFC00105D7BE8B55085142010AAD157545F7AEA8B55A2FBFF",
INIT_39 => X"EAB45080015410007FEAA0055517DE00A2AA955FFFF80020BAAAAA9754508000",
INIT_3A => X"AA8B555D557FE00A280020BAAAD140000A2AEBFFEF082A82010F7802AABA5D7F",
INIT_3B => X"803DE00FFD557400AAD56AB455D5140145007BE8B55087BEAB555D04001EFF7A",
INIT_3C => X"82EBFFEF007BE8BFF5D2ABDF55F7AABDEAAF784154BA08557FEAAA284000AAFF",
INIT_3D => X"FF80174AA557FC21EF082A80145F780020105D7BEAB45557BE8B45082EBFEBA0",
INIT_3E => X"0000000000000000000000000000000000000A2FFD54105D7FC21EFFFD16AA10",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(14),        -- Port A data input
DOA(0)   => data_read_a_hi_256(14),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(14),        -- Port B data input
DOB(0)   => data_read_b_hi_256(14),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_15_13 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000A000000000284000280000001800020030000000033022000000180002",
INIT_01 => X"8000080000000048000000000000026040000000080000080200000000110200",
INIT_02 => X"0020042004010E60004C0080000800000410000000020090020000300245E005",
INIT_03 => X"0000010000080400000000408400480111000000610008000000C00000E54400",
INIT_04 => X"980000010000000088C2550080000040000040000008A00028C8100000120000",
INIT_05 => X"020004012E025000000001322000000A28008000011000000220004D41000000",
INIT_06 => X"819588000800101000011008040000100001060418800510000A620000000092",
INIT_07 => X"0000000800044004010C20008440810284020002102220002000340800062480",
INIT_08 => X"0000000001140800002C0A001214050540C800400406180000002DF004000244",
INIT_09 => X"1E00400900000000000016041044400440000000000042008001000000000022",
INIT_0A => X"0000000000000220000000000000080C00000081000045901118000040000000",
INIT_0B => X"0000000200404000010500004000000114000009000000000000004200000000",
INIT_0C => X"0000000000000000000040001000040001000000000000000001000020000800",
INIT_0D => X"000000000000001001208000180800000000030200000180800C400030002000",
INIT_0E => X"0000000000002600020800000000001080004000000000000002000000000000",
INIT_0F => X"A400000000000000000008000000000000000000000014800000000000000052",
INIT_10 => X"0000000000000000000000010240000000000000000000290000000000000000",
INIT_11 => X"2001C05838120800000000000000000000010000000000000000000000001804",
INIT_12 => X"081004000000000000A010000000000000902000000000180010002020000000",
INIT_13 => X"6600000000000000000024080000000000000000280400000000000000000000",
INIT_14 => X"0000000000200801000000000000000000501001920000000000000000000A40",
INIT_15 => X"0000020000000000000000003000000000000000000A101C3614000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000080000120980000000010",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000400200000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"28BEF00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"5555555D2AAAABAAAD1420BAFF8000010082A954BA00003DFEF085155400F784",
INIT_29 => X"AE95555A2FBE8BEFA2843DE00AA8015400FF84001EFA2FBE8B55A2AE80000F7D",
INIT_2A => X"2FBEAB45F7D56AABAAAD5554BA087FFFF55557BD54AAF7FBC01FFA2802ABEFF7",
INIT_2B => X"A28402000AAAE955455500155EF0804155EFFFFBE8BFF0800174AA557BFDE10A",
INIT_2C => X"A00557DE10F7D1574AAA2D16AB55FFD568BEF087FE8A1055003FE00A2AA801FF",
INIT_2D => X"00AA802AA00AAAE800BA5D0015545AA843FE0008557DFFF0800020105D557FEA",
INIT_2E => X"00000516AA00A2AE800BAFFFFC20BAF7AEA8B45080417400FFFFC21450800154",
INIT_2F => X"8FD7005150438F78A2DBFF000000000000000000000000000000000000000000",
INIT_30 => X"EDB55B6A080038E3DB50555412AA8ABAAADB40092E38E070280024904AA1C043",
INIT_31 => X"1C71C7BE8A2ABD7E3AA9257DA2FFE8BC7BE8E38E10A28017400E38A051FFA2FF",
INIT_32 => X"00124AA557FFDE10A2FBEDB6DF7D16AABAA2DB50482147FFAF554971D0492E3F",
INIT_33 => X"10038E38A2AE851FFB68402038AAAA955554900105FF0800175D7E3FFEFBD700",
INIT_34 => X"000005010495B7AE921C517DE10FFDF50482A2DB6AB45FFD56DBD7087BEAA384",
INIT_35 => X"0FFF1C017D140410400BE8E28A10AAA085082550A1057DBE803AE38145B78FD7",
INIT_36 => X"000000000000000000001C556FA00A2A0800BAE3F1C0092EBAAADB6D080A1241",
INIT_37 => X"4AA0800020BA550028B550855400AAF7AEBDFEF0000000000000000000000000",
INIT_38 => X"7400AAAE975EFA2FBFFF55FF84000AAAAFBC0145002AA8AAAAAFFC2000AAAA97",
INIT_39 => X"E8B55085142010AAD157545F7AEA8B55AAAE821EFAAFBEAB55F7AAA8A00AA841",
INIT_3A => X"417555AAFFFDF450804020AA557BFFE10A2FFFFFEFF7D568ABAA2FFC00105D7B",
INIT_3B => X"D17DF45007FE8AAA08002AAAAA2AA955FFFF80020BAAAAA975450800001EF080",
INIT_3C => X"7802AABA5D7FEAB45080015410007FEAA0055517DE00FFFBC2000AAFBE8B55F7",
INIT_3D => X"A2AEBFFEF082A82010FFD5421EF5D0000010F7AAA8A10AA8017400552A801EFF",
INIT_3E => X"00000000000000000000000000000000000005D557FE00A280020BAAAD140000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(15),        -- Port A data input
DOA(0)   => data_read_a_hi_256(15),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(15),        -- Port B data input
DOB(0)   => data_read_b_hi_256(15),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_16_13 : RAMB16_S1_S1
generic map (
INIT_00 => X"DA22C618B1000482B688B186588884862A400438255FC38381441205BA803003",
INIT_01 => X"7045A80028404C211203A952A90341080B173340412000E1005D628000820484",
INIT_02 => X"428406A4000850848330118D0AAC55001349B108818005460229044001C01784",
INIT_03 => X"092C4020000500020000500986812C405000001A48202050000A214AC0650115",
INIT_04 => X"4804A55440256F504025E003A054F46415A4E62B6FE3307943965A00001A1152",
INIT_05 => X"0000001C40A5B950ADB8EA097057ECE14C86D2B7F85AAD17F4B100000B88148C",
INIT_06 => X"415401DCDCF2C0A8030140BCB0820A200342A1C641C1E8782F508F2B00003584",
INIT_07 => X"002701881A3202080AE00480A2002840BE1480FA004342AA6F12000054004867",
INIT_08 => X"08C54828091002000002B32A8C19064E486A8001510000014140C1E2A14891E0",
INIT_09 => X"015452B103020814004088B64102680B6596594800400413CAC0208944800000",
INIT_0A => X"96AA000484094C000000000000012C9000A0000D0A80000BF8028E87C1B99270",
INIT_0B => X"014808A02004200E540480212000A448C0082024AE50064B44000000000002A2",
INIT_0C => X"0004000D5846256AAEA811150445411150445411150445411150422A088A8200",
INIT_0D => X"00000004010042A204A0C5817D00005034052E40000817D00440004004AD3240",
INIT_0E => X"632B2673FA4587978A2004102800809225545155121740000004900090000000",
INIT_0F => X"00C6564CE7F4EA4B940076D296D003030800462CBD320018CAAAACFE9164C800",
INIT_10 => X"28834ADB1440A114793A4A30A40839AA14910D08DCB2640031955559FD3AC990",
INIT_11 => X"594AB0B1A025371CA0E034E8443C097A800EB090D4AAC91208ED2FA0CE5E09B1",
INIT_12 => X"7B50446083001B94BB38C540EBE61284BB304880E3E4579EDC00992980D58033",
INIT_13 => X"5511121840E7A2CD952ECC12ABC3E6ACB3DFB12ECE315000F61FF1727A85FDBC",
INIT_14 => X"75DEB07F6F2E7084517F126F8395CB2BEFBAB8BA8AF698228CC5E2F08ECA5159",
INIT_15 => X"5580A840A8009F8B108C80A1021B080AFC0DF6422C6077F4A77F20D0C0E21084",
INIT_16 => X"0000000000000000000000000000000000044000102A0001148442A110810359",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"558D11544C690DA64C1C4F68A360400000000000000000000000000000000000",
INIT_1A => X"14D14D14D14D14D14D14D14D14D14D14D14514514514514529E5F87869E79E78",
INIT_1B => X"D1E8F47A3D1E8F47A7D3E9F4FA7D3E9F4FA7D3E9F47A7D1E9F47A7D1E9F4D14D",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000007D3E9F4FA7D3E8F47A3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"C00AA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"03DFEF085155400F78428BEF087FFFFEFF7D168B55AAD17FFFF552EBFE00007F",
INIT_29 => X"2E975EFF7D568BFFFF80175EF0004000BA552A821FFFF8000010082A954BA000",
INIT_2A => X"55540000082EAABFFA2FBE8B55A2AE80000F7D5555555D2AAAABAAAD1420BA5D",
INIT_2B => X"A2FBE8BEFA2843DE00AA8015400FF84001EF0000020AA5D00154005D043FF455",
INIT_2C => X"FA2802ABEF557BEABEF5D0415410087FD74BAAAAEBFFEF557FC00AAF7AE95555",
INIT_2D => X"FFFFAABFEAAFF84001FF002A821FFAAD5554BA087FFFF55557BD54AAF7FBC01F",
INIT_2E => X"000FFFBE8BFF0800174AA557BFDE10A2FBEAB45F7D56AABA082A97545F7D16AB",
INIT_2F => X"FFEF552AB8E38087FC2092000000000000000000000000000000000000000000",
INIT_30 => X"070280024904AA1C0438FD7005150438F78A2DBFF0871F8FC7E3D56AB6DBEDB7",
INIT_31 => X"AA8ABAAADB400924920925EFF7D16ABFFE38E175EF1400000BA412E871FFE38E",
INIT_32 => X"0A1240055003FF6D5551420101C2EAFBD7A2FFEDB55B6A080038E3DB50555412",
INIT_33 => X"57FC00BAE3AA9257DA2FFE8BC7BE8E38E10A28017400E38A051FF0804050BA41",
INIT_34 => X"4971D0492E3F1C71C7BE8A2ABD74975EDBC7550E12410087FD74AAB6AABFFC75",
INIT_35 => X"A08249756DF7D168BC7F7AABAEAAF780051C70824851D7A2DB50482147FFAF55",
INIT_36 => X"00000000000000000000E3FFEFBD70000124AA557FFDE10A2FBEDB6DF7D16AAB",
INIT_37 => X"B55A2D16ABEFFFFBFDFFF552AAAAAA007BC00000000000000000000000000000",
INIT_38 => X"20AA002A955EFAAAA974AA0800020BA550028B550855400AAF7AEBDFEF08516A",
INIT_39 => X"000AAAAFBC0145002AA8AAAAAFFC20000000021EFF7D568BFFA2AA955FF5D040",
INIT_3A => X"E975EF0800174BA002E820105D003DFEF5D51420005D2ABFF45A2FBFFF55FF84",
INIT_3B => X"7BD74AAF7AEBDF455D7BC20BAAAAE821EFAAFBEAB55F7AAA8A00AA8417400AAA",
INIT_3C => X"2FFC00105D7BE8B55085142010AAD157545F7AEA8B5500557DF45552A8200000",
INIT_3D => X"A2FFFFFEFF7D568ABA0804155FFF7D568B55FFAAAAABAFF8415545000015555A",
INIT_3E => X"0000000000000000000000000000000000000AAFFFDF450804020AA557BFFE10",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(16),        -- Port A data input
DOA(0)   => data_read_a_hi_256(16),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(16),        -- Port B data input
DOB(0)   => data_read_b_hi_256(16),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_17_13 : RAMB16_S1_S1
generic map (
INIT_00 => X"5284CE4FB7BD2C8994A13392DBD02E14006B82AC7E800D44D3DD2FD5F9B961C0",
INIT_01 => X"2EACD01F7E03FC6793F2199B39FC233C11D93AE6F3BB92B32091DBC339B24542",
INIT_02 => X"E63CCCC00A82C08092A2AFAE667033DB50853379C10BFDC5C6F4044443C817C6",
INIT_03 => X"7FF183635AEF9E3635AEF9E18E237040404446965C0607EE6DB7854AC4DE060C",
INIT_04 => X"D78AC33FB604488B000892EF17BE6D84196482236FE100294152E294350FB697",
INIT_05 => X"081B5F9B409420D0CDB47A05403F6CE0C08A4AB7F840EDB6F48100DFC8081081",
INIT_06 => X"768465354781CBC30316367077B4BDB50646E8D87100A8201ED01C19C020F71A",
INIT_07 => X"4002A110C922480A82D0841147162C48EBB9537A0022DC67987042EE976ABEA7",
INIT_08 => X"DB931BFEF91C00002CC0E019C0C82A4E4820C15A2330E004401891181168C4D1",
INIT_09 => X"09F3A1BC11EFBC66DB65307071477FF1030C397C060B4254064302042F803A69",
INIT_0A => X"3F330802162F3B7EE3F3EC7C7DEF207000F00059D2ED56D7EED2ED3C9A867DC0",
INIT_0B => X"185C44B91BC1740B7605040BE0018CFC7429F326B9E822FFC00074D5A0AB033A",
INIT_0C => X"00367A28FC1B7F7FEFFCFBFF3EFFCFBFF3EFFCFBFF3EFFCFBFF3EFFE7DFF9E00",
INIT_0D => X"0000000008004BA78428C7AD7FC94B533F5B4FFBD2FAD7FCCA786D43FE67C218",
INIT_0E => X"BA494CEBFD4F2667ABB6F68B29760593F33FA0CF170F40006001B1A05C000000",
INIT_0F => X"7F749299D7FAEB237DFE5865B6D2BF23265CBACE542A6FEE92333AFF33E0A9BF",
INIT_10 => X"F6C24B6D18C3C9F8E2881F3F787D776B5DB94A09955054DFDD246675FE7AC153",
INIT_11 => X"BFB349E08FF9A27EDE9FA8AEFD9E7467BFCB195CFEB56A1A70D34D1706FFFA3E",
INIT_12 => X"6FE219CA80725B875EED723FF7FCB2875EDAAFEAF7FD929BFD55BBC71D79F639",
INIT_13 => X"546670D018E7A6E581D7B6AB75FDFCECA6E581D7BB5DDFC6FF0EB7D7E859FDB5",
INIT_14 => X"B978177F6D6AF5ECDB5FB76A5F5FA165B456E0FB308710C49FCFB741598B9C7E",
INIT_15 => X"CFDAAB00AC00A8BBFC8B501CF7A0FED9A540EA1952586CEB54D143ACFF9A3BA9",
INIT_16 => X"000000000000000000000000000000000026E100002F382DBD9ECFE117805F20",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"4372003009EDCC4052E917114F981800C0000000000000000000000000000000",
INIT_1A => X"BA69A69AEBA69AEBA69A69AEBA69AEBA69A69A69A69A69A68698686981D75D74",
INIT_1B => X"6A351A8D46A351A8D068341A0D068341A0D068341A0D46A341A0D46A341A69AE",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000000000046A351A8D46A351A8D4",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"7FEAA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"17FFFF552EBFE00007FC00AA087FFFFFFFFFFFFFEFF7FBEAB450804001EFAAD5",
INIT_29 => X"D168A000004020AA5D7BE8B450051401EF087FD74AA087FFFFEFF7D168B55AAD",
INIT_2A => X"D7FEAB55FF80175EFFF8000010082A954BA00003DFEF085155400F78428BEFAA",
INIT_2B => X"F7D568BFFFF80175EF0004000BA552A821FF5D00020BA552A82000552A821555",
INIT_2C => X"AAAD1420BAFFFFFDF45AAD17FFFFAAFBC01EF5D0015555557BFDEBA5D2E975EF",
INIT_2D => X"BA007FEABEF005555555A2D1554BAA2FBE8B55A2AE80000F7D5555555D2AAAAB",
INIT_2E => X"0000000020AA5D00154005D043FF45555540000082EAABFF00516AA10552E820",
INIT_2F => X"8B550000071EFB6DF7AE92000000000000000000000000000000000000000000",
INIT_30 => X"F8FC7E3D56AB6DBEDB7FFEF552AB8E38087FC2092147FFFFFFFFFBFDFC7EBF5E",
INIT_31 => X"150438F78A2DBFFBED16AA381C0A07082497FEFB6D1451471EF007BD04920871",
INIT_32 => X"2A850105D2A80155417BEFB6DEB8E175FFE38E070280024904AA1C0438FD7005",
INIT_33 => X"D7BFAEBA4920925EFF7D16ABFFE38E175EF1400000BA412E871FF550A0009249",
INIT_34 => X"E3DB50555412AA8ABAAADB40092FFF5FFF6DAADF7FFD7B6F1C71EF55001756D5",
INIT_35 => X"7145B6AA28492487082007FEDBD700515556DA2DF50492A2FFEDB55B6A080038",
INIT_36 => X"000000000000000000000804050BA410A1240055003FF6D5551420101C2EAFBD",
INIT_37 => X"FEFF7FBFFF55A2D16AB550000175EFFFFBEAA000000000000000000000000000",
INIT_38 => X"55EF087FC200008516AB55A2D16ABEFFFFBFDFFF552AAAAAA007BC0000557FFD",
INIT_39 => X"020BA550028B550855400AAF7AEBDFEFF7D568AAA5D2A97410007BFFFFF55515",
INIT_3A => X"A955EF5D2E80010002A954005D2A82155087FFFFEFAAAA975EFAAAA974AA0800",
INIT_3B => X"D1575FF5504175EF5D7FEAAAA0000021EFF7D568BFFA2AA955FF5D04020AA002",
INIT_3C => X"2FBFFF55FF84000AAAAFBC0145002AA8AAAAAFFC2000FFD57DFFFAAFFFDF55FF",
INIT_3D => X"5D51420005D2ABFF45557FE8AAA000415410007BFFF450051555EFA2FBC0000A",
INIT_3E => X"00000000000000000000000000000000000000800174BA002E820105D003DFEF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(17),        -- Port A data input
DOA(0)   => data_read_a_hi_256(17),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(17),        -- Port B data input
DOB(0)   => data_read_b_hi_256(17),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_18_13 : RAMB16_S1_S1
generic map (
INIT_00 => X"69844019080000A21A611406840014122A641074155FC28A2024001001801003",
INIT_01 => X"7443D920034004180005E9E3C90360C0041C0181002001602025800008440084",
INIT_02 => X"E2DCCCE61D5C008103F2000781FC0FEDEAC2161B0B8FB0008620044443006010",
INIT_03 => X"884E300802006900802006995C896D605200000856E24A040000640052141103",
INIT_04 => X"480520FC026125AC0025C9122644E3E40EC8E2001001302281841A009038A86A",
INIT_05 => X"432000040089983070019400F01010004C8DB841405A80A100B586200FAC24AE",
INIT_06 => X"09044359DC7040000000002C109B0E0A00A1104641C0803804000707284600E1",
INIT_07 => X"400D10100400481D5EB08501620000007500CE801241021FE78E404860140060",
INIT_08 => X"00880C0106A0528020019307CC082A0A4A6A01ED725021400040D028000A9729",
INIT_09 => X"00117063038000282081402E4106400B6186128040600C10C1C0200950508110",
INIT_0A => X"C0C30C2E21580C874004008080003C32A10A19090C02010E1022944061688000",
INIT_0B => X"0180A8062026000DC425C0301311324AA2373088479105D044A1022000001835",
INIT_0C => X"0D89844703649000000200000000000000000000000000000000000000000010",
INIT_0D => X"0D8306C182701404C1973010802020404084001E00010802046092B5001FB365",
INIT_0E => X"528EB314068AB8B803DB00002900800400FC503F08180050942E4200020C1B06",
INIT_0F => X"40A51D66280D6032C5F96D3C51555D5D7D5AA87285820814A3CCC501C2A60820",
INIT_10 => X"8B35A3FEBF1FEDFD9C2B30E0468AAAD5D48F37E8FC1304102947998A03984C10",
INIT_11 => X"440FE1DD772D37A0A321BC6968F32658BF2D4F2A80BF8FE3F9FE3AC362080529",
INIT_12 => X"5487910D7E5A6D961A28456A1832E5161A100DD5182BC54020EA67A189C6ED36",
INIT_13 => X"AA444CAF91EDD1B725868403BE06323551B725868A100ABD119753B70964122B",
INIT_14 => X"EDC259048ACD868EE3803D65CEDC258A8F80D55E007C3F8EBB56F4C5362C978F",
INIT_15 => X"3F240014BE84370001B6922070440556B15F7FABBC0031BCF2257C41634B14D4",
INIT_16 => X"C1B06C1B06C1B06C1B06C1B06C1B06C1B0491069068000004060300A005A0118",
INIT_17 => X"1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06",
INIT_18 => X"B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C",
INIT_19 => X"B28BBECEB80EE173C2300F7DF16000000000000000000000000041B06C1B06C1",
INIT_1A => X"8A28A28AAAAAAA28A28A28AAAAAAA28A28A28A28A28A28A2910591505C104104",
INIT_1B => X"28944A25128944A25128944A25128944A25128944A2552A954AA5128944AAAA2",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000128944A25128944A251",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"9540000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"BEAB450804001EFAAD57FEAA087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974BA082E",
INIT_29 => X"7FFFFFFFFFBFDF45AAD568B55080028B55002E82000087FFFFFFFFFFFFFEFF7F",
INIT_2A => X"0043DE10AA843DE00087FFFFEFF7D168B55AAD17FFFF552EBFE00007FC00AA08",
INIT_2B => X"0004020AA5D7BE8B450051401EF087FD74AAAAFFFDF45A2D16AB55F7FFFFFFF0",
INIT_2C => X"0F78428BEFAA80000000804154BA55042ABEF5D7FD75FFAAD540145AAD168A00",
INIT_2D => X"00082E95555085168A10557FD7545FF8000010082A954BA00003DFEF08515540",
INIT_2E => X"0005D00020BA552A82000552A821555D7FEAB55FF80175EF5D00020105D2A974",
INIT_2F => X"DFFF5D2A954AA082A92428000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFBFDFC7EBF5E8B550000071EFB6DF7AE921C7FFFFFFFFFFFFFFFF7FBF",
INIT_31 => X"AB8E38087FC2092087FFDFC7E3F1FAF55A2DF6DB7D1C002AB7D002A82028147F",
INIT_32 => X"DF6DB7DE3F5FAFC708003DE28B68E38E280871F8FC7E3D56AB6DBEDB7FFEF552",
INIT_33 => X"ADF4516DBED16AA381C0A07082497FEFB6D1451471EF007BD0492B6F1F8F55AA",
INIT_34 => X"1C0438FD7005150438F78A2DBFFA28407038140410492550A2ABC7497BD25FFA",
INIT_35 => X"F5D0E05000492097428002E9557D1C516FA28417BD5545E38E070280024904AA",
INIT_36 => X"00000000000000000000550A00092492A850105D2A80155417BEFB6DEB8E175F",
INIT_37 => X"FFFFFFFFDFEFF7FBFFFEF552E974AA082A820AA0000000000000000000000000",
INIT_38 => X"ABEF002A800AA557FFDFEFF7FBFFF55A2D16AB550000175EFFFFBEAA00557FFF",
INIT_39 => X"6ABEFFFFBFDFFF552AAAAAA007BC0000087BFDF45AAD568B55AAFBFDFEF55042",
INIT_3A => X"FC2000FFD56AB45A2FFFDFFFAAD16AB4500043DEAAFFAEAAAAA08516AB55A2D1",
INIT_3B => X"2AA8B45087FC01EFA2FFD55EFF7D568AAA5D2A97410007BFFFFF5551555EF087",
INIT_3C => X"AAA974AA0800020BA550028B550855400AAF7AEBDFEFA280154BA55040000055",
INIT_3D => X"087FFFFEFAAAA975EF5D2E974000804154BA082A975EF5D517DEAA007BD5545A",
INIT_3E => X"00000000000000000000000000000000000005D2E80010002A954005D2A82155",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(18),        -- Port A data input
DOA(0)   => data_read_a_hi_256(18),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(18),        -- Port B data input
DOB(0)   => data_read_b_hi_256(18),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_19_13 : RAMB16_S1_S1
generic map (
INIT_00 => X"042200000000000041088001001AA00000000000000000000000500802000003",
INIT_01 => X"040048000024000000000404000000000A22000800000800004A200000000001",
INIT_02 => X"200C8840085EB00480060000001C008002489E0F000405EA0004040404000000",
INIT_03 => X"24004000000000000000000900002C4050000000000069500208400002E14100",
INIT_04 => X"4800200C0000000044002000C80020E40000E200000130200188000000800100",
INIT_05 => X"000000000080181000000000701000004C8000000058800000B1000009880480",
INIT_06 => X"80500081081040000000002C100040400000004641C080380400070100000000",
INIT_07 => X"4020109801A4CE005C00048380142810010564C4100114012002402028044808",
INIT_08 => X"0070700000000000000083004C3902420062000020E0000100004082A140102B",
INIT_09 => X"001150200000000000000026400000016186100000000010C04002C000000000",
INIT_0A => X"007C00008082C0002000000000002C3000000004050001030102040000000000",
INIT_0B => X"0000000000000000000000000000010000800011000000000000000000000BC0",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"000000000000000000000000000000042000760000000000000000010004B200",
INIT_0E => X"0D74002280300F0002FB069040000060000C5003000800000000000000000000",
INIT_0F => X"C01AE8004500744C780687DBA828008080A5FC0D385598035D0008A00C015660",
INIT_10 => X"39D8140040201BF861F0E7D693E6170022408116DFE0AB3006BA0011401D02AC",
INIT_11 => X"5412E4997F5249FD005043B8680CC98F00D0F2DD0140100406FE053A98F6ECC7",
INIT_12 => X"7418663001858040E153888000010840E165D0000000285C246A181C03FE4662",
INIT_13 => X"8199830066F0020858385974000001260208583854E2200000660208D6B1423F",
INIT_14 => X"8235AC508FCE8811042040F008235AE04420C040CF00C031C80009B8F224978B",
INIT_15 => X"030004E00000C220010808C10D9A92A74CD7CF4A09051110AD5A3C9200B7F280",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000118",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"07208BBA3F0C7010C660C7441920000000000000000000000000000000000000",
INIT_1A => X"861869A61861861861869A61861861861861861861861861A8208C4C1534D34C",
INIT_1B => X"984C26130984C26130984C26130984C26130984D26930984C26130984C261861",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000984C26130984C26130",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"174BA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFDFEF5D2A974BA082E95400F7FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0004",
INIT_29 => X"FFFFFFFFFFFFFFFFF7FBFDFFF552E974BAA2FFFFE10087FFFFFFFFFFFFFFFFFF",
INIT_2A => X"004001EFAAAEA8ABA087FFFFFFFFFFFFFEFF7FBEAB450804001EFAAD57FEAAF7",
INIT_2B => X"FFFBFDF45AAD568B55080028B55002E82000F7FFFFFFFFFFFFDFEFA2D568B550",
INIT_2C => X"0007FC00AAF7FFFFFFFF7FBE8B55AAD16ABEF5D2ABFF55080402010087FFFFFF",
INIT_2D => X"55A2FFFDFEF5D2EBFE00AAFFFFEBA087FFFFEFF7D168B55AAD17FFFF552EBFE0",
INIT_2E => X"000AAFFFDF45A2D16AB55F7FFFFFFF00043DE10AA843DE00557FFDFEFA2D16AB",
INIT_2F => X"FFEF552A974AA0000104AA000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFF7FBFDFFF5D2A954AA082A92428E3FFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"0071EFB6DF7AE92EBFFFFFFFFFFFFDFEFF7F5FAFC7492A974AAB6F5F8E101C7F",
INIT_32 => X"F1F8FD7AAD16AB450000001FFBEA4A8AAA147FFFFFFFFFBFDFC7EBF5E8B55000",
INIT_33 => X"00000010087FFDFC7E3F1FAF55A2DF6DB7D1C002AB7D002A82028FFFFFFFEFF7",
INIT_34 => X"BEDB7FFEF552AB8E38087FC2092F7FBF8FC7E3F5EAB45B6DF6FBEF5D2AB8F7D0",
INIT_35 => X"84971F8FC7AAD56DB6DBEF5F8FD7412ABFE28B6F5F8E820871F8FC7E3D56AB6D",
INIT_36 => X"00000000000000000000B6F1F8F55AADF6DB7DE3F5FAFC708003DE28B68E38E2",
INIT_37 => X"FFFFFFFFFFFFFFFFFDFEF552E954AA0004000AA0000000000000000000000000",
INIT_38 => X"54AAF7D568A00557FFFFFFFFFFFDFEFF7FBFFFEF552E974AA082A820AAA2FFFF",
INIT_39 => X"FFF55A2D16AB550000175EFFFFBEAA00A2FFFFFFFF7FBFDFFFFFD568B55002A9",
INIT_3A => X"A800AAF7FBFDFEFF7D56AB45AAD56AB450004001EFFF842AAAA557FFDFEFF7FB",
INIT_3B => X"FFFFFFF552AA8BEF080402000087BFDF45AAD568B55AAFBFDFEF55042ABEF002",
INIT_3C => X"8516AB55A2D16ABEFFFFBFDFFF552AAAAAA007BC0000FFFBE8B55AAD168B55F7",
INIT_3D => X"00043DEAAFFAEAAAAA08556AB55A2D57FFFFF7D568B45002ABDEAAFFD16AA000",
INIT_3E => X"0000000000000000000000000000000000000FFD56AB45A2FFFDFFFAAD16AB45",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(19),        -- Port A data input
DOA(0)   => data_read_a_hi_256(19),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(19),        -- Port B data input
DOB(0)   => data_read_b_hi_256(19),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_20_13 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000003",
INIT_01 => X"F55FF80000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"E05022020800008400F655001FFCFF80018FA804400000000000004400000001",
INIT_03 => X"00000000000000000000000900002CC07000000000000000000000000000013F",
INIT_04 => X"68002FFE40900010000180000001FFEC0012EE0C001370F40780000000000000",
INIT_05 => X"0840000880FCBBF0100E204DF0F88311DD8005080679800000F3000029980580",
INIT_06 => X"001000030817C8E8840155FDF9001001050023F6C3C3D0F87FA19F7F011000E4",
INIT_07 => X"000000090492260800008000EE00000000000000002101FF2002C00000004018",
INIT_08 => X"2A040001071004000013FF7FCA302C0C0008214800002101554031F800000000",
INIT_09 => X"801F57F200000090000489FEC0000001EFBEF0040008023FDFC0000000004006",
INIT_0A => X"0000000008000000000000000000ADF000000200000008000008028300110230",
INIT_0B => X"0000000000000800080000000000000000000000000000000800800A40000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"000000040900005C848538000020000000800000080000020000800101FFB600",
INIT_0E => X"00800000003A010003000000000000600FFC53FF001800000002004080000000",
INIT_0F => X"0001000000007408040000004000000004E9000008020000200000000E800800",
INIT_10 => X"00200000000313100010002000008000000000129600040000400000001D0010",
INIT_11 => X"81C012060000000000218F7840000100800004000000000066C0000080080000",
INIT_12 => X"800000000017C000100000000001A800080000000001A8040000002840008185",
INIT_13 => X"0000000006F00000100200000000012600001004000000000066000000801040",
INIT_14 => X"0000200410100000000005F00000020080090A0000000085C800002000586000",
INIT_15 => X"FF00400000000000020020020001000040283024E4F2860400008000030ED080",
INIT_16 => X"00000000000000000000000000000004010201001003020200000000000127DB",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"A0700030038200010089120104D2040020000000000000000000000000000000",
INIT_1A => X"2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2C30C30C30C30C306982121A1E79E79",
INIT_1B => X"32190C86432190C86432190C86432190C86432190C86432190C86432190CB2CB",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000432190C86432190C864",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0201000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF552A974AA0004174BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA0804",
INIT_29 => X"7FFFFFFFFFFFFFFFFFFFFFFEF552E954AA000400000F7FFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E954BA007FC00BA087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974BA082E9540000",
INIT_2B => X"FFFFFFFFFF7FBFDFFF552E974BAA2FFFFE10FFFFFFFFFFFFFFFFFFFFFBFDFFF5",
INIT_2C => X"FAAD57FEAA007FFFFFFFFFFFFFEFF7FBFFF550800020BAAAD56AAAAF7FFFFFFF",
INIT_2D => X"EFF7D56AB450000021EFA2D57DE10087FFFFFFFFFFFFFEFF7FBEAB450804001E",
INIT_2E => X"000F7FFFFFFFFFFFFDFEFA2D568B550004001EFAAAEA8ABA5D7FFFFFFFFFFFDF",
INIT_2F => X"FFFF5D2E954AA080005000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFEF552A974AA0000104AAFFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"A954AA082A92428087FFFFFFFFFFFFFFFFFFBFDFEF5D2E974AA000A07000E3FF",
INIT_32 => X"FFFFFEFF7FBFFFFF552E974AA0071C50BA1C7FFFFFFFFFFFFFFFF7FBFDFFF5D2",
INIT_33 => X"EDF6FABAEBFFFFFFFFFFFFDFEFF7F5FAFC7492A974AAB6F5F8E10E3FFFFFFFFF",
INIT_34 => X"EBF5E8B550000071EFB6DF7AE921C7FFFFFFFFFBFDFEFE3F5F8F450004050AAB",
INIT_35 => X"A497FFFFFFF7FBF8FC7EBD168B450804021FFB6D57DE28147FFFFFFFFFBFDFC7",
INIT_36 => X"00000000000000000000FFFFFFFEFF7F1F8FD7AAD16AB450000001FFBEA4A8AA",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2A954AA0800174100000000000000000000000000",
INIT_38 => X"74AA002E95410A2FFFFFFFFFFFFFFFFFFFFFDFEF552E954AA0004000AAFFFFFF",
INIT_39 => X"FDFEFF7FBFFFEF552E974AA082A820AA087FFFFFFFFFFFFFEFF7FBFDFFF5D2A9",
INIT_3A => X"568A00AAFFFFFFFFFFBFDFEFFFFFFDFEF5D2E954AA0051554BA557FFFFFFFFFF",
INIT_3B => X"D16AB450804174AAFFFFFFEBAA2FFFFFFFF7FBFDFFFFFD568B55002A954AAF7D",
INIT_3C => X"57FFDFEFF7FBFFF55A2D16AB550000175EFFFFBEAA005D7FFFFEFF7FBFDFFFAA",
INIT_3D => X"0004001EFFF842AAAA087BFDFEFF7FFEAB45A2D568B550804001EFF7D57DEBA5",
INIT_3E => X"0000000000000000000000000000000000000F7FBFDFEFF7D56AB45AAD56AB45",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(20),        -- Port A data input
DOA(0)   => data_read_a_hi_256(20),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(20),        -- Port B data input
DOB(0)   => data_read_b_hi_256(20),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_21_13 : RAMB16_S1_S1
generic map (
INIT_00 => X"4A302428B824900A128C090A5C1800261500213C005FE812D10420054085A202",
INIT_01 => X"001FFE3440B609703B0427F801A40B8115BC4F655300340288A40D30040E4DD8",
INIT_02 => X"E00424256888D8819801000F9FFFFFFFF149FF1FCA448046C60A0D2437C517F9",
INIT_03 => X"20030640003250640003250F06002CC1740002019824E001CD357832440001FF",
INIT_04 => X"EA2C3FFD400006E04401A8837001FFFC004AEF00080B70E08FB5789421007C5C",
INIT_05 => X"00011A0C40F9FFF80920954FF0F00809DF84A0202879800000F3000029980780",
INIT_06 => X"0805984B7A1FC0A0000101FFF0480080002281F7C3C381F87C03DFFF00009004",
INIT_07 => X"B424068086A205481A60A19000908204A855B000A08A61FF20C3D004D331D340",
INIT_08 => X"1BFA0001600802000023F7FFC08D234B40C2028253000040114200000D0226C0",
INIT_09 => X"EF1F5FF054096C6ADBA169FFC202B1C1FFBEF0440021083DFFCE22DC2880E24D",
INIT_0A => X"45FF0C004041D84862A28C54518DBFF00020004C0A6044901112A0908AA0A300",
INIT_0B => X"018C241102068006C620C03882019480E63180855A492712CC01C49C20201BFE",
INIT_0C => X"08A9464116544302C02D92236488D92236488D92236488D922366446C911B210",
INIT_0D => X"08800444021048034004001890000806002804A0822189000900D80621FFBE00",
INIT_0E => X"060580261013813A2CC396506102C4053FFD5BFF00A04A00200602CA52001100",
INIT_0F => X"080C0B004C202621A85C09411500135844C196D3606941018150098404C1A304",
INIT_10 => X"B02901013416181C96C2C9C600890A2028172192C460D1820302A0130809834A",
INIT_11 => X"9C5E803408250180AC268D185DB3F4350B811068C00049A0A4AA68F05C96A001",
INIT_12 => X"002C006560138F032B1804101244C883052208209040CC849063A747512B7678",
INIT_13 => X"41401E240665750440C9488280254530314080C2C601040420352148A00501B1",
INIT_14 => X"500811204D000700114204A70422016149916011008CAA8858850B00C32591C0",
INIT_15 => X"FFC06E60AC0496022300233104663040808E991765205000070121D41D18D098",
INIT_16 => X"40100401004010040100401004010040102090010008000001C0E010020007DF",
INIT_17 => X"0100401004010040100401004010040100401004010040100401004010040100",
INIT_18 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_19 => X"FFEF9FEEFF7FFDF7FF3E3DFDF7E0000000000000000000000000401004010040",
INIT_1A => X"BEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBFFDFDFFFCF3CF3F",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFEFF7FBFDFEFF7FBFDFEFBEF",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000FFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0001000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E954AA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0004",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA0004154BAFFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"52E974BA0804000AAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0004174BAFF",
INIT_2B => X"FFFFFFFFFFFFFFFFEF552E954AA000400000007FFFFFFFFFFFFFFFFFFFFFFEF5",
INIT_2C => X"A082E95400007FFFFFFFFFFFFFFFFFFFFDFEF5D2E974BA002E97400007FFFFFF",
INIT_2D => X"FFFFFBFDFEF5D2A954AA002E974BA087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFBFDFFF5D2E954BA007FC00BA5D7FFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA000002000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080005000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"A974AA0000104AAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974BA0000174AAFFFF",
INIT_32 => X"FFFFFFFFFFFFDFEF552E954BA080A000AAE3FFFFFFFFFFFFFFFFFFFFFFFEF552",
INIT_33 => X"02A95400087FFFFFFFFFFFFFFFFFFBFDFEF5D2E974AA000A07000007FFFFFFFF",
INIT_34 => X"F7FBFDFFF5D2A954AA082A924281C7FFFFFFFFFFFFFFFFFFBFDFEF5D2A974BA0",
INIT_35 => X"A557FFFFFFFFFFFFFFFF7FBFDFFF552E974BA0020924BA1C7FFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000E3FFFFFFFFFFFFFFEFF7FBFFFFF552E974AA0071C50B",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0000020000000000000000000000000000",
INIT_38 => X"74BA0000174BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954AA080017410FFFFFF",
INIT_39 => X"FFFFFFFFFFDFEF552E954AA0004000AAF7FFFFFFFFFFFFFFFFFFFFFFFEF552A9",
INIT_3A => X"E95410087FFFFFFFFFFFFFFFF7FBFDFEF5D2A954BA082E800AAA2FFFFFFFFFFF",
INIT_3B => X"FBFFFFF552E954BA002E97410087FFFFFFFFFFFFFEFF7FBFDFFF5D2A974AA002",
INIT_3C => X"57FFFFFFFFFFFDFEFF7FBFFFEF552E974AA082A820AA557FFFFFFFFFFFFFEFF7",
INIT_3D => X"5D2E954AA0051554BA5D7FFFFFFFFFBFDFEFF7FFFFFEF5D2A974BA0000020AA5",
INIT_3E => X"0000000000000000000000000000000000000AAFFFFFFFFFFBFDFEFFFFFFDFEF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(21),        -- Port A data input
DOA(0)   => data_read_a_hi_256(21),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(21),        -- Port B data input
DOB(0)   => data_read_b_hi_256(21),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_22_13 : RAMB16_S1_S1
generic map (
INIT_00 => X"5290F4CDE914905A14A43D33F488243E17122300F55FEB189B343A1140548380",
INIT_01 => X"A54007B259F6A975386262000C344BA9573C6FF57B18A5FB0ABFCD3C2C5F4F0C",
INIT_02 => X"021DFF8C38B3C009D203551040030071869D0040180AA2DC53DB89BEA8204001",
INIT_03 => X"2603475A969D0475A969D0460EAA401005111011BD506954EDB40F5EF41434C0",
INIT_04 => X"922D9002100ED69E443D988B0D5400103E48003D0800011E803B06B5B9125A15",
INIT_05 => X"281B5A0C06000408F4DF9422010D8802022F2124A8022492580040440002021C",
INIT_06 => X"F780C4C052881ADA0E05440205DA50930FA182010004700083E220800440B588",
INIT_07 => X"049D028B93FB561833D8094A02F5EA92FD7247E10305C40040D136E6A023F7FC",
INIT_08 => X"00028241680A0E002A9400803A884B5B5206B7C2E53CA25144009007A64EBD64",
INIT_09 => X"41008810240240C6694008010392354010000560141801002028A83D2A08E06D",
INIT_0A => X"34000000848BCA6902A29C54539C020E11810098D4067EFF9FF284D483E2AB41",
INIT_0B => X"500001840000C80B410014088040F4A944B1AA313C0022AA0011C0DC00028001",
INIT_0C => X"80B14004D158C8CA24A1C2A870AA1C2A870AA1C2A870AA1C2A872550E1543800",
INIT_0D => X"80A14050A01509E050854498B5281A1C34E506A2C6898B52A154DAC6B6000850",
INIT_0E => X"0B03001A483A4146603050080410089180008800143D83888281A2034A850142",
INIT_0F => X"A4160600349075238473F1210006133835E92273612B3482C090068A0E84AC56",
INIT_10 => X"30060181BA1B13959DC08DA902458870201970B29602562B0581200D141D0959",
INIT_11 => X"E042021C040D0152C8058B3840F044708E7E1C20A0106EA166C13AFC14AA3804",
INIT_12 => X"080E004B0C17C1439A9838301DC1A8438EA32C009DC1A8255300650458A1D588",
INIT_13 => X"018010E186F110A908E3A8CB0026C9A610A908E6A60F0807626610E160589C4C",
INIT_14 => X"2A701667334005800B1605F043858125E0D04110408D2485CA034681E43A1E40",
INIT_15 => X"00646002304244A91102C93A2D608D2A258DF8034188200C050171A41108F084",
INIT_16 => X"110441104411044110441104411044110466C440446CA06951D4EA8010009804",
INIT_17 => X"0040100401004411044110441104411044110441104411044110441104411044",
INIT_18 => X"0401004010040100401004010040100401004010040100401004010040100401",
INIT_19 => X"F7DFBFDEFE8FF1F7DEBDDF7DF7D05122890000000003FFFFFFFF900401004010",
INIT_1A => X"9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7BFFDFD7DDDF7DF7D",
INIT_1B => X"F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE79E7",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000003F9FCFE7F3F9FCFE7F3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA000400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0800",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000002000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2A954BA000015400FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080402010FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2A954BA0004154BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A0004174BAFFFFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0800154AAFFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF552A974AA0000174BAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974A",
INIT_2E => X"000007FFFFFFFFFFFFFFFFFFFFFFEF552E974BA0804000AAA2FFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080400010000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E954AA080005000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000402010FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2A954BA000417410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"804154BAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974BA0000174AAFFFFFFFFFFF",
INIT_34 => X"FFFFFFFEF552A974AA0000104AAE3FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0",
INIT_35 => X"AA2FFFFFFFFFFFFFFFFFFFFFFFEF552E954BA000E124BAE3FFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000007FFFFFFFFFFFFFFFFFFFFDFEF552E954BA080A000A",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804000100000000000000000000000000",
INIT_38 => X"54AA000400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2A954AA080017410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"0174BAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A954BA000415400FFFFFFFFFFFFF",
INIT_3B => X"FFFDFEF552E974AA0804174AAF7FFFFFFFFFFFFFFFFFFFFFFFEF552A974BA000",
INIT_3C => X"2FFFFFFFFFFFFFFFFFFFFFDFEF552E954AA0004000AAA2FFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2A954BA082E800AAAAFFFFFFFFFFFFFFFFFFFBFDFEF5D2E954BA002A820BAA",
INIT_3E => X"0000000000000000000000000000000000000087FFFFFFFFFFFFFFFF7FBFDFEF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(22),        -- Port A data input
DOA(0)   => data_read_a_hi_256(22),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(22),        -- Port B data input
DOB(0)   => data_read_b_hi_256(22),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_23_13 : RAMB16_S1_S1
generic map (
INIT_00 => X"EF20906D902424807BC8241BC81801B97D38AD3C0800103362A6741C80A12A02",
INIT_01 => X"001FFF8409F089003B4422000D80C80106804A7951C5B9D1C828043EA28838F9",
INIT_02 => X"E01CEE21649C82C40800000F9FFEFF8E72CA7F5FC2E22809925A0D3611C877F8",
INIT_03 => X"24000400402670400402670D48222DC1764446838624000080007460C40001BF",
INIT_04 => X"68403FFC020560E0443E21037C01FFFC0002EE00628BF0E02FAD781014085014",
INIT_05 => X"0112000202FBFFF00920017FF0F0628BFF8488890979800002F702002BB807A0",
INIT_06 => X"EF85788B681FC000000001FFF0010000000001F7CBC385F87C0BFFFF20040001",
INIT_07 => X"F6E200000000C1440E3AE408009120071070FA07A1CB23FFA403F0C4D23BF7C0",
INIT_08 => X"0BF87CA400804000003FF7FFD8880A034AC09662305AB10555421006891A1089",
INIT_09 => X"BE1F5FEA10092C0896A243FFC0008087FFBEF2000000001DFFC612C0C0400100",
INIT_0A => X"41FF0C2060501000600000000001BFFA800808189A657EF81DD0C00079CC8001",
INIT_0B => X"018C24110A860006C620C0312241C482B20400CC52492710CC80060020A81BFE",
INIT_0C => X"0C08866907048320C20C10030400C10030400C10030400C10030400608018210",
INIT_0D => X"040002000041500300100040000500C000801000C02400000952800001FFBF04",
INIT_0E => X"FC850015385380380CDB86106502C5043FFD5FFF00A04BC010A7724B10000800",
INIT_0F => X"89F90A002A70A710A51C01C05904014861433602A1CAF13F2110055614C72FC0",
INIT_10 => X"E02D02001C1E14981B43253EE50C8220180F1082E06397E07E42200AAC298E57",
INIT_11 => X"8421802400A90022B0070FAE18019214A380344920080B21A58B02AC60BACDF0",
INIT_12 => X"0A2A000C480B0704B54028101AC49C84BB4100009AC49C80857A82D20CE8CB22",
INIT_13 => X"01E00C8103416445C12ED0400027C5292445C12D500B0005A62D344CB241D095",
INIT_14 => X"132C907425604680038706A35132C94BDD011010404428886AC91B11311C8280",
INIT_15 => X"FF000470BE0692020328CA0028042054A92771C50FC070110001C1680809591D",
INIT_16 => X"00802008020080200802008020080200800800200200000000000008004807DF",
INIT_17 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_18 => X"8020080200802008020080200802008020080200802008020080200802008020",
INIT_19 => X"0000000000000000000000000000000000000000000000000000008020080200",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080002010FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974AA000400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000400010FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974AA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080000010FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E954AA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954A",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA000015400FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080002010FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974AA000400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000402010FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E954AA080005000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA080407000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA00041741",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080000010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000402010FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2A954AA080002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954AA080017410FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"552A954BA000415400F7FFFFFFFFFFFFFFFFFFFFFFFFF552A954BA080015410F",
INIT_3E => X"0000000000000000000000000000000000000F7FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(23),        -- Port A data input
DOA(0)   => data_read_a_hi_256(23),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(23),        -- Port B data input
DOB(0)   => data_read_b_hi_256(23),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_24_13 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100600007FFF000080108004000800020000840041000080808",
INIT_02 => X"FC5CA803400EB8209000000F9FFEFF8E7240FF1FC22409EA04018E50074017F0",
INIT_03 => X"11100400000000400000000D00002CC07400000090C080019001010A000001BF",
INIT_04 => X"68003FFC00040000000000008001FFFC0002EE00000370E007A100000000E468",
INIT_05 => X"0000000000F8BFF00920004DF0F00001DF8000000079800000F3000029980780",
INIT_06 => X"6E461803081FC000000001FFF0000000000001F7C3C380F87C019FFF00000000",
INIT_07 => X"600C2400013649609C8000980040814210254000A00B21FF2003F2A80D500000",
INIT_08 => X"0BF80000000000000003F7FFD88D2B4A02C0940062EC2804001610020408178B",
INIT_09 => X"8E1F5FE010092C0892A041FFC0000001FFBEF0000000001DFFC002C000000000",
INIT_0A => X"41FF0C0000000000600000000001BFFA0000005501AA00000CE2000009400000",
INIT_0B => X"018C0411020600048620C030020502000200000400490510CC00040020201BF4",
INIT_0C => X"0808064106040300C00C10030400C10030400C10030400C10030400608018210",
INIT_0D => X"0000000000004003000000000000001200580000000000000000000001FFBE00",
INIT_0E => X"0086C022005381380FDB96516140C6043FFD5BFF000041000000004110000000",
INIT_0F => X"80010D804400A7240C840C201D0210840043B4804012500021E0088014C04940",
INIT_10 => X"4109038041021C980200D06410C1924030008142E06024A00043C01100298092",
INIT_11 => X"587CC200002100C14428090A1D02348190814C09C010104025AA40041A0D8005",
INIT_12 => X"022E0030300B0E46177004208000D8C61D7004300000D884817B00011306B2D9",
INIT_13 => X"01E003060344710009875C018100013831000985DC000C20003C310006143B70",
INIT_14 => X"4001850EDC004780144806A64400186CBF8961104000C3807884000846EB9500",
INIT_15 => X"FF0006E08C063C0220002201490418082010A57263E0100008000290161E711C",
INIT_16 => X"00000000000000000000000000000000000000000000000000000000000007DF",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"F2D0AEEAF6E7CC1132CDB4441990000000000000000000000000000000000000",
INIT_1A => X"BEFBE79E79E79E79E79EFBEFBEFBEFBEFBEF9EF9EF9EF9EFA69861219575D75F",
INIT_1B => X"783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1EFBEF",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000783C1E0F0783C1E0F0",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0201000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A000400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA000400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000400000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402010000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"00002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080002010FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000400010FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA00040000",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020100000000000000000000000000",
INIT_38 => X"74BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"000010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA000002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974AA000402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000002010F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(24),        -- Port A data input
DOA(0)   => data_read_a_hi_256(24),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(24),        -- Port B data input
DOB(0)   => data_read_b_hi_256(24),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_25_13 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100200002000000080100004000000020000800041000080808",
INIT_02 => X"FC400086000000800000000F9FFEFF8E738FFF1FC204010000000111568DD7F8",
INIT_03 => X"00000400000000400000000D00002CC4740000008000000080000000000001BF",
INIT_04 => X"68003FFF64A564AC000000000001FFFE0082EF00010370E007A1000000004000",
INIT_05 => X"0A00040148F8BFF80920804DF0F00101DFC040000079C92484F30499299837C1",
INIT_06 => X"66041803081FC0E0801101FFFD000E41002299F7E3C380F87C019FFF81200096",
INIT_07 => X"000000080480AE00000080000000000000000000A00B21FF2003E00000000000",
INIT_08 => X"1BF80000400A02000003F7FFFA0008000200A0400008A0000014100200081000",
INIT_09 => X"8E1F5FFA53EFBCACB2E369FFE0010001FFBEF80C40630C7DFFEEBAF000800202",
INIT_0A => X"41FF0C0600000000600000000001BFFE00301000000000000CC020000140000C",
INIT_0B => X"01DCCC31222730A49620C030020100000200000400490D10EC00040220201BF4",
INIT_0C => X"0808064106240300C00C10030400C10030400C10030400C10030400608018210",
INIT_0D => X"0883044582114013412080000000000000000000000000000012800001FFBE00",
INIT_0E => X"00040020000180380FC386106140C6043FFD5BFF00A04B80608003CB120C1106",
INIT_0F => X"0000080040000200040400000100000000009480000240000100080000400900",
INIT_10 => X"0001000000000808000000240000020000000100006004800002001000008012",
INIT_11 => X"0001001808220000002004001900000080800008000000000022400000088000",
INIT_12 => X"0010000000000E00110000000000408009000000000040808063004000008200",
INIT_13 => X"6000000000046100000240000000001021000004400000000010210000001010",
INIT_14 => X"4000000404000800000000060400000088000001800000001084000000088000",
INIT_15 => X"FF800C608C041002000002000006100000002100000000180600000000100018",
INIT_16 => X"4110441104411044110441104411044510629041040D180400000010028047DF",
INIT_17 => X"1104411044110441104411044110441104411044110441104411044110441104",
INIT_18 => X"1044110441104411044110441104411044110441104411044110441104411044",
INIT_19 => X"FBA2894A196A8C5A2932EC15DA080800002FFFFFFFFFFFFFFFFFC11044110441",
INIT_1A => X"2492492492492492492410410410410410410492410492412000531215A69A6B",
INIT_1B => X"158AC562B158AC562B158AC562B158AC562B1588C46231188C46231188C49249",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000B158AC562B158AC562B",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080000010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000010FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08000000",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(25),        -- Port A data input
DOA(0)   => data_read_a_hi_256(25),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(25),        -- Port B data input
DOB(0)   => data_read_b_hi_256(25),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_26_13 : RAMB16_S1_S1
generic map (
INIT_00 => X"E9264EAB20190CA3BA4997AA9002AE9C001006B0778015CFA17E0811039879C7",
INIT_01 => X"2FFFF9BB1F773C7F9BB07DFFFDD863FC5FFF3FEFFBBF9FFB22FFFBC7B9F30686",
INIT_02 => X"E06CCC62052E708180F6FFBFFFFCFFFFF9C7FF7FC24332E642090000074037F6",
INIT_03 => X"428003739CD9863739CD9869FE2B7DEAF300029E4E300DFE69A6E644E6FF473F",
INIT_04 => X"7C2FEFFFF5BA124F003DD31EAFFFFFEE9FF7EE6F4C0770FFD7DC7CA53997B2B1",
INIT_05 => X"DFFB5421C1F8BBFAFDBFFACDF0FFCC05DDDBFF3690F9EDB7F5F7AFF639BD7DE3",
INIT_06 => X"EFD044ABC817C3E3A74667FDFFB6FF5727CC3BFEF7C3FAF87FF59F7FFBFEF69F",
INIT_07 => X"00003002132462052E708180EF060C18E5BEFB051225CDFF7002C4EEDE77F6E0",
INIT_08 => X"3FFF7D5000EC75088ED3FF7FC8790E46426CE06CB1F8E041051831FA3068D77E",
INIT_09 => X"C05FD7FF9BEFBDCEFBEE59FEF44F6603EFBEFAFCC2E35E7FDFD147CCF3F583FA",
INIT_0A => X"67FF1C7FBFADEB31E35768E8ED6BFDF3EB3EBF9DDBCE7FDC1DF8A760F3EACC02",
INIT_0B => X"5BDDCC3B336F7C548667D47B7737AF3FD62601EDC25B3533DCEB07F262213FFC",
INIT_0C => X"5F9A06E19F4D93A0EA0F78C35E30D78C35E30D78C35E30D78C35E986BC61AE31",
INIT_0D => X"5FD7AFEFDFFAF59B6FF28FE1D80D73D840607307DCFE1D80EF69A004DFFFF7FF",
INIT_0E => X"0004001F8041897B2FFFC6D86D70CE04FFFFF3FF1F5F5475BD7F72E4D75EBFAF",
INIT_0F => X"F60008003F008237B0040A00010003E020023E0201F45EC0010007E01047D17B",
INIT_10 => X"00010001DC0004C81003DE050A700200001DC0006863E8BD8002000FC0208FA2",
INIT_11 => X"2200E400002801E1A00004C21C0206F60081800800007B00010F02007EC09A0E",
INIT_12 => X"0880007E000807C7C1A612001E0015C7C19C22001E0015C59DFE82011A311AA0",
INIT_13 => X"00001BC00101F60409F0670840070809760409F06984800780097604067D0010",
INIT_14 => X"81019F40042100001F800203D81019EC085614000085C80023D81009CF008A74",
INIT_15 => X"FF802FFDFFAFD082003B032FB987E04021D481D4000819060801E0D00001231D",
INIT_16 => X"EBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEFFBFBFBFBBFCFBB0FFDFEFFEF2DFFFFFB",
INIT_17 => X"BFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAF",
INIT_18 => X"FAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFE",
INIT_19 => X"475B15BCF491E166CC8553F86EDB5C88646FFFFFFFFFFFFFFFFFEBFAFEBFAFEB",
INIT_1A => X"861861861861861861861861861861861861869A69A61861AFBD54D5F871C71D",
INIT_1B => X"984C26130984C26130984C26130984C26130984C26130984C26130984C261861",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000984C26130984C26130",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040201",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(26),        -- Port A data input
DOA(0)   => data_read_a_hi_256(26),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(26),        -- Port B data input
DOB(0)   => data_read_b_hi_256(26),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_27_13 : RAMB16_S1_S1
generic map (
INIT_00 => X"00080A40000A41248002029000050A088000008242A0004404480002000A1155",
INIT_01 => X"2FFFF1C11F781C129C107DFFFE0860941E81258CA2B71C2220EC1B86E1A00002",
INIT_02 => X"E1000000810000014400FF6FFFF0FFFFF8007F1FC21110005080200000221FF0",
INIT_03 => X"4080026318C18226318C1821302232EAE00002BE001115FE48620040840A863F",
INIT_04 => X"643D4FFC2530000F003D821C0BFFFF8E9EF79E6D440748FED70060842105B0B0",
INIT_05 => X"D6F39020D1F8A3FAFDBFBACDC8FDC405D1DB7F1490E5EDB7D5CBADB2385D79C3",
INIT_06 => X"6FE000A38007C3032646EFF1F0B6FF46A78C39F8E723F2E47FE59C7F9ADA2612",
INIT_07 => X"00002820000000810000014401060C180190310540118DFF1000C0849673F6C0",
INIT_08 => X"3FF779100062B12A8EC3F47FC80208808210880C00082050000110023068D030",
INIT_09 => X"005F07E09BFFBD07FBAC09F8E42922038F7DF8BEC2E39C5F1FD047CEF1B582D8",
INIT_0A => X"63FF5D5F9FADE911E81C09818109E1F16B16B71092CE7ED81CF403601228C402",
INIT_0B => X"1BFDCC39732F3554866AD57C37BEAF1C152201A4C05B7531D56B05B06A213FF8",
INIT_0C => X"5BCA06F18FC59380F00E34430D10C34430D10C34430D10C34430F0861A2186B5",
INIT_0D => X"5B56ADAB5FAAE58B2F628EA0C80FA3F04040510768EA0C80CC61A0044DFFC6EB",
INIT_0E => X"0004001D800188792CE79715710AE4047FFD23FF315D54358D593474955AB6AD",
INIT_0F => X"520008003B000297B0040200010003E020001F0201E44A400100076000579129",
INIT_10 => X"00010001DC00004A10035E0408300200001DC000086BC8948002000EC000AF22",
INIT_11 => X"02002400002801E1A00000C01E0202F60080800800007B00000782006EC0820A",
INIT_12 => X"0080007E000006A7C10602001E0001A7C10C02001E0001C18DE282010A311AA0",
INIT_13 => X"00001BC00000FE0401F04300400708007E0401F04180800780007E04047D0010",
INIT_14 => X"81011F40040100001F800002F81011EC080604000085C80001F810094F008034",
INIT_15 => X"FF800C6DDDAFD082001B03249887E04001D481D4000009020801E0D00001021F",
INIT_16 => X"AB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6BF1EBDABD8E270BF84A25C6ACB777E3",
INIT_17 => X"B6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6AD",
INIT_18 => X"6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADA",
INIT_19 => X"490E2168100481CA860402104A471688747FFFFFFFFFFFFFFFFFAB6ADAB6ADAB",
INIT_1A => X"000000000000000000000000000000000008200000000000200072F210000001",
INIT_1B => X"05028140A05028140A05028140A05028140A0500804020100804020100800000",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000A05028140A05028140A",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040201",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(27),        -- Port A data input
DOA(0)   => data_read_a_hi_256(27),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(27),        -- Port B data input
DOB(0)   => data_read_b_hi_256(27),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_28_13 : RAMB16_S1_S1
generic map (
INIT_00 => X"02200AA400180030808802A900002A08001280A08A801044104A1000001818C3",
INIT_01 => X"0AA00011460214428114180000882214413D0A71592A01D92213D28005210202",
INIT_02 => X"0451110A012100884000AA30200000000C100040104112101100008888200000",
INIT_03 => X"448000318C52A20318C52A20148810200111100C211004AA00034204200A2200",
INIT_04 => X"04004001001A90110000121402AA0000003C00000500000040080421080D0080",
INIT_05 => X"4060000C8001000000002E000000050000001610300000010000802202040012",
INIT_06 => X"1000002080001111001222000425A1040026A008000000000000000009328280",
INIT_07 => X"2491008A00491201210088400122448908A20402000408001000040820000000",
INIT_08 => X"20058310402A160026500000028040101004200C840082115554000112244814",
INIT_09 => X"4140000800000060000720000102028000000490160801020002200011100010",
INIT_0A => X"020000081B34211082B694D4D294000020020381040000000200032040004400",
INIT_0B => X"4800210C19808400500010009110091500020B408810000100200020408B0000",
INIT_0C => X"01028000080118020023604858121604858121604858121604858090B0242C00",
INIT_0D => X"010000800920040804020A6058003108402043058C460580653020005A004039",
INIT_0E => X"00000002800008014004104104420A00C000200005000010040A0020CC000200",
INIT_0F => X"520000000500000010000200000000000000280000040A40000000A000001029",
INIT_10 => X"00000000000000C0000002000830000000000000480008148000000140000020",
INIT_11 => X"020024000000000000000440000000020000800000000000000C00000040020A",
INIT_12 => X"00800000000001804006020000000500400C0200000005400A90000000100000",
INIT_13 => X"0000000000018200001003004000000142000010018080000001420000200000",
INIT_14 => X"8000080000010000000000018800008000060400000000000310000008000034",
INIT_15 => X"000002040080000000110006B081400000400000000009020000000000002200",
INIT_16 => X"802008020080200802008020080200802101210810C39A66A90A85420413A820",
INIT_17 => X"0200802008020080200802008020080200802008020080200802008020080200",
INIT_18 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_19 => X"DE21102C110A00246972BD89A40A0C22E1000000000000000000002008020080",
INIT_1A => X"2082082082082082082082082082082082082082082082080D35050758C30C31",
INIT_1B => X"0582C160B0582C160B0582C160B0582C160B0580C06030180C06030180C08208",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000B0582C160B0582C160B",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(28),        -- Port A data input
DOA(0)   => data_read_a_hi_256(28),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(28),        -- Port B data input
DOB(0)   => data_read_b_hi_256(28),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_29_13 : RAMB16_S1_S1
generic map (
INIT_00 => X"79964E4BA01DACAB9E659792D00AAE160002829C7FDFEFCEE97C2815039D70C3",
INIT_01 => X"0ABFF9AB0775343F9AB01DF80D5821FC0FFF3FEFD1AF9FF1207FFBC7B9720586",
INIT_02 => X"002CCC60050E700080F6AAA7BFFC007189C7FF2FC00330E602800000074037F6",
INIT_03 => X"468003210868A63210868A68DA017D207200021C4E200CAA6186A40042FF4300",
INIT_04 => X"7C2FE002F0900001003C5316A6ABFFE21F36E02F0D03701F47D41800109FB281",
INIT_05 => X"4979440580F9B808F49F6A4DF00F8D01DC4B97369078249370F482E62BA41462",
INIT_06 => X"B250442BC81001E1870223FC0BF7F11507C423FE33C078F803F19F00E936721D",
INIT_07 => X"00011080012460050E700080EF020408EC8CFA01122149FF700200665A35D260",
INIT_08 => X"2BFD055040A452000443FF00007906464068406C31F84000000831FA1028575A",
INIT_09 => X"805FD017102690AA694551FE30444681E0820AD40201423FC00122C493500172",
INIT_0A => X"0600002AFFBE2330815568A8AD6ABC02A02A0B0CCB463B4C0748A720B1EA4C00",
INIT_0B => X"0850400A11414C005005000B51158936D20601A98A10200308A002E240010BFC",
INIT_0C => X"05928020194918A22A2268C81A32068C81A32068C81A32068C81A99034640C00",
INIT_0D => X"058102C48970541944B20FA1580561D040406305587A158046282000DBFFF13D",
INIT_0E => X"000000028040890327DCD28928324400DFFFF0001F1F0050342D42A086040B02",
INIT_0F => X"F60000000500802010000A000000000000022A0000141EC0000000A01000507B",
INIT_10 => X"00000000000004C0000082010A700000000000006800283D80000001402000A0",
INIT_11 => X"2200E4000000000000000442040004020001800000000000010D000010401A0E",
INIT_12 => X"08800000000801C040A6120000001540409C2200000015441DAC800010100000",
INIT_13 => X"0000000001019600081027084000000956000810298480000009560002200000",
INIT_14 => X"800088000021000000000201D800088000561400000000002358000088000A74",
INIT_15 => X"00802594A282C0000033010FB181E00020400000000819060000000000002305",
INIT_16 => X"C0B02C0B02C0B02C0B02C0B02C0B02C4B12B312912831A27FCFE7FFB175B6FF8",
INIT_17 => X"0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02",
INIT_18 => X"B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C",
INIT_19 => X"BBCF9F96EE7FFDF7FE783FFDFFEA0C00602FFFFFFFFFFFFFFFFFC0B02C0B02C0",
INIT_1A => X"EFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEEBAEBAEBAEBAEBBFFDF9FBEFFFFFFE",
INIT_1B => X"BFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFBEFB",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000FBFDFEFF7FBFDFEFF7F",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(29),        -- Port A data input
DOA(0)   => data_read_a_hi_256(29),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(29),        -- Port B data input
DOB(0)   => data_read_b_hi_256(29),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_30_13 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"F7FFBFFEFF9FE1F7FFBFFFFDFFD0000000000000000000000000000000000000",
INIT_1A => X"9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7AFBD75F5FDF7DF7F",
INIT_1B => X"F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE79E7",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000003F9FCFE7F3F9FCFE7F3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(30),        -- Port A data input
DOA(0)   => data_read_a_hi_256(30),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(30),        -- Port B data input
DOB(0)   => data_read_b_hi_256(30),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_31_13 : RAMB16_S1_S1
generic map (
INIT_00 => X"129000008004A00804A40000400800020000000C005FEA005800200400050100",
INIT_01 => X"255FF18019700810180065FFFC0040801E80258CA2951C2200EC0906A0804140",
INIT_02 => X"E0000000000000011000550FDFF0FFFFF0007F1FC200000044000000000817F0",
INIT_03 => X"0000024210A30024210A3001002220C06044469200040154482000408400043F",
INIT_04 => X"602D0FFC2420000E003D80080955FF8E1ECA8E2D400340FE870060842100B030",
INIT_05 => X"0213100040F8A3F8FDBF944DC0FDC001D1CB6904A061EDB6D4C30490281831C1",
INIT_06 => X"6FC000830007C202060445F1F0D25E4207A099F0E303F0E07FE19C7F80402412",
INIT_07 => X"0000200000000000000001100004081001103107000185FF0000C0849673F6C0",
INIT_08 => X"1BF27A00000000000883F47FC800080002008000000820440000100220489020",
INIT_09 => X"011F07E013EFBC06FBA009F8E00120038F3CF82C44630C5D1FC002CCE0808248",
INIT_0A => X"61FF0C06C48BC801600000000001A1F00110101092CE7ED81CF0004012288000",
INIT_0B => X"11DCCC31222730048620C4382204A608142002A440492530C401049020221BF8",
INIT_0C => X"0888066187448380E00C10030400C10030400C10030400C10030600608018210",
INIT_0D => X"080204010200418301208480800D02D00040100240A808008840800405FF8640",
INIT_0E => X"0004001D000180780CE386106100C4043FFD03FF101D40008001304018081004",
INIT_0F => X"000008003A000217A0040000010003E02000160201E040000100074000478100",
INIT_10 => X"00010001DC00000810035C0400000200001DC0000063C0800002000E80008F02",
INIT_11 => X"00000000002801E1A00000801C0202F40080000800007B00000302006E808000",
INIT_12 => X"0000007E00000607810000001E000087810000001E000081846282010A211AA0",
INIT_13 => X"00001BC00000740401E0400000070800340401E04000000780003404045D0010",
INIT_14 => X"01011740040000001F8000025010116C080000000085C80000C8100947008000",
INIT_15 => X"FF800C609C06D082000A03200806A040019481D4000000000801E0D00001001D",
INIT_16 => X"010040100401004010040100401004010060C040040C200950402090128057C3",
INIT_17 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_18 => X"0040100401004010040100401004010040100401004010040100401004010040",
INIT_19 => X"00000000000000000000000000001000802FFFFFFFFFFFFFFFFF810040100401",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(31),        -- Port A data input
DOA(0)   => data_read_a_hi_256(31),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(31),        -- Port B data input
DOB(0)   => data_read_b_hi_256(31),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_0_12 : RAMB16_S1_S1
generic map (
INIT_00 => X"ED39BA795990D275FB4A6E96ACC4731DEA4598B0AFB54867F6EE4618C3749803",
INIT_01 => X"8AA0047D8607944AC7DA180001ECA2444042106208408208C20022E9173734B3",
INIT_02 => X"1A7DDD79F9A73E6CCA7DAAF00001000008478020113D98E382FEDF333027C80F",
INIT_03 => X"75D341110C58F31110C58F32A208921F8051500147A0E4AB3493FB3A01EBE240",
INIT_04 => X"86424001531009B100425A97B2AA0001E03501D0A39C8F0078420001106D0C4C",
INIT_05 => X"BCC8CA2EBF03400700402BB20F00239E20341699198600000B08694B16434804",
INIT_06 => X"103FB860B2800161F8432200012DA185F80F24081C3C0707800E600056881308",
INIT_07 => X"B24197ABCDA467F9A73E6CCAFDC3870EEEEC44E2BDFE220094D03022210C011C",
INIT_08 => X"240581B5695EAA80262C080032BF07C7C1FC3F8E94F65B11555EAFFC1C306758",
INIT_09 => X"7E40000BEC004170040DB60017FED1CC0001045002984202003DB931192D60A5",
INIT_0A => X"120071411A74315881A28C141118000C5A85A60444210123820B43B40804674D",
INIT_0B => X"0820008E514045BB514F0106D1D8599581D3A958BC104A89215AC14C48898403",
INIT_0C => X"C261C01C48B1584A0CA3E2687A9A1E2687A9A1E2687A9A1E26870CD061343885",
INIT_0D => X"D274E93A758FA8683AC54B287522E10A74AF4AA59C568752662F5AC218000002",
INIT_0E => X"FF83C002783A0904231C70470C7E0B92800224008AE09FAD4BD48D1FC5D3A4E9",
INIT_0F => X"5BFF078004F075885DFBF7E15C06101C55E921F1F80FAB7FE0F0009E0E903EAD",
INIT_10 => X"F12E0380231F13978FF023FAFDBD9870380230F2D6081F56FFC1E0013C1D207D",
INIT_11 => X"DE7F263C0C8700125C0F8F3C43F1F10BBF7EFC61E01804E1E6C8F8FE807F67FB",
INIT_12 => X"02BE00017C17C1007E5E2E3081C5AC007E6F0E3081C5AC44418D65FE45DEE55B",
INIT_13 => X"61E0042786F103E9F01F9BC3C120C5A703E9F01F978B8C20666703E9F8A0FFED",
INIT_14 => X"FA7E283FFB414F80005F05F10FA7E283F78F6511C048278DCA174FF038FF15B4",
INIT_15 => X"0066A20B61692F293185D8D724E15D3FCC6B7C236FE0691B0700132C1F0EF880",
INIT_16 => X"3A4E93A4E93A4E93A4E93A4E93A4E93A4F942F92E9628540AD2A91442525A000",
INIT_17 => X"A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E9",
INIT_18 => X"4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93",
INIT_19 => X"55F3898E09B56C74DAB15D1CF13501AA495000000000000000003A4E93A4E93A",
INIT_1A => X"082082082082082082082082082082082082082082082082082084E41DC71C71",
INIT_1B => X"E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F82082",
INIT_1C => X"FFFFFFFFFFFFFFF94A5294A5294A5294A5294A52800003E1F0F87C3E1F0F87C3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"3060C183060C187FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"BDEBA0000000000000000000000000000000000000000000003060C183060C18",
INIT_28 => X"168ABA002E82145085155545F7AA975EFFFAABDE00FFAEBDFFF5D2EAAAAAF7AE",
INIT_29 => X"7FFFE10005542145557FD5545FF8000155087FC0155F7D168B55007BFDF45085",
INIT_2A => X"7FFC0010080017555555568AAAFFFFD7545AA8028A00A2802AABAFF8028BEF5D",
INIT_2B => X"FF842AABAA2AE95545FFD168ABAF7AEAAAAAA2FFFDF4500043FE105D2E954BAF",
INIT_2C => X"5007FD7400550415410002E974BA5D5168A00A2D142155005142010FFAE820AA",
INIT_2D => X"FFF780000BA007FE8AAAFF803FFFF5D2A821550000000BA007FD55FF5D7FC014",
INIT_2E => X"000AAFBEAA00007BFDFFF082EBDF455D5142000082E82145FFD17DFEFFFD168B",
INIT_2F => X"DFD75D2AA8A80EA8E2FE3F000000000000000000000000000000000000000000",
INIT_30 => X"68B551475FAF6D1C556F0AA1C24AABEA495FC716F002A975FFE3AA95E00EBAEB",
INIT_31 => X"42A0070071C50BAFEF1FAE0016D56A16D557BC257D415E0216FA3F1E8FC0145B",
INIT_32 => X"8010E004924874825D7FEAA85487FD24AFE3D02DAAAE12BD5545A2803AA00005",
INIT_33 => X"120155EA568E870BAEB8A05A2AEA8B50F55A2F150005A3A438BD04AFAB8F550A",
INIT_34 => X"545E055FFBE81D0BE8EA8A3AA05A2A5504001C74BA42A1571E8028E3DB7816D0",
INIT_35 => X"A5C7E3DFFFE90B45B47ABA497A82FFAFD2A82485FD2415A105C21451ED42A002",
INIT_36 => X"00000000000000000000B55EAAA100AA1D0F6F480B6A555A2A57A002A3D5FDB6",
INIT_37 => X"5EFAAAAB5E1AF3AABFF45592E88A0AFE80A8B0A0000000000000000000000000",
INIT_38 => X"65F520EBE9EF67D7BEA1FD5D556ABEF5D557FEBA55022A3F70C6B405F4D2AE97",
INIT_39 => X"C114728007521170821CE0FDE69411A8DED57CE1055555E5F58EFFC01FE2CACB",
INIT_3A => X"42341D5DEEBEF55080034E0A592A4AD0079C75D6070CC5CBB0280C029ABAA3EB",
INIT_3B => X"7F353AAF6C77F7F20D968BF57812A95E02A2AAB5EB0F280800EFAEE9F5D18F31",
INIT_3C => X"C91565455C141E41887D58AC448B69C30E02116220415A9540AA854140A0A204",
INIT_3D => X"DE6BE93172D7D625B556EEAB157ABEBE1B4D792A4AD1183454180DD3FDCAAAB7",
INIT_3E => X"F0000001FF0000001FF0000001FF0000001FF01EABC4B8014174FF7DA80F52FE",
INIT_3F => X"FF0000001FF0000001FF0000001FF0000001FF0000001FF0000001FF0000001F")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(0),               -- Port A write enable input
DIA(0)   => data_write_a(0),        -- Port A data input
DOA(0)   => data_read_a_lo_512(0),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(0),               -- Port B write enable input
DIB(0)   => data_write_b(0),        -- Port B data input
DOB(0)   => data_read_b_lo_512(0),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_1_12 : RAMB16_S1_S1
generic map (
INIT_00 => X"212C001411984004084D000508C53810A03D1450E839B003342114428A000803",
INIT_01 => X"00000019400B100A8196000000CC004400400002000000000000028001340000",
INIT_02 => X"052137AE8031800C0044009000000000061800001CD4019802AD04CCCFC20004",
INIT_03 => X"04514108C60C21008C6042108400000201440020505100000043C30E10E9F000",
INIT_04 => X"02104001011DEFE088805681920000008000004001900800004002108C280008",
INIT_05 => X"040002340105000200000000080001900010000108040000000008411600401C",
INIT_06 => X"1034001042800808201000000001000820020000102000040000000000800180",
INIT_07 => X"64BF81A15EDFDE8031800C00843060C19E030022103600000450020800040004",
INIT_08 => X"00008004691687AA840008000090248CC84E000046000311555521F183060AC5",
INIT_09 => X"0820800D08100171000DB000154440C800400500000852020011200201012021",
INIT_0A => X"02000040001000880A2A04445004000102002041000001008208001440004140",
INIT_0B => X"4820018A1140440078050040511000102000A008183000010002404400000000",
INIT_0C => X"1000C80008000C030030880C2A030A00C28030A80C2A030A00C28018D4061401",
INIT_0D => X"10040802050080200284401C0022880F009E08008205C0020118088018000000",
INIT_0E => X"0F03C00280000000420860C60C0C0B92C0000000004000010042000040102008",
INIT_0F => X"001E078005000108400005E11C0610000000288058000003C0F000A000100000",
INIT_10 => X"F10E0380000000C202300000008D187038000000480800000781E00140002000",
INIT_11 => X"806302380C870010000004400100110800007861E0180000000C400680000001",
INIT_12 => X"023E00000000018000580C308000050000610C30800005000215006800000101",
INIT_13 => X"61E0000000018100B0001843812000014100B00016030C20000141002880026D",
INIT_14 => X"400A20009B404F80000000018400A20044096111C04000000304026000501580",
INIT_15 => X"0046820040082300218450C2800010094000482141E060190700100000002200",
INIT_16 => X"020080200802008020080200802008020080008008600500A82A1100A8000000",
INIT_17 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_18 => X"0080200802008020080200802008020080200802008020080200802008020080",
INIT_19 => X"81328A46BABEFC54A0810C7452B4428A14000000000000000000020080200802",
INIT_1A => X"AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA28A28A28A28A2A8218D2C0C924925",
INIT_1B => X"E974BA5D2E974BA5D2E974BA5D2E974BA5D2E975BADD6EB75BADD6EB75BAAAAA",
INIT_1C => X"FFFFFFFFFFFFFFFD8C6318C6318C6318C6318C63000002E974BA5D2E974BA5D2",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"70E1C3870E1C387FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"5555500000000000000000000000000000000000000000000070E1C3870E1C38",
INIT_28 => X"EBDF455D2EAABEFF7FFE8BFF5D0002155557FFFFFF007FC21EFA2FFD74AAAAD5",
INIT_29 => X"AA95400552AAAABAFFD1574105D7FD75FFAAAA800AAF7AA974BAFFFBE8B45F7A",
INIT_2A => X"0517DF555D2EAAA1055000015500557DF45AAD1400BAA2AE801550051555EFF7",
INIT_2B => X"FFD540155557FD5400F78028BFFFFFBEAB55F780020AAAA80020AA082EAAB550",
INIT_2C => X"AFF842ABEF5D517DF55552A974AAF7AE820AA0851574BAA2D1574AA5D7BFDEBA",
INIT_2D => X"EFAAD1575EF557FFFE10557FFFFFFFFD56AAAAFFFFD7555AAD168B45AAAEAAAB",
INIT_2E => X"0005D7FFDF4500043FE105D2E954BAF7AE80010082A97410557FEABFFAAFBE8B",
INIT_2F => X"51C7A2FBD5490BFD1C056A000000000000000000000000000000000000000000",
INIT_30 => X"974BAF7FFEFB45FFAABDF55492AA8BC2EBDFEAF7F1F840017D4975D2FEF147FC",
INIT_31 => X"080BEF495FC71D54124924385FAAA8AAAE3D145410F7F1D55D71C002DABAEBAA",
INIT_32 => X"002D082082AB8B6DBEDB7DF7F540E2AE85028B40155145F7AF6DBED5450AA1C2",
INIT_33 => X"78E021FF1471FDEAAFFD56F16D5571D2E28E38E0216FA2D1E8E80140F45082B4",
INIT_34 => X"A2DA3FB7DAAD4AAAAF487BC70BFA97F7AF6D417E92482BF84020BA495557E3FF",
INIT_35 => X"55554ADBD7A2FFC7BEFF6FFD7FC7002FD74951D71EDFFABFD16FAAAE92BD5545",
INIT_36 => X"00000000000000000000547AB8F550A8010E00492487482FFFE82A85EBAE2FFC",
INIT_37 => X"1EF005162BEF047FD5545AAFBF7400FBF9424F70000000000000000000000000",
INIT_38 => X"714F8338AAAA1D0AE974AAF7FFFDF55F7AABFF55082CA8B4DF6C1E8F5E540002",
INIT_39 => X"EABEF75550ACBB7582225FF5843404547184164AA5D2EBEEB0A2D555410D3555",
INIT_3A => X"FEAAEB083BC1000FF8409000512AEABFFDF79DCBF755962010BDCBBC21455D7F",
INIT_3B => X"801F8BA0C57740BDAA0688E5405D57D412F7D55F5E50C7F401BAAE8403CF5A3F",
INIT_3C => X"5D16BABAA3EBC3157ABD5FFE55F2AA9FEAFDF7F431A9F7FFE81FF013A8001AFF",
INIT_3D => X"FB863550229BCABEB7DA403FFFDA2FBF7FED2C7F955445079E280A00C56145EF",
INIT_3E => X"0000000000000000000000000000000000000596EBEF55080034E0A592A4AD00",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(0),               -- Port A write enable input
DIA(0)   => data_write_a(1),        -- Port A data input
DOA(0)   => data_read_a_lo_512(1),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(0),               -- Port B write enable input
DIB(0)   => data_write_b(1),        -- Port B data input
DOB(0)   => data_read_b_lo_512(1),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_2_12 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10E006600180111284380310006289800480032283E000A34301002001A0817",
INIT_01 => X"0005A00810790848048044A54E404350404000720885800802000906E4910200",
INIT_02 => X"407004208400408044C600C50AA055254010541A110222841200000002402544",
INIT_03 => X"0600011004182401004102408C28414043101000408118000145840440F5C415",
INIT_04 => X"5035855703A2900A000CD3088400F40688C9844409060850925E58A4081A0221",
INIT_05 => X"0200840D1021A15AC50494894850890540D1E12020C6E510818500440A280090",
INIT_06 => X"113044094002801020440090A8011A1224AB9380552102442884882A20004097",
INIT_07 => X"000100880004428400408044860000008C022402102100AA40004404B5075460",
INIT_08 => X"15C23440408C862A2A12382A8A5244145048C06085008010141521F000001240",
INIT_09 => X"400582B9033AA0E7AA4110B0506744810554542450694E710A836188C2C00222",
INIT_0A => X"443518360012C2210B020414109130A28038188096A06B8C120CA440A9C00802",
INIT_0B => X"1345E53300EC68005605002964AF222A5704004D080211121C80024200821780",
INIT_0C => X"181080C1110C882202211488452213C88472213C88472213488441109A442231",
INIT_0D => X"008204440210091341208041000810C00000300220201800A908000038AD0284",
INIT_0E => X"00040002804180300E88D28D206A40000554815500481440300000C44A081100",
INIT_0F => X"000008000500828700000000010000000002380000A00000010000A010050000",
INIT_10 => X"00010000000004CA000214000000020000000000684280000002000140200500",
INIT_11 => X"000000000020000000000442100002840000000800000000010C000026000000",
INIT_12 => X"00000000000805A4800000000000152300000000000015801272000100210020",
INIT_13 => X"000000000101C00000C000000000000940000120000000000009600004050000",
INIT_14 => X"0000130000000000000002018000106000000000000000002380000141000000",
INIT_15 => X"55000190000000000002000280000000011080C0000000000000000000002310",
INIT_16 => X"40902409064190641906419024090244902A9003004800415120D4A190804241",
INIT_17 => X"0900409004090641906419064190240902409024090641906419064190240902",
INIT_18 => X"9044090040900409004190441904419044090040900409004190441904419044",
INIT_19 => X"75960040138D70C030B51C50C7D100A2052F81F81F83F03F03F0419044190441",
INIT_1A => X"0410410410410410410410410410410410410410410410410248602081659659",
INIT_1B => X"5128944A25128944A25128944A25128944A25128944A25128944A25128941041",
INIT_1C => X"FFFFFFFFFFFFFFFE1084210842108421084210843FFF825128944A25128944A2",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"7FD5FF555815607FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"2AA000000000000000000000000000000000000000000000007FD5FF55581560",
INIT_28 => X"FC21EFA2FFD75EFAA8415410AA8415555087BFFF55A2AA800BAFFAE954000800",
INIT_29 => X"84155EFA2AEBDEAAA2FBEAABA5D7FE8B555551421455D0002145552EBFEBA007",
INIT_2A => X"2AEBDF555D2E954BAA2AA974BAFFFFE8B45552EBDF45FFAEAABFFF7FFE8B55F7",
INIT_2B => X"AAAAAAAAAFFD1574105D7FFFF555D2AAAAAA5D2E820BAA2FBEAB5555557DF55A",
INIT_2C => X"50055575EFFF84021555D043DEAA5D04021EF557FC21FFAA8428BFFAAAA954AA",
INIT_2D => X"10085568A00FF80175FFA2D17DFEFF7800215500557DF55AA80001FFAA800015",
INIT_2E => X"0005D00020AAAA80020AA082EAAB5500517DF555D042AA10A284154005D00154",
INIT_2F => X"00AAFFAA9543A080038A2A000000000000000000000000000000000000000000",
INIT_30 => X"0017D5D20B8EAA007FC51C7A2FBD55D2BE800042AFE8E1557D0075D2F45BEAA8",
INIT_31 => X"AA8BC7EBDFEAFEFFD00105FFBC20BDEAAA2FBF8AAA557BE8B6D5D5FFABEF4904",
INIT_32 => X"FFEFB6D555578F7DB6A0BDF7D480E174BFA02A974BAF7F5EFB455D2ABDF55492",
INIT_33 => X"ED1FDE90E3A497492B6AAADAAAE3D155E105571D55D71C002DABA5524820BAB6",
INIT_34 => X"BE8F401D7B6A0001470155C51D0092A071555D5E3AE821D00001FF0871C016DB",
INIT_35 => X"5BE8555400550A38428007FED000E3DA3DFD5E3DFFFBD5A38A021551C5F7AF6D",
INIT_36 => X"00000000000000000000410F45082B4002D082082AB8B6D1C5B7DF7FF78E075C",
INIT_37 => X"5EF005560B55F7AA800AAF7AA954AA00042AAA20000000000000000000000000",
INIT_38 => X"ABEF057D68F5F5A00021EF55042AAAA007FD5555AAFBD7545FBB8020A3F7AE97",
INIT_39 => X"7DF55D7AABFF5428ACA8F45A6C1E8F5EFF84165EFF7802BAB0A2FFEAABA557BE",
INIT_3A => X"CA8AA80800020AAF7FBFFFEF04552ABFFFF841FFE75CA882108202E974AAF7D5",
INIT_3B => X"00151FF0C57401E5F3D1E00A1A884174A8FFAEBFEB0A2D55541051555694F002",
INIT_3C => X"2AA801455D7FE8BFFF680800FFF7AAA155F595542455512A975455D3AA8A0055",
INIT_3D => X"5D79FCAF774AE005BE7895554005D2A8A0B882FFFFE10AAAAAB755A66B6AF56A",
INIT_3E => X"00000000000000000000000000000000000000C3BC1000FF8409000512AEABFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(0),               -- Port A write enable input
DIA(0)   => data_write_a(2),        -- Port A data input
DOA(0)   => data_read_a_lo_512(2),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(0),               -- Port B write enable input
DIB(0)   => data_write_b(2),        -- Port B data input
DOB(0)   => data_read_b_lo_512(2),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_3_12 : RAMB16_S1_S1
generic map (
INIT_00 => X"210C00A20020000108430020001600B8156021104940741B3530400E02B92203",
INIT_01 => X"014C9BCA58B1296D24A402C992500B69404040028804A0080A000416A8D90A08",
INIT_02 => X"C12026A484318004404405C9C66E331352180D468B8203980300204442E02B34",
INIT_03 => X"04000748D60D24648D60524C88804D0215011020D15018148040C10A70E1D58C",
INIT_04 => X"18283333240FE41244187308C9104D70944852640901083801750EB0A418C220",
INIT_05 => X"0613142D01912CC2A1B4140528348900C612A104201C689044340ED413A07649",
INIT_06 => X"119000034019881822104C5E68035250A222829710A0A02C18C01A9920842413",
INIT_07 => X"402F00AB0016CA0431800444841020509D038B021230C1990001C644C8273200",
INIT_08 => X"16905000408482088290E8E64010248C4A5AA840C2000110001521F0810A92E7",
INIT_09 => X"0003CE6581BD016342A951AB146C4480530C3B2A8088D3542651670200C1826A",
INIT_0A => X"00735D36209A8A20020894004284B660821030C8990467401218004041020002",
INIT_0B => X"512445B740457154562F957CC08B00093700080D0A4851001D8302D20A0A1530",
INIT_0C => X"00508650008008021021A40861021840869021A408610218C0869810D6043095",
INIT_0D => X"1C8508438450801043A08090380A8834207007022209038080190000999C8F84",
INIT_0E => X"000400200000C0002A48A206204C4205F3304B33004C0041006240140A1C310A",
INIT_0F => X"0000080040000083800400000100000000008400018040000100080000510100",
INIT_10 => X"0001000000000800000244040000020000000100002A0080000200100000A702",
INIT_11 => X"000000000020000000200000080002C000800008000000000022000006808000",
INIT_12 => X"0000000000000A2281000000000040A3810000000000402001400000022002A0",
INIT_13 => X"000000000004200001C0400000000010200001C0400000000010000004490010",
INIT_14 => X"0001070004000000000000060000104C08000000000000001000000903008000",
INIT_15 => X"CC004050CA0C00020220200070040000010401C4000000000000000000100008",
INIT_16 => X"4310E4310A4210A4210A4210A4210A4210A8D0830A68010001B4DA881048061C",
INIT_17 => X"21084290A4210A4210A4210A4210A4210A4210A4210E4310E4310E4310E4310E",
INIT_18 => X"90A421084290A421084390E4310C4390E4310C4390E4310C4290A421084290A4",
INIT_19 => X"015303C0C78C706428A14C586291000A044001FFE000003FFC004290A4210842",
INIT_1A => X"2492492492492492492492492492492492410410410410412821600001249249",
INIT_1B => X"51A8D46A351A8D46A351A8D46A351A8D46A351A9D4EA753A9D4EA753A9D49249",
INIT_1C => X"FFFFFFFFFFFFFFFC00000000000000000000000038F56351A8D46A351A8D46A3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"55AB02055AB0207FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"420000000000000000000000000000000000000000000000007FFFAB57FFFAB5",
INIT_28 => X"A800BAFFAE9554508002AA00AA843DF55FFAA955EFA2D168B55557BEAA000055",
INIT_29 => X"002AB55AAAA955EF005568A00087BE8BFFA2D155410AA8415555087BFFF55A2A",
INIT_2A => X"AAABFF5508003FF555D0002145552ABFEBA007FC21EF007FD75FFAA841541008",
INIT_2B => X"082EBDEAAA2FBEAABA5D7FC0155005168B455D042AB45F7FFD741000042AA10A",
INIT_2C => X"FF7FBEAB55F7AABDEBA5D7FC2010A2D1575FFF7AA975555D2E80145F78415545",
INIT_2D => X"EF5555554AA087BC01FFFFAAAAB55552A954BAFFFFE8B55552EBDE00F7AEAABF",
INIT_2E => X"000082E820BAA2FBEAB5555557DF55A2AEBDF555D2E954BA002EAAABA002A821",
INIT_2F => X"FB7D5D7FEAA3808554203A000000000000000000000000000000000000000000",
INIT_30 => X"1557D1475FAF45BEAA800AAFFAA95578080038A2AA28E3AF55E3A0BA5D7AADB6",
INIT_31 => X"BD55D7BE80004AA1E8E2AB55B6A0925D7085F6AA10087FEABD7AAD57AEBAB68E",
INIT_32 => X"F5D0438140E2FA38B6AEBFF6D1D04AAFFA41040017D5D20B8EAA007FC51C7A2F",
INIT_33 => X"D0A901FFFF801557D1C20B8EAAA2FBE80AA557BE8B6D5D5FFABEF49002FB55FF",
INIT_34 => X"5D20BDE00EBAAA8BC7EBDFEAFEFAB8ABAE925D21C7010EADB525D7FFAE975C75",
INIT_35 => X"F002EADA921420871D74971D24820875C21D5EB8AA8FFF012A954BAFFF5EFB45",
INIT_36 => X"000000000000000000001C24820BAB6FFEFB6D555578F7DB6A0BDF7DEB8E125F",
INIT_37 => X"B55A28408145AAFFFFFFF5D7FEAABA0051400A20000000000000000000000000",
INIT_38 => X"AB55FAD568AA2AFAE975EF555168B55F7AA800BAF7AA955EF00042AAA2A2AEAA",
INIT_39 => X"2AAAA007FD55558A7BD7145FBB8020A35D2ABEF55F7800015F087FEAA00007FE",
INIT_3A => X"968F575D003FF55F7D5420BA5D2ABFEAAF7AE9DFF759A82AEF70800021EF5504",
INIT_3B => X"FFD5145FBAC9755F05040255FFD84175EF55002AAB0A2FFEAABA557BEA3EF057",
INIT_3C => X"82E974AAF7D57DF45552A3FF10AA8429F45A7D5EAF5FFBAEAAA10554155400AA",
INIT_3D => X"FF843FFE77C80825BC052ABFE10550415557085540000005156155FE90A8F5C0",
INIT_3E => X"00000000000000000000000000000000000005500020AAF7FBFFFEF04552ABFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(0),               -- Port A write enable input
DIA(0)   => data_write_a(3),        -- Port A data input
DOA(0)   => data_read_a_lo_512(3),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(0),               -- Port B write enable input
DIB(0)   => data_write_b(3),        -- Port B data input
DOB(0)   => data_read_b_lo_512(3),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_4_12 : RAMB16_S1_S1
generic map (
INIT_00 => X"A108400020612C80284210081034849800A00030300004833522C82D04A16002",
INIT_01 => X"2043998A1839284D1CA0650E1E504368403008418984014902030806A0D10200",
INIT_02 => X"C120042200000000044441CE01E80F00A49043118680008002000000026208E4",
INIT_03 => X"040001020019200020011209CC0164C060000000690111040144800042F5C403",
INIT_04 => X"7029AF0F81A00010CCA47700CC513CAC0D0B8E02010740E19754080108988021",
INIT_05 => X"02139405007133C0712244CD20F20105D583000020E9892201D304D42A9835E1",
INIT_06 => X"9190440300078002014405D9EE814C0284A883B6D7038AE079059B7800048092",
INIT_07 => X"000100AA0004408000000004840400008D200102503000782000C00C8025C000",
INIT_08 => X"00728A00408403220811991E02120C044058080004000001101121F220000260",
INIT_09 => X"811001E1185B38AD23C3707AD46440818F3CF80EC423CA7D01D123C80200816A",
INIT_0A => X"45810810A01B40216361056D6150F41200280001900439001FD8A00041400000",
INIT_0B => X"11FC88076266E800D605402962A820211500024808010512C40106D222223B14",
INIT_0C => X"0408804116040B02C02C500B0C02C100B0C02C100B0402C300B0401618058611",
INIT_0D => X"040200050200501301208482200D00D0A0408402C4282200A84800009B878680",
INIT_0E => X"00000020000100024AC88300300060090F0D830F00025400300204D018000804",
INIT_0F => X"8000000040000206A2000800000000000000950002E010000000080000588040",
INIT_10 => X"0000000000000808000554000200000000000100006D0020000000100000BB00",
INIT_11 => X"0000400000000000002000001A0002504001000000000000002280000D800800",
INIT_12 => X"0800000000000E2C802000000000408D801000000000408012440000200110A0",
INIT_13 => X"000000000004680003A0040000000010280003800800000000102800000B0000",
INIT_14 => X"000005C0002000000000000620000158000010000000000010A0000B00000200",
INIT_15 => X"C30146200400104002602600400000000294004000000004000000000010001A",
INIT_16 => X"0080200000008020000000802000000080080000004090014134DA101288C6DB",
INIT_17 => X"0802000000000401806010040180601004018060100000802000000080200000",
INIT_18 => X"8060180601004010040080200802000000000000802008020000000000008020",
INIT_19 => X"C0A28A063807E0500014063450404882846FFE000003FFC00000010040100401",
INIT_1A => X"AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA28A28A28A28A2934C8D0CCD145144",
INIT_1B => X"68341A0D068341A0D068341A0D068341A0D068351A8D46A351A8D46A351AAAAA",
INIT_1C => X"FFFFFFFFFFFFFFFC0000000000000000000000001FE32068341A0D068341A0D0",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"408102040810207FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"800AA00000000000000000000000000000000000000000000040810204081020",
INIT_28 => X"168B55557BEAB4500554200000557FE10FFFBEAA10007FD7410FFAA97555082A",
INIT_29 => X"55574105D2A800AA00043FEBA5D7FEAA00007BE8AAAAA843DF55FFAA955EFA2D",
INIT_2A => X"57BC00AAA2FFEAAAAAA8415555087BFFF55A2AA800BAFFAE9555508002AA0000",
INIT_2B => X"A2AA955EF005568A00087BE8BFFA2D17DE1000517FE10AAAAA8AAA002E975455",
INIT_2C => X"FAA8417410A2D140000F7FBC2010A2D157400AAAE974AAAAAA974BA08002AB55",
INIT_2D => X"EFA2AABDEAA087BEAAAAA2FBD54BA080002145552ABFEAA007FC21EF007FD75F",
INIT_2E => X"00055042AB45F7FFD741000042AA10AAAABFF5508003FF55F7D568A00552EA8B",
INIT_2F => X"5400F7A49057D0824850B8000000000000000000000000000000000000000000",
INIT_30 => X"3AF55F7A0925D7AADB6FB7D5D7FEAB7808554203A145178E00FFFBE8A101475D",
INIT_31 => X"A9557D080038AAA145157428492E8008200043FE925571EFA380871C7028A28E",
INIT_32 => X"AEA8A9200249056D4175C5092AAF5FDA38BE8E1557D1475FAF45BEAA800AAFFA",
INIT_33 => X"AA4954281C0E2FB55B6A0925D7085F6AA10087FEABD7AAD57AEBA08517DE00AA",
INIT_34 => X"007FC51C7007BD55D7BE80004AAFEDB42028EBFBC2028BED152438AAA092492A",
INIT_35 => X"AF7DF6AA00412EAABFFAA803DEBA0875EDA80BEF1C743840040017D5520B8EAA",
INIT_36 => X"0000000000000000000041002FB55FFF5D0438140E2FA38B6AEBFF6DBE84AAEB",
INIT_37 => X"A00FFFFEAA105D5155410FF84021EF0800154B20000000000000000000000000",
INIT_38 => X"DEBA0851574B2AAAEAAB55F78400145AAFFFFFEF5D7FEABFF0051400A25D5568",
INIT_39 => X"68B55F7AA800BAF7AA955EF00042AAA25555410BA082E8201000043FE005D517",
INIT_3A => X"568AA200557DE00AAAAAAA000804001FF005575408AA557FEB2FFAE975EF5551",
INIT_3B => X"D1550AAAA8002010F2AC154B25F2ABFF55F7800015F087FEAA00007FEAB55FAD",
INIT_3C => X"800021EF55042AAAA007FD5555087BD6145FAAC000A2A6FBC00BAAAFBC00BAF7",
INIT_3D => X"F7AEBDFF779A82AA43F7FBE8A00082EA8BFFAA843FEBA08517DE00F3F9574B30",
INIT_3E => X"000000000000000000000000000000000000008003FF55F7D5420BA5D2ABFEAA",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(0),               -- Port A write enable input
DIA(0)   => data_write_a(4),        -- Port A data input
DOA(0)   => data_read_a_lo_512(4),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(0),               -- Port B write enable input
DIB(0)   => data_write_b(4),        -- Port B data input
DOB(0)   => data_read_b_lo_512(4),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_5_12 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50DF4A0791B3FCB694379283C81FD996A091832102004A336A20E03C040C002",
INIT_01 => X"805FBDC69830A84D5C6A60000C34C26841280A00084000C8C212892EEAD53235",
INIT_02 => X"3B2026B578918E640A4F01CF8011FF0002080000082CA9998276DF7772C7C80D",
INIT_03 => X"37134108420D700084205702A4008A1D9100002171C0E0051554D93A11F5D140",
INIT_04 => X"8A41A0FC03A56DA000425A819410E3816C086198A388B702A8CA1210844A0C4C",
INIT_05 => X"B1808A062E8BC835F5E84532D708238A282F00A9291224800A2861490343082C",
INIT_06 => X"903FB8483A90581859050424100940825C6184401CDC451B860A6507160C4100",
INIT_07 => X"D26F068BCC96CDF8918E640E96D1A3469D6300E2FFEA27F8E4D23248130E259C",
INIT_08 => X"0BFA82E568442B2A082C0A7E3014250D49DA37A2420619000002AFF48D1222E5",
INIT_09 => X"3F005001E40969289429360416DCD1C46083030604B1CA20C03DF83B0A2C60A5",
INIT_0A => X"14613C71005A10492B888120288F480D58858449026145B3830F449449062B4F",
INIT_0B => X"11AC04934AC648BFD727C031E64170A137D5AA5C3E4B0F8A3C58C34C002290E3",
INIT_0C => X"CA29C6CC50384B6AC6AC86AB31AACA6AB39AAC86AB39AACA6AB3055643559C31",
INIT_0D => X"C673E33CF28F38603855401985228A0614BD30A0A2819852011E5AC2B87F9182",
INIT_0E => X"FF87C002F87A803E460B2516510CA594FF0044FFA4B08BAC4BB2CD0F09CF84E3",
INIT_0F => X"0DFF0F8005F0F5100DFFF5E15D06101C55EB29F1E00BE53FE1F000BE1E802F94",
INIT_10 => X"F12F0380231F17D78FC029FFF58D9A70380230F2FE0017C37FC3E0017C3D005F",
INIT_11 => X"FC7F023C0CA700125C0F8F7E43F1F001BFFE7C69E01804E1E7CCF8FC003FF5F1",
INIT_12 => X"023E00017C1FC1A4BFD82C3081C5BD27BFE30C3081C5BD00C02365D645CEEF5B",
INIT_13 => X"61E0042787F181E9C1EFD8CB8120C5AF41E9C18FD60F0C20666F41E9F009FFFD",
INIT_14 => X"7A7C077FFF404F80005F07F187A7D14BFFC96111C048278DEB074F9930FF9D80",
INIT_15 => X"C064014B8B652E2B3120C81284641D3E8DBF7D636FE860190700132C1F0EFB80",
INIT_16 => X"38CE1384E3384E338CE138CE1384E33C4E3ECE32E128882551349A1CBAA44103",
INIT_17 => X"84E3384E3384E3384E338CE138CE1384E3384E338CE138CE1384E3384E338CE1",
INIT_18 => X"CE138CE138CE138CE1384E3384E3384E3384E338CE138CE138CE138CE1384E33",
INIT_19 => X"F5E5BB4E7F7B9DB7FF3A1B6DB7E8410A8C000000000000000000384E3384E338",
INIT_1A => X"BEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEF9F7CFDFDDCF3CF3D",
INIT_1B => X"BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEFBEF",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000001711C7BBDDEEF77BBDDEEF77",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"FDFFF00000000000000000000000000000000000000000000080000000000000",
INIT_28 => X"FD7410FFAA97410082A800AAAAAE955450055421FFFFFBC0010AAD5574BA557F",
INIT_29 => X"7FD74000055574BA5D7FD7555A2D5575EF55517FF5500557FE10FFFBEAA10007",
INIT_2A => X"0002AABA5D2ABFFFFAA843DF55FFAA955EFA2D168B55557BEAB5500554200000",
INIT_2B => X"5D2A800AA00043FEBA5D7FEAA00007BC00AAAAAEBDF45A28428B45FFD168BFF0",
INIT_2C => X"5080028A00A2FFFDE00F7D57FEBAFF80174BAAAD1555EF555555555005557410",
INIT_2D => X"BA5D2E821FFA2D5554BA557BD75FFAA8415555087BFFF55A2AA800BAFFAE9555",
INIT_2E => X"00000517FE10AAAAA8AAA002E97545557BC00AAA2FFEAAAA082A97545F7D5420",
INIT_2F => X"7010BEDF524AA5571FDFEF000000000000000000000000000000000000000000",
INIT_30 => X"78E00EBFBE8A101475D5400F7A49043D0824850B8A2AE9756D145B401FFFFFFC",
INIT_31 => X"FEAB7D0855420BA1471D74380851524BA5571D757DB6D5525EF555178F6D1451",
INIT_32 => X"8A28B6DEBDF6DBEF1C0A28AAA5524BFFFFA28E3AF55F7A0925D7AADB6FB7D5D7",
INIT_33 => X"5555057D145152428492E8008200043FE925571EFA380871C7028B6AEBDF45B6",
INIT_34 => X"BEAA800AAFFAA9557D080038AAAA2FBF8E10EBD578EAAFF8415482BED1555EF5",
INIT_35 => X"81C209256DFFDF420BA552A821FFB6DF574A85575C55EFBE8E1557D1475FAF45",
INIT_36 => X"0000000000000000000008517DE00AAAEA8A9200249056D4175C50920875FDA3",
INIT_37 => X"5FF5D7BC21EFF7FBD7400F7FBC00BA55557DFF70000000000000000000000000",
INIT_38 => X"01FF5D5568BE7555568A00AAFFEAA105D5155410FF84020AA0800154B2AAAA97",
INIT_39 => X"00145AAFFFFFEF5D7FEABFF0051400A25551554BA0051400BA5551575EFF7D14",
INIT_3A => X"1574B2FFAABFF45FFAAAABFFAAFFFDFFF552EA8AAA55043DFF7AAAEAAB55F784",
INIT_3B => X"8002410FFD5575EF5555421E75555400BA082E8201000043FE005D517DEBA085",
INIT_3C => X"FAE975EF555168B55F7AA800BAF7AA955EF00002AAA2A2FBE8A00A2D16AAAAFF",
INIT_3D => X"0055554088A557FEB25D00021FFFFFFC00BA552A821EFFFFFD74BA5D51575F7F",
INIT_3E => X"000000000000000000000000000000000000000557DE00AAAAAAA000804001FF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(0),               -- Port A write enable input
DIA(0)   => data_write_a(5),        -- Port A data input
DOA(0)   => data_read_a_lo_512(5),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(0),               -- Port B write enable input
DIB(0)   => data_write_b(5),        -- Port B data input
DOB(0)   => data_read_b_lo_512(5),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_6_12 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10800B0061A01002840002C03002818000402322520070B313301C4389B2082",
INIT_01 => X"250041CA3839684D18A160000C52426841000000090800090210080008110200",
INIT_02 => X"0020042080010000044654C0000C008010000000001020900200200002620814",
INIT_03 => X"060881021088200021080200E4000A0891000020610111500104C00000F14400",
INIT_04 => X"0880000100000002000052288144004281C050400100280000C8100000080001",
INIT_05 => X"928080840001100A08009000280201000850E022401400002028214043410820",
INIT_06 => X"10100518090012122100C808049310002040000410A0001400000200120840D2",
INIT_07 => X"000100800004400001000000860408108C22000A502010074120044800040001",
INIT_08 => X"50000040D0C4E2088003FD01C01004044058082004000000000121F020408244",
INIT_09 => X"00BF17E9001205A5204911F814444080400100020000D200DFD16400C2A40AA0",
INIT_0A => X"04611C17849000022862A1596C8B5DF04834948900000100220C244840000880",
INIT_0B => X"03AD0413424E4044D665C070C22602291504400D084915020448114080201000",
INIT_0C => X"5E08864011088B22D22C008B0022C408B1022C208B0822C608B1111600458010",
INIT_0D => X"4251A12CD28A300429688001000800000020280204001000A00804309A002182",
INIT_0E => X"0000000280402400420800000000006200FC10002442042429324294014E8CA7",
INIT_0F => X"A40000000500800840000800000000000002280018001480000000A010100052",
INIT_10 => X"00000000000004C2003000010240000000000000680800290000000140202000",
INIT_11 => X"2000C0000000000000000442000001080001000000000000010C000280001804",
INIT_12 => X"08000000000801C300A010000000156000902000000015101200002800000000",
INIT_13 => X"000000000101800038002408000000094000386028040000000940000ED40000",
INIT_14 => X"0003B000002000000000020180002A24005010000000000023000060C7000A40",
INIT_15 => X"3F0280090321000040A410C28108000160008094000810040000000000002300",
INIT_16 => X"284A5284A728CA5284A528CA728CA52C4A5A0A32A300940101349A0408240818",
INIT_17 => X"9CA1294A329CA5284A728CA7284A5284A728CA5284A528CA728CA5284A728CA7",
INIT_18 => X"CA3294A129CA3294A129CA1294A329CA1294A3294A129CA3294A129CA3294A32",
INIT_19 => X"F5F78BCE7F8FF0F4FA955F7CF7F40A80145D55555556AAAAAAAAA94A329CA129",
INIT_1A => X"8E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E39B6CEDECDDF7DF7D",
INIT_1B => X"F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE38E3",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000001A1A33F9FCFE7F3F9FCFE7F3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"555FF00000000000000000000000000000000000000000000080000000000000",
INIT_28 => X"BC0010AAD5574BA557FFDFFF087BFDF45F7AA974AAAAAA97555F784174BAF7D5",
INIT_29 => X"515555508043FE00F7AA97555A2FBD7410AA8428AAAAAAE955450055421FFFFF",
INIT_2A => X"7D1575EFFFAA9555500557FE10FFFBEAA10007FD7410FFAA97400082A800AA08",
INIT_2B => X"0055574BA5D7FD7555A2D5575EF55517FF55A2AA97400552AAAB45082E80155F",
INIT_2C => X"500554200000003DE10FFD5401FFF7AAA8A10082EAAB45A2FFC2000007FD7400",
INIT_2D => X"10AA803FE105D516AABAFF843FFFFAA843DF55FFAA955EFA2D168B55557BEAB5",
INIT_2E => X"000AAAEBDF45A28428B45FFD168BFF00002AABA5D2ABFFFF087BD5545007BFDE",
INIT_2F => X"256DEB84104BAFFD1525FF000000000000000000000000000000000000000000",
INIT_30 => X"9756D145B401FFFFFFC7010BEDF524AA5571FDFEF1C7BFFF55FFA095482B6A49",
INIT_31 => X"4904380824850381C5B5057D1C003DE28F7A49057DAAF5D2428A2842AAAAA2AE",
INIT_32 => X"2AAFB451C2A8017DE3DF525FFFFA49756D145178E00EBFBE8A101475D5400F7A",
INIT_33 => X"2F1C50381471D74380851524BA5571D757DB6D5525EF555178F6DAAA49542841",
INIT_34 => X"AADB6FB7D5D7FEAB7D0855420BA1C0E3FE00E3DB471EFE3AAAAA00082EA8B6DA",
INIT_35 => X"F1C7BD057D1C71FFE10A28038E1049516AAB8FF8428FEFA28E3AF55F7A0925D7",
INIT_36 => X"00000000000000000000B6AEBDF45B68A28B6DEBDF6DBEF1C0A28AAA5524BFFF",
INIT_37 => X"F55F78017400F780001FFAA84000AAFFD1401E70000000000000000000000000",
INIT_38 => X"20BAAA8428AA2AAAA975FF5D7BC21EFF7FBD7400F7FBC00BA55557DFF7557BFD",
INIT_39 => X"EAA105D5155410FF84020AA0800154B2557FC01EF55043FEAAFF80021EFA2D14",
INIT_3A => X"568BE7AA80174AA082ABDF555D2A821EFAAFBC01FFF780155F7555568A00AAFF",
INIT_3B => X"AEA8A10082EA8BEFAAD5554B25551554BA0051400BA5551575EFF7D1401FF5D5",
INIT_3C => X"AAEAAB55F78400145AAFFFFFEF5D7FEABFF0051400A25D2EBFE10AAFFD55EFA2",
INIT_3D => X"552EA8AAA55043DFF7557BC01EF55557DE00AA842AA0000516AABAFF8428BE7A",
INIT_3E => X"0000000000000000000000000000000000000FFAABFF45FFAAAABFFAAFFFDFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(0),               -- Port A write enable input
DIA(0)   => data_write_a(6),        -- Port A data input
DOA(0)   => data_read_a_lo_512(6),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(0),               -- Port B write enable input
DIB(0)   => data_write_b(6),        -- Port B data input
DOB(0)   => data_read_b_lo_512(6),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_7_12 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10844B00482258A2842112C02450418800002300500030B313300C418992002",
INIT_01 => X"000009CA3839684D1CA0E0000E51424840000000080000080200080008510204",
INIT_02 => X"0120042086010000044600C00008000004100000000260900200000002402004",
INIT_03 => X"8628A10000082400000002408400080011000000610008000208C00000E14400",
INIT_04 => X"0911800100A000000000524084000040000050001140200100C8100000080102",
INIT_05 => X"0300812401011000000000002000114008008060441000000020024093000000",
INIT_06 => X"9190431C0D4010100000880804010010800000041080081000000200010424B2",
INIT_07 => X"000100AA0004408601000004860000008C02000A103010006928040800062481",
INIT_08 => X"84000048D484C20888000A0002120484C048007004000000000021F000000244",
INIT_09 => X"00A06009881201A520491004106C48A04040002400A15A208001650004001020",
INIT_0A => X"C99E1060201002044809C1040140A001004808810000459033189C0A400118A0",
INIT_0B => X"102000024040484050050041648A0041140C500B08821054C000264120000400",
INIT_0C => X"0404A083260E0832132011880462011880462051881462051881D31018C40620",
INIT_0D => X"0001000080001000813094801A8F80F00A600B52602801A88848011118003700",
INIT_0E => X"000003C007C002808228010410082042C000C000000004001002000400040002",
INIT_0F => X"A4000007800F80C840000800009864038A1200081C0014800000F001F0200052",
INIT_10 => X"00002C0E00E0E4004038000102400002C0E00E0D20100029000001E003E04000",
INIT_11 => X"2000C04031100E0403D0700300080908000100000661801E1900040380001804",
INIT_12 => X"0840878083E8003780A01043203A101780902043203A10082410082880000000",
INIT_13 => X"0601E0187900181035E0240806483248181035E0280410C8198818100DDD0000",
INIT_14 => X"0403774000201021E020FA006040376C00501022131210722060806D47000A40",
INIT_15 => X"00928A0002000110888600C032128201519480D40009902430160403E0E00506",
INIT_16 => X"01000000020080601802000000000405000A0020020081014134928820480010",
INIT_17 => X"0802018040000000006018020080200804010000000000806018020080000004",
INIT_18 => X"0000000001806008020000001006008020080001004008020080201004000020",
INIT_19 => X"0000000000000000000000000000400A004618618618C30C30C3000020180600",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000000B0840000000000000000000",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"1555500000000000000000000000000000000000000000000080000000000000",
INIT_28 => X"A97555F784174BAF7D5555FFF780155EFAAAEA8ABAAAFBFDE0055556AA005D04",
INIT_29 => X"55555EFAAFFFDFEFAAAAAAB455D556AA00FFAE95555087BFDF45F7AA974AAAAA",
INIT_2A => X"02EAAAAA082EA8A00AAAE955450055421FFFFFBC0010AAD5574BA557FFDFFF55",
INIT_2B => X"08043FE00F7AA97555A2FBD7410AA8428AAA557BFDFFF55003DFFFF7FBEAA000",
INIT_2C => X"0082A800AAF7AE975FFA28000010552EBDE00007BEAAAAA2D140000085155555",
INIT_2D => X"45087FEAB455D516AB55557BD55FF00557FE10FFFBEAA10007FD7410FFAA9740",
INIT_2E => X"000A2AA97400552AAAB45082E80155F7D1575EFFFAA955555D51574AAAAFFD55",
INIT_2F => X"AE105D556AA10410E17555000000000000000000000000000000000000000000",
INIT_30 => X"FFF55FFA095482B6A49256DEB84104BAFFD1525FFFF8E175C7A2AAAAA82A2F1F",
INIT_31 => X"F524AA5571FDFEF415B575D7AAF1FFFD7AAAAAFB7D495F6AA10E3AE905551C7B",
INIT_32 => X"003AFEFEBFBEAA001C2EA8A821C2EAAA00A2AE9756D145B401FFFFFFC7010BED",
INIT_33 => X"EDB470101C5B5057D1C003DE28F7A49057DAAF5D2428A2842AAAA497BFAFFF49",
INIT_34 => X"1475D5400F7A490438082485038F7A4905C7A28A070384120BDE100075EAA82B",
INIT_35 => X"D495150492BEF1D2555087BE8B7D555F6AB57417BC05D7145178E00EBFBE8A10",
INIT_36 => X"00000000000000000000AAA495428412AAFB451C2A8017DE3DF525FFFFA49756",
INIT_37 => X"555A2AEA8A10AAD568A00555168A10002E9754D0000000000000000000000000",
INIT_38 => X"8A10AAAE8215D557BFDF55F78017400F780001FFAA84000AAFFD1401E7FFAA97",
INIT_39 => X"C21EFF7FBD7400F7FBC00BA55557DFF7007BD5555AAD57DF55AAAEBDFEF007BE",
INIT_3A => X"428AA2007FE8BFF080028BFFAAFFEAA105D2EAAA005D2AAAA18AAAA975FF5D7B",
INIT_3B => X"043DE0000516AA10F7FBD7408557FC01EF55043FEAAFF80021EFA2D1420BAAA8",
INIT_3C => X"55568A00AAFFEAA105D5155410FF84020AA0800154B2FF8402145A2AA954AA00",
INIT_3D => X"AAFBC01FFF780155F7005140000FFD140145007FE8BEF557BEAB55087FC215D5",
INIT_3E => X"0000000000000000000000000000000000000AA80174AA082ABDF555D2A821EF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(0),               -- Port A write enable input
DIA(0)   => data_write_a(7),        -- Port A data input
DOA(0)   => data_read_a_lo_512(7),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(0),               -- Port B write enable input
DIB(0)   => data_write_b(7),        -- Port B data input
DOB(0)   => data_read_b_lo_512(7),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_8_12 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00000648E2840112C00000418000002700500030B3132000400812082",
INIT_01 => X"100008480009004C04A100000252024840000000180800080200010040110204",
INIT_02 => X"0020042000490000004600804008000005100000000024900200000002400004",
INIT_03 => X"0A0C33400008082400000080A4004B0891000020610112000040C00000E5C000",
INIT_04 => X"18800001000000000000512080000040800150400824280110C8100000120200",
INIT_05 => X"908084A10100100200004080280008240810802206940000012C214451610800",
INIT_06 => X"81B000080860109021400008040000202048020414A0021400040200322824C1",
INIT_07 => X"000000080004408049000004860000008402001A50208000630C040800062483",
INIT_08 => X"440000428644212280800A00021004044048002124000000000021F000000244",
INIT_09 => X"00004009001001010008100414644410400102228000D20080114502006409A2",
INIT_0A => X"000051312000042200294429148A4801C80C8C81000045907118040340020832",
INIT_0B => X"4020000240404140004D0544C4AA0001150410090302500011C813428A000400",
INIT_0C => X"46501090008820240240409000240009000240009000240009000120204808A5",
INIT_0D => X"42D1A168D09A301468402480004780F00140080860280004085904309A002196",
INIT_0E => X"00783FC00044340242280000000000020000C0000442106419120004034685A3",
INIT_0F => X"8000F07F800088A80000081EA2F9EC0000064004081010001E0FF00011104040",
INIT_10 => X"0ED0FC7E00000422201080000202658FC7E0000021882020003C1FE000222080",
INIT_11 => X"018059C3F350FE0C00000002A0040500000103961FE780000110010090000800",
INIT_12 => X"FD41FF80000830200021C1CF600012200010D1CF600012121600100810000004",
INIT_13 => X"9E1FE000010A1802100004343ED8000898021000087073D80008980200800002",
INIT_14 => X"0080200000BEB07FE00002086008020000209AEE3F300000246020200000620B",
INIT_15 => X"0088881903210000440610C8000A808040000208901786E4F0FE0C0000000166",
INIT_16 => X"685A1685A769DA368DA368DA769DA36CDA121A11A141800011309284002C0810",
INIT_17 => X"95A5685A1685A5695A368DA368DA769DA368DA368DA7695A1685A1685A5695A1",
INIT_18 => X"5A1695A568DA368DA369DA768DA1685A1695A5685A168DA369DA768DA368DA16",
INIT_19 => X"A4028A0A543EBC57A10A1E75D64108080468618618630C30C30C69DA5685A168",
INIT_1A => X"9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7BF3CCD8DF5B2DB2C",
INIT_1B => X"F87D3E1F4F87D3E1F4F87D3E1F4F87D3E1F4F87C3E1F0F87C3E1F0F87C3E79E7",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000006A6D4F87D3E1F4F87D3E1F4",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"155FF00000000000000000000000000000000000000000000080000000000000",
INIT_28 => X"BFDE0055556AA005D0415555080000000087BEAA10F7803DE00FFAEBFFFF0800",
INIT_29 => X"2AA8AAA557FC0010F780154105D7FC2145005155555F780155EFAAAEA8ABAAAF",
INIT_2A => X"7FFFFF55AA80155FF087BFDF45F7AA974AAAAAA97555F784174BAF7D5555FF55",
INIT_2B => X"AAFFFDFEFAAAAAAB455D556AA00FFAE95555AAFFE8A00552EBFE00F7D17FF45F",
INIT_2C => X"A557FFDFFF5504000AAAAAAA8B55F7D140010552E821EFAAAABDF555555555EF",
INIT_2D => X"55AA8028A00A2D57FF45557BE8A00AAAE955450055421FFFFFBC0010AAD5574B",
INIT_2E => X"000557BFDFFF55003DFFFF7FBEAA00002EAAAAA082EA8A00002AA8A10F784021",
INIT_2F => X"FE10F7AEBAFFF080A175D7000000000000000000000000000000000000000000",
INIT_30 => X"175C7A2AAAAA82A2F1FAE105D556AA10410E17555080E000280071E8A00EB8E3",
INIT_31 => X"4104BAFFD1525FF492EA8AAA5571C2000FF8A17400557FC015514555757DFF8E",
INIT_32 => X"2ABDE10EBDF7AF6DE3FFF8F7DB68A105D71C7BFFF55FFA095482B6A49256DEB8",
INIT_33 => X"AA0BDF6D415B575D7AAF1FFFD7AAAAAFB7D495F6AA10E3AE90555A2FBE8A3849",
INIT_34 => X"FFFFC7010BEDF524AA5571FDFEF550E00082B6A0AFB55F7D1420104124821D7A",
INIT_35 => X"01C2EA8A00F7800017DA2842FA00B6D578F6D557FFDA00A2AE9756D145B401FF",
INIT_36 => X"00000000000000000000497BFAFFF49003AFEFEBFBEAA001C2EA8A821C2EAAA0",
INIT_37 => X"0BA08556AA00AAAABFE00F7AEAABEF082E955450000000000000000000000000",
INIT_38 => X"21555D51575EFFFAA97555A2AEA8A10AAD568A00555168A10002E9754D082E82",
INIT_39 => X"17400F780001FFAA84000AAFFD1401E7082EAAABA5D5140010F7AE974105D7BC",
INIT_3A => X"E8215DA2FFE8ABA082ABFE00AAFBEABFFAAFBEABFFF7AA80145557BFDF55F780",
INIT_3B => X"D540000000402145AA843FFFF007BD5555AAD57DF55AAAEBDFEF007BE8A10AAA",
INIT_3C => X"AAA975FF5D7BC21EFF7FBD7400F7FBC00BA55557DFF75D2E82010F7843DF45FF",
INIT_3D => X"5D2EAAA005D2AAAA185D2AAAA10F780021FFA2803DE10FFD16ABFF5D7BFDE10A",
INIT_3E => X"0000000000000000000000000000000000000007FE8BFF080028BFFAAFFEAA10",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(1),               -- Port A write enable input
DIA(0)   => data_write_a(8),        -- Port A data input
DOA(0)   => data_read_a_lo_512(8),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(1),               -- Port B write enable input
DIB(0)   => data_write_b(8),        -- Port B data input
DOB(0)   => data_read_b_lo_512(8),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_9_12 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00018248A2840112C00002C18000002300500030B3132000400812006",
INIT_01 => X"400008000000004C0020000000100248413C0A61590001D90213C10008110204",
INIT_02 => X"01A0042080010000054600C04008000004100000001020900200200002420804",
INIT_03 => X"024003400008012400000010E4004B0891000020610310000144C00000F5C000",
INIT_04 => X"1801800100E000000000510084000040010050020810200000C8900000320200",
INIT_05 => X"918004311104100000000000200008100800002000100000002C234415610820",
INIT_06 => X"81B00008080010100000980804000008800042041080001000100200322C2481",
INIT_07 => X"0000811800044080010000058600000086020002502080006000040800062C80",
INIT_08 => X"0000004001D4618008800A00061004044048002004000000000061F000000244",
INIT_09 => X"000040090802009420409004104444084001022400214A2080014400026401A2",
INIT_0A => X"04000071200000A003CA294140200800C80C8C8100004590111C040040120800",
INIT_0B => X"12210002404848502847040164880021150400080222000200C8034200000000",
INIT_0C => X"4610088010080421021040841021000841021000841021000841010800420820",
INIT_0D => X"42D0A16C529A321068500484000500D10042080040284000084900001A002196",
INIT_0E => X"00000002804000004228010410082002C000C0002400046419120410034285A1",
INIT_0F => X"A00000000500800800000800000000000002290008001080000000A010100042",
INIT_10 => X"00000000000004C2001000000240000000000000680800280000000140202000",
INIT_11 => X"0000C0000000000000000442020001000001000000000000010C800080000804",
INIT_12 => X"08000000000801A7802010000000152780102000000015000600000800000000",
INIT_13 => X"000000000101900011E0240000000009500011E0280000000009500004DD0000",
INIT_14 => X"000137400020000000000201C000136C00101000000000002340002947000240",
INIT_15 => X"0080881901210000000600C280028000419480D4000010040000000000002304",
INIT_16 => X"68DA368DA1685A1685A1685A1685A16C5A121A13A141950051309284A82C0010",
INIT_17 => X"85A1685A1685A1685A368DA368DA368DA368DA368DA368DA368DA368DA368DA3",
INIT_18 => X"5A1685A168DA368DA368DA368DA368DA368DA368DA3685A1685A1685A1685A16",
INIT_19 => X"0157344CCCF48DE68A895C38E2540A8010100000000000000000685A1685A168",
INIT_1A => X"14514514514514514514514514514514514D34D34D34D34D28E1004039248209",
INIT_1B => X"D268341A4D268341A0D069349A0D069349A0D068341A0D068341A0D068345145",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000014D490D069349A0D068341A4",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"EAABA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"03DE00FFAEBFFFF0800155FFAAFBE8B45002A974AAAA803DFFFAA843DF45FFFF",
INIT_29 => X"7BFDE00A2FBD7400F7FBFDFFFA2AEBDE00AAFBEAABA080000000087BEAA10F78",
INIT_2A => X"055401FFF7AEAAA10F780155EFAAAEA8ABAAAFBFDE0055556AA005D041555508",
INIT_2B => X"557FC0010F780154105D7FC2145005155555557BE8BEF007FFDEAAAAD1555EF0",
INIT_2C => X"AF7D5555FFF780154AA5D2AA8A10F7AA974AA082E80010A2AAAAA10552AA8AAA",
INIT_2D => X"BAF7D17FEBAA2AEBDF45002EAAABA087BFDF45F7AA974AAAAAA97555F784174B",
INIT_2E => X"000AAFFE8A00552EBFE00F7D17FF45F7FFFFF55AA80155FF080400145FFFBEAA",
INIT_2F => X"8FC7BE8A3DF7DF7F5E8A92000000000000000000000000000000000000000000",
INIT_30 => X"000280071E8A00EB8E3FE10F7AEBAFFF080A175D7BEF1E8B6D002090482B68E3",
INIT_31 => X"56AA10410E175550871FFE00A2FBD0400FFF5FDFC7B6A0BDE38B6F5E8A92080E",
INIT_32 => X"7BFAE82A2DB555C71C5B451D7FFAAA8A38FF8E175C7A2AAAAA82A2F1FAE105D5",
INIT_33 => X"2AEADA38492EA8AAA5571C2000FF8A17400557FC015514555757D5D71E8BEF14",
INIT_34 => X"B6A49256DEB84104BAFFD1525FFFF84174BA5D20AAA00E3AA904BA142A87010A",
INIT_35 => X"7000400155FFFBEDA82FFD57DEBAAAA0BFF7D0024ADA921C7BFFF55FFA095482",
INIT_36 => X"00000000000000000000A2FBE8A38492ABDE10EBDF7AF6DE3FFF8F7DB68A105D",
INIT_37 => X"BEF080402000F7AAA8B55FFAABDFEFF7D16AA000000000000000000000000000",
INIT_38 => X"FEAAFFD16AA00082E820BA08556AA00AAAABFE00F7AEAABEF082E95545F7D568",
INIT_39 => X"A8A10AAD568A00555168A10002E9754D00517DE00A2FFC2000F7D17FF55FF803",
INIT_3A => X"1575EF555568BEF5D7FE8A10AAFFD55555D7FD5555FFAAA8AAAFFAA97555A2AE",
INIT_3B => X"AE800AA552A97400A2AEBDEAA082EAAABA5D5140010F7AE974105D7BC21555D5",
INIT_3C => X"57BFDF55F78017400F780001FFAA84000AAFFD1401E7FF80174AA5D0028A00AA",
INIT_3D => X"AAFBEABFFF7AA80145080002145F7FBFFE00FFD17FEAAA2803DFEF08043FE005",
INIT_3E => X"0000000000000000000000000000000000000A2FFE8ABA082ABFE00AAFBEABFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(1),               -- Port A write enable input
DIA(0)   => data_write_a(9),        -- Port A data input
DOA(0)   => data_read_a_lo_512(9),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(1),               -- Port B write enable input
DIB(0)   => data_write_b(9),        -- Port B data input
DOB(0)   => data_read_b_lo_512(9),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_10_12 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00018248A2840112C00002C18000202300500030B3132000400992006",
INIT_01 => X"254008000000004C002000000010026840000000080000080200010008110204",
INIT_02 => X"0020042000010000004455800008000004100000000000900200000002400004",
INIT_03 => X"020001021089000021081000C400090011000000610001540104C00000F14400",
INIT_04 => X"0811800101A00002000050088554004200C840000000200080C8100000000001",
INIT_05 => X"030080001000100800009400200000000840E020201000000024024001200020",
INIT_06 => X"81B00008080012120004CC080492500280208004148000100000020020042493",
INIT_07 => X"0000000800044080010000048404081085020002502000006000040800062480",
INIT_08 => X"100202400084410808000A00021004044048000004000000000021F020408264",
INIT_09 => X"010040090002008420401004144440004040022484214A2080110108C2C00320",
INIT_0A => X"04004166A48A0001080000000000080080181881000045901118044040020800",
INIT_0B => X"1201000200484910000F0105602622291404020902005002018002400A022000",
INIT_0C => X"0440001011808020120004801120044800120004801120044800110002400884",
INIT_0D => X"008000440210100041308480800F82F00040180260A808008848000018002104",
INIT_0E => X"000000028040000002280104100820020000400020000440100204100A000100",
INIT_0F => X"040000000500800800000000000000000002280008000400000000A010100010",
INIT_10 => X"00000000000004C2001000010000000000000000680800010000000140202000",
INIT_11 => X"200000000000000000000442000001000000000000000000010C000080001000",
INIT_12 => X"00000000000801C0008000000000154000800000000015000410000800000000",
INIT_13 => X"0000000001019800180000080000000958001800000400000009580002800000",
INIT_14 => X"0000A0000000000000000201E0000A0000400000000000002360002080000800",
INIT_15 => X"0080881000000000000600C28102800060000000000800000000000000002306",
INIT_16 => X"401004010040100401004010040100441020D0030008840051309A90BA884010",
INIT_17 => X"0902409024090240900401004010040100401004010040100401004010040100",
INIT_18 => X"1004010040902409024090240902409024090240902409024090240902409024",
INIT_19 => X"F546890A940FE0D3971243555205428290100000000000000000401004010040",
INIT_1A => X"8A28A28A28A28A28A28A28A28A28A28A28A28A28A28A28A29554199854514514",
INIT_1B => X"2B95CAE532994CA6532995CAE572B94CA6532994CA6532994CA6532994CA28A2",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000002718E72B94CA6532994CA657",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"FDE1000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"03DFFFAA843DF45FFFFEAABA007FC2155F7D155545AA80001EFAAFBEAB45557F",
INIT_29 => X"042AB55FFD168B55AA8000010FFFBE8BFFF78402155AAFBE8B45002A974AAAA8",
INIT_2A => X"AD16AABA002ABDE10080000000087BEAA10F7803DE00FFAEBFFFF0800155FF00",
INIT_2B => X"A2FBD7400F7FBFDFFFA2AEBDE00AAFBEAABAA2FFD741055003DFEFF7AA801FFA",
INIT_2C => X"05D0415555007FD74105555555EFF7FBC0145F78028A00A2D142155087BFDE00",
INIT_2D => X"55AAD168ABA002A975FFF7AEBDEBAF780155EFAAAEA8ABAAAFBFDE0055556AA0",
INIT_2E => X"000557BE8BEF007FFDEAAAAD1555EF0055401FFF7AEAAA105D042ABFF5D556AB",
INIT_2F => X"71D7AAFBEFB455D71F8E00000000000000000000000000000000000000000000",
INIT_30 => X"E8B6D002090482B68E38FC7BE8A3DF7DF7F5E8A92007BC217DEBDB55555AA8E0",
INIT_31 => X"EBAFFF080A175D700042AB7DEBDB6DB55BE8E05000EBFFE8BC7E38E07145BEF1",
INIT_32 => X"0A3DFD7F7A4821D7A2D16FA82142EB8E00080E000280071E8A00EB8E3FE10F7A",
INIT_33 => X"ED1421450871FFE00A2FBD0400FFF5FDFC7B6A0BDE38B6F5E8A92B6FBD541049",
INIT_34 => X"A2F1FAE105D556AA10410E175550071D54104951555D7EBF5C5155E3842AA00B",
INIT_35 => X"8410E2ABD749516FB55BED16FA820820955EFE3AEBDEAAFF8E175C7A2AAAAA82",
INIT_36 => X"000000000000000000005D71E8BEF147BFAE82A2DB555C71C5B451D7FFAAA8A3",
INIT_37 => X"1EFA2FFD7545AAAE97555A2FBFDF455D556AA000000000000000000000000000",
INIT_38 => X"8B45AAAA95545F7D568BEF080402000F7AAA8B55FFAABDFEFF7D16AA00087FC0",
INIT_39 => X"6AA00AAAABFE00F7AEAABEF082E9554500042ABFFA2FFFFF45F7AE97400AAFFE",
INIT_3A => X"16AA00FFFBD5400082EBFF45F78400155A2D57FE00552EA8A00082E820BA0855",
INIT_3B => X"D557555A2802AA10FFD54214500517DE00A2FFC2000F7D17FF55FF803FEAAFFD",
INIT_3C => X"FAA97555A2AEA8A10AAD568A00555168A10002E9754D085155410085557555AA",
INIT_3D => X"5D7FD5555FFAAA8AAA002AAAB4508557DF55F7D17FE000804155FFAAAABDEAAF",
INIT_3E => X"0000000000000000000000000000000000000555568BEF5D7FE8A10AAFFD5555",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(1),               -- Port A write enable input
DIA(0)   => data_write_a(10),        -- Port A data input
DOA(0)   => data_read_a_lo_512(10),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(1),               -- Port B write enable input
DIB(0)   => data_write_b(10),        -- Port B data input
DOB(0)   => data_read_b_lo_512(10),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_11_12 : RAMB16_S1_S1
generic map (
INIT_00 => X"A101C4B05A0034CA2840712C2D001419000002300500030B31B20084EC992002",
INIT_01 => X"90000986B83028491800E0000C26426040000000080000088200080802512224",
INIT_02 => X"1A2004205E010640024D00800008000004100000040EC090820018003241A00C",
INIT_03 => X"28639100000C5C00000045C08400C8001100000061806A001618C03001E54400",
INIT_04 => X"1A800001000009A0804059A190000040400040008058220008C8100000120D4E",
INIT_05 => X"02000E81080250010000002022000058080400000E1200000020004401000004",
INIT_06 => X"819435143F20101010001008040800B8100102041088011100022200000024B2",
INIT_07 => X"90640D280884453E01064002944180008402001295BA100022E4340800062D82",
INIT_08 => X"400000093204802200280A0012160585C1D808D004000000000323F40C102244",
INIT_09 => X"380040098010001100009204107C5950400000220080C200800900020C006827",
INIT_0A => X"80007100004016EA080801010000080D00200081000045B0511D289940103399",
INIT_0B => X"002000024040410A000D0104408810C115D9C008050042400100D04E88000002",
INIT_0C => X"00655010009264201200C7B421ED0C7B421ED0C7B431ED087B43176843DA1085",
INIT_0D => X"0401020080400A10012494881A4F80F209500BB2602881A488485C1318002000",
INIT_0E => X"6619A540124814800228010410082022C00040002020090020220C9600040802",
INIT_0F => X"ACCC334A802491600C587949B6D0141B4CC600D5761B1599865A500490B86A56",
INIT_10 => X"BAC845542056A61686EC81E3A6CB68AA2C622C9A251C352B330CB4A0092170D8",
INIT_11 => X"BCCAD0B5A81536080CC6B21A21B1FC09CB0F1076D4A200B2AD4068F4101639B5",
INIT_12 => X"4D2CC281E31AA0103AB8D5514066380804B268A2E060901204112566F10AC418",
INIT_13 => X"D551443C47281002540B2C9AAAA8662A1152B202AE3554403028115AA88201A1",
INIT_14 => X"548A20A0492A2724A0621620402A020141F172FB182A32AB6845AB6200251BC9",
INIT_15 => X"00C00A000200074044E6801832728080D00A380B753952C4877E0104DDE4D124",
INIT_16 => X"0080200802008020080200802008020480080022020081010124988800400010",
INIT_17 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_18 => X"0000000000802008020080200802008020080200802008020080200802008020",
INIT_19 => X"55062608804180C0B10A42104201400204000000000000000000000000000000",
INIT_1A => X"00000000000000000000000000000000000820820820820801C4149470000000",
INIT_1B => X"0000000000000000040200000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000007E0F0000000000000100800",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"000AA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0001EFAAFBEAB45557FFDE10082ABDF5508557DF45002ABDFFFF7803DE10AA80",
INIT_29 => X"AEBFF45FFAEBFEAA002A801FFF7FFE8A10A28000000007FC2155F7D155545AA8",
INIT_2A => X"2AABFE10082ABFFEFAAFBE8B45002A974AAAA803DFFFAA843DF45FFFFEAABAA2",
INIT_2B => X"FFD168B55AA8000010FFFBE8BFFF78402155AAD155555A28428BFF002ABDE00A",
INIT_2C => X"F0800155FF00557FF45557FC2010002A80010A2842AAAA007BFFF4500042AB55",
INIT_2D => X"FF5D00154BAF7FBE8BEFFFD540000080000000087BEAA10F7803DE00FFAEBFFF",
INIT_2E => X"000A2FFD741055003DFEFF7AA801FFAAD16AABA002ABDE10A2D168A10A284021",
INIT_2F => X"DFC7F78E3FE28B684070AA000000000000000000000000000000000000000000",
INIT_30 => X"C217DEBDB55555AA8E071D7AAFBEFB455D71F8E00002EBDF6D005B78F7D142AB",
INIT_31 => X"A3DF7DF7F5E8A92BEAEBFF7DEBA0BDEAA1C2A801C7E3FFEFA10B68407038007B",
INIT_32 => X"8A28BFF082ABAE10B6AAB8E280820B8FEFBEF1E8B6D002090482B68E38FC7BE8",
INIT_33 => X"07FF8F7D00042AB7DEBDB6DB55BE8E05000EBFFE8BC7E38E07145B6D15756DA2",
INIT_34 => X"EB8E3FE10F7AEBAFFF080A175D708517DF7D497BC5028142A87000A28A2AA920",
INIT_35 => X"0B6DB6AA28A280001FF5D0A10482FFFFEFBC7E3DF42028080E000280071E8A00",
INIT_36 => X"00000000000000000000B6FBD5410490A3DFD7F7A4821D7A2D16FA82142EB8E0",
INIT_37 => X"FEF007BE8BFF5D2ABDF55F7AABDEAAF784154BA0000000000000000000000000",
INIT_38 => X"DE00FF84154BA087FC01EFA2FFD7545AAAE97555A2FBFDF455D556AA00082EBF",
INIT_39 => X"02000F7AAA8B55FFAABDFEFF7D16AA00FFAEBFFEFAA803DEBA5D2E82155A2FBF",
INIT_3A => X"A95545F7D5555FFAAAAA8BFF002AAAA00FFAAA8AAA080028BFFF7D568BEF0804",
INIT_3B => X"2E95400A2AEA8A00007FEABFF00042ABFFA2FFFFF45F7AE97400AAFFE8B45AAA",
INIT_3C => X"82E820BA08556AA00AAAABFE00F7AEAABEF082E9554508557DFFF007BD54BA5D",
INIT_3D => X"A2D57FE00552EA8A00FFFFE8AAAAA80001FF5D2E82000F7FFFFF45AAFFC20BA0",
INIT_3E => X"0000000000000000000000000000000000000FFFBD5400082EBFF45F78400155",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(1),               -- Port A write enable input
DIA(0)   => data_write_a(11),        -- Port A data input
DOA(0)   => data_read_a_lo_512(11),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(1),               -- Port B write enable input
DIB(0)   => data_write_b(11),        -- Port B data input
DOB(0)   => data_read_b_lo_512(11),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_12_12 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50080B01BC002006940202C0DE041196A83183000000023322287E0FC000006",
INIT_01 => X"75400D849830C84C5823E0000C17424840000000080000088200002802153231",
INIT_02 => X"18A026B43ED180040147558040090000061800000C06ED9802768F4472C52005",
INIT_03 => X"2A67E34A528D0524A52850528400C8001100000171C02B550618C91A10E55440",
INIT_04 => X"1BC0000100056C8280825DE98154004300C840800850240080CA921084520A07",
INIT_05 => X"02000F832000500C0000941024000852084060202E100001002000448100000C",
INIT_06 => X"819A1D1C3FE01A1A40045408049A50BA4020C6041090001200006200000000F2",
INIT_07 => X"C26A0719CC96CC6ED18A64019695A854870300FA3968B20068FC06080106249F",
INIT_08 => X"D002024B3E040800008C0A002610240D494A06F3460409000000E3F0AD5282E5",
INIT_09 => X"27A06009200040000400120412445D78400001000410420080218029CC807A27",
INIT_0A => X"18000006848A026F000000000000080000F010C100204593F11A6CDF48003BF8",
INIT_0B => X"000000820040402B28050400400432C9349DF21A31A00ACC0000F04F80020001",
INIT_0C => X"00357804611AE45D05D0833430CD0833420CD0C33420CD0833430668619A1000",
INIT_0D => X"0000000000000A74812DF00E87E80A079F9F90FA0280E87E800C7FF3B8002000",
INIT_0E => X"3B6B0E404D26160682082002000401EA0000C40000800A006002818808000000",
INIT_0F => X"A476D61C809A4DA84272592D6246FC1B17B541F97E1B348EDA93900B2B286C56",
INIT_10 => X"30C669E622DBC325CFD881A962454CFBE5403AB99594362B1DB52720165650D9",
INIT_11 => X"F8D2D39A3745261E4A95A110A3F855000E4B1D32BAB504BB7490FCFF912A3834",
INIT_12 => X"B90E9B018C7530200AB8F8BF41F9A22006B37DC8E1F9A21A70116D4C5080651C",
INIT_13 => X"118780319CCA08AB1001ACDF34B8F1C688AB1002AE3F7B807B6289F368828C4C",
INIT_14 => X"2AF020233376A5ECC016B1A827CDA21160F051DE610A34C50427E6E220323E4A",
INIT_15 => X"0077020000000439FDC05C5806781FAB46095A0B5199B0AC55521524F1864022",
INIT_16 => X"000000000000000000000000000000000026C000002884000130921092804010",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"8020080200000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0051B946088881360A95090CB054420290100000000000000000008020080200",
INIT_1A => X"041041041041041041041041041041041049249249249249200100002D451451",
INIT_1B => X"92C964B2592C964B2592C964B2592C964B2592C86432190C86432190C8641041",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000003800F592C964B2592C964B25",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"7DE1000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"ABDFFFF7803DE10AA80000AAAA843FE0008557DFFF0800020105D557FEAA0055",
INIT_29 => X"D5420000051555FFA2AA8200000557DFFFF7AA80000082ABDF5508557DF45002",
INIT_2A => X"82AA8AAAAAFFC00BA007FC2155F7D155545AA80001EFAAFBEAB45557FFDE10AA",
INIT_2B => X"FFAEBFEAA002A801FFF7FFE8A10A28000000A2D155410F7FFFFEBA08003FE000",
INIT_2C => X"5FFFFEAABA000028A105D2ABFE10A2AABFE1055516ABEF5D517DEAAA2AEBFF45",
INIT_2D => X"55002A820AA08557DFFFF7AA82155AAFBE8B45002A974AAAA803DFFFAA843DF4",
INIT_2E => X"000AAD155555A28428BFF002ABDE00A2AABFE10082ABFFEF0855420000004175",
INIT_2F => X"5010495B7AE921C517DE10000000000000000000000000000000000000000000",
INIT_30 => X"BDF6D005B78F7D142ABDFC7F78E3FE28B684070AABE803AE38145B78FD700000",
INIT_31 => X"BEFB455D71F8E00BED547038145B505FFB6A487000005F7AFD7F7A482038002E",
INIT_32 => X"F1FDE821C003FE001C2EAAAAAB6F5C2082007BC217DEBDB55555AA8E071D7AAF",
INIT_33 => X"D517DEAABEAEBFF7DEBA0BDEAA1C2A801C7E3FFEFA10B68407038B6D550428FF",
INIT_34 => X"B68E38FC7BE8A3DF7DF7F5E8A9200002FA285D20BDE28A2A4B8E10555B68BEF5",
INIT_35 => X"F085F47038140010555142082082005F7DFD7F7A482155BEF1E8B6D002090482",
INIT_36 => X"00000000000000000000B6D15756DA28A28BFF082ABAE10B6AAB8E280820B8FE",
INIT_37 => X"ABA5D7FEAB45080015410007FEAA0055517DE000000000000000000000000000",
INIT_38 => X"AB45F780020BA082EBFFEF007BE8BFF5D2ABDF55F7AABDEAAF784154BAF7802A",
INIT_39 => X"D7545AAAE97555A2FBFDF455D556AA00F7D1554BA5D7BC01FFFF8015410007FE",
INIT_3A => X"4154BAF7D1400BAFFD57FE005D043FE10552EAAAAAFFD140000087FC01EFA2FF",
INIT_3B => X"8428A105D7FEABEF55557DEBAFFAEBFFEFAA803DEBA5D2E82155A2FBFDE00FF8",
INIT_3C => X"7D568BEF080402000F7AAA8B55FFAABDFEFF7D16AA0008003FEBA55003DEBAA2",
INIT_3D => X"FFAAA8AAA080028BFF087BD54AA550402145550000010087FFFF45F78402145F",
INIT_3E => X"0000000000000000000000000000000000000F7D5555FFAAAAA8BFF002AAAA00",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(1),               -- Port A write enable input
DIA(0)   => data_write_a(12),        -- Port A data input
DOA(0)   => data_read_a_lo_512(12),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(1),               -- Port B write enable input
DIB(0)   => data_write_b(12),        -- Port B data input
DOB(0)   => data_read_b_lo_512(12),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_13_12 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10154A0441836CA2840512822007C18000E02700500030B31B300040081A042",
INIT_01 => X"00000804A000C04800020000000002404001000008220008A200100802110204",
INIT_02 => X"02200430000104000A4700804008000004100000000420918204D3033240400D",
INIT_03 => X"AA4003400008592400000590C40009141100000C6180C0000000C00001E14000",
INIT_04 => X"0800000102400120088054019000004160004190BAA0270000C8100000600206",
INIT_05 => X"21000012040610050040000227003AA0082400E94C1200000824424005220020",
INIT_06 => X"81963B180C001010580000080400000058000004109C00138000020024142581",
INIT_07 => X"002C8008000441600106400A9600010494020002B8AAA000EF003408000E2580",
INIT_08 => X"000000E48194408000A00A001210040441C80320040210000002ABF004102244",
INIT_09 => X"2A004009640040100400940412D4C4004000022000104200802D983000480120",
INIT_0A => X"8000202020401480000000000000080C90090881000145B0111A14004015080D",
INIT_0B => X"00000002004040AA08050400404040C11444000805200A402090024000008002",
INIT_0C => X"8410000A00280020020040800020040800020000801020000800010020400000",
INIT_0D => X"84A14250A055100050100490000500D00040080040290000084E4000B800610C",
INIT_0E => X"DCD13042BEDA36820228000000000000C000400081A08BC812A2092B02850942",
INIT_0F => X"89B9A260857DB400431969CA985D480949D32804A40AB137341C10B7D6A02EC0",
INIT_10 => X"E6ACA678001CE7D0296C213A460CA4271CA2168AEC1017606E6838216FAD4055",
INIT_11 => X"84AD4961C281B20213073C5FC0058008632D30D522CE80239DCC01AB013A4D20",
INIT_12 => X"2E6B13804A4B01D83461299900F6BD583A519104A0EEBD1A141010B2A4C8E116",
INIT_13 => X"89E5E40913419151EE0E94641828F72B5151EE0D184B321037AF5158BB02D085",
INIT_14 => X"562EC0B42162D68EE0073AE1C562EC13D521921A4170300B2B458B56B01C2280",
INIT_15 => X"00888A120240034000E6DC8285028014B82372011FC1E4F5E0A00929684EAF84",
INIT_16 => X"50942509425094250942509425094254940A1421420082020120908800480030",
INIT_17 => X"0942509425094250942509425094250942509425094250942509425094250942",
INIT_18 => X"9425094250942509425094250942509425094250942509425094250942509425",
INIT_19 => X"F7EFBBEEFF3F7DF7FF3E9F7DF7E2450228000000000000000000509425094250",
INIT_1A => X"BAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBF7DFDFDDD555555",
INIT_1B => X"EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAEBAE",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000000000F7EBF5FAFD7EBF5FAFD7",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"2ABEF00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0020105D557FEAA00557DE10AAD5554BA087FFFF55557BD54AAF7FBC01FFA280",
INIT_29 => X"7BD75EF087FFFFEF557BEAB45552E80155AA802AB45AA843FE0008557DFFF080",
INIT_2A => X"FAE820AA5D5557555082ABDF5508557DF45002ABDFFFF7803DE10AA80000AA08",
INIT_2B => X"0051555FFA2AA8200000557DFFFF7AA80000AAD1420AA087BD7555FFD168AAAF",
INIT_2C => X"5557FFDE10AAAEA8BFFA2FBD7545FFD157555085140010F7AEAABFFAAD542000",
INIT_2D => X"BA557BE8A10A284154BAFFAAAAB45007FC2155F7D155545AA80001EFAAFBEAB4",
INIT_2E => X"000A2D155410F7FFFFEBA08003FE00082AA8AAAAAFFC00BA00002AAAAF7D5574",
INIT_2F => X"0492E3F1C71C7BE8A2ABD7000000000000000000000000000000000000000000",
INIT_30 => X"3AE38145B78FD7000005010495B7AE921C517DE10A2DB50482147FFAF554971D",
INIT_31 => X"E3FE28B684070AA1C71D25D7007FFAFD7497BE8B5555208217DBE8A2AB45BE80",
INIT_32 => X"7FD257DFFD568A82FFA4870BA555F5056D002EBDF6D005B78F7D142ABDFC7F78",
INIT_33 => X"FAAAFBFFBED547038145B505FFB6A487000005F7AFD7F7A482038AADF4709214",
INIT_34 => X"AA8E071D7AAFBEFB455D71F8E00A2A0ADBC7A2FFD257DE3DF52555085142000F",
INIT_35 => X"21C002AA92FFDF574824171EAA10B680124BAFFAAAFB45007BC217DEBDB55555",
INIT_36 => X"00000000000000000000B6D550428FFF1FDE821C003FE001C2EAAAAAB6F5C208",
INIT_37 => X"0105D7BE8B55085142010AAD157545F7AEA8B550000000000000000000000000",
INIT_38 => X"01EFF7AAA8B55F7802AABA5D7FEAB45080015410007FEAA0055517DE00A2FFC0",
INIT_39 => X"E8BFF5D2ABDF55F7AABDEAAF784154BA5D5140145007BE8B55087BEAB555D040",
INIT_3A => X"0020BAA2FFD54105D7FC21EFFFD16AA10FF80174AA557FC21EF082EBFFEF007B",
INIT_3B => X"FBC0155085540000FFAEBFFEFF7D1554BA5D7BC01FFFF8015410007FEAB45F78",
INIT_3C => X"87FC01EFA2FFD7545AAAE97555A2FBFDF455D556AA00A2803FF45AAFFC21EFAA",
INIT_3D => X"552EAAAAAFFD1400005D042AA00F7FBD5410085568A10FF80020AAFFAABFF550",
INIT_3E => X"0000000000000000000000000000000000000F7D1400BAFFD57FE005D043FE10",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(1),               -- Port A write enable input
DIA(0)   => data_write_a(13),        -- Port A data input
DOA(0)   => data_read_a_lo_512(13),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(1),               -- Port B write enable input
DIB(0)   => data_write_b(13),        -- Port B data input
DOB(0)   => data_read_b_lo_512(13),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_14_12 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10020A000180000284008280000281800000030000000033022000000580002",
INIT_01 => X"000008020000204D006800000030824840000000084000084200090008510200",
INIT_02 => X"0220043170010A600A4D008040080000041000000028009002000F333240800C",
INIT_03 => X"111813400008002400000000C400090011000000610200001104D83000F14000",
INIT_04 => X"0801800100A000000000540084000040000040000800200000C8100000000748",
INIT_05 => X"0100000000001000000000002000080008000000001000000024024001200020",
INIT_06 => X"819EB84028001010000000080400000000000004108000100000020020040081",
INIT_07 => X"92040608000440100102400A94810206844200021DA2A0002000340800062C80",
INIT_08 => X"000000000084400008800A001214040441481500040000000000A7F408002244",
INIT_09 => X"0A0040090002008420401004104444004000020400214A208001000002400120",
INIT_0A => X"0400002020000000000000000000080C8008088100004590111B480040120000",
INIT_0B => X"1000000200404800000504016000002114000008020000020080024000000000",
INIT_0C => X"0410000010000000000040001000000000000040000000000001000000000000",
INIT_0D => X"04810244825010004010000000000000000000000000000000080000B8002104",
INIT_0E => X"0002C38280001202020800000000001000004000000000401022000002040902",
INIT_0F => X"20000587050001404E8084341CBA3404800828805200008000E0E0A000080002",
INIT_10 => X"4D18178E012010C00224004091C3514072C000444A0400080001C1C140001000",
INIT_11 => X"51709A07424142084458476001003809D0104B01C5710044020C4006010500C5",
INIT_12 => X"C26EE3803180C18006519462A00005001460E4730000050A1011004001060049",
INIT_13 => X"01F9E00660318000000538318740000140000001B4600CE80001400000002B62",
INIT_14 => X"0000000AD89857B0E0684411800000003799EB764D000330C300000000E3554B",
INIT_15 => X"0000021002002C000024008284001A0902000422E3F5960080480A0216A07240",
INIT_16 => X"4090240902409024090240902409024090081021020080015134920800480010",
INIT_17 => X"0902409024090240902409024090240902409024090240902409024090240902",
INIT_18 => X"9024090240902409024090240902409024090240902409024090240902409024",
INIT_19 => X"F5579B4E5C8FF0F7BE9D5F7DF650400200000000000000000000409024090240",
INIT_1A => X"9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7BF7DDDDDFCF3CF3D",
INIT_1B => X"F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE79E7",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000003FFF03F9FCFE7F3F9FCFE7F3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"420BA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"BD54AAF7FBC01FFA2802ABEFA2FBE8B55A2AE80000F7D5555555D2AAAABAAAD1",
INIT_29 => X"AA801FFA28402000AAAE955455500155EF0804155EFAAD5554BA087FFFF55557",
INIT_2A => X"7AEA8B45080417400AA843FE0008557DFFF0800020105D557FEAA00557DE10A2",
INIT_2B => X"087FFFFEF557BEAB45552E80155AA802AB4500516AA00A2AE800BAFFFFC20BAF",
INIT_2C => X"0AA80000AA005568ABAA28402010A2843FEBAFFFBD7410A2D168BFF087BD75EF",
INIT_2D => X"005D7FFDF4555517DFEF00043FEAA082ABDF5508557DF45002ABDFFFF7803DE1",
INIT_2E => X"000AAD1420AA087BD7555FFD168AAAFFAE820AA5D5557555002E80155A280000",
INIT_2F => X"0555412AA8ABAAADB40092000000000000000000000000000000000000000000",
INIT_30 => X"50482147FFAF554971D0492E3F1C71C7BE8A2ABD7A2FFEDB55B6A080038E3DB5",
INIT_31 => X"B7AE921C517DE10A2AE851FFB68402038AAAA955554900105FF0800175D7A2DB",
INIT_32 => X"A0800BAE3F1C0092EBAAADB6D080A12410BE803AE38145B78FD7000005010495",
INIT_33 => X"2D568BC71C71D25D7007FFAFD7497BE8B5555208217DBE8A2AB451C556FA00A2",
INIT_34 => X"142ABDFC7F78E3FE28B684070AA00516DABAA28402038B6803DE82F7F5D5410A",
INIT_35 => X"D002A80155B680000105D7FF8F455D5F78FD7000E3FEAA002EBDF6D005B78F7D",
INIT_36 => X"00000000000000000000AADF47092147FD257DFFD568A82FFA4870BA555F5056",
INIT_37 => X"F55FF84000AAAAFBC0145002AA8AAAAAFFC20000000000000000000000000000",
INIT_38 => X"01EF080417555A2FFC00105D7BE8B55085142010AAD157545F7AEA8B55A2FBFF",
INIT_39 => X"EAB45080015410007FEAA0055517DE00A2AA955FFFF80020BAAAAA9754508000",
INIT_3A => X"AA8B555D557FE00A280020BAAAD140000A2AEBFFEF082A82010F7802AABA5D7F",
INIT_3B => X"803DE00FFD557400AAD56AB455D5140145007BE8B55087BEAB555D04001EFF7A",
INIT_3C => X"82EBFFEF007BE8BFF5D2ABDF55F7AABDEAAF784154BA08557FEAAA284000AAFF",
INIT_3D => X"FF80174AA557FC21EF082A80145F780020105D7BEAB45557BE8B45082EBFEBA0",
INIT_3E => X"0000000000000000000000000000000000000A2FFD54105D7FC21EFFFD16AA10",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(1),               -- Port A write enable input
DIA(0)   => data_write_a(14),        -- Port A data input
DOA(0)   => data_read_a_lo_512(14),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(1),               -- Port B write enable input
DIB(0)   => data_write_b(14),        -- Port B data input
DOB(0)   => data_read_b_lo_512(14),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_15_12 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000A000000000284000280000001800020030000000033022000000180002",
INIT_01 => X"8000080000000048000000000000026040000000080000080200000000110200",
INIT_02 => X"0020042004010E60004C0080000800000410000000020090020000300245E005",
INIT_03 => X"0000010000080400000000408400480111000000610008000000C00000E54400",
INIT_04 => X"980000010000000088C2550080000040000040000008A00028C8100000120000",
INIT_05 => X"020004012E025000000001322000000A28008000011000000220004D41000000",
INIT_06 => X"819588000800101000011008040000100001060418800510000A620000000092",
INIT_07 => X"0000000800044004010C20008440810284020002102220002000340800062480",
INIT_08 => X"0000000001140800002C0A001214050540C800400406180000002DF004000244",
INIT_09 => X"1E00400900000000000016041044400440000000000042008001000000000022",
INIT_0A => X"0000000000000220000000000000080C00000081000045901118000040000000",
INIT_0B => X"0000000200404000010500004000000114000009000000000000004200000000",
INIT_0C => X"0000000000000000000040001000040001000000000000000001000020000800",
INIT_0D => X"000000000000001001208000180800000000030200000180800C400030002000",
INIT_0E => X"0000000000002600020800000000001080004000000000000002000000000000",
INIT_0F => X"A400000000000000000008000000000000000000000014800000000000000052",
INIT_10 => X"0000000000000000000000010240000000000000000000290000000000000000",
INIT_11 => X"2001C05838120800000000000000000000010000000000000000000000001804",
INIT_12 => X"081004000000000000A010000000000000902000000000180010002020000000",
INIT_13 => X"6600000000000000000024080000000000000000280400000000000000000000",
INIT_14 => X"0000000000200801000000000000000000501001920000000000000000000A40",
INIT_15 => X"0000020000000000000000003000000000000000000A101C3614000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000080000120980000000010",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000400200000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"28BEF00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"5555555D2AAAABAAAD1420BAFF8000010082A954BA00003DFEF085155400F784",
INIT_29 => X"AE95555A2FBE8BEFA2843DE00AA8015400FF84001EFA2FBE8B55A2AE80000F7D",
INIT_2A => X"2FBEAB45F7D56AABAAAD5554BA087FFFF55557BD54AAF7FBC01FFA2802ABEFF7",
INIT_2B => X"A28402000AAAE955455500155EF0804155EFFFFBE8BFF0800174AA557BFDE10A",
INIT_2C => X"A00557DE10F7D1574AAA2D16AB55FFD568BEF087FE8A1055003FE00A2AA801FF",
INIT_2D => X"00AA802AA00AAAE800BA5D0015545AA843FE0008557DFFF0800020105D557FEA",
INIT_2E => X"00000516AA00A2AE800BAFFFFC20BAF7AEA8B45080417400FFFFC21450800154",
INIT_2F => X"8FD7005150438F78A2DBFF000000000000000000000000000000000000000000",
INIT_30 => X"EDB55B6A080038E3DB50555412AA8ABAAADB40092E38E070280024904AA1C043",
INIT_31 => X"1C71C7BE8A2ABD7E3AA9257DA2FFE8BC7BE8E38E10A28017400E38A051FFA2FF",
INIT_32 => X"00124AA557FFDE10A2FBEDB6DF7D16AABAA2DB50482147FFAF554971D0492E3F",
INIT_33 => X"10038E38A2AE851FFB68402038AAAA955554900105FF0800175D7E3FFEFBD700",
INIT_34 => X"000005010495B7AE921C517DE10FFDF50482A2DB6AB45FFD56DBD7087BEAA384",
INIT_35 => X"0FFF1C017D140410400BE8E28A10AAA085082550A1057DBE803AE38145B78FD7",
INIT_36 => X"000000000000000000001C556FA00A2A0800BAE3F1C0092EBAAADB6D080A1241",
INIT_37 => X"4AA0800020BA550028B550855400AAF7AEBDFEF0000000000000000000000000",
INIT_38 => X"7400AAAE975EFA2FBFFF55FF84000AAAAFBC0145002AA8AAAAAFFC2000AAAA97",
INIT_39 => X"E8B55085142010AAD157545F7AEA8B55AAAE821EFAAFBEAB55F7AAA8A00AA841",
INIT_3A => X"417555AAFFFDF450804020AA557BFFE10A2FFFFFEFF7D568ABAA2FFC00105D7B",
INIT_3B => X"D17DF45007FE8AAA08002AAAAA2AA955FFFF80020BAAAAA975450800001EF080",
INIT_3C => X"7802AABA5D7FEAB45080015410007FEAA0055517DE00FFFBC2000AAFBE8B55F7",
INIT_3D => X"A2AEBFFEF082A82010FFD5421EF5D0000010F7AAA8A10AA8017400552A801EFF",
INIT_3E => X"00000000000000000000000000000000000005D557FE00A280020BAAAD140000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(1),               -- Port A write enable input
DIA(0)   => data_write_a(15),        -- Port A data input
DOA(0)   => data_read_a_lo_512(15),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(1),               -- Port B write enable input
DIB(0)   => data_write_b(15),        -- Port B data input
DOB(0)   => data_read_b_lo_512(15),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_16_12 : RAMB16_S1_S1
generic map (
INIT_00 => X"DA22C618B1000482B688B186588884862A400438255FC38381441205BA803003",
INIT_01 => X"7045A80028404C211203A952A90341080B173340412000E1005D628000820484",
INIT_02 => X"428406A4000850848330118D0AAC55001349B108818005460229044001C01784",
INIT_03 => X"092C4020000500020000500986812C405000001A48202050000A214AC0650115",
INIT_04 => X"4804A55440256F504025E003A054F46415A4E62B6FE3307943965A00001A1152",
INIT_05 => X"0000001C40A5B950ADB8EA097057ECE14C86D2B7F85AAD17F4B100000B88148C",
INIT_06 => X"415401DCDCF2C0A8030140BCB0820A200342A1C641C1E8782F508F2B00003584",
INIT_07 => X"002701881A3202080AE00480A2002840BE1480FA004342AA6F12000054004867",
INIT_08 => X"08C54828091002000002B32A8C19064E486A8001510000014140C1E2A14891E0",
INIT_09 => X"015452B103020814004088B64102680B6596594800400413CAC0208944800000",
INIT_0A => X"96AA000484094C000000000000012C9000A0000D0A80000BF8028E87C1B99270",
INIT_0B => X"014808A02004200E540480212000A448C0082024AE50064B44000000000002A2",
INIT_0C => X"0004000D5846256AAEA811150445411150445411150445411150422A088A8200",
INIT_0D => X"00000004010042A204A0C5817D00005034052E40000817D00440004004AD3240",
INIT_0E => X"632B2673FA4587978A2004102800809225545155121740000004900090000000",
INIT_0F => X"00C6564CE7F4EA4B940076D296D003030800462CBD320018CAAAACFE9164C800",
INIT_10 => X"28834ADB1440A114793A4A30A40839AA14910D08DCB2640031955559FD3AC990",
INIT_11 => X"594AB0B1A025371CA0E034E8443C097A800EB090D4AAC91208ED2FA0CE5E09B1",
INIT_12 => X"7B50446083001B94BB38C540EBE61284BB304880E3E4579EDC00992980D58033",
INIT_13 => X"5511121840E7A2CD952ECC12ABC3E6ACB3DFB12ECE315000F61FF1727A85FDBC",
INIT_14 => X"75DEB07F6F2E7084517F126F8395CB2BEFBAB8BA8AF698228CC5E2F08ECA5159",
INIT_15 => X"5580A840A8009F8B108C80A1021B080AFC0DF6422C6077F4A77F20D0C0E21084",
INIT_16 => X"0000000000000000000000000000000000044000102A0001148442A110810359",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"558D11544C690DA64C1C4F68A360400000000000000000000000000000000000",
INIT_1A => X"14D14D14D14D14D14D14D14D14D14D14D14514514514514529E5F87869E79E78",
INIT_1B => X"D1E8F47A3D1E8F47A7D3E9F4FA7D3E9F4FA7D3E9F47A7D1E9F47A7D1E9F4D14D",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000007D3E9F4FA7D3E8F47A3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"C00AA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"03DFEF085155400F78428BEF087FFFFEFF7D168B55AAD17FFFF552EBFE00007F",
INIT_29 => X"2E975EFF7D568BFFFF80175EF0004000BA552A821FFFF8000010082A954BA000",
INIT_2A => X"55540000082EAABFFA2FBE8B55A2AE80000F7D5555555D2AAAABAAAD1420BA5D",
INIT_2B => X"A2FBE8BEFA2843DE00AA8015400FF84001EF0000020AA5D00154005D043FF455",
INIT_2C => X"FA2802ABEF557BEABEF5D0415410087FD74BAAAAEBFFEF557FC00AAF7AE95555",
INIT_2D => X"FFFFAABFEAAFF84001FF002A821FFAAD5554BA087FFFF55557BD54AAF7FBC01F",
INIT_2E => X"000FFFBE8BFF0800174AA557BFDE10A2FBEAB45F7D56AABA082A97545F7D16AB",
INIT_2F => X"FFEF552AB8E38087FC2092000000000000000000000000000000000000000000",
INIT_30 => X"070280024904AA1C0438FD7005150438F78A2DBFF0871F8FC7E3D56AB6DBEDB7",
INIT_31 => X"AA8ABAAADB400924920925EFF7D16ABFFE38E175EF1400000BA412E871FFE38E",
INIT_32 => X"0A1240055003FF6D5551420101C2EAFBD7A2FFEDB55B6A080038E3DB50555412",
INIT_33 => X"57FC00BAE3AA9257DA2FFE8BC7BE8E38E10A28017400E38A051FF0804050BA41",
INIT_34 => X"4971D0492E3F1C71C7BE8A2ABD74975EDBC7550E12410087FD74AAB6AABFFC75",
INIT_35 => X"A08249756DF7D168BC7F7AABAEAAF780051C70824851D7A2DB50482147FFAF55",
INIT_36 => X"00000000000000000000E3FFEFBD70000124AA557FFDE10A2FBEDB6DF7D16AAB",
INIT_37 => X"B55A2D16ABEFFFFBFDFFF552AAAAAA007BC00000000000000000000000000000",
INIT_38 => X"20AA002A955EFAAAA974AA0800020BA550028B550855400AAF7AEBDFEF08516A",
INIT_39 => X"000AAAAFBC0145002AA8AAAAAFFC20000000021EFF7D568BFFA2AA955FF5D040",
INIT_3A => X"E975EF0800174BA002E820105D003DFEF5D51420005D2ABFF45A2FBFFF55FF84",
INIT_3B => X"7BD74AAF7AEBDF455D7BC20BAAAAE821EFAAFBEAB55F7AAA8A00AA8417400AAA",
INIT_3C => X"2FFC00105D7BE8B55085142010AAD157545F7AEA8B5500557DF45552A8200000",
INIT_3D => X"A2FFFFFEFF7D568ABA0804155FFF7D568B55FFAAAAABAFF8415545000015555A",
INIT_3E => X"0000000000000000000000000000000000000AAFFFDF450804020AA557BFFE10",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(2),               -- Port A write enable input
DIA(0)   => data_write_a(16),        -- Port A data input
DOA(0)   => data_read_a_lo_512(16),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(2),               -- Port B write enable input
DIB(0)   => data_write_b(16),        -- Port B data input
DOB(0)   => data_read_b_lo_512(16),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_17_12 : RAMB16_S1_S1
generic map (
INIT_00 => X"5284CE4FB7BD2C8994A13392DBD02E14006B82AC7E800D44D3DD2FD5F9B961C0",
INIT_01 => X"2EACD01F7E03FC6793F2199B39FC233C11D93AE6F3BB92B32091DBC339B24542",
INIT_02 => X"E63CCCC00A82C08092A2AFAE667033DB50853379C10BFDC5C6F4044443C817C6",
INIT_03 => X"7FF183635AEF9E3635AEF9E18E237040404446965C0607EE6DB7854AC4DE060C",
INIT_04 => X"D78AC33FB604488B000892EF17BE6D84196482236FE100294152E294350FB697",
INIT_05 => X"081B5F9B409420D0CDB47A05403F6CE0C08A4AB7F840EDB6F48100DFC8081081",
INIT_06 => X"768465354781CBC30316367077B4BDB50646E8D87100A8201ED01C19C020F71A",
INIT_07 => X"4002A110C922480A82D0841147162C48EBB9537A0022DC67987042EE976ABEA7",
INIT_08 => X"DB931BFEF91C00002CC0E019C0C82A4E4820C15A2330E004401891181168C4D1",
INIT_09 => X"09F3A1BC11EFBC66DB65307071477FF1030C397C060B4254064302042F803A69",
INIT_0A => X"3F330802162F3B7EE3F3EC7C7DEF207000F00059D2ED56D7EED2ED3C9A867DC0",
INIT_0B => X"185C44B91BC1740B7605040BE0018CFC7429F326B9E822FFC00074D5A0AB033A",
INIT_0C => X"00367A28FC1B7F7FEFFCFBFF3EFFCFBFF3EFFCFBFF3EFFCFBFF3EFFE7DFF9E00",
INIT_0D => X"0000000008004BA78428C7AD7FC94B533F5B4FFBD2FAD7FCCA786D43FE67C218",
INIT_0E => X"BA494CEBFD4F2667ABB6F68B29760593F33FA0CF170F40006001B1A05C000000",
INIT_0F => X"7F749299D7FAEB237DFE5865B6D2BF23265CBACE542A6FEE92333AFF33E0A9BF",
INIT_10 => X"F6C24B6D18C3C9F8E2881F3F787D776B5DB94A09955054DFDD246675FE7AC153",
INIT_11 => X"BFB349E08FF9A27EDE9FA8AEFD9E7467BFCB195CFEB56A1A70D34D1706FFFA3E",
INIT_12 => X"6FE219CA80725B875EED723FF7FCB2875EDAAFEAF7FD929BFD55BBC71D79F639",
INIT_13 => X"546670D018E7A6E581D7B6AB75FDFCECA6E581D7BB5DDFC6FF0EB7D7E859FDB5",
INIT_14 => X"B978177F6D6AF5ECDB5FB76A5F5FA165B456E0FB308710C49FCFB741598B9C7E",
INIT_15 => X"CFDAAB00AC00A8BBFC8B501CF7A0FED9A540EA1952586CEB54D143ACFF9A3BA9",
INIT_16 => X"000000000000000000000000000000000026E100002F382DBD9ECFE117805F20",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"4372003009EDCC4052E917114F981800C0000000000000000000000000000000",
INIT_1A => X"BA69A69AEBA69AEBA69A69AEBA69AEBA69A69A69A69A69A68698686981D75D74",
INIT_1B => X"6A351A8D46A351A8D068341A0D068341A0D068341A0D46A341A0D46A341A69AE",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000000000046A351A8D46A351A8D4",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"7FEAA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"17FFFF552EBFE00007FC00AA087FFFFFFFFFFFFFEFF7FBEAB450804001EFAAD5",
INIT_29 => X"D168A000004020AA5D7BE8B450051401EF087FD74AA087FFFFEFF7D168B55AAD",
INIT_2A => X"D7FEAB55FF80175EFFF8000010082A954BA00003DFEF085155400F78428BEFAA",
INIT_2B => X"F7D568BFFFF80175EF0004000BA552A821FF5D00020BA552A82000552A821555",
INIT_2C => X"AAAD1420BAFFFFFDF45AAD17FFFFAAFBC01EF5D0015555557BFDEBA5D2E975EF",
INIT_2D => X"BA007FEABEF005555555A2D1554BAA2FBE8B55A2AE80000F7D5555555D2AAAAB",
INIT_2E => X"0000000020AA5D00154005D043FF45555540000082EAABFF00516AA10552E820",
INIT_2F => X"8B550000071EFB6DF7AE92000000000000000000000000000000000000000000",
INIT_30 => X"F8FC7E3D56AB6DBEDB7FFEF552AB8E38087FC2092147FFFFFFFFFBFDFC7EBF5E",
INIT_31 => X"150438F78A2DBFFBED16AA381C0A07082497FEFB6D1451471EF007BD04920871",
INIT_32 => X"2A850105D2A80155417BEFB6DEB8E175FFE38E070280024904AA1C0438FD7005",
INIT_33 => X"D7BFAEBA4920925EFF7D16ABFFE38E175EF1400000BA412E871FF550A0009249",
INIT_34 => X"E3DB50555412AA8ABAAADB40092FFF5FFF6DAADF7FFD7B6F1C71EF55001756D5",
INIT_35 => X"7145B6AA28492487082007FEDBD700515556DA2DF50492A2FFEDB55B6A080038",
INIT_36 => X"000000000000000000000804050BA410A1240055003FF6D5551420101C2EAFBD",
INIT_37 => X"FEFF7FBFFF55A2D16AB550000175EFFFFBEAA000000000000000000000000000",
INIT_38 => X"55EF087FC200008516AB55A2D16ABEFFFFBFDFFF552AAAAAA007BC0000557FFD",
INIT_39 => X"020BA550028B550855400AAF7AEBDFEFF7D568AAA5D2A97410007BFFFFF55515",
INIT_3A => X"A955EF5D2E80010002A954005D2A82155087FFFFEFAAAA975EFAAAA974AA0800",
INIT_3B => X"D1575FF5504175EF5D7FEAAAA0000021EFF7D568BFFA2AA955FF5D04020AA002",
INIT_3C => X"2FBFFF55FF84000AAAAFBC0145002AA8AAAAAFFC2000FFD57DFFFAAFFFDF55FF",
INIT_3D => X"5D51420005D2ABFF45557FE8AAA000415410007BFFF450051555EFA2FBC0000A",
INIT_3E => X"00000000000000000000000000000000000000800174BA002E820105D003DFEF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(2),               -- Port A write enable input
DIA(0)   => data_write_a(17),        -- Port A data input
DOA(0)   => data_read_a_lo_512(17),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(2),               -- Port B write enable input
DIB(0)   => data_write_b(17),        -- Port B data input
DOB(0)   => data_read_b_lo_512(17),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_18_12 : RAMB16_S1_S1
generic map (
INIT_00 => X"69844019080000A21A611406840014122A641074155FC28A2024001001801003",
INIT_01 => X"7443D920034004180005E9E3C90360C0041C0181002001602025800008440084",
INIT_02 => X"E2DCCCE61D5C008103F2000781FC0FEDEAC2161B0B8FB0008620044443006010",
INIT_03 => X"884E300802006900802006995C896D605200000856E24A040000640052141103",
INIT_04 => X"480520FC026125AC0025C9122644E3E40EC8E2001001302281841A009038A86A",
INIT_05 => X"432000040089983070019400F01010004C8DB841405A80A100B586200FAC24AE",
INIT_06 => X"09044359DC7040000000002C109B0E0A00A1104641C0803804000707284600E1",
INIT_07 => X"400D10100400481D5EB08501620000007500CE801241021FE78E404860140060",
INIT_08 => X"00880C0106A0528020019307CC082A0A4A6A01ED725021400040D028000A9729",
INIT_09 => X"00117063038000282081402E4106400B6186128040600C10C1C0200950508110",
INIT_0A => X"C0C30C2E21580C874004008080003C32A10A19090C02010E1022944061688000",
INIT_0B => X"0180A8062026000DC425C0301311324AA2373088479105D044A1022000001835",
INIT_0C => X"0D89844703649000000200000000000000000000000000000000000000000010",
INIT_0D => X"0D8306C182701404C1973010802020404084001E00010802046092B5001FB365",
INIT_0E => X"528EB314068AB8B803DB00002900800400FC503F08180050942E4200020C1B06",
INIT_0F => X"40A51D66280D6032C5F96D3C51555D5D7D5AA87285820814A3CCC501C2A60820",
INIT_10 => X"8B35A3FEBF1FEDFD9C2B30E0468AAAD5D48F37E8FC1304102947998A03984C10",
INIT_11 => X"440FE1DD772D37A0A321BC6968F32658BF2D4F2A80BF8FE3F9FE3AC362080529",
INIT_12 => X"5487910D7E5A6D961A28456A1832E5161A100DD5182BC54020EA67A189C6ED36",
INIT_13 => X"AA444CAF91EDD1B725868403BE06323551B725868A100ABD119753B70964122B",
INIT_14 => X"EDC259048ACD868EE3803D65CEDC258A8F80D55E007C3F8EBB56F4C5362C978F",
INIT_15 => X"3F240014BE84370001B6922070440556B15F7FABBC0031BCF2257C41634B14D4",
INIT_16 => X"C1B06C1B06C1B06C1B06C1B06C1B06C1B0491069068000004060300A005A0118",
INIT_17 => X"1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06",
INIT_18 => X"B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C",
INIT_19 => X"B28BBECEB80EE173C2300F7DF16000000000000000000000000041B06C1B06C1",
INIT_1A => X"8A28A28AAAAAAA28A28A28AAAAAAA28A28A28A28A28A28A2910591505C104104",
INIT_1B => X"28944A25128944A25128944A25128944A25128944A2552A954AA5128944AAAA2",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000128944A25128944A251",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"9540000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"BEAB450804001EFAAD57FEAA087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974BA082E",
INIT_29 => X"7FFFFFFFFFBFDF45AAD568B55080028B55002E82000087FFFFFFFFFFFFFEFF7F",
INIT_2A => X"0043DE10AA843DE00087FFFFEFF7D168B55AAD17FFFF552EBFE00007FC00AA08",
INIT_2B => X"0004020AA5D7BE8B450051401EF087FD74AAAAFFFDF45A2D16AB55F7FFFFFFF0",
INIT_2C => X"0F78428BEFAA80000000804154BA55042ABEF5D7FD75FFAAD540145AAD168A00",
INIT_2D => X"00082E95555085168A10557FD7545FF8000010082A954BA00003DFEF08515540",
INIT_2E => X"0005D00020BA552A82000552A821555D7FEAB55FF80175EF5D00020105D2A974",
INIT_2F => X"DFFF5D2A954AA082A92428000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFBFDFC7EBF5E8B550000071EFB6DF7AE921C7FFFFFFFFFFFFFFFF7FBF",
INIT_31 => X"AB8E38087FC2092087FFDFC7E3F1FAF55A2DF6DB7D1C002AB7D002A82028147F",
INIT_32 => X"DF6DB7DE3F5FAFC708003DE28B68E38E280871F8FC7E3D56AB6DBEDB7FFEF552",
INIT_33 => X"ADF4516DBED16AA381C0A07082497FEFB6D1451471EF007BD0492B6F1F8F55AA",
INIT_34 => X"1C0438FD7005150438F78A2DBFFA28407038140410492550A2ABC7497BD25FFA",
INIT_35 => X"F5D0E05000492097428002E9557D1C516FA28417BD5545E38E070280024904AA",
INIT_36 => X"00000000000000000000550A00092492A850105D2A80155417BEFB6DEB8E175F",
INIT_37 => X"FFFFFFFFDFEFF7FBFFFEF552E974AA082A820AA0000000000000000000000000",
INIT_38 => X"ABEF002A800AA557FFDFEFF7FBFFF55A2D16AB550000175EFFFFBEAA00557FFF",
INIT_39 => X"6ABEFFFFBFDFFF552AAAAAA007BC0000087BFDF45AAD568B55AAFBFDFEF55042",
INIT_3A => X"FC2000FFD56AB45A2FFFDFFFAAD16AB4500043DEAAFFAEAAAAA08516AB55A2D1",
INIT_3B => X"2AA8B45087FC01EFA2FFD55EFF7D568AAA5D2A97410007BFFFFF5551555EF087",
INIT_3C => X"AAA974AA0800020BA550028B550855400AAF7AEBDFEFA280154BA55040000055",
INIT_3D => X"087FFFFEFAAAA975EF5D2E974000804154BA082A975EF5D517DEAA007BD5545A",
INIT_3E => X"00000000000000000000000000000000000005D2E80010002A954005D2A82155",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(2),               -- Port A write enable input
DIA(0)   => data_write_a(18),        -- Port A data input
DOA(0)   => data_read_a_lo_512(18),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(2),               -- Port B write enable input
DIB(0)   => data_write_b(18),        -- Port B data input
DOB(0)   => data_read_b_lo_512(18),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_19_12 : RAMB16_S1_S1
generic map (
INIT_00 => X"042200000000000041088001001AA00000000000000000000000500802000003",
INIT_01 => X"040048000024000000000404000000000A22000800000800004A200000000001",
INIT_02 => X"200C8840085EB00480060000001C008002489E0F000405EA0004040404000000",
INIT_03 => X"24004000000000000000000900002C4050000000000069500208400002E14100",
INIT_04 => X"4800200C0000000044002000C80020E40000E200000130200188000000800100",
INIT_05 => X"000000000080181000000000701000004C8000000058800000B1000009880480",
INIT_06 => X"80500081081040000000002C100040400000004641C080380400070100000000",
INIT_07 => X"4020109801A4CE005C00048380142810010564C4100114012002402028044808",
INIT_08 => X"0070700000000000000083004C3902420062000020E0000100004082A140102B",
INIT_09 => X"001150200000000000000026400000016186100000000010C04002C000000000",
INIT_0A => X"007C00008082C0002000000000002C3000000004050001030102040000000000",
INIT_0B => X"0000000000000000000000000000010000800011000000000000000000000BC0",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"000000000000000000000000000000042000760000000000000000010004B200",
INIT_0E => X"0D74002280300F0002FB069040000060000C5003000800000000000000000000",
INIT_0F => X"C01AE8004500744C780687DBA828008080A5FC0D385598035D0008A00C015660",
INIT_10 => X"39D8140040201BF861F0E7D693E6170022408116DFE0AB3006BA0011401D02AC",
INIT_11 => X"5412E4997F5249FD005043B8680CC98F00D0F2DD0140100406FE053A98F6ECC7",
INIT_12 => X"7418663001858040E153888000010840E165D0000000285C246A181C03FE4662",
INIT_13 => X"8199830066F0020858385974000001260208583854E2200000660208D6B1423F",
INIT_14 => X"8235AC508FCE8811042040F008235AE04420C040CF00C031C80009B8F224978B",
INIT_15 => X"030004E00000C220010808C10D9A92A74CD7CF4A09051110AD5A3C9200B7F280",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000118",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"07208BBA3F0C7010C660C7441920000000000000000000000000000000000000",
INIT_1A => X"861869A61861861861869A61861861861861861861861861A8208C4C1534D34C",
INIT_1B => X"984C26130984C26130984C26130984C26130984D26930984C26130984C261861",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000984C26130984C26130",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"174BA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFDFEF5D2A974BA082E95400F7FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0004",
INIT_29 => X"FFFFFFFFFFFFFFFFF7FBFDFFF552E974BAA2FFFFE10087FFFFFFFFFFFFFFFFFF",
INIT_2A => X"004001EFAAAEA8ABA087FFFFFFFFFFFFFEFF7FBEAB450804001EFAAD57FEAAF7",
INIT_2B => X"FFFBFDF45AAD568B55080028B55002E82000F7FFFFFFFFFFFFDFEFA2D568B550",
INIT_2C => X"0007FC00AAF7FFFFFFFF7FBE8B55AAD16ABEF5D2ABFF55080402010087FFFFFF",
INIT_2D => X"55A2FFFDFEF5D2EBFE00AAFFFFEBA087FFFFEFF7D168B55AAD17FFFF552EBFE0",
INIT_2E => X"000AAFFFDF45A2D16AB55F7FFFFFFF00043DE10AA843DE00557FFDFEFA2D16AB",
INIT_2F => X"FFEF552A974AA0000104AA000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFF7FBFDFFF5D2A954AA082A92428E3FFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"0071EFB6DF7AE92EBFFFFFFFFFFFFDFEFF7F5FAFC7492A974AAB6F5F8E101C7F",
INIT_32 => X"F1F8FD7AAD16AB450000001FFBEA4A8AAA147FFFFFFFFFBFDFC7EBF5E8B55000",
INIT_33 => X"00000010087FFDFC7E3F1FAF55A2DF6DB7D1C002AB7D002A82028FFFFFFFEFF7",
INIT_34 => X"BEDB7FFEF552AB8E38087FC2092F7FBF8FC7E3F5EAB45B6DF6FBEF5D2AB8F7D0",
INIT_35 => X"84971F8FC7AAD56DB6DBEF5F8FD7412ABFE28B6F5F8E820871F8FC7E3D56AB6D",
INIT_36 => X"00000000000000000000B6F1F8F55AADF6DB7DE3F5FAFC708003DE28B68E38E2",
INIT_37 => X"FFFFFFFFFFFFFFFFFDFEF552E954AA0004000AA0000000000000000000000000",
INIT_38 => X"54AAF7D568A00557FFFFFFFFFFFDFEFF7FBFFFEF552E974AA082A820AAA2FFFF",
INIT_39 => X"FFF55A2D16AB550000175EFFFFBEAA00A2FFFFFFFF7FBFDFFFFFD568B55002A9",
INIT_3A => X"A800AAF7FBFDFEFF7D56AB45AAD56AB450004001EFFF842AAAA557FFDFEFF7FB",
INIT_3B => X"FFFFFFF552AA8BEF080402000087BFDF45AAD568B55AAFBFDFEF55042ABEF002",
INIT_3C => X"8516AB55A2D16ABEFFFFBFDFFF552AAAAAA007BC0000FFFBE8B55AAD168B55F7",
INIT_3D => X"00043DEAAFFAEAAAAA08556AB55A2D57FFFFF7D568B45002ABDEAAFFD16AA000",
INIT_3E => X"0000000000000000000000000000000000000FFD56AB45A2FFFDFFFAAD16AB45",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(2),               -- Port A write enable input
DIA(0)   => data_write_a(19),        -- Port A data input
DOA(0)   => data_read_a_lo_512(19),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(2),               -- Port B write enable input
DIB(0)   => data_write_b(19),        -- Port B data input
DOB(0)   => data_read_b_lo_512(19),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_20_12 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000003",
INIT_01 => X"F55FF80000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"E05022020800008400F655001FFCFF80018FA804400000000000004400000001",
INIT_03 => X"00000000000000000000000900002CC07000000000000000000000000000013F",
INIT_04 => X"68002FFE40900010000180000001FFEC0012EE0C001370F40780000000000000",
INIT_05 => X"0840000880FCBBF0100E204DF0F88311DD8005080679800000F3000029980580",
INIT_06 => X"001000030817C8E8840155FDF9001001050023F6C3C3D0F87FA19F7F011000E4",
INIT_07 => X"000000090492260800008000EE00000000000000002101FF2002C00000004018",
INIT_08 => X"2A040001071004000013FF7FCA302C0C0008214800002101554031F800000000",
INIT_09 => X"801F57F200000090000489FEC0000001EFBEF0040008023FDFC0000000004006",
INIT_0A => X"0000000008000000000000000000ADF000000200000008000008028300110230",
INIT_0B => X"0000000000000800080000000000000000000000000000000800800A40000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"000000040900005C848538000020000000800000080000020000800101FFB600",
INIT_0E => X"00800000003A010003000000000000600FFC53FF001800000002004080000000",
INIT_0F => X"0001000000007408040000004000000004E9000008020000200000000E800800",
INIT_10 => X"00200000000313100010002000008000000000129600040000400000001D0010",
INIT_11 => X"81C012060000000000218F7840000100800004000000000066C0000080080000",
INIT_12 => X"800000000017C000100000000001A800080000000001A8040000002840008185",
INIT_13 => X"0000000006F00000100200000000012600001004000000000066000000801040",
INIT_14 => X"0000200410100000000005F00000020080090A0000000085C800002000586000",
INIT_15 => X"FF00400000000000020020020001000040283024E4F2860400008000030ED080",
INIT_16 => X"00000000000000000000000000000004010201001003020200000000000127DB",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"A0700030038200010089120104D2040020000000000000000000000000000000",
INIT_1A => X"2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2C30C30C30C30C306982121A1E79E79",
INIT_1B => X"32190C86432190C86432190C86432190C86432190C86432190C86432190CB2CB",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000432190C86432190C864",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0201000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF552A974AA0004174BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA0804",
INIT_29 => X"7FFFFFFFFFFFFFFFFFFFFFFEF552E954AA000400000F7FFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E954BA007FC00BA087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974BA082E9540000",
INIT_2B => X"FFFFFFFFFF7FBFDFFF552E974BAA2FFFFE10FFFFFFFFFFFFFFFFFFFFFBFDFFF5",
INIT_2C => X"FAAD57FEAA007FFFFFFFFFFFFFEFF7FBFFF550800020BAAAD56AAAAF7FFFFFFF",
INIT_2D => X"EFF7D56AB450000021EFA2D57DE10087FFFFFFFFFFFFFEFF7FBEAB450804001E",
INIT_2E => X"000F7FFFFFFFFFFFFDFEFA2D568B550004001EFAAAEA8ABA5D7FFFFFFFFFFFDF",
INIT_2F => X"FFFF5D2E954AA080005000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFEF552A974AA0000104AAFFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"A954AA082A92428087FFFFFFFFFFFFFFFFFFBFDFEF5D2E974AA000A07000E3FF",
INIT_32 => X"FFFFFEFF7FBFFFFF552E974AA0071C50BA1C7FFFFFFFFFFFFFFFF7FBFDFFF5D2",
INIT_33 => X"EDF6FABAEBFFFFFFFFFFFFDFEFF7F5FAFC7492A974AAB6F5F8E10E3FFFFFFFFF",
INIT_34 => X"EBF5E8B550000071EFB6DF7AE921C7FFFFFFFFFBFDFEFE3F5F8F450004050AAB",
INIT_35 => X"A497FFFFFFF7FBF8FC7EBD168B450804021FFB6D57DE28147FFFFFFFFFBFDFC7",
INIT_36 => X"00000000000000000000FFFFFFFEFF7F1F8FD7AAD16AB450000001FFBEA4A8AA",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2A954AA0800174100000000000000000000000000",
INIT_38 => X"74AA002E95410A2FFFFFFFFFFFFFFFFFFFFFDFEF552E954AA0004000AAFFFFFF",
INIT_39 => X"FDFEFF7FBFFFEF552E974AA082A820AA087FFFFFFFFFFFFFEFF7FBFDFFF5D2A9",
INIT_3A => X"568A00AAFFFFFFFFFFBFDFEFFFFFFDFEF5D2E954AA0051554BA557FFFFFFFFFF",
INIT_3B => X"D16AB450804174AAFFFFFFEBAA2FFFFFFFF7FBFDFFFFFD568B55002A954AAF7D",
INIT_3C => X"57FFDFEFF7FBFFF55A2D16AB550000175EFFFFBEAA005D7FFFFEFF7FBFDFFFAA",
INIT_3D => X"0004001EFFF842AAAA087BFDFEFF7FFEAB45A2D568B550804001EFF7D57DEBA5",
INIT_3E => X"0000000000000000000000000000000000000F7FBFDFEFF7D56AB45AAD56AB45",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(2),               -- Port A write enable input
DIA(0)   => data_write_a(20),        -- Port A data input
DOA(0)   => data_read_a_lo_512(20),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(2),               -- Port B write enable input
DIB(0)   => data_write_b(20),        -- Port B data input
DOB(0)   => data_read_b_lo_512(20),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_21_12 : RAMB16_S1_S1
generic map (
INIT_00 => X"4A302428B824900A128C090A5C1800261500213C005FE812D10420054085A202",
INIT_01 => X"001FFE3440B609703B0427F801A40B8115BC4F655300340288A40D30040E4DD8",
INIT_02 => X"E00424256888D8819801000F9FFFFFFFF149FF1FCA448046C60A0D2437C517F9",
INIT_03 => X"20030640003250640003250F06002CC1740002019824E001CD357832440001FF",
INIT_04 => X"EA2C3FFD400006E04401A8837001FFFC004AEF00080B70E08FB5789421007C5C",
INIT_05 => X"00011A0C40F9FFF80920954FF0F00809DF84A0202879800000F3000029980780",
INIT_06 => X"0805984B7A1FC0A0000101FFF0480080002281F7C3C381F87C03DFFF00009004",
INIT_07 => X"B424068086A205481A60A19000908204A855B000A08A61FF20C3D004D331D340",
INIT_08 => X"1BFA0001600802000023F7FFC08D234B40C2028253000040114200000D0226C0",
INIT_09 => X"EF1F5FF054096C6ADBA169FFC202B1C1FFBEF0440021083DFFCE22DC2880E24D",
INIT_0A => X"45FF0C004041D84862A28C54518DBFF00020004C0A6044901112A0908AA0A300",
INIT_0B => X"018C241102068006C620C03882019480E63180855A492712CC01C49C20201BFE",
INIT_0C => X"08A9464116544302C02D92236488D92236488D92236488D922366446C911B210",
INIT_0D => X"08800444021048034004001890000806002804A0822189000900D80621FFBE00",
INIT_0E => X"060580261013813A2CC396506102C4053FFD5BFF00A04A00200602CA52001100",
INIT_0F => X"080C0B004C202621A85C09411500135844C196D3606941018150098404C1A304",
INIT_10 => X"B02901013416181C96C2C9C600890A2028172192C460D1820302A0130809834A",
INIT_11 => X"9C5E803408250180AC268D185DB3F4350B811068C00049A0A4AA68F05C96A001",
INIT_12 => X"002C006560138F032B1804101244C883052208209040CC849063A747512B7678",
INIT_13 => X"41401E240665750440C9488280254530314080C2C601040420352148A00501B1",
INIT_14 => X"500811204D000700114204A70422016149916011008CAA8858850B00C32591C0",
INIT_15 => X"FFC06E60AC0496022300233104663040808E991765205000070121D41D18D098",
INIT_16 => X"40100401004010040100401004010040102090010008000001C0E010020007DF",
INIT_17 => X"0100401004010040100401004010040100401004010040100401004010040100",
INIT_18 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_19 => X"FFEF9FEEFF7FFDF7FF3E3DFDF7E0000000000000000000000000401004010040",
INIT_1A => X"BEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBFFDFDFFFCF3CF3F",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFEFF7FBFDFEFF7FBFDFEFBEF",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000FFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0001000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E954AA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0004",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA0004154BAFFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"52E974BA0804000AAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0004174BAFF",
INIT_2B => X"FFFFFFFFFFFFFFFFEF552E954AA000400000007FFFFFFFFFFFFFFFFFFFFFFEF5",
INIT_2C => X"A082E95400007FFFFFFFFFFFFFFFFFFFFDFEF5D2E974BA002E97400007FFFFFF",
INIT_2D => X"FFFFFBFDFEF5D2A954AA002E974BA087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFBFDFFF5D2E954BA007FC00BA5D7FFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA000002000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080005000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"A974AA0000104AAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974BA0000174AAFFFF",
INIT_32 => X"FFFFFFFFFFFFDFEF552E954BA080A000AAE3FFFFFFFFFFFFFFFFFFFFFFFEF552",
INIT_33 => X"02A95400087FFFFFFFFFFFFFFFFFFBFDFEF5D2E974AA000A07000007FFFFFFFF",
INIT_34 => X"F7FBFDFFF5D2A954AA082A924281C7FFFFFFFFFFFFFFFFFFBFDFEF5D2A974BA0",
INIT_35 => X"A557FFFFFFFFFFFFFFFF7FBFDFFF552E974BA0020924BA1C7FFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000E3FFFFFFFFFFFFFFEFF7FBFFFFF552E974AA0071C50B",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0000020000000000000000000000000000",
INIT_38 => X"74BA0000174BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954AA080017410FFFFFF",
INIT_39 => X"FFFFFFFFFFDFEF552E954AA0004000AAF7FFFFFFFFFFFFFFFFFFFFFFFEF552A9",
INIT_3A => X"E95410087FFFFFFFFFFFFFFFF7FBFDFEF5D2A954BA082E800AAA2FFFFFFFFFFF",
INIT_3B => X"FBFFFFF552E954BA002E97410087FFFFFFFFFFFFFEFF7FBFDFFF5D2A974AA002",
INIT_3C => X"57FFFFFFFFFFFDFEFF7FBFFFEF552E974AA082A820AA557FFFFFFFFFFFFFEFF7",
INIT_3D => X"5D2E954AA0051554BA5D7FFFFFFFFFBFDFEFF7FFFFFEF5D2A974BA0000020AA5",
INIT_3E => X"0000000000000000000000000000000000000AAFFFFFFFFFFBFDFEFFFFFFDFEF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(2),               -- Port A write enable input
DIA(0)   => data_write_a(21),        -- Port A data input
DOA(0)   => data_read_a_lo_512(21),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(2),               -- Port B write enable input
DIB(0)   => data_write_b(21),        -- Port B data input
DOB(0)   => data_read_b_lo_512(21),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_22_12 : RAMB16_S1_S1
generic map (
INIT_00 => X"5290F4CDE914905A14A43D33F488243E17122300F55FEB189B343A1140548380",
INIT_01 => X"A54007B259F6A975386262000C344BA9573C6FF57B18A5FB0ABFCD3C2C5F4F0C",
INIT_02 => X"021DFF8C38B3C009D203551040030071869D0040180AA2DC53DB89BEA8204001",
INIT_03 => X"2603475A969D0475A969D0460EAA401005111011BD506954EDB40F5EF41434C0",
INIT_04 => X"922D9002100ED69E443D988B0D5400103E48003D0800011E803B06B5B9125A15",
INIT_05 => X"281B5A0C06000408F4DF9422010D8802022F2124A8022492580040440002021C",
INIT_06 => X"F780C4C052881ADA0E05440205DA50930FA182010004700083E220800440B588",
INIT_07 => X"049D028B93FB561833D8094A02F5EA92FD7247E10305C40040D136E6A023F7FC",
INIT_08 => X"00028241680A0E002A9400803A884B5B5206B7C2E53CA25144009007A64EBD64",
INIT_09 => X"41008810240240C6694008010392354010000560141801002028A83D2A08E06D",
INIT_0A => X"34000000848BCA6902A29C54539C020E11810098D4067EFF9FF284D483E2AB41",
INIT_0B => X"500001840000C80B410014088040F4A944B1AA313C0022AA0011C0DC00028001",
INIT_0C => X"80B14004D158C8CA24A1C2A870AA1C2A870AA1C2A870AA1C2A872550E1543800",
INIT_0D => X"80A14050A01509E050854498B5281A1C34E506A2C6898B52A154DAC6B6000850",
INIT_0E => X"0B03001A483A4146603050080410089180008800143D83888281A2034A850142",
INIT_0F => X"A4160600349075238473F1210006133835E92273612B3482C090068A0E84AC56",
INIT_10 => X"30060181BA1B13959DC08DA902458870201970B29602562B0581200D141D0959",
INIT_11 => X"E042021C040D0152C8058B3840F044708E7E1C20A0106EA166C13AFC14AA3804",
INIT_12 => X"080E004B0C17C1439A9838301DC1A8438EA32C009DC1A8255300650458A1D588",
INIT_13 => X"018010E186F110A908E3A8CB0026C9A610A908E6A60F0807626610E160589C4C",
INIT_14 => X"2A701667334005800B1605F043858125E0D04110408D2485CA034681E43A1E40",
INIT_15 => X"00646002304244A91102C93A2D608D2A258DF8034188200C050171A41108F084",
INIT_16 => X"110441104411044110441104411044110466C440446CA06951D4EA8010009804",
INIT_17 => X"0040100401004411044110441104411044110441104411044110441104411044",
INIT_18 => X"0401004010040100401004010040100401004010040100401004010040100401",
INIT_19 => X"F7DFBFDEFE8FF1F7DEBDDF7DF7D05122890000000003FFFFFFFF900401004010",
INIT_1A => X"9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7BFFDFD7DDDF7DF7D",
INIT_1B => X"F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE79E7",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000003F9FCFE7F3F9FCFE7F3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA000400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0800",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000002000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2A954BA000015400FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080402010FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2A954BA0004154BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A0004174BAFFFFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0800154AAFFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF552A974AA0000174BAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974A",
INIT_2E => X"000007FFFFFFFFFFFFFFFFFFFFFFEF552E974BA0804000AAA2FFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080400010000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E954AA080005000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000402010FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2A954BA000417410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"804154BAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974BA0000174AAFFFFFFFFFFF",
INIT_34 => X"FFFFFFFEF552A974AA0000104AAE3FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0",
INIT_35 => X"AA2FFFFFFFFFFFFFFFFFFFFFFFEF552E954BA000E124BAE3FFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000007FFFFFFFFFFFFFFFFFFFFDFEF552E954BA080A000A",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804000100000000000000000000000000",
INIT_38 => X"54AA000400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2A954AA080017410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"0174BAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A954BA000415400FFFFFFFFFFFFF",
INIT_3B => X"FFFDFEF552E974AA0804174AAF7FFFFFFFFFFFFFFFFFFFFFFFEF552A974BA000",
INIT_3C => X"2FFFFFFFFFFFFFFFFFFFFFDFEF552E954AA0004000AAA2FFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2A954BA082E800AAAAFFFFFFFFFFFFFFFFFFFBFDFEF5D2E954BA002A820BAA",
INIT_3E => X"0000000000000000000000000000000000000087FFFFFFFFFFFFFFFF7FBFDFEF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(2),               -- Port A write enable input
DIA(0)   => data_write_a(22),        -- Port A data input
DOA(0)   => data_read_a_lo_512(22),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(2),               -- Port B write enable input
DIB(0)   => data_write_b(22),        -- Port B data input
DOB(0)   => data_read_b_lo_512(22),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_23_12 : RAMB16_S1_S1
generic map (
INIT_00 => X"EF20906D902424807BC8241BC81801B97D38AD3C0800103362A6741C80A12A02",
INIT_01 => X"001FFF8409F089003B4422000D80C80106804A7951C5B9D1C828043EA28838F9",
INIT_02 => X"E01CEE21649C82C40800000F9FFEFF8E72CA7F5FC2E22809925A0D3611C877F8",
INIT_03 => X"24000400402670400402670D48222DC1764446838624000080007460C40001BF",
INIT_04 => X"68403FFC020560E0443E21037C01FFFC0002EE00628BF0E02FAD781014085014",
INIT_05 => X"0112000202FBFFF00920017FF0F0628BFF8488890979800002F702002BB807A0",
INIT_06 => X"EF85788B681FC000000001FFF0010000000001F7CBC385F87C0BFFFF20040001",
INIT_07 => X"F6E200000000C1440E3AE408009120071070FA07A1CB23FFA403F0C4D23BF7C0",
INIT_08 => X"0BF87CA400804000003FF7FFD8880A034AC09662305AB10555421006891A1089",
INIT_09 => X"BE1F5FEA10092C0896A243FFC0008087FFBEF2000000001DFFC612C0C0400100",
INIT_0A => X"41FF0C2060501000600000000001BFFA800808189A657EF81DD0C00079CC8001",
INIT_0B => X"018C24110A860006C620C0312241C482B20400CC52492710CC80060020A81BFE",
INIT_0C => X"0C08866907048320C20C10030400C10030400C10030400C10030400608018210",
INIT_0D => X"040002000041500300100040000500C000801000C02400000952800001FFBF04",
INIT_0E => X"FC850015385380380CDB86106502C5043FFD5FFF00A04BC010A7724B10000800",
INIT_0F => X"89F90A002A70A710A51C01C05904014861433602A1CAF13F2110055614C72FC0",
INIT_10 => X"E02D02001C1E14981B43253EE50C8220180F1082E06397E07E42200AAC298E57",
INIT_11 => X"8421802400A90022B0070FAE18019214A380344920080B21A58B02AC60BACDF0",
INIT_12 => X"0A2A000C480B0704B54028101AC49C84BB4100009AC49C80857A82D20CE8CB22",
INIT_13 => X"01E00C8103416445C12ED0400027C5292445C12D500B0005A62D344CB241D095",
INIT_14 => X"132C907425604680038706A35132C94BDD011010404428886AC91B11311C8280",
INIT_15 => X"FF000470BE0692020328CA0028042054A92771C50FC070110001C1680809591D",
INIT_16 => X"00802008020080200802008020080200800800200200000000000008004807DF",
INIT_17 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_18 => X"8020080200802008020080200802008020080200802008020080200802008020",
INIT_19 => X"0000000000000000000000000000000000000000000000000000008020080200",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080002010FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974AA000400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000400010FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974AA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080000010FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E954AA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954A",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA000015400FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080002010FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974AA000400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000402010FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E954AA080005000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA080407000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA00041741",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080000010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000402010FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2A954AA080002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954AA080017410FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"552A954BA000415400F7FFFFFFFFFFFFFFFFFFFFFFFFF552A954BA080015410F",
INIT_3E => X"0000000000000000000000000000000000000F7FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(2),               -- Port A write enable input
DIA(0)   => data_write_a(23),        -- Port A data input
DOA(0)   => data_read_a_lo_512(23),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(2),               -- Port B write enable input
DIB(0)   => data_write_b(23),        -- Port B data input
DOB(0)   => data_read_b_lo_512(23),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_24_12 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100600007FFF000080108004000800020000840041000080808",
INIT_02 => X"FC5CA803400EB8209000000F9FFEFF8E7240FF1FC22409EA04018E50074017F0",
INIT_03 => X"11100400000000400000000D00002CC07400000090C080019001010A000001BF",
INIT_04 => X"68003FFC00040000000000008001FFFC0002EE00000370E007A100000000E468",
INIT_05 => X"0000000000F8BFF00920004DF0F00001DF8000000079800000F3000029980780",
INIT_06 => X"6E461803081FC000000001FFF0000000000001F7C3C380F87C019FFF00000000",
INIT_07 => X"600C2400013649609C8000980040814210254000A00B21FF2003F2A80D500000",
INIT_08 => X"0BF80000000000000003F7FFD88D2B4A02C0940062EC2804001610020408178B",
INIT_09 => X"8E1F5FE010092C0892A041FFC0000001FFBEF0000000001DFFC002C000000000",
INIT_0A => X"41FF0C0000000000600000000001BFFA0000005501AA00000CE2000009400000",
INIT_0B => X"018C0411020600048620C030020502000200000400490510CC00040020201BF4",
INIT_0C => X"0808064106040300C00C10030400C10030400C10030400C10030400608018210",
INIT_0D => X"0000000000004003000000000000001200580000000000000000000001FFBE00",
INIT_0E => X"0086C022005381380FDB96516140C6043FFD5BFF000041000000004110000000",
INIT_0F => X"80010D804400A7240C840C201D0210840043B4804012500021E0088014C04940",
INIT_10 => X"4109038041021C980200D06410C1924030008142E06024A00043C01100298092",
INIT_11 => X"587CC200002100C14428090A1D02348190814C09C010104025AA40041A0D8005",
INIT_12 => X"022E0030300B0E46177004208000D8C61D7004300000D884817B00011306B2D9",
INIT_13 => X"01E003060344710009875C018100013831000985DC000C20003C310006143B70",
INIT_14 => X"4001850EDC004780144806A64400186CBF8961104000C3807884000846EB9500",
INIT_15 => X"FF0006E08C063C0220002201490418082010A57263E0100008000290161E711C",
INIT_16 => X"00000000000000000000000000000000000000000000000000000000000007DF",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"F2D0AEEAF6E7CC1132CDB4441990000000000000000000000000000000000000",
INIT_1A => X"BEFBE79E79E79E79E79EFBEFBEFBEFBEFBEF9EF9EF9EF9EFA69861219575D75F",
INIT_1B => X"783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1EFBEF",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000783C1E0F0783C1E0F0",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0201000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A000400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA000400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000400000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402010000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"00002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080002010FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000400010FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA00040000",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020100000000000000000000000000",
INIT_38 => X"74BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"000010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA000002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974AA000402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000002010F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(3),               -- Port A write enable input
DIA(0)   => data_write_a(24),        -- Port A data input
DOA(0)   => data_read_a_lo_512(24),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(3),               -- Port B write enable input
DIB(0)   => data_write_b(24),        -- Port B data input
DOB(0)   => data_read_b_lo_512(24),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_25_12 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100200002000000080100004000000020000800041000080808",
INIT_02 => X"FC400086000000800000000F9FFEFF8E738FFF1FC204010000000111568DD7F8",
INIT_03 => X"00000400000000400000000D00002CC4740000008000000080000000000001BF",
INIT_04 => X"68003FFF64A564AC000000000001FFFE0082EF00010370E007A1000000004000",
INIT_05 => X"0A00040148F8BFF80920804DF0F00101DFC040000079C92484F30499299837C1",
INIT_06 => X"66041803081FC0E0801101FFFD000E41002299F7E3C380F87C019FFF81200096",
INIT_07 => X"000000080480AE00000080000000000000000000A00B21FF2003E00000000000",
INIT_08 => X"1BF80000400A02000003F7FFFA0008000200A0400008A0000014100200081000",
INIT_09 => X"8E1F5FFA53EFBCACB2E369FFE0010001FFBEF80C40630C7DFFEEBAF000800202",
INIT_0A => X"41FF0C0600000000600000000001BFFE00301000000000000CC020000140000C",
INIT_0B => X"01DCCC31222730A49620C030020100000200000400490D10EC00040220201BF4",
INIT_0C => X"0808064106240300C00C10030400C10030400C10030400C10030400608018210",
INIT_0D => X"0883044582114013412080000000000000000000000000000012800001FFBE00",
INIT_0E => X"00040020000180380FC386106140C6043FFD5BFF00A04B80608003CB120C1106",
INIT_0F => X"0000080040000200040400000100000000009480000240000100080000400900",
INIT_10 => X"0001000000000808000000240000020000000100006004800002001000008012",
INIT_11 => X"0001001808220000002004001900000080800008000000000022400000088000",
INIT_12 => X"0010000000000E00110000000000408009000000000040808063004000008200",
INIT_13 => X"6000000000046100000240000000001021000004400000000010210000001010",
INIT_14 => X"4000000404000800000000060400000088000001800000001084000000088000",
INIT_15 => X"FF800C608C041002000002000006100000002100000000180600000000100018",
INIT_16 => X"4110441104411044110441104411044510629041040D180400000010028047DF",
INIT_17 => X"1104411044110441104411044110441104411044110441104411044110441104",
INIT_18 => X"1044110441104411044110441104411044110441104411044110441104411044",
INIT_19 => X"FBA2894A196A8C5A2932EC15DA080800002FFFFFFFFFFFFFFFFFC11044110441",
INIT_1A => X"2492492492492492492410410410410410410492410492412000531215A69A6B",
INIT_1B => X"158AC562B158AC562B158AC562B158AC562B1588C46231188C46231188C49249",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000B158AC562B158AC562B",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080000010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000010FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08000000",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(3),               -- Port A write enable input
DIA(0)   => data_write_a(25),        -- Port A data input
DOA(0)   => data_read_a_lo_512(25),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(3),               -- Port B write enable input
DIB(0)   => data_write_b(25),        -- Port B data input
DOB(0)   => data_read_b_lo_512(25),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_26_12 : RAMB16_S1_S1
generic map (
INIT_00 => X"E9264EAB20190CA3BA4997AA9002AE9C001006B0778015CFA17E0811039879C7",
INIT_01 => X"2FFFF9BB1F773C7F9BB07DFFFDD863FC5FFF3FEFFBBF9FFB22FFFBC7B9F30686",
INIT_02 => X"E06CCC62052E708180F6FFBFFFFCFFFFF9C7FF7FC24332E642090000074037F6",
INIT_03 => X"428003739CD9863739CD9869FE2B7DEAF300029E4E300DFE69A6E644E6FF473F",
INIT_04 => X"7C2FEFFFF5BA124F003DD31EAFFFFFEE9FF7EE6F4C0770FFD7DC7CA53997B2B1",
INIT_05 => X"DFFB5421C1F8BBFAFDBFFACDF0FFCC05DDDBFF3690F9EDB7F5F7AFF639BD7DE3",
INIT_06 => X"EFD044ABC817C3E3A74667FDFFB6FF5727CC3BFEF7C3FAF87FF59F7FFBFEF69F",
INIT_07 => X"00003002132462052E708180EF060C18E5BEFB051225CDFF7002C4EEDE77F6E0",
INIT_08 => X"3FFF7D5000EC75088ED3FF7FC8790E46426CE06CB1F8E041051831FA3068D77E",
INIT_09 => X"C05FD7FF9BEFBDCEFBEE59FEF44F6603EFBEFAFCC2E35E7FDFD147CCF3F583FA",
INIT_0A => X"67FF1C7FBFADEB31E35768E8ED6BFDF3EB3EBF9DDBCE7FDC1DF8A760F3EACC02",
INIT_0B => X"5BDDCC3B336F7C548667D47B7737AF3FD62601EDC25B3533DCEB07F262213FFC",
INIT_0C => X"5F9A06E19F4D93A0EA0F78C35E30D78C35E30D78C35E30D78C35E986BC61AE31",
INIT_0D => X"5FD7AFEFDFFAF59B6FF28FE1D80D73D840607307DCFE1D80EF69A004DFFFF7FF",
INIT_0E => X"0004001F8041897B2FFFC6D86D70CE04FFFFF3FF1F5F5475BD7F72E4D75EBFAF",
INIT_0F => X"F60008003F008237B0040A00010003E020023E0201F45EC0010007E01047D17B",
INIT_10 => X"00010001DC0004C81003DE050A700200001DC0006863E8BD8002000FC0208FA2",
INIT_11 => X"2200E400002801E1A00004C21C0206F60081800800007B00010F02007EC09A0E",
INIT_12 => X"0880007E000807C7C1A612001E0015C7C19C22001E0015C59DFE82011A311AA0",
INIT_13 => X"00001BC00101F60409F0670840070809760409F06984800780097604067D0010",
INIT_14 => X"81019F40042100001F800203D81019EC085614000085C80023D81009CF008A74",
INIT_15 => X"FF802FFDFFAFD082003B032FB987E04021D481D4000819060801E0D00001231D",
INIT_16 => X"EBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEFFBFBFBFBBFCFBB0FFDFEFFEF2DFFFFFB",
INIT_17 => X"BFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAF",
INIT_18 => X"FAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFE",
INIT_19 => X"475B15BCF491E166CC8553F86EDB5C88646FFFFFFFFFFFFFFFFFEBFAFEBFAFEB",
INIT_1A => X"861861861861861861861861861861861861869A69A61861AFBD54D5F871C71D",
INIT_1B => X"984C26130984C26130984C26130984C26130984C26130984C26130984C261861",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000984C26130984C26130",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040201",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(3),               -- Port A write enable input
DIA(0)   => data_write_a(26),        -- Port A data input
DOA(0)   => data_read_a_lo_512(26),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(3),               -- Port B write enable input
DIB(0)   => data_write_b(26),        -- Port B data input
DOB(0)   => data_read_b_lo_512(26),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_27_12 : RAMB16_S1_S1
generic map (
INIT_00 => X"00080A40000A41248002029000050A088000008242A0004404480002000A1155",
INIT_01 => X"2FFFF1C11F781C129C107DFFFE0860941E81258CA2B71C2220EC1B86E1A00002",
INIT_02 => X"E1000000810000014400FF6FFFF0FFFFF8007F1FC21110005080200000221FF0",
INIT_03 => X"4080026318C18226318C1821302232EAE00002BE001115FE48620040840A863F",
INIT_04 => X"643D4FFC2530000F003D821C0BFFFF8E9EF79E6D440748FED70060842105B0B0",
INIT_05 => X"D6F39020D1F8A3FAFDBFBACDC8FDC405D1DB7F1490E5EDB7D5CBADB2385D79C3",
INIT_06 => X"6FE000A38007C3032646EFF1F0B6FF46A78C39F8E723F2E47FE59C7F9ADA2612",
INIT_07 => X"00002820000000810000014401060C180190310540118DFF1000C0849673F6C0",
INIT_08 => X"3FF779100062B12A8EC3F47FC80208808210880C00082050000110023068D030",
INIT_09 => X"005F07E09BFFBD07FBAC09F8E42922038F7DF8BEC2E39C5F1FD047CEF1B582D8",
INIT_0A => X"63FF5D5F9FADE911E81C09818109E1F16B16B71092CE7ED81CF403601228C402",
INIT_0B => X"1BFDCC39732F3554866AD57C37BEAF1C152201A4C05B7531D56B05B06A213FF8",
INIT_0C => X"5BCA06F18FC59380F00E34430D10C34430D10C34430D10C34430F0861A2186B5",
INIT_0D => X"5B56ADAB5FAAE58B2F628EA0C80FA3F04040510768EA0C80CC61A0044DFFC6EB",
INIT_0E => X"0004001D800188792CE79715710AE4047FFD23FF315D54358D593474955AB6AD",
INIT_0F => X"520008003B000297B0040200010003E020001F0201E44A400100076000579129",
INIT_10 => X"00010001DC00004A10035E0408300200001DC000086BC8948002000EC000AF22",
INIT_11 => X"02002400002801E1A00000C01E0202F60080800800007B00000782006EC0820A",
INIT_12 => X"0080007E000006A7C10602001E0001A7C10C02001E0001C18DE282010A311AA0",
INIT_13 => X"00001BC00000FE0401F04300400708007E0401F04180800780007E04047D0010",
INIT_14 => X"81011F40040100001F800002F81011EC080604000085C80001F810094F008034",
INIT_15 => X"FF800C6DDDAFD082001B03249887E04001D481D4000009020801E0D00001021F",
INIT_16 => X"AB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6BF1EBDABD8E270BF84A25C6ACB777E3",
INIT_17 => X"B6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6AD",
INIT_18 => X"6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADA",
INIT_19 => X"490E2168100481CA860402104A471688747FFFFFFFFFFFFFFFFFAB6ADAB6ADAB",
INIT_1A => X"000000000000000000000000000000000008200000000000200072F210000001",
INIT_1B => X"05028140A05028140A05028140A05028140A0500804020100804020100800000",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000A05028140A05028140A",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040201",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(3),               -- Port A write enable input
DIA(0)   => data_write_a(27),        -- Port A data input
DOA(0)   => data_read_a_lo_512(27),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(3),               -- Port B write enable input
DIB(0)   => data_write_b(27),        -- Port B data input
DOB(0)   => data_read_b_lo_512(27),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_28_12 : RAMB16_S1_S1
generic map (
INIT_00 => X"02200AA400180030808802A900002A08001280A08A801044104A1000001818C3",
INIT_01 => X"0AA00011460214428114180000882214413D0A71592A01D92213D28005210202",
INIT_02 => X"0451110A012100884000AA30200000000C100040104112101100008888200000",
INIT_03 => X"448000318C52A20318C52A20148810200111100C211004AA00034204200A2200",
INIT_04 => X"04004001001A90110000121402AA0000003C00000500000040080421080D0080",
INIT_05 => X"4060000C8001000000002E000000050000001610300000010000802202040012",
INIT_06 => X"1000002080001111001222000425A1040026A008000000000000000009328280",
INIT_07 => X"2491008A00491201210088400122448908A20402000408001000040820000000",
INIT_08 => X"20058310402A160026500000028040101004200C840082115554000112244814",
INIT_09 => X"4140000800000060000720000102028000000490160801020002200011100010",
INIT_0A => X"020000081B34211082B694D4D294000020020381040000000200032040004400",
INIT_0B => X"4800210C19808400500010009110091500020B408810000100200020408B0000",
INIT_0C => X"01028000080118020023604858121604858121604858121604858090B0242C00",
INIT_0D => X"010000800920040804020A6058003108402043058C460580653020005A004039",
INIT_0E => X"00000002800008014004104104420A00C000200005000010040A0020CC000200",
INIT_0F => X"520000000500000010000200000000000000280000040A40000000A000001029",
INIT_10 => X"00000000000000C0000002000830000000000000480008148000000140000020",
INIT_11 => X"020024000000000000000440000000020000800000000000000C00000040020A",
INIT_12 => X"00800000000001804006020000000500400C0200000005400A90000000100000",
INIT_13 => X"0000000000018200001003004000000142000010018080000001420000200000",
INIT_14 => X"8000080000010000000000018800008000060400000000000310000008000034",
INIT_15 => X"000002040080000000110006B081400000400000000009020000000000002200",
INIT_16 => X"802008020080200802008020080200802101210810C39A66A90A85420413A820",
INIT_17 => X"0200802008020080200802008020080200802008020080200802008020080200",
INIT_18 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_19 => X"DE21102C110A00246972BD89A40A0C22E1000000000000000000002008020080",
INIT_1A => X"2082082082082082082082082082082082082082082082080D35050758C30C31",
INIT_1B => X"0582C160B0582C160B0582C160B0582C160B0580C06030180C06030180C08208",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000B0582C160B0582C160B",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(3),               -- Port A write enable input
DIA(0)   => data_write_a(28),        -- Port A data input
DOA(0)   => data_read_a_lo_512(28),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(3),               -- Port B write enable input
DIB(0)   => data_write_b(28),        -- Port B data input
DOB(0)   => data_read_b_lo_512(28),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_29_12 : RAMB16_S1_S1
generic map (
INIT_00 => X"79964E4BA01DACAB9E659792D00AAE160002829C7FDFEFCEE97C2815039D70C3",
INIT_01 => X"0ABFF9AB0775343F9AB01DF80D5821FC0FFF3FEFD1AF9FF1207FFBC7B9720586",
INIT_02 => X"002CCC60050E700080F6AAA7BFFC007189C7FF2FC00330E602800000074037F6",
INIT_03 => X"468003210868A63210868A68DA017D207200021C4E200CAA6186A40042FF4300",
INIT_04 => X"7C2FE002F0900001003C5316A6ABFFE21F36E02F0D03701F47D41800109FB281",
INIT_05 => X"4979440580F9B808F49F6A4DF00F8D01DC4B97369078249370F482E62BA41462",
INIT_06 => X"B250442BC81001E1870223FC0BF7F11507C423FE33C078F803F19F00E936721D",
INIT_07 => X"00011080012460050E700080EF020408EC8CFA01122149FF700200665A35D260",
INIT_08 => X"2BFD055040A452000443FF00007906464068406C31F84000000831FA1028575A",
INIT_09 => X"805FD017102690AA694551FE30444681E0820AD40201423FC00122C493500172",
INIT_0A => X"0600002AFFBE2330815568A8AD6ABC02A02A0B0CCB463B4C0748A720B1EA4C00",
INIT_0B => X"0850400A11414C005005000B51158936D20601A98A10200308A002E240010BFC",
INIT_0C => X"05928020194918A22A2268C81A32068C81A32068C81A32068C81A99034640C00",
INIT_0D => X"058102C48970541944B20FA1580561D040406305587A158046282000DBFFF13D",
INIT_0E => X"000000028040890327DCD28928324400DFFFF0001F1F0050342D42A086040B02",
INIT_0F => X"F60000000500802010000A000000000000022A0000141EC0000000A01000507B",
INIT_10 => X"00000000000004C0000082010A700000000000006800283D80000001402000A0",
INIT_11 => X"2200E4000000000000000442040004020001800000000000010D000010401A0E",
INIT_12 => X"08800000000801C040A6120000001540409C2200000015441DAC800010100000",
INIT_13 => X"0000000001019600081027084000000956000810298480000009560002200000",
INIT_14 => X"800088000021000000000201D800088000561400000000002358000088000A74",
INIT_15 => X"00802594A282C0000033010FB181E00020400000000819060000000000002305",
INIT_16 => X"C0B02C0B02C0B02C0B02C0B02C0B02C4B12B312912831A27FCFE7FFB175B6FF8",
INIT_17 => X"0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02",
INIT_18 => X"B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C",
INIT_19 => X"BBCF9F96EE7FFDF7FE783FFDFFEA0C00602FFFFFFFFFFFFFFFFFC0B02C0B02C0",
INIT_1A => X"EFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEEBAEBAEBAEBAEBBFFDF9FBEFFFFFFE",
INIT_1B => X"BFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFBEFB",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000FBFDFEFF7FBFDFEFF7F",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(3),               -- Port A write enable input
DIA(0)   => data_write_a(29),        -- Port A data input
DOA(0)   => data_read_a_lo_512(29),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(3),               -- Port B write enable input
DIB(0)   => data_write_b(29),        -- Port B data input
DOB(0)   => data_read_b_lo_512(29),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_30_12 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"F7FFBFFEFF9FE1F7FFBFFFFDFFD0000000000000000000000000000000000000",
INIT_1A => X"9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7AFBD75F5FDF7DF7F",
INIT_1B => X"F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE79E7",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000003F9FCFE7F3F9FCFE7F3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(3),               -- Port A write enable input
DIA(0)   => data_write_a(30),        -- Port A data input
DOA(0)   => data_read_a_lo_512(30),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(3),               -- Port B write enable input
DIB(0)   => data_write_b(30),        -- Port B data input
DOB(0)   => data_read_b_lo_512(30),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_31_12 : RAMB16_S1_S1
generic map (
INIT_00 => X"129000008004A00804A40000400800020000000C005FEA005800200400050100",
INIT_01 => X"255FF18019700810180065FFFC0040801E80258CA2951C2200EC0906A0804140",
INIT_02 => X"E0000000000000011000550FDFF0FFFFF0007F1FC200000044000000000817F0",
INIT_03 => X"0000024210A30024210A3001002220C06044469200040154482000408400043F",
INIT_04 => X"602D0FFC2420000E003D80080955FF8E1ECA8E2D400340FE870060842100B030",
INIT_05 => X"0213100040F8A3F8FDBF944DC0FDC001D1CB6904A061EDB6D4C30490281831C1",
INIT_06 => X"6FC000830007C202060445F1F0D25E4207A099F0E303F0E07FE19C7F80402412",
INIT_07 => X"0000200000000000000001100004081001103107000185FF0000C0849673F6C0",
INIT_08 => X"1BF27A00000000000883F47FC800080002008000000820440000100220489020",
INIT_09 => X"011F07E013EFBC06FBA009F8E00120038F3CF82C44630C5D1FC002CCE0808248",
INIT_0A => X"61FF0C06C48BC801600000000001A1F00110101092CE7ED81CF0004012288000",
INIT_0B => X"11DCCC31222730048620C4382204A608142002A440492530C401049020221BF8",
INIT_0C => X"0888066187448380E00C10030400C10030400C10030400C10030600608018210",
INIT_0D => X"080204010200418301208480800D02D00040100240A808008840800405FF8640",
INIT_0E => X"0004001D000180780CE386106100C4043FFD03FF101D40008001304018081004",
INIT_0F => X"000008003A000217A0040000010003E02000160201E040000100074000478100",
INIT_10 => X"00010001DC00000810035C0400000200001DC0000063C0800002000E80008F02",
INIT_11 => X"00000000002801E1A00000801C0202F40080000800007B00000302006E808000",
INIT_12 => X"0000007E00000607810000001E000087810000001E000081846282010A211AA0",
INIT_13 => X"00001BC00000740401E0400000070800340401E04000000780003404045D0010",
INIT_14 => X"01011740040000001F8000025010116C080000000085C80000C8100947008000",
INIT_15 => X"FF800C609C06D082000A03200806A040019481D4000000000801E0D00001001D",
INIT_16 => X"010040100401004010040100401004010060C040040C200950402090128057C3",
INIT_17 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_18 => X"0040100401004010040100401004010040100401004010040100401004010040",
INIT_19 => X"00000000000000000000000000001000802FFFFFFFFFFFFFFFFF810040100401",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(3),               -- Port A write enable input
DIA(0)   => data_write_a(31),        -- Port A data input
DOA(0)   => data_read_a_lo_512(31),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(3),               -- Port B write enable input
DIB(0)   => data_write_b(31),        -- Port B data input
DOB(0)   => data_read_b_lo_512(31),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_0_11 : RAMB16_S1_S1
generic map (
INIT_00 => X"ED39BA795990D275FB4A6E96ACC4731DEA4598B0AFB54867F6EE4618C3749803",
INIT_01 => X"8AA0047D8607944AC7DA180001ECA2444042106208408208C20022E9173734B3",
INIT_02 => X"1A7DDD79F9A73E6CCA7DAAF00001000008478020113D98E382FEDF333027C80F",
INIT_03 => X"75D341110C58F31110C58F32A208921F8051500147A0E4AB3493FB3A01EBE240",
INIT_04 => X"86424001531009B100425A97B2AA0001E03501D0A39C8F0078420001106D0C4C",
INIT_05 => X"BCC8CA2EBF03400700402BB20F00239E20341699198600000B08694B16434804",
INIT_06 => X"103FB860B2800161F8432200012DA185F80F24081C3C0707800E600056881308",
INIT_07 => X"B24197ABCDA467F9A73E6CCAFDC3870EEEEC44E2BDFE220094D03022210C011C",
INIT_08 => X"240581B5695EAA80262C080032BF07C7C1FC3F8E94F65B11555EAFFC1C306758",
INIT_09 => X"7E40000BEC004170040DB60017FED1CC0001045002984202003DB931192D60A5",
INIT_0A => X"120071411A74315881A28C141118000C5A85A60444210123820B43B40804674D",
INIT_0B => X"0820008E514045BB514F0106D1D8599581D3A958BC104A89215AC14C48898403",
INIT_0C => X"C261C01C48B1584A0CA3E2687A9A1E2687A9A1E2687A9A1E26870CD061343885",
INIT_0D => X"D274E93A758FA8683AC54B287522E10A74AF4AA59C568752662F5AC218000002",
INIT_0E => X"FF83C002783A0904231C70470C7E0B92800224008AE09FAD4BD48D1FC5D3A4E9",
INIT_0F => X"5BFF078004F075885DFBF7E15C06101C55E921F1F80FAB7FE0F0009E0E903EAD",
INIT_10 => X"F12E0380231F13978FF023FAFDBD9870380230F2D6081F56FFC1E0013C1D207D",
INIT_11 => X"DE7F263C0C8700125C0F8F3C43F1F10BBF7EFC61E01804E1E6C8F8FE807F67FB",
INIT_12 => X"02BE00017C17C1007E5E2E3081C5AC007E6F0E3081C5AC44418D65FE45DEE55B",
INIT_13 => X"61E0042786F103E9F01F9BC3C120C5A703E9F01F978B8C20666703E9F8A0FFED",
INIT_14 => X"FA7E283FFB414F80005F05F10FA7E283F78F6511C048278DCA174FF038FF15B4",
INIT_15 => X"0066A20B61692F293185D8D724E15D3FCC6B7C236FE0691B0700132C1F0EF880",
INIT_16 => X"3A4E93A4E93A4E93A4E93A4E93A4E93A4F942F92E9628540AD2A91442525A000",
INIT_17 => X"A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E9",
INIT_18 => X"4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93",
INIT_19 => X"55F3898E09B56C74DAB15D1CF13501AA495000000000000000003A4E93A4E93A",
INIT_1A => X"082082082082082082082082082082082082082082082082082084E41DC71C71",
INIT_1B => X"E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F82082",
INIT_1C => X"FFFFFFFFFFFFFFF94A5294A5294A5294A5294A52800003E1F0F87C3E1F0F87C3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"3060C183060C187FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"BDEBA0000000000000000000000000000000000000000000003060C183060C18",
INIT_28 => X"168ABA002E82145085155545F7AA975EFFFAABDE00FFAEBDFFF5D2EAAAAAF7AE",
INIT_29 => X"7FFFE10005542145557FD5545FF8000155087FC0155F7D168B55007BFDF45085",
INIT_2A => X"7FFC0010080017555555568AAAFFFFD7545AA8028A00A2802AABAFF8028BEF5D",
INIT_2B => X"FF842AABAA2AE95545FFD168ABAF7AEAAAAAA2FFFDF4500043FE105D2E954BAF",
INIT_2C => X"5007FD7400550415410002E974BA5D5168A00A2D142155005142010FFAE820AA",
INIT_2D => X"FFF780000BA007FE8AAAFF803FFFF5D2A821550000000BA007FD55FF5D7FC014",
INIT_2E => X"000AAFBEAA00007BFDFFF082EBDF455D5142000082E82145FFD17DFEFFFD168B",
INIT_2F => X"DFD75D2AA8A80EA8E2FE3F000000000000000000000000000000000000000000",
INIT_30 => X"68B551475FAF6D1C556F0AA1C24AABEA495FC716F002A975FFE3AA95E00EBAEB",
INIT_31 => X"42A0070071C50BAFEF1FAE0016D56A16D557BC257D415E0216FA3F1E8FC0145B",
INIT_32 => X"8010E004924874825D7FEAA85487FD24AFE3D02DAAAE12BD5545A2803AA00005",
INIT_33 => X"120155EA568E870BAEB8A05A2AEA8B50F55A2F150005A3A438BD04AFAB8F550A",
INIT_34 => X"545E055FFBE81D0BE8EA8A3AA05A2A5504001C74BA42A1571E8028E3DB7816D0",
INIT_35 => X"A5C7E3DFFFE90B45B47ABA497A82FFAFD2A82485FD2415A105C21451ED42A002",
INIT_36 => X"00000000000000000000B55EAAA100AA1D0F6F480B6A555A2A57A002A3D5FDB6",
INIT_37 => X"5EFAAAAB5E1AF3AABFF45592E88A0AFE80A8B0A0000000000000000000000000",
INIT_38 => X"65F520EBE9EF67D7BEA1FD5D556ABEF5D557FEBA55022A3F70C6B405F4D2AE97",
INIT_39 => X"C114728007521170821CE0FDE69411A8DED57CE1055555E5F58EFFC01FE2CACB",
INIT_3A => X"42341D5DEEBEF55080034E0A592A4AD0079C75D6070CC5CBB0280C029ABAA3EB",
INIT_3B => X"7F353AAF6C77F7F20D968BF57812A95E02A2AAB5EB0F280800EFAEE9F5D18F31",
INIT_3C => X"C91565455C141E41887D58AC448B69C30E02116220415A9540AA854140A0A204",
INIT_3D => X"DE6BE93172D7D625B556EEAB157ABEBE1B4D792A4AD1183454180DD3FDCAAAB7",
INIT_3E => X"F0000001FF0000001FF0000001FF0000001FF01EABC4B8014174FF7DA80F52FE",
INIT_3F => X"FF0000001FF0000001FF0000001FF0000001FF0000001FF0000001FF0000001F")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(0),               -- Port A write enable input
DIA(0)   => data_write_a(0),        -- Port A data input
DOA(0)   => data_read_a_hi_512(0),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(0),               -- Port B write enable input
DIB(0)   => data_write_b(0),        -- Port B data input
DOB(0)   => data_read_b_hi_512(0),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_1_11 : RAMB16_S1_S1
generic map (
INIT_00 => X"212C001411984004084D000508C53810A03D1450E839B003342114428A000803",
INIT_01 => X"00000019400B100A8196000000CC004400400002000000000000028001340000",
INIT_02 => X"052137AE8031800C0044009000000000061800001CD4019802AD04CCCFC20004",
INIT_03 => X"04514108C60C21008C6042108400000201440020505100000043C30E10E9F000",
INIT_04 => X"02104001011DEFE088805681920000008000004001900800004002108C280008",
INIT_05 => X"040002340105000200000000080001900010000108040000000008411600401C",
INIT_06 => X"1034001042800808201000000001000820020000102000040000000000800180",
INIT_07 => X"64BF81A15EDFDE8031800C00843060C19E030022103600000450020800040004",
INIT_08 => X"00008004691687AA840008000090248CC84E000046000311555521F183060AC5",
INIT_09 => X"0820800D08100171000DB000154440C800400500000852020011200201012021",
INIT_0A => X"02000040001000880A2A04445004000102002041000001008208001440004140",
INIT_0B => X"4820018A1140440078050040511000102000A008183000010002404400000000",
INIT_0C => X"1000C80008000C030030880C2A030A00C28030A80C2A030A00C28018D4061401",
INIT_0D => X"10040802050080200284401C0022880F009E08008205C0020118088018000000",
INIT_0E => X"0F03C00280000000420860C60C0C0B92C0000000004000010042000040102008",
INIT_0F => X"001E078005000108400005E11C0610000000288058000003C0F000A000100000",
INIT_10 => X"F10E0380000000C202300000008D187038000000480800000781E00140002000",
INIT_11 => X"806302380C870010000004400100110800007861E0180000000C400680000001",
INIT_12 => X"023E00000000018000580C308000050000610C30800005000215006800000101",
INIT_13 => X"61E0000000018100B0001843812000014100B00016030C20000141002880026D",
INIT_14 => X"400A20009B404F80000000018400A20044096111C04000000304026000501580",
INIT_15 => X"0046820040082300218450C2800010094000482141E060190700100000002200",
INIT_16 => X"020080200802008020080200802008020080008008600500A82A1100A8000000",
INIT_17 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_18 => X"0080200802008020080200802008020080200802008020080200802008020080",
INIT_19 => X"81328A46BABEFC54A0810C7452B4428A14000000000000000000020080200802",
INIT_1A => X"AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA28A28A28A28A2A8218D2C0C924925",
INIT_1B => X"E974BA5D2E974BA5D2E974BA5D2E974BA5D2E975BADD6EB75BADD6EB75BAAAAA",
INIT_1C => X"FFFFFFFFFFFFFFFD8C6318C6318C6318C6318C63000002E974BA5D2E974BA5D2",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"70E1C3870E1C387FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"5555500000000000000000000000000000000000000000000070E1C3870E1C38",
INIT_28 => X"EBDF455D2EAABEFF7FFE8BFF5D0002155557FFFFFF007FC21EFA2FFD74AAAAD5",
INIT_29 => X"AA95400552AAAABAFFD1574105D7FD75FFAAAA800AAF7AA974BAFFFBE8B45F7A",
INIT_2A => X"0517DF555D2EAAA1055000015500557DF45AAD1400BAA2AE801550051555EFF7",
INIT_2B => X"FFD540155557FD5400F78028BFFFFFBEAB55F780020AAAA80020AA082EAAB550",
INIT_2C => X"AFF842ABEF5D517DF55552A974AAF7AE820AA0851574BAA2D1574AA5D7BFDEBA",
INIT_2D => X"EFAAD1575EF557FFFE10557FFFFFFFFD56AAAAFFFFD7555AAD168B45AAAEAAAB",
INIT_2E => X"0005D7FFDF4500043FE105D2E954BAF7AE80010082A97410557FEABFFAAFBE8B",
INIT_2F => X"51C7A2FBD5490BFD1C056A000000000000000000000000000000000000000000",
INIT_30 => X"974BAF7FFEFB45FFAABDF55492AA8BC2EBDFEAF7F1F840017D4975D2FEF147FC",
INIT_31 => X"080BEF495FC71D54124924385FAAA8AAAE3D145410F7F1D55D71C002DABAEBAA",
INIT_32 => X"002D082082AB8B6DBEDB7DF7F540E2AE85028B40155145F7AF6DBED5450AA1C2",
INIT_33 => X"78E021FF1471FDEAAFFD56F16D5571D2E28E38E0216FA2D1E8E80140F45082B4",
INIT_34 => X"A2DA3FB7DAAD4AAAAF487BC70BFA97F7AF6D417E92482BF84020BA495557E3FF",
INIT_35 => X"55554ADBD7A2FFC7BEFF6FFD7FC7002FD74951D71EDFFABFD16FAAAE92BD5545",
INIT_36 => X"00000000000000000000547AB8F550A8010E00492487482FFFE82A85EBAE2FFC",
INIT_37 => X"1EF005162BEF047FD5545AAFBF7400FBF9424F70000000000000000000000000",
INIT_38 => X"714F8338AAAA1D0AE974AAF7FFFDF55F7AABFF55082CA8B4DF6C1E8F5E540002",
INIT_39 => X"EABEF75550ACBB7582225FF5843404547184164AA5D2EBEEB0A2D555410D3555",
INIT_3A => X"FEAAEB083BC1000FF8409000512AEABFFDF79DCBF755962010BDCBBC21455D7F",
INIT_3B => X"801F8BA0C57740BDAA0688E5405D57D412F7D55F5E50C7F401BAAE8403CF5A3F",
INIT_3C => X"5D16BABAA3EBC3157ABD5FFE55F2AA9FEAFDF7F431A9F7FFE81FF013A8001AFF",
INIT_3D => X"FB863550229BCABEB7DA403FFFDA2FBF7FED2C7F955445079E280A00C56145EF",
INIT_3E => X"0000000000000000000000000000000000000596EBEF55080034E0A592A4AD00",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(0),               -- Port A write enable input
DIA(0)   => data_write_a(1),        -- Port A data input
DOA(0)   => data_read_a_hi_512(1),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(0),               -- Port B write enable input
DIB(0)   => data_write_b(1),        -- Port B data input
DOB(0)   => data_read_b_hi_512(1),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_2_11 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10E006600180111284380310006289800480032283E000A34301002001A0817",
INIT_01 => X"0005A00810790848048044A54E404350404000720885800802000906E4910200",
INIT_02 => X"407004208400408044C600C50AA055254010541A110222841200000002402544",
INIT_03 => X"0600011004182401004102408C28414043101000408118000145840440F5C415",
INIT_04 => X"5035855703A2900A000CD3088400F40688C9844409060850925E58A4081A0221",
INIT_05 => X"0200840D1021A15AC50494894850890540D1E12020C6E510818500440A280090",
INIT_06 => X"113044094002801020440090A8011A1224AB9380552102442884882A20004097",
INIT_07 => X"000100880004428400408044860000008C022402102100AA40004404B5075460",
INIT_08 => X"15C23440408C862A2A12382A8A5244145048C06085008010141521F000001240",
INIT_09 => X"400582B9033AA0E7AA4110B0506744810554542450694E710A836188C2C00222",
INIT_0A => X"443518360012C2210B020414109130A28038188096A06B8C120CA440A9C00802",
INIT_0B => X"1345E53300EC68005605002964AF222A5704004D080211121C80024200821780",
INIT_0C => X"181080C1110C882202211488452213C88472213C88472213488441109A442231",
INIT_0D => X"008204440210091341208041000810C00000300220201800A908000038AD0284",
INIT_0E => X"00040002804180300E88D28D206A40000554815500481440300000C44A081100",
INIT_0F => X"000008000500828700000000010000000002380000A00000010000A010050000",
INIT_10 => X"00010000000004CA000214000000020000000000684280000002000140200500",
INIT_11 => X"000000000020000000000442100002840000000800000000010C000026000000",
INIT_12 => X"00000000000805A4800000000000152300000000000015801272000100210020",
INIT_13 => X"000000000101C00000C000000000000940000120000000000009600004050000",
INIT_14 => X"0000130000000000000002018000106000000000000000002380000141000000",
INIT_15 => X"55000190000000000002000280000000011080C0000000000000000000002310",
INIT_16 => X"40902409064190641906419024090244902A9003004800415120D4A190804241",
INIT_17 => X"0900409004090641906419064190240902409024090641906419064190240902",
INIT_18 => X"9044090040900409004190441904419044090040900409004190441904419044",
INIT_19 => X"75960040138D70C030B51C50C7D100A2052F81F81F83F03F03F0419044190441",
INIT_1A => X"0410410410410410410410410410410410410410410410410248602081659659",
INIT_1B => X"5128944A25128944A25128944A25128944A25128944A25128944A25128941041",
INIT_1C => X"FFFFFFFFFFFFFFFE1084210842108421084210843FFF825128944A25128944A2",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"7FD5FF555815607FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"2AA000000000000000000000000000000000000000000000007FD5FF55581560",
INIT_28 => X"FC21EFA2FFD75EFAA8415410AA8415555087BFFF55A2AA800BAFFAE954000800",
INIT_29 => X"84155EFA2AEBDEAAA2FBEAABA5D7FE8B555551421455D0002145552EBFEBA007",
INIT_2A => X"2AEBDF555D2E954BAA2AA974BAFFFFE8B45552EBDF45FFAEAABFFF7FFE8B55F7",
INIT_2B => X"AAAAAAAAAFFD1574105D7FFFF555D2AAAAAA5D2E820BAA2FBEAB5555557DF55A",
INIT_2C => X"50055575EFFF84021555D043DEAA5D04021EF557FC21FFAA8428BFFAAAA954AA",
INIT_2D => X"10085568A00FF80175FFA2D17DFEFF7800215500557DF55AA80001FFAA800015",
INIT_2E => X"0005D00020AAAA80020AA082EAAB5500517DF555D042AA10A284154005D00154",
INIT_2F => X"00AAFFAA9543A080038A2A000000000000000000000000000000000000000000",
INIT_30 => X"0017D5D20B8EAA007FC51C7A2FBD55D2BE800042AFE8E1557D0075D2F45BEAA8",
INIT_31 => X"AA8BC7EBDFEAFEFFD00105FFBC20BDEAAA2FBF8AAA557BE8B6D5D5FFABEF4904",
INIT_32 => X"FFEFB6D555578F7DB6A0BDF7D480E174BFA02A974BAF7F5EFB455D2ABDF55492",
INIT_33 => X"ED1FDE90E3A497492B6AAADAAAE3D155E105571D55D71C002DABA5524820BAB6",
INIT_34 => X"BE8F401D7B6A0001470155C51D0092A071555D5E3AE821D00001FF0871C016DB",
INIT_35 => X"5BE8555400550A38428007FED000E3DA3DFD5E3DFFFBD5A38A021551C5F7AF6D",
INIT_36 => X"00000000000000000000410F45082B4002D082082AB8B6D1C5B7DF7FF78E075C",
INIT_37 => X"5EF005560B55F7AA800AAF7AA954AA00042AAA20000000000000000000000000",
INIT_38 => X"ABEF057D68F5F5A00021EF55042AAAA007FD5555AAFBD7545FBB8020A3F7AE97",
INIT_39 => X"7DF55D7AABFF5428ACA8F45A6C1E8F5EFF84165EFF7802BAB0A2FFEAABA557BE",
INIT_3A => X"CA8AA80800020AAF7FBFFFEF04552ABFFFF841FFE75CA882108202E974AAF7D5",
INIT_3B => X"00151FF0C57401E5F3D1E00A1A884174A8FFAEBFEB0A2D55541051555694F002",
INIT_3C => X"2AA801455D7FE8BFFF680800FFF7AAA155F595542455512A975455D3AA8A0055",
INIT_3D => X"5D79FCAF774AE005BE7895554005D2A8A0B882FFFFE10AAAAAB755A66B6AF56A",
INIT_3E => X"00000000000000000000000000000000000000C3BC1000FF8409000512AEABFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(0),               -- Port A write enable input
DIA(0)   => data_write_a(2),        -- Port A data input
DOA(0)   => data_read_a_hi_512(2),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(0),               -- Port B write enable input
DIB(0)   => data_write_b(2),        -- Port B data input
DOB(0)   => data_read_b_hi_512(2),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_3_11 : RAMB16_S1_S1
generic map (
INIT_00 => X"210C00A20020000108430020001600B8156021104940741B3530400E02B92203",
INIT_01 => X"014C9BCA58B1296D24A402C992500B69404040028804A0080A000416A8D90A08",
INIT_02 => X"C12026A484318004404405C9C66E331352180D468B8203980300204442E02B34",
INIT_03 => X"04000748D60D24648D60524C88804D0215011020D15018148040C10A70E1D58C",
INIT_04 => X"18283333240FE41244187308C9104D70944852640901083801750EB0A418C220",
INIT_05 => X"0613142D01912CC2A1B4140528348900C612A104201C689044340ED413A07649",
INIT_06 => X"119000034019881822104C5E68035250A222829710A0A02C18C01A9920842413",
INIT_07 => X"402F00AB0016CA0431800444841020509D038B021230C1990001C644C8273200",
INIT_08 => X"16905000408482088290E8E64010248C4A5AA840C2000110001521F0810A92E7",
INIT_09 => X"0003CE6581BD016342A951AB146C4480530C3B2A8088D3542651670200C1826A",
INIT_0A => X"00735D36209A8A20020894004284B660821030C8990467401218004041020002",
INIT_0B => X"512445B740457154562F957CC08B00093700080D0A4851001D8302D20A0A1530",
INIT_0C => X"00508650008008021021A40861021840869021A408610218C0869810D6043095",
INIT_0D => X"1C8508438450801043A08090380A8834207007022209038080190000999C8F84",
INIT_0E => X"000400200000C0002A48A206204C4205F3304B33004C0041006240140A1C310A",
INIT_0F => X"0000080040000083800400000100000000008400018040000100080000510100",
INIT_10 => X"0001000000000800000244040000020000000100002A0080000200100000A702",
INIT_11 => X"000000000020000000200000080002C000800008000000000022000006808000",
INIT_12 => X"0000000000000A2281000000000040A3810000000000402001400000022002A0",
INIT_13 => X"000000000004200001C0400000000010200001C0400000000010000004490010",
INIT_14 => X"0001070004000000000000060000104C08000000000000001000000903008000",
INIT_15 => X"CC004050CA0C00020220200070040000010401C4000000000000000000100008",
INIT_16 => X"4310E4310A4210A4210A4210A4210A4210A8D0830A68010001B4DA881048061C",
INIT_17 => X"21084290A4210A4210A4210A4210A4210A4210A4210E4310E4310E4310E4310E",
INIT_18 => X"90A421084290A421084390E4310C4390E4310C4390E4310C4290A421084290A4",
INIT_19 => X"015303C0C78C706428A14C586291000A044001FFE000003FFC004290A4210842",
INIT_1A => X"2492492492492492492492492492492492410410410410412821600001249249",
INIT_1B => X"51A8D46A351A8D46A351A8D46A351A8D46A351A9D4EA753A9D4EA753A9D49249",
INIT_1C => X"FFFFFFFFFFFFFFFC00000000000000000000000038F56351A8D46A351A8D46A3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"55AB02055AB0207FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"420000000000000000000000000000000000000000000000007FFFAB57FFFAB5",
INIT_28 => X"A800BAFFAE9554508002AA00AA843DF55FFAA955EFA2D168B55557BEAA000055",
INIT_29 => X"002AB55AAAA955EF005568A00087BE8BFFA2D155410AA8415555087BFFF55A2A",
INIT_2A => X"AAABFF5508003FF555D0002145552ABFEBA007FC21EF007FD75FFAA841541008",
INIT_2B => X"082EBDEAAA2FBEAABA5D7FC0155005168B455D042AB45F7FFD741000042AA10A",
INIT_2C => X"FF7FBEAB55F7AABDEBA5D7FC2010A2D1575FFF7AA975555D2E80145F78415545",
INIT_2D => X"EF5555554AA087BC01FFFFAAAAB55552A954BAFFFFE8B55552EBDE00F7AEAABF",
INIT_2E => X"000082E820BAA2FBEAB5555557DF55A2AEBDF555D2E954BA002EAAABA002A821",
INIT_2F => X"FB7D5D7FEAA3808554203A000000000000000000000000000000000000000000",
INIT_30 => X"1557D1475FAF45BEAA800AAFFAA95578080038A2AA28E3AF55E3A0BA5D7AADB6",
INIT_31 => X"BD55D7BE80004AA1E8E2AB55B6A0925D7085F6AA10087FEABD7AAD57AEBAB68E",
INIT_32 => X"F5D0438140E2FA38B6AEBFF6D1D04AAFFA41040017D5D20B8EAA007FC51C7A2F",
INIT_33 => X"D0A901FFFF801557D1C20B8EAAA2FBE80AA557BE8B6D5D5FFABEF49002FB55FF",
INIT_34 => X"5D20BDE00EBAAA8BC7EBDFEAFEFAB8ABAE925D21C7010EADB525D7FFAE975C75",
INIT_35 => X"F002EADA921420871D74971D24820875C21D5EB8AA8FFF012A954BAFFF5EFB45",
INIT_36 => X"000000000000000000001C24820BAB6FFEFB6D555578F7DB6A0BDF7DEB8E125F",
INIT_37 => X"B55A28408145AAFFFFFFF5D7FEAABA0051400A20000000000000000000000000",
INIT_38 => X"AB55FAD568AA2AFAE975EF555168B55F7AA800BAF7AA955EF00042AAA2A2AEAA",
INIT_39 => X"2AAAA007FD55558A7BD7145FBB8020A35D2ABEF55F7800015F087FEAA00007FE",
INIT_3A => X"968F575D003FF55F7D5420BA5D2ABFEAAF7AE9DFF759A82AEF70800021EF5504",
INIT_3B => X"FFD5145FBAC9755F05040255FFD84175EF55002AAB0A2FFEAABA557BEA3EF057",
INIT_3C => X"82E974AAF7D57DF45552A3FF10AA8429F45A7D5EAF5FFBAEAAA10554155400AA",
INIT_3D => X"FF843FFE77C80825BC052ABFE10550415557085540000005156155FE90A8F5C0",
INIT_3E => X"00000000000000000000000000000000000005500020AAF7FBFFFEF04552ABFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(0),               -- Port A write enable input
DIA(0)   => data_write_a(3),        -- Port A data input
DOA(0)   => data_read_a_hi_512(3),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(0),               -- Port B write enable input
DIB(0)   => data_write_b(3),        -- Port B data input
DOB(0)   => data_read_b_hi_512(3),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_4_11 : RAMB16_S1_S1
generic map (
INIT_00 => X"A108400020612C80284210081034849800A00030300004833522C82D04A16002",
INIT_01 => X"2043998A1839284D1CA0650E1E504368403008418984014902030806A0D10200",
INIT_02 => X"C120042200000000044441CE01E80F00A49043118680008002000000026208E4",
INIT_03 => X"040001020019200020011209CC0164C060000000690111040144800042F5C403",
INIT_04 => X"7029AF0F81A00010CCA47700CC513CAC0D0B8E02010740E19754080108988021",
INIT_05 => X"02139405007133C0712244CD20F20105D583000020E9892201D304D42A9835E1",
INIT_06 => X"9190440300078002014405D9EE814C0284A883B6D7038AE079059B7800048092",
INIT_07 => X"000100AA0004408000000004840400008D200102503000782000C00C8025C000",
INIT_08 => X"00728A00408403220811991E02120C044058080004000001101121F220000260",
INIT_09 => X"811001E1185B38AD23C3707AD46440818F3CF80EC423CA7D01D123C80200816A",
INIT_0A => X"45810810A01B40216361056D6150F41200280001900439001FD8A00041400000",
INIT_0B => X"11FC88076266E800D605402962A820211500024808010512C40106D222223B14",
INIT_0C => X"0408804116040B02C02C500B0C02C100B0C02C100B0402C300B0401618058611",
INIT_0D => X"040200050200501301208482200D00D0A0408402C4282200A84800009B878680",
INIT_0E => X"00000020000100024AC88300300060090F0D830F00025400300204D018000804",
INIT_0F => X"8000000040000206A2000800000000000000950002E010000000080000588040",
INIT_10 => X"0000000000000808000554000200000000000100006D0020000000100000BB00",
INIT_11 => X"0000400000000000002000001A0002504001000000000000002280000D800800",
INIT_12 => X"0800000000000E2C802000000000408D801000000000408012440000200110A0",
INIT_13 => X"000000000004680003A0040000000010280003800800000000102800000B0000",
INIT_14 => X"000005C0002000000000000620000158000010000000000010A0000B00000200",
INIT_15 => X"C30146200400104002602600400000000294004000000004000000000010001A",
INIT_16 => X"0080200000008020000000802000000080080000004090014134DA101288C6DB",
INIT_17 => X"0802000000000401806010040180601004018060100000802000000080200000",
INIT_18 => X"8060180601004010040080200802000000000000802008020000000000008020",
INIT_19 => X"C0A28A063807E0500014063450404882846FFE000003FFC00000010040100401",
INIT_1A => X"AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA28A28A28A28A2934C8D0CCD145144",
INIT_1B => X"68341A0D068341A0D068341A0D068341A0D068351A8D46A351A8D46A351AAAAA",
INIT_1C => X"FFFFFFFFFFFFFFFC0000000000000000000000001FE32068341A0D068341A0D0",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"408102040810207FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"800AA00000000000000000000000000000000000000000000040810204081020",
INIT_28 => X"168B55557BEAB4500554200000557FE10FFFBEAA10007FD7410FFAA97555082A",
INIT_29 => X"55574105D2A800AA00043FEBA5D7FEAA00007BE8AAAAA843DF55FFAA955EFA2D",
INIT_2A => X"57BC00AAA2FFEAAAAAA8415555087BFFF55A2AA800BAFFAE9555508002AA0000",
INIT_2B => X"A2AA955EF005568A00087BE8BFFA2D17DE1000517FE10AAAAA8AAA002E975455",
INIT_2C => X"FAA8417410A2D140000F7FBC2010A2D157400AAAE974AAAAAA974BA08002AB55",
INIT_2D => X"EFA2AABDEAA087BEAAAAA2FBD54BA080002145552ABFEAA007FC21EF007FD75F",
INIT_2E => X"00055042AB45F7FFD741000042AA10AAAABFF5508003FF55F7D568A00552EA8B",
INIT_2F => X"5400F7A49057D0824850B8000000000000000000000000000000000000000000",
INIT_30 => X"3AF55F7A0925D7AADB6FB7D5D7FEAB7808554203A145178E00FFFBE8A101475D",
INIT_31 => X"A9557D080038AAA145157428492E8008200043FE925571EFA380871C7028A28E",
INIT_32 => X"AEA8A9200249056D4175C5092AAF5FDA38BE8E1557D1475FAF45BEAA800AAFFA",
INIT_33 => X"AA4954281C0E2FB55B6A0925D7085F6AA10087FEABD7AAD57AEBA08517DE00AA",
INIT_34 => X"007FC51C7007BD55D7BE80004AAFEDB42028EBFBC2028BED152438AAA092492A",
INIT_35 => X"AF7DF6AA00412EAABFFAA803DEBA0875EDA80BEF1C743840040017D5520B8EAA",
INIT_36 => X"0000000000000000000041002FB55FFF5D0438140E2FA38B6AEBFF6DBE84AAEB",
INIT_37 => X"A00FFFFEAA105D5155410FF84021EF0800154B20000000000000000000000000",
INIT_38 => X"DEBA0851574B2AAAEAAB55F78400145AAFFFFFEF5D7FEABFF0051400A25D5568",
INIT_39 => X"68B55F7AA800BAF7AA955EF00042AAA25555410BA082E8201000043FE005D517",
INIT_3A => X"568AA200557DE00AAAAAAA000804001FF005575408AA557FEB2FFAE975EF5551",
INIT_3B => X"D1550AAAA8002010F2AC154B25F2ABFF55F7800015F087FEAA00007FEAB55FAD",
INIT_3C => X"800021EF55042AAAA007FD5555087BD6145FAAC000A2A6FBC00BAAAFBC00BAF7",
INIT_3D => X"F7AEBDFF779A82AA43F7FBE8A00082EA8BFFAA843FEBA08517DE00F3F9574B30",
INIT_3E => X"000000000000000000000000000000000000008003FF55F7D5420BA5D2ABFEAA",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(0),               -- Port A write enable input
DIA(0)   => data_write_a(4),        -- Port A data input
DOA(0)   => data_read_a_hi_512(4),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(0),               -- Port B write enable input
DIB(0)   => data_write_b(4),        -- Port B data input
DOB(0)   => data_read_b_hi_512(4),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_5_11 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50DF4A0791B3FCB694379283C81FD996A091832102004A336A20E03C040C002",
INIT_01 => X"805FBDC69830A84D5C6A60000C34C26841280A00084000C8C212892EEAD53235",
INIT_02 => X"3B2026B578918E640A4F01CF8011FF0002080000082CA9998276DF7772C7C80D",
INIT_03 => X"37134108420D700084205702A4008A1D9100002171C0E0051554D93A11F5D140",
INIT_04 => X"8A41A0FC03A56DA000425A819410E3816C086198A388B702A8CA1210844A0C4C",
INIT_05 => X"B1808A062E8BC835F5E84532D708238A282F00A9291224800A2861490343082C",
INIT_06 => X"903FB8483A90581859050424100940825C6184401CDC451B860A6507160C4100",
INIT_07 => X"D26F068BCC96CDF8918E640E96D1A3469D6300E2FFEA27F8E4D23248130E259C",
INIT_08 => X"0BFA82E568442B2A082C0A7E3014250D49DA37A2420619000002AFF48D1222E5",
INIT_09 => X"3F005001E40969289429360416DCD1C46083030604B1CA20C03DF83B0A2C60A5",
INIT_0A => X"14613C71005A10492B888120288F480D58858449026145B3830F449449062B4F",
INIT_0B => X"11AC04934AC648BFD727C031E64170A137D5AA5C3E4B0F8A3C58C34C002290E3",
INIT_0C => X"CA29C6CC50384B6AC6AC86AB31AACA6AB39AAC86AB39AACA6AB3055643559C31",
INIT_0D => X"C673E33CF28F38603855401985228A0614BD30A0A2819852011E5AC2B87F9182",
INIT_0E => X"FF87C002F87A803E460B2516510CA594FF0044FFA4B08BAC4BB2CD0F09CF84E3",
INIT_0F => X"0DFF0F8005F0F5100DFFF5E15D06101C55EB29F1E00BE53FE1F000BE1E802F94",
INIT_10 => X"F12F0380231F17D78FC029FFF58D9A70380230F2FE0017C37FC3E0017C3D005F",
INIT_11 => X"FC7F023C0CA700125C0F8F7E43F1F001BFFE7C69E01804E1E7CCF8FC003FF5F1",
INIT_12 => X"023E00017C1FC1A4BFD82C3081C5BD27BFE30C3081C5BD00C02365D645CEEF5B",
INIT_13 => X"61E0042787F181E9C1EFD8CB8120C5AF41E9C18FD60F0C20666F41E9F009FFFD",
INIT_14 => X"7A7C077FFF404F80005F07F187A7D14BFFC96111C048278DEB074F9930FF9D80",
INIT_15 => X"C064014B8B652E2B3120C81284641D3E8DBF7D636FE860190700132C1F0EFB80",
INIT_16 => X"38CE1384E3384E338CE138CE1384E33C4E3ECE32E128882551349A1CBAA44103",
INIT_17 => X"84E3384E3384E3384E338CE138CE1384E3384E338CE138CE1384E3384E338CE1",
INIT_18 => X"CE138CE138CE138CE1384E3384E3384E3384E338CE138CE138CE138CE1384E33",
INIT_19 => X"F5E5BB4E7F7B9DB7FF3A1B6DB7E8410A8C000000000000000000384E3384E338",
INIT_1A => X"BEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEF9F7CFDFDDCF3CF3D",
INIT_1B => X"BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEFBEF",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000001711C7BBDDEEF77BBDDEEF77",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"FDFFF00000000000000000000000000000000000000000000080000000000000",
INIT_28 => X"FD7410FFAA97410082A800AAAAAE955450055421FFFFFBC0010AAD5574BA557F",
INIT_29 => X"7FD74000055574BA5D7FD7555A2D5575EF55517FF5500557FE10FFFBEAA10007",
INIT_2A => X"0002AABA5D2ABFFFFAA843DF55FFAA955EFA2D168B55557BEAB5500554200000",
INIT_2B => X"5D2A800AA00043FEBA5D7FEAA00007BC00AAAAAEBDF45A28428B45FFD168BFF0",
INIT_2C => X"5080028A00A2FFFDE00F7D57FEBAFF80174BAAAD1555EF555555555005557410",
INIT_2D => X"BA5D2E821FFA2D5554BA557BD75FFAA8415555087BFFF55A2AA800BAFFAE9555",
INIT_2E => X"00000517FE10AAAAA8AAA002E97545557BC00AAA2FFEAAAA082A97545F7D5420",
INIT_2F => X"7010BEDF524AA5571FDFEF000000000000000000000000000000000000000000",
INIT_30 => X"78E00EBFBE8A101475D5400F7A49043D0824850B8A2AE9756D145B401FFFFFFC",
INIT_31 => X"FEAB7D0855420BA1471D74380851524BA5571D757DB6D5525EF555178F6D1451",
INIT_32 => X"8A28B6DEBDF6DBEF1C0A28AAA5524BFFFFA28E3AF55F7A0925D7AADB6FB7D5D7",
INIT_33 => X"5555057D145152428492E8008200043FE925571EFA380871C7028B6AEBDF45B6",
INIT_34 => X"BEAA800AAFFAA9557D080038AAAA2FBF8E10EBD578EAAFF8415482BED1555EF5",
INIT_35 => X"81C209256DFFDF420BA552A821FFB6DF574A85575C55EFBE8E1557D1475FAF45",
INIT_36 => X"0000000000000000000008517DE00AAAEA8A9200249056D4175C50920875FDA3",
INIT_37 => X"5FF5D7BC21EFF7FBD7400F7FBC00BA55557DFF70000000000000000000000000",
INIT_38 => X"01FF5D5568BE7555568A00AAFFEAA105D5155410FF84020AA0800154B2AAAA97",
INIT_39 => X"00145AAFFFFFEF5D7FEABFF0051400A25551554BA0051400BA5551575EFF7D14",
INIT_3A => X"1574B2FFAABFF45FFAAAABFFAAFFFDFFF552EA8AAA55043DFF7AAAEAAB55F784",
INIT_3B => X"8002410FFD5575EF5555421E75555400BA082E8201000043FE005D517DEBA085",
INIT_3C => X"FAE975EF555168B55F7AA800BAF7AA955EF00002AAA2A2FBE8A00A2D16AAAAFF",
INIT_3D => X"0055554088A557FEB25D00021FFFFFFC00BA552A821EFFFFFD74BA5D51575F7F",
INIT_3E => X"000000000000000000000000000000000000000557DE00AAAAAAA000804001FF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(0),               -- Port A write enable input
DIA(0)   => data_write_a(5),        -- Port A data input
DOA(0)   => data_read_a_hi_512(5),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(0),               -- Port B write enable input
DIB(0)   => data_write_b(5),        -- Port B data input
DOB(0)   => data_read_b_hi_512(5),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_6_11 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10800B0061A01002840002C03002818000402322520070B313301C4389B2082",
INIT_01 => X"250041CA3839684D18A160000C52426841000000090800090210080008110200",
INIT_02 => X"0020042080010000044654C0000C008010000000001020900200200002620814",
INIT_03 => X"060881021088200021080200E4000A0891000020610111500104C00000F14400",
INIT_04 => X"0880000100000002000052288144004281C050400100280000C8100000080001",
INIT_05 => X"928080840001100A08009000280201000850E022401400002028214043410820",
INIT_06 => X"10100518090012122100C808049310002040000410A0001400000200120840D2",
INIT_07 => X"000100800004400001000000860408108C22000A502010074120044800040001",
INIT_08 => X"50000040D0C4E2088003FD01C01004044058082004000000000121F020408244",
INIT_09 => X"00BF17E9001205A5204911F814444080400100020000D200DFD16400C2A40AA0",
INIT_0A => X"04611C17849000022862A1596C8B5DF04834948900000100220C244840000880",
INIT_0B => X"03AD0413424E4044D665C070C22602291504400D084915020448114080201000",
INIT_0C => X"5E08864011088B22D22C008B0022C408B1022C208B0822C608B1111600458010",
INIT_0D => X"4251A12CD28A300429688001000800000020280204001000A00804309A002182",
INIT_0E => X"0000000280402400420800000000006200FC10002442042429324294014E8CA7",
INIT_0F => X"A40000000500800840000800000000000002280018001480000000A010100052",
INIT_10 => X"00000000000004C2003000010240000000000000680800290000000140202000",
INIT_11 => X"2000C0000000000000000442000001080001000000000000010C000280001804",
INIT_12 => X"08000000000801C300A010000000156000902000000015101200002800000000",
INIT_13 => X"000000000101800038002408000000094000386028040000000940000ED40000",
INIT_14 => X"0003B000002000000000020180002A24005010000000000023000060C7000A40",
INIT_15 => X"3F0280090321000040A410C28108000160008094000810040000000000002300",
INIT_16 => X"284A5284A728CA5284A528CA728CA52C4A5A0A32A300940101349A0408240818",
INIT_17 => X"9CA1294A329CA5284A728CA7284A5284A728CA5284A528CA728CA5284A728CA7",
INIT_18 => X"CA3294A129CA3294A129CA1294A329CA1294A3294A129CA3294A129CA3294A32",
INIT_19 => X"F5F78BCE7F8FF0F4FA955F7CF7F40A80145D55555556AAAAAAAAA94A329CA129",
INIT_1A => X"8E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E39B6CEDECDDF7DF7D",
INIT_1B => X"F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE38E3",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000001A1A33F9FCFE7F3F9FCFE7F3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"555FF00000000000000000000000000000000000000000000080000000000000",
INIT_28 => X"BC0010AAD5574BA557FFDFFF087BFDF45F7AA974AAAAAA97555F784174BAF7D5",
INIT_29 => X"515555508043FE00F7AA97555A2FBD7410AA8428AAAAAAE955450055421FFFFF",
INIT_2A => X"7D1575EFFFAA9555500557FE10FFFBEAA10007FD7410FFAA97400082A800AA08",
INIT_2B => X"0055574BA5D7FD7555A2D5575EF55517FF55A2AA97400552AAAB45082E80155F",
INIT_2C => X"500554200000003DE10FFD5401FFF7AAA8A10082EAAB45A2FFC2000007FD7400",
INIT_2D => X"10AA803FE105D516AABAFF843FFFFAA843DF55FFAA955EFA2D168B55557BEAB5",
INIT_2E => X"000AAAEBDF45A28428B45FFD168BFF00002AABA5D2ABFFFF087BD5545007BFDE",
INIT_2F => X"256DEB84104BAFFD1525FF000000000000000000000000000000000000000000",
INIT_30 => X"9756D145B401FFFFFFC7010BEDF524AA5571FDFEF1C7BFFF55FFA095482B6A49",
INIT_31 => X"4904380824850381C5B5057D1C003DE28F7A49057DAAF5D2428A2842AAAAA2AE",
INIT_32 => X"2AAFB451C2A8017DE3DF525FFFFA49756D145178E00EBFBE8A101475D5400F7A",
INIT_33 => X"2F1C50381471D74380851524BA5571D757DB6D5525EF555178F6DAAA49542841",
INIT_34 => X"AADB6FB7D5D7FEAB7D0855420BA1C0E3FE00E3DB471EFE3AAAAA00082EA8B6DA",
INIT_35 => X"F1C7BD057D1C71FFE10A28038E1049516AAB8FF8428FEFA28E3AF55F7A0925D7",
INIT_36 => X"00000000000000000000B6AEBDF45B68A28B6DEBDF6DBEF1C0A28AAA5524BFFF",
INIT_37 => X"F55F78017400F780001FFAA84000AAFFD1401E70000000000000000000000000",
INIT_38 => X"20BAAA8428AA2AAAA975FF5D7BC21EFF7FBD7400F7FBC00BA55557DFF7557BFD",
INIT_39 => X"EAA105D5155410FF84020AA0800154B2557FC01EF55043FEAAFF80021EFA2D14",
INIT_3A => X"568BE7AA80174AA082ABDF555D2A821EFAAFBC01FFF780155F7555568A00AAFF",
INIT_3B => X"AEA8A10082EA8BEFAAD5554B25551554BA0051400BA5551575EFF7D1401FF5D5",
INIT_3C => X"AAEAAB55F78400145AAFFFFFEF5D7FEABFF0051400A25D2EBFE10AAFFD55EFA2",
INIT_3D => X"552EA8AAA55043DFF7557BC01EF55557DE00AA842AA0000516AABAFF8428BE7A",
INIT_3E => X"0000000000000000000000000000000000000FFAABFF45FFAAAABFFAAFFFDFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(0),               -- Port A write enable input
DIA(0)   => data_write_a(6),        -- Port A data input
DOA(0)   => data_read_a_hi_512(6),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(0),               -- Port B write enable input
DIB(0)   => data_write_b(6),        -- Port B data input
DOB(0)   => data_read_b_hi_512(6),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_7_11 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10844B00482258A2842112C02450418800002300500030B313300C418992002",
INIT_01 => X"000009CA3839684D1CA0E0000E51424840000000080000080200080008510204",
INIT_02 => X"0120042086010000044600C00008000004100000000260900200000002402004",
INIT_03 => X"8628A10000082400000002408400080011000000610008000208C00000E14400",
INIT_04 => X"0911800100A000000000524084000040000050001140200100C8100000080102",
INIT_05 => X"0300812401011000000000002000114008008060441000000020024093000000",
INIT_06 => X"9190431C0D4010100000880804010010800000041080081000000200010424B2",
INIT_07 => X"000100AA0004408601000004860000008C02000A103010006928040800062481",
INIT_08 => X"84000048D484C20888000A0002120484C048007004000000000021F000000244",
INIT_09 => X"00A06009881201A520491004106C48A04040002400A15A208001650004001020",
INIT_0A => X"C99E1060201002044809C1040140A001004808810000459033189C0A400118A0",
INIT_0B => X"102000024040484050050041648A0041140C500B08821054C000264120000400",
INIT_0C => X"0404A083260E0832132011880462011880462051881462051881D31018C40620",
INIT_0D => X"0001000080001000813094801A8F80F00A600B52602801A88848011118003700",
INIT_0E => X"000003C007C002808228010410082042C000C000000004001002000400040002",
INIT_0F => X"A4000007800F80C840000800009864038A1200081C0014800000F001F0200052",
INIT_10 => X"00002C0E00E0E4004038000102400002C0E00E0D20100029000001E003E04000",
INIT_11 => X"2000C04031100E0403D0700300080908000100000661801E1900040380001804",
INIT_12 => X"0840878083E8003780A01043203A101780902043203A10082410082880000000",
INIT_13 => X"0601E0187900181035E0240806483248181035E0280410C8198818100DDD0000",
INIT_14 => X"0403774000201021E020FA006040376C00501022131210722060806D47000A40",
INIT_15 => X"00928A0002000110888600C032128201519480D40009902430160403E0E00506",
INIT_16 => X"01000000020080601802000000000405000A0020020081014134928820480010",
INIT_17 => X"0802018040000000006018020080200804010000000000806018020080000004",
INIT_18 => X"0000000001806008020000001006008020080001004008020080201004000020",
INIT_19 => X"0000000000000000000000000000400A004618618618C30C30C3000020180600",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000000B0840000000000000000000",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"1555500000000000000000000000000000000000000000000080000000000000",
INIT_28 => X"A97555F784174BAF7D5555FFF780155EFAAAEA8ABAAAFBFDE0055556AA005D04",
INIT_29 => X"55555EFAAFFFDFEFAAAAAAB455D556AA00FFAE95555087BFDF45F7AA974AAAAA",
INIT_2A => X"02EAAAAA082EA8A00AAAE955450055421FFFFFBC0010AAD5574BA557FFDFFF55",
INIT_2B => X"08043FE00F7AA97555A2FBD7410AA8428AAA557BFDFFF55003DFFFF7FBEAA000",
INIT_2C => X"0082A800AAF7AE975FFA28000010552EBDE00007BEAAAAA2D140000085155555",
INIT_2D => X"45087FEAB455D516AB55557BD55FF00557FE10FFFBEAA10007FD7410FFAA9740",
INIT_2E => X"000A2AA97400552AAAB45082E80155F7D1575EFFFAA955555D51574AAAAFFD55",
INIT_2F => X"AE105D556AA10410E17555000000000000000000000000000000000000000000",
INIT_30 => X"FFF55FFA095482B6A49256DEB84104BAFFD1525FFFF8E175C7A2AAAAA82A2F1F",
INIT_31 => X"F524AA5571FDFEF415B575D7AAF1FFFD7AAAAAFB7D495F6AA10E3AE905551C7B",
INIT_32 => X"003AFEFEBFBEAA001C2EA8A821C2EAAA00A2AE9756D145B401FFFFFFC7010BED",
INIT_33 => X"EDB470101C5B5057D1C003DE28F7A49057DAAF5D2428A2842AAAA497BFAFFF49",
INIT_34 => X"1475D5400F7A490438082485038F7A4905C7A28A070384120BDE100075EAA82B",
INIT_35 => X"D495150492BEF1D2555087BE8B7D555F6AB57417BC05D7145178E00EBFBE8A10",
INIT_36 => X"00000000000000000000AAA495428412AAFB451C2A8017DE3DF525FFFFA49756",
INIT_37 => X"555A2AEA8A10AAD568A00555168A10002E9754D0000000000000000000000000",
INIT_38 => X"8A10AAAE8215D557BFDF55F78017400F780001FFAA84000AAFFD1401E7FFAA97",
INIT_39 => X"C21EFF7FBD7400F7FBC00BA55557DFF7007BD5555AAD57DF55AAAEBDFEF007BE",
INIT_3A => X"428AA2007FE8BFF080028BFFAAFFEAA105D2EAAA005D2AAAA18AAAA975FF5D7B",
INIT_3B => X"043DE0000516AA10F7FBD7408557FC01EF55043FEAAFF80021EFA2D1420BAAA8",
INIT_3C => X"55568A00AAFFEAA105D5155410FF84020AA0800154B2FF8402145A2AA954AA00",
INIT_3D => X"AAFBC01FFF780155F7005140000FFD140145007FE8BEF557BEAB55087FC215D5",
INIT_3E => X"0000000000000000000000000000000000000AA80174AA082ABDF555D2A821EF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(0),               -- Port A write enable input
DIA(0)   => data_write_a(7),        -- Port A data input
DOA(0)   => data_read_a_hi_512(7),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(0),               -- Port B write enable input
DIB(0)   => data_write_b(7),        -- Port B data input
DOB(0)   => data_read_b_hi_512(7),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_8_11 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00000648E2840112C00000418000002700500030B3132000400812082",
INIT_01 => X"100008480009004C04A100000252024840000000180800080200010040110204",
INIT_02 => X"0020042000490000004600804008000005100000000024900200000002400004",
INIT_03 => X"0A0C33400008082400000080A4004B0891000020610112000040C00000E5C000",
INIT_04 => X"18800001000000000000512080000040800150400824280110C8100000120200",
INIT_05 => X"908084A10100100200004080280008240810802206940000012C214451610800",
INIT_06 => X"81B000080860109021400008040000202048020414A0021400040200322824C1",
INIT_07 => X"000000080004408049000004860000008402001A50208000630C040800062483",
INIT_08 => X"440000428644212280800A00021004044048002124000000000021F000000244",
INIT_09 => X"00004009001001010008100414644410400102228000D20080114502006409A2",
INIT_0A => X"000051312000042200294429148A4801C80C8C81000045907118040340020832",
INIT_0B => X"4020000240404140004D0544C4AA0001150410090302500011C813428A000400",
INIT_0C => X"46501090008820240240409000240009000240009000240009000120204808A5",
INIT_0D => X"42D1A168D09A301468402480004780F00140080860280004085904309A002196",
INIT_0E => X"00783FC00044340242280000000000020000C0000442106419120004034685A3",
INIT_0F => X"8000F07F800088A80000081EA2F9EC0000064004081010001E0FF00011104040",
INIT_10 => X"0ED0FC7E00000422201080000202658FC7E0000021882020003C1FE000222080",
INIT_11 => X"018059C3F350FE0C00000002A0040500000103961FE780000110010090000800",
INIT_12 => X"FD41FF80000830200021C1CF600012200010D1CF600012121600100810000004",
INIT_13 => X"9E1FE000010A1802100004343ED8000898021000087073D80008980200800002",
INIT_14 => X"0080200000BEB07FE00002086008020000209AEE3F300000246020200000620B",
INIT_15 => X"0088881903210000440610C8000A808040000208901786E4F0FE0C0000000166",
INIT_16 => X"685A1685A769DA368DA368DA769DA36CDA121A11A141800011309284002C0810",
INIT_17 => X"95A5685A1685A5695A368DA368DA769DA368DA368DA7695A1685A1685A5695A1",
INIT_18 => X"5A1695A568DA368DA369DA768DA1685A1695A5685A168DA369DA768DA368DA16",
INIT_19 => X"A4028A0A543EBC57A10A1E75D64108080468618618630C30C30C69DA5685A168",
INIT_1A => X"9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7BF3CCD8DF5B2DB2C",
INIT_1B => X"F87D3E1F4F87D3E1F4F87D3E1F4F87D3E1F4F87C3E1F0F87C3E1F0F87C3E79E7",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000006A6D4F87D3E1F4F87D3E1F4",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"155FF00000000000000000000000000000000000000000000080000000000000",
INIT_28 => X"BFDE0055556AA005D0415555080000000087BEAA10F7803DE00FFAEBFFFF0800",
INIT_29 => X"2AA8AAA557FC0010F780154105D7FC2145005155555F780155EFAAAEA8ABAAAF",
INIT_2A => X"7FFFFF55AA80155FF087BFDF45F7AA974AAAAAA97555F784174BAF7D5555FF55",
INIT_2B => X"AAFFFDFEFAAAAAAB455D556AA00FFAE95555AAFFE8A00552EBFE00F7D17FF45F",
INIT_2C => X"A557FFDFFF5504000AAAAAAA8B55F7D140010552E821EFAAAABDF555555555EF",
INIT_2D => X"55AA8028A00A2D57FF45557BE8A00AAAE955450055421FFFFFBC0010AAD5574B",
INIT_2E => X"000557BFDFFF55003DFFFF7FBEAA00002EAAAAA082EA8A00002AA8A10F784021",
INIT_2F => X"FE10F7AEBAFFF080A175D7000000000000000000000000000000000000000000",
INIT_30 => X"175C7A2AAAAA82A2F1FAE105D556AA10410E17555080E000280071E8A00EB8E3",
INIT_31 => X"4104BAFFD1525FF492EA8AAA5571C2000FF8A17400557FC015514555757DFF8E",
INIT_32 => X"2ABDE10EBDF7AF6DE3FFF8F7DB68A105D71C7BFFF55FFA095482B6A49256DEB8",
INIT_33 => X"AA0BDF6D415B575D7AAF1FFFD7AAAAAFB7D495F6AA10E3AE90555A2FBE8A3849",
INIT_34 => X"FFFFC7010BEDF524AA5571FDFEF550E00082B6A0AFB55F7D1420104124821D7A",
INIT_35 => X"01C2EA8A00F7800017DA2842FA00B6D578F6D557FFDA00A2AE9756D145B401FF",
INIT_36 => X"00000000000000000000497BFAFFF49003AFEFEBFBEAA001C2EA8A821C2EAAA0",
INIT_37 => X"0BA08556AA00AAAABFE00F7AEAABEF082E955450000000000000000000000000",
INIT_38 => X"21555D51575EFFFAA97555A2AEA8A10AAD568A00555168A10002E9754D082E82",
INIT_39 => X"17400F780001FFAA84000AAFFD1401E7082EAAABA5D5140010F7AE974105D7BC",
INIT_3A => X"E8215DA2FFE8ABA082ABFE00AAFBEABFFAAFBEABFFF7AA80145557BFDF55F780",
INIT_3B => X"D540000000402145AA843FFFF007BD5555AAD57DF55AAAEBDFEF007BE8A10AAA",
INIT_3C => X"AAA975FF5D7BC21EFF7FBD7400F7FBC00BA55557DFF75D2E82010F7843DF45FF",
INIT_3D => X"5D2EAAA005D2AAAA185D2AAAA10F780021FFA2803DE10FFD16ABFF5D7BFDE10A",
INIT_3E => X"0000000000000000000000000000000000000007FE8BFF080028BFFAAFFEAA10",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(1),               -- Port A write enable input
DIA(0)   => data_write_a(8),        -- Port A data input
DOA(0)   => data_read_a_hi_512(8),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(1),               -- Port B write enable input
DIB(0)   => data_write_b(8),        -- Port B data input
DOB(0)   => data_read_b_hi_512(8),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_9_11 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00018248A2840112C00002C18000002300500030B3132000400812006",
INIT_01 => X"400008000000004C0020000000100248413C0A61590001D90213C10008110204",
INIT_02 => X"01A0042080010000054600C04008000004100000001020900200200002420804",
INIT_03 => X"024003400008012400000010E4004B0891000020610310000144C00000F5C000",
INIT_04 => X"1801800100E000000000510084000040010050020810200000C8900000320200",
INIT_05 => X"918004311104100000000000200008100800002000100000002C234415610820",
INIT_06 => X"81B00008080010100000980804000008800042041080001000100200322C2481",
INIT_07 => X"0000811800044080010000058600000086020002502080006000040800062C80",
INIT_08 => X"0000004001D4618008800A00061004044048002004000000000061F000000244",
INIT_09 => X"000040090802009420409004104444084001022400214A2080014400026401A2",
INIT_0A => X"04000071200000A003CA294140200800C80C8C8100004590111C040040120800",
INIT_0B => X"12210002404848502847040164880021150400080222000200C8034200000000",
INIT_0C => X"4610088010080421021040841021000841021000841021000841010800420820",
INIT_0D => X"42D0A16C529A321068500484000500D10042080040284000084900001A002196",
INIT_0E => X"00000002804000004228010410082002C000C0002400046419120410034285A1",
INIT_0F => X"A00000000500800800000800000000000002290008001080000000A010100042",
INIT_10 => X"00000000000004C2001000000240000000000000680800280000000140202000",
INIT_11 => X"0000C0000000000000000442020001000001000000000000010C800080000804",
INIT_12 => X"08000000000801A7802010000000152780102000000015000600000800000000",
INIT_13 => X"000000000101900011E0240000000009500011E0280000000009500004DD0000",
INIT_14 => X"000137400020000000000201C000136C00101000000000002340002947000240",
INIT_15 => X"0080881901210000000600C280028000419480D4000010040000000000002304",
INIT_16 => X"68DA368DA1685A1685A1685A1685A16C5A121A13A141950051309284A82C0010",
INIT_17 => X"85A1685A1685A1685A368DA368DA368DA368DA368DA368DA368DA368DA368DA3",
INIT_18 => X"5A1685A168DA368DA368DA368DA368DA368DA368DA3685A1685A1685A1685A16",
INIT_19 => X"0157344CCCF48DE68A895C38E2540A8010100000000000000000685A1685A168",
INIT_1A => X"14514514514514514514514514514514514D34D34D34D34D28E1004039248209",
INIT_1B => X"D268341A4D268341A0D069349A0D069349A0D068341A0D068341A0D068345145",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000014D490D069349A0D068341A4",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"EAABA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"03DE00FFAEBFFFF0800155FFAAFBE8B45002A974AAAA803DFFFAA843DF45FFFF",
INIT_29 => X"7BFDE00A2FBD7400F7FBFDFFFA2AEBDE00AAFBEAABA080000000087BEAA10F78",
INIT_2A => X"055401FFF7AEAAA10F780155EFAAAEA8ABAAAFBFDE0055556AA005D041555508",
INIT_2B => X"557FC0010F780154105D7FC2145005155555557BE8BEF007FFDEAAAAD1555EF0",
INIT_2C => X"AF7D5555FFF780154AA5D2AA8A10F7AA974AA082E80010A2AAAAA10552AA8AAA",
INIT_2D => X"BAF7D17FEBAA2AEBDF45002EAAABA087BFDF45F7AA974AAAAAA97555F784174B",
INIT_2E => X"000AAFFE8A00552EBFE00F7D17FF45F7FFFFF55AA80155FF080400145FFFBEAA",
INIT_2F => X"8FC7BE8A3DF7DF7F5E8A92000000000000000000000000000000000000000000",
INIT_30 => X"000280071E8A00EB8E3FE10F7AEBAFFF080A175D7BEF1E8B6D002090482B68E3",
INIT_31 => X"56AA10410E175550871FFE00A2FBD0400FFF5FDFC7B6A0BDE38B6F5E8A92080E",
INIT_32 => X"7BFAE82A2DB555C71C5B451D7FFAAA8A38FF8E175C7A2AAAAA82A2F1FAE105D5",
INIT_33 => X"2AEADA38492EA8AAA5571C2000FF8A17400557FC015514555757D5D71E8BEF14",
INIT_34 => X"B6A49256DEB84104BAFFD1525FFFF84174BA5D20AAA00E3AA904BA142A87010A",
INIT_35 => X"7000400155FFFBEDA82FFD57DEBAAAA0BFF7D0024ADA921C7BFFF55FFA095482",
INIT_36 => X"00000000000000000000A2FBE8A38492ABDE10EBDF7AF6DE3FFF8F7DB68A105D",
INIT_37 => X"BEF080402000F7AAA8B55FFAABDFEFF7D16AA000000000000000000000000000",
INIT_38 => X"FEAAFFD16AA00082E820BA08556AA00AAAABFE00F7AEAABEF082E95545F7D568",
INIT_39 => X"A8A10AAD568A00555168A10002E9754D00517DE00A2FFC2000F7D17FF55FF803",
INIT_3A => X"1575EF555568BEF5D7FE8A10AAFFD55555D7FD5555FFAAA8AAAFFAA97555A2AE",
INIT_3B => X"AE800AA552A97400A2AEBDEAA082EAAABA5D5140010F7AE974105D7BC21555D5",
INIT_3C => X"57BFDF55F78017400F780001FFAA84000AAFFD1401E7FF80174AA5D0028A00AA",
INIT_3D => X"AAFBEABFFF7AA80145080002145F7FBFFE00FFD17FEAAA2803DFEF08043FE005",
INIT_3E => X"0000000000000000000000000000000000000A2FFE8ABA082ABFE00AAFBEABFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(1),               -- Port A write enable input
DIA(0)   => data_write_a(9),        -- Port A data input
DOA(0)   => data_read_a_hi_512(9),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(1),               -- Port B write enable input
DIB(0)   => data_write_b(9),        -- Port B data input
DOB(0)   => data_read_b_hi_512(9),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_10_11 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00018248A2840112C00002C18000202300500030B3132000400992006",
INIT_01 => X"254008000000004C002000000010026840000000080000080200010008110204",
INIT_02 => X"0020042000010000004455800008000004100000000000900200000002400004",
INIT_03 => X"020001021089000021081000C400090011000000610001540104C00000F14400",
INIT_04 => X"0811800101A00002000050088554004200C840000000200080C8100000000001",
INIT_05 => X"030080001000100800009400200000000840E020201000000024024001200020",
INIT_06 => X"81B00008080012120004CC080492500280208004148000100000020020042493",
INIT_07 => X"0000000800044080010000048404081085020002502000006000040800062480",
INIT_08 => X"100202400084410808000A00021004044048000004000000000021F020408264",
INIT_09 => X"010040090002008420401004144440004040022484214A2080110108C2C00320",
INIT_0A => X"04004166A48A0001080000000000080080181881000045901118044040020800",
INIT_0B => X"1201000200484910000F0105602622291404020902005002018002400A022000",
INIT_0C => X"0440001011808020120004801120044800120004801120044800110002400884",
INIT_0D => X"008000440210100041308480800F82F00040180260A808008848000018002104",
INIT_0E => X"000000028040000002280104100820020000400020000440100204100A000100",
INIT_0F => X"040000000500800800000000000000000002280008000400000000A010100010",
INIT_10 => X"00000000000004C2001000010000000000000000680800010000000140202000",
INIT_11 => X"200000000000000000000442000001000000000000000000010C000080001000",
INIT_12 => X"00000000000801C0008000000000154000800000000015000410000800000000",
INIT_13 => X"0000000001019800180000080000000958001800000400000009580002800000",
INIT_14 => X"0000A0000000000000000201E0000A0000400000000000002360002080000800",
INIT_15 => X"0080881000000000000600C28102800060000000000800000000000000002306",
INIT_16 => X"401004010040100401004010040100441020D0030008840051309A90BA884010",
INIT_17 => X"0902409024090240900401004010040100401004010040100401004010040100",
INIT_18 => X"1004010040902409024090240902409024090240902409024090240902409024",
INIT_19 => X"F546890A940FE0D3971243555205428290100000000000000000401004010040",
INIT_1A => X"8A28A28A28A28A28A28A28A28A28A28A28A28A28A28A28A29554199854514514",
INIT_1B => X"2B95CAE532994CA6532995CAE572B94CA6532994CA6532994CA6532994CA28A2",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000002718E72B94CA6532994CA657",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"FDE1000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"03DFFFAA843DF45FFFFEAABA007FC2155F7D155545AA80001EFAAFBEAB45557F",
INIT_29 => X"042AB55FFD168B55AA8000010FFFBE8BFFF78402155AAFBE8B45002A974AAAA8",
INIT_2A => X"AD16AABA002ABDE10080000000087BEAA10F7803DE00FFAEBFFFF0800155FF00",
INIT_2B => X"A2FBD7400F7FBFDFFFA2AEBDE00AAFBEAABAA2FFD741055003DFEFF7AA801FFA",
INIT_2C => X"05D0415555007FD74105555555EFF7FBC0145F78028A00A2D142155087BFDE00",
INIT_2D => X"55AAD168ABA002A975FFF7AEBDEBAF780155EFAAAEA8ABAAAFBFDE0055556AA0",
INIT_2E => X"000557BE8BEF007FFDEAAAAD1555EF0055401FFF7AEAAA105D042ABFF5D556AB",
INIT_2F => X"71D7AAFBEFB455D71F8E00000000000000000000000000000000000000000000",
INIT_30 => X"E8B6D002090482B68E38FC7BE8A3DF7DF7F5E8A92007BC217DEBDB55555AA8E0",
INIT_31 => X"EBAFFF080A175D700042AB7DEBDB6DB55BE8E05000EBFFE8BC7E38E07145BEF1",
INIT_32 => X"0A3DFD7F7A4821D7A2D16FA82142EB8E00080E000280071E8A00EB8E3FE10F7A",
INIT_33 => X"ED1421450871FFE00A2FBD0400FFF5FDFC7B6A0BDE38B6F5E8A92B6FBD541049",
INIT_34 => X"A2F1FAE105D556AA10410E175550071D54104951555D7EBF5C5155E3842AA00B",
INIT_35 => X"8410E2ABD749516FB55BED16FA820820955EFE3AEBDEAAFF8E175C7A2AAAAA82",
INIT_36 => X"000000000000000000005D71E8BEF147BFAE82A2DB555C71C5B451D7FFAAA8A3",
INIT_37 => X"1EFA2FFD7545AAAE97555A2FBFDF455D556AA000000000000000000000000000",
INIT_38 => X"8B45AAAA95545F7D568BEF080402000F7AAA8B55FFAABDFEFF7D16AA00087FC0",
INIT_39 => X"6AA00AAAABFE00F7AEAABEF082E9554500042ABFFA2FFFFF45F7AE97400AAFFE",
INIT_3A => X"16AA00FFFBD5400082EBFF45F78400155A2D57FE00552EA8A00082E820BA0855",
INIT_3B => X"D557555A2802AA10FFD54214500517DE00A2FFC2000F7D17FF55FF803FEAAFFD",
INIT_3C => X"FAA97555A2AEA8A10AAD568A00555168A10002E9754D085155410085557555AA",
INIT_3D => X"5D7FD5555FFAAA8AAA002AAAB4508557DF55F7D17FE000804155FFAAAABDEAAF",
INIT_3E => X"0000000000000000000000000000000000000555568BEF5D7FE8A10AAFFD5555",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(1),               -- Port A write enable input
DIA(0)   => data_write_a(10),        -- Port A data input
DOA(0)   => data_read_a_hi_512(10),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(1),               -- Port B write enable input
DIB(0)   => data_write_b(10),        -- Port B data input
DOB(0)   => data_read_b_hi_512(10),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_11_11 : RAMB16_S1_S1
generic map (
INIT_00 => X"A101C4B05A0034CA2840712C2D001419000002300500030B31B20084EC992002",
INIT_01 => X"90000986B83028491800E0000C26426040000000080000088200080802512224",
INIT_02 => X"1A2004205E010640024D00800008000004100000040EC090820018003241A00C",
INIT_03 => X"28639100000C5C00000045C08400C8001100000061806A001618C03001E54400",
INIT_04 => X"1A800001000009A0804059A190000040400040008058220008C8100000120D4E",
INIT_05 => X"02000E81080250010000002022000058080400000E1200000020004401000004",
INIT_06 => X"819435143F20101010001008040800B8100102041088011100022200000024B2",
INIT_07 => X"90640D280884453E01064002944180008402001295BA100022E4340800062D82",
INIT_08 => X"400000093204802200280A0012160585C1D808D004000000000323F40C102244",
INIT_09 => X"380040098010001100009204107C5950400000220080C200800900020C006827",
INIT_0A => X"80007100004016EA080801010000080D00200081000045B0511D289940103399",
INIT_0B => X"002000024040410A000D0104408810C115D9C008050042400100D04E88000002",
INIT_0C => X"00655010009264201200C7B421ED0C7B421ED0C7B431ED087B43176843DA1085",
INIT_0D => X"0401020080400A10012494881A4F80F209500BB2602881A488485C1318002000",
INIT_0E => X"6619A540124814800228010410082022C00040002020090020220C9600040802",
INIT_0F => X"ACCC334A802491600C587949B6D0141B4CC600D5761B1599865A500490B86A56",
INIT_10 => X"BAC845542056A61686EC81E3A6CB68AA2C622C9A251C352B330CB4A0092170D8",
INIT_11 => X"BCCAD0B5A81536080CC6B21A21B1FC09CB0F1076D4A200B2AD4068F4101639B5",
INIT_12 => X"4D2CC281E31AA0103AB8D5514066380804B268A2E060901204112566F10AC418",
INIT_13 => X"D551443C47281002540B2C9AAAA8662A1152B202AE3554403028115AA88201A1",
INIT_14 => X"548A20A0492A2724A0621620402A020141F172FB182A32AB6845AB6200251BC9",
INIT_15 => X"00C00A000200074044E6801832728080D00A380B753952C4877E0104DDE4D124",
INIT_16 => X"0080200802008020080200802008020480080022020081010124988800400010",
INIT_17 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_18 => X"0000000000802008020080200802008020080200802008020080200802008020",
INIT_19 => X"55062608804180C0B10A42104201400204000000000000000000000000000000",
INIT_1A => X"00000000000000000000000000000000000820820820820801C4149470000000",
INIT_1B => X"0000000000000000040200000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000007E0F0000000000000100800",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"000AA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0001EFAAFBEAB45557FFDE10082ABDF5508557DF45002ABDFFFF7803DE10AA80",
INIT_29 => X"AEBFF45FFAEBFEAA002A801FFF7FFE8A10A28000000007FC2155F7D155545AA8",
INIT_2A => X"2AABFE10082ABFFEFAAFBE8B45002A974AAAA803DFFFAA843DF45FFFFEAABAA2",
INIT_2B => X"FFD168B55AA8000010FFFBE8BFFF78402155AAD155555A28428BFF002ABDE00A",
INIT_2C => X"F0800155FF00557FF45557FC2010002A80010A2842AAAA007BFFF4500042AB55",
INIT_2D => X"FF5D00154BAF7FBE8BEFFFD540000080000000087BEAA10F7803DE00FFAEBFFF",
INIT_2E => X"000A2FFD741055003DFEFF7AA801FFAAD16AABA002ABDE10A2D168A10A284021",
INIT_2F => X"DFC7F78E3FE28B684070AA000000000000000000000000000000000000000000",
INIT_30 => X"C217DEBDB55555AA8E071D7AAFBEFB455D71F8E00002EBDF6D005B78F7D142AB",
INIT_31 => X"A3DF7DF7F5E8A92BEAEBFF7DEBA0BDEAA1C2A801C7E3FFEFA10B68407038007B",
INIT_32 => X"8A28BFF082ABAE10B6AAB8E280820B8FEFBEF1E8B6D002090482B68E38FC7BE8",
INIT_33 => X"07FF8F7D00042AB7DEBDB6DB55BE8E05000EBFFE8BC7E38E07145B6D15756DA2",
INIT_34 => X"EB8E3FE10F7AEBAFFF080A175D708517DF7D497BC5028142A87000A28A2AA920",
INIT_35 => X"0B6DB6AA28A280001FF5D0A10482FFFFEFBC7E3DF42028080E000280071E8A00",
INIT_36 => X"00000000000000000000B6FBD5410490A3DFD7F7A4821D7A2D16FA82142EB8E0",
INIT_37 => X"FEF007BE8BFF5D2ABDF55F7AABDEAAF784154BA0000000000000000000000000",
INIT_38 => X"DE00FF84154BA087FC01EFA2FFD7545AAAE97555A2FBFDF455D556AA00082EBF",
INIT_39 => X"02000F7AAA8B55FFAABDFEFF7D16AA00FFAEBFFEFAA803DEBA5D2E82155A2FBF",
INIT_3A => X"A95545F7D5555FFAAAAA8BFF002AAAA00FFAAA8AAA080028BFFF7D568BEF0804",
INIT_3B => X"2E95400A2AEA8A00007FEABFF00042ABFFA2FFFFF45F7AE97400AAFFE8B45AAA",
INIT_3C => X"82E820BA08556AA00AAAABFE00F7AEAABEF082E9554508557DFFF007BD54BA5D",
INIT_3D => X"A2D57FE00552EA8A00FFFFE8AAAAA80001FF5D2E82000F7FFFFF45AAFFC20BA0",
INIT_3E => X"0000000000000000000000000000000000000FFFBD5400082EBFF45F78400155",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(1),               -- Port A write enable input
DIA(0)   => data_write_a(11),        -- Port A data input
DOA(0)   => data_read_a_hi_512(11),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(1),               -- Port B write enable input
DIB(0)   => data_write_b(11),        -- Port B data input
DOB(0)   => data_read_b_hi_512(11),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_12_11 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50080B01BC002006940202C0DE041196A83183000000023322287E0FC000006",
INIT_01 => X"75400D849830C84C5823E0000C17424840000000080000088200002802153231",
INIT_02 => X"18A026B43ED180040147558040090000061800000C06ED9802768F4472C52005",
INIT_03 => X"2A67E34A528D0524A52850528400C8001100000171C02B550618C91A10E55440",
INIT_04 => X"1BC0000100056C8280825DE98154004300C840800850240080CA921084520A07",
INIT_05 => X"02000F832000500C0000941024000852084060202E100001002000448100000C",
INIT_06 => X"819A1D1C3FE01A1A40045408049A50BA4020C6041090001200006200000000F2",
INIT_07 => X"C26A0719CC96CC6ED18A64019695A854870300FA3968B20068FC06080106249F",
INIT_08 => X"D002024B3E040800008C0A002610240D494A06F3460409000000E3F0AD5282E5",
INIT_09 => X"27A06009200040000400120412445D78400001000410420080218029CC807A27",
INIT_0A => X"18000006848A026F000000000000080000F010C100204593F11A6CDF48003BF8",
INIT_0B => X"000000820040402B28050400400432C9349DF21A31A00ACC0000F04F80020001",
INIT_0C => X"00357804611AE45D05D0833430CD0833420CD0C33420CD0833430668619A1000",
INIT_0D => X"0000000000000A74812DF00E87E80A079F9F90FA0280E87E800C7FF3B8002000",
INIT_0E => X"3B6B0E404D26160682082002000401EA0000C40000800A006002818808000000",
INIT_0F => X"A476D61C809A4DA84272592D6246FC1B17B541F97E1B348EDA93900B2B286C56",
INIT_10 => X"30C669E622DBC325CFD881A962454CFBE5403AB99594362B1DB52720165650D9",
INIT_11 => X"F8D2D39A3745261E4A95A110A3F855000E4B1D32BAB504BB7490FCFF912A3834",
INIT_12 => X"B90E9B018C7530200AB8F8BF41F9A22006B37DC8E1F9A21A70116D4C5080651C",
INIT_13 => X"118780319CCA08AB1001ACDF34B8F1C688AB1002AE3F7B807B6289F368828C4C",
INIT_14 => X"2AF020233376A5ECC016B1A827CDA21160F051DE610A34C50427E6E220323E4A",
INIT_15 => X"0077020000000439FDC05C5806781FAB46095A0B5199B0AC55521524F1864022",
INIT_16 => X"000000000000000000000000000000000026C000002884000130921092804010",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"8020080200000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0051B946088881360A95090CB054420290100000000000000000008020080200",
INIT_1A => X"041041041041041041041041041041041049249249249249200100002D451451",
INIT_1B => X"92C964B2592C964B2592C964B2592C964B2592C86432190C86432190C8641041",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000003800F592C964B2592C964B25",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"7DE1000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"ABDFFFF7803DE10AA80000AAAA843FE0008557DFFF0800020105D557FEAA0055",
INIT_29 => X"D5420000051555FFA2AA8200000557DFFFF7AA80000082ABDF5508557DF45002",
INIT_2A => X"82AA8AAAAAFFC00BA007FC2155F7D155545AA80001EFAAFBEAB45557FFDE10AA",
INIT_2B => X"FFAEBFEAA002A801FFF7FFE8A10A28000000A2D155410F7FFFFEBA08003FE000",
INIT_2C => X"5FFFFEAABA000028A105D2ABFE10A2AABFE1055516ABEF5D517DEAAA2AEBFF45",
INIT_2D => X"55002A820AA08557DFFFF7AA82155AAFBE8B45002A974AAAA803DFFFAA843DF4",
INIT_2E => X"000AAD155555A28428BFF002ABDE00A2AABFE10082ABFFEF0855420000004175",
INIT_2F => X"5010495B7AE921C517DE10000000000000000000000000000000000000000000",
INIT_30 => X"BDF6D005B78F7D142ABDFC7F78E3FE28B684070AABE803AE38145B78FD700000",
INIT_31 => X"BEFB455D71F8E00BED547038145B505FFB6A487000005F7AFD7F7A482038002E",
INIT_32 => X"F1FDE821C003FE001C2EAAAAAB6F5C2082007BC217DEBDB55555AA8E071D7AAF",
INIT_33 => X"D517DEAABEAEBFF7DEBA0BDEAA1C2A801C7E3FFEFA10B68407038B6D550428FF",
INIT_34 => X"B68E38FC7BE8A3DF7DF7F5E8A9200002FA285D20BDE28A2A4B8E10555B68BEF5",
INIT_35 => X"F085F47038140010555142082082005F7DFD7F7A482155BEF1E8B6D002090482",
INIT_36 => X"00000000000000000000B6D15756DA28A28BFF082ABAE10B6AAB8E280820B8FE",
INIT_37 => X"ABA5D7FEAB45080015410007FEAA0055517DE000000000000000000000000000",
INIT_38 => X"AB45F780020BA082EBFFEF007BE8BFF5D2ABDF55F7AABDEAAF784154BAF7802A",
INIT_39 => X"D7545AAAE97555A2FBFDF455D556AA00F7D1554BA5D7BC01FFFF8015410007FE",
INIT_3A => X"4154BAF7D1400BAFFD57FE005D043FE10552EAAAAAFFD140000087FC01EFA2FF",
INIT_3B => X"8428A105D7FEABEF55557DEBAFFAEBFFEFAA803DEBA5D2E82155A2FBFDE00FF8",
INIT_3C => X"7D568BEF080402000F7AAA8B55FFAABDFEFF7D16AA0008003FEBA55003DEBAA2",
INIT_3D => X"FFAAA8AAA080028BFF087BD54AA550402145550000010087FFFF45F78402145F",
INIT_3E => X"0000000000000000000000000000000000000F7D5555FFAAAAA8BFF002AAAA00",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(1),               -- Port A write enable input
DIA(0)   => data_write_a(12),        -- Port A data input
DOA(0)   => data_read_a_hi_512(12),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(1),               -- Port B write enable input
DIB(0)   => data_write_b(12),        -- Port B data input
DOB(0)   => data_read_b_hi_512(12),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_13_11 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10154A0441836CA2840512822007C18000E02700500030B31B300040081A042",
INIT_01 => X"00000804A000C04800020000000002404001000008220008A200100802110204",
INIT_02 => X"02200430000104000A4700804008000004100000000420918204D3033240400D",
INIT_03 => X"AA4003400008592400000590C40009141100000C6180C0000000C00001E14000",
INIT_04 => X"0800000102400120088054019000004160004190BAA0270000C8100000600206",
INIT_05 => X"21000012040610050040000227003AA0082400E94C1200000824424005220020",
INIT_06 => X"81963B180C001010580000080400000058000004109C00138000020024142581",
INIT_07 => X"002C8008000441600106400A9600010494020002B8AAA000EF003408000E2580",
INIT_08 => X"000000E48194408000A00A001210040441C80320040210000002ABF004102244",
INIT_09 => X"2A004009640040100400940412D4C4004000022000104200802D983000480120",
INIT_0A => X"8000202020401480000000000000080C90090881000145B0111A14004015080D",
INIT_0B => X"00000002004040AA08050400404040C11444000805200A402090024000008002",
INIT_0C => X"8410000A00280020020040800020040800020000801020000800010020400000",
INIT_0D => X"84A14250A055100050100490000500D00040080040290000084E4000B800610C",
INIT_0E => X"DCD13042BEDA36820228000000000000C000400081A08BC812A2092B02850942",
INIT_0F => X"89B9A260857DB400431969CA985D480949D32804A40AB137341C10B7D6A02EC0",
INIT_10 => X"E6ACA678001CE7D0296C213A460CA4271CA2168AEC1017606E6838216FAD4055",
INIT_11 => X"84AD4961C281B20213073C5FC0058008632D30D522CE80239DCC01AB013A4D20",
INIT_12 => X"2E6B13804A4B01D83461299900F6BD583A519104A0EEBD1A141010B2A4C8E116",
INIT_13 => X"89E5E40913419151EE0E94641828F72B5151EE0D184B321037AF5158BB02D085",
INIT_14 => X"562EC0B42162D68EE0073AE1C562EC13D521921A4170300B2B458B56B01C2280",
INIT_15 => X"00888A120240034000E6DC8285028014B82372011FC1E4F5E0A00929684EAF84",
INIT_16 => X"50942509425094250942509425094254940A1421420082020120908800480030",
INIT_17 => X"0942509425094250942509425094250942509425094250942509425094250942",
INIT_18 => X"9425094250942509425094250942509425094250942509425094250942509425",
INIT_19 => X"F7EFBBEEFF3F7DF7FF3E9F7DF7E2450228000000000000000000509425094250",
INIT_1A => X"BAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBF7DFDFDDD555555",
INIT_1B => X"EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAEBAE",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000000000F7EBF5FAFD7EBF5FAFD7",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"2ABEF00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0020105D557FEAA00557DE10AAD5554BA087FFFF55557BD54AAF7FBC01FFA280",
INIT_29 => X"7BD75EF087FFFFEF557BEAB45552E80155AA802AB45AA843FE0008557DFFF080",
INIT_2A => X"FAE820AA5D5557555082ABDF5508557DF45002ABDFFFF7803DE10AA80000AA08",
INIT_2B => X"0051555FFA2AA8200000557DFFFF7AA80000AAD1420AA087BD7555FFD168AAAF",
INIT_2C => X"5557FFDE10AAAEA8BFFA2FBD7545FFD157555085140010F7AEAABFFAAD542000",
INIT_2D => X"BA557BE8A10A284154BAFFAAAAB45007FC2155F7D155545AA80001EFAAFBEAB4",
INIT_2E => X"000A2D155410F7FFFFEBA08003FE00082AA8AAAAAFFC00BA00002AAAAF7D5574",
INIT_2F => X"0492E3F1C71C7BE8A2ABD7000000000000000000000000000000000000000000",
INIT_30 => X"3AE38145B78FD7000005010495B7AE921C517DE10A2DB50482147FFAF554971D",
INIT_31 => X"E3FE28B684070AA1C71D25D7007FFAFD7497BE8B5555208217DBE8A2AB45BE80",
INIT_32 => X"7FD257DFFD568A82FFA4870BA555F5056D002EBDF6D005B78F7D142ABDFC7F78",
INIT_33 => X"FAAAFBFFBED547038145B505FFB6A487000005F7AFD7F7A482038AADF4709214",
INIT_34 => X"AA8E071D7AAFBEFB455D71F8E00A2A0ADBC7A2FFD257DE3DF52555085142000F",
INIT_35 => X"21C002AA92FFDF574824171EAA10B680124BAFFAAAFB45007BC217DEBDB55555",
INIT_36 => X"00000000000000000000B6D550428FFF1FDE821C003FE001C2EAAAAAB6F5C208",
INIT_37 => X"0105D7BE8B55085142010AAD157545F7AEA8B550000000000000000000000000",
INIT_38 => X"01EFF7AAA8B55F7802AABA5D7FEAB45080015410007FEAA0055517DE00A2FFC0",
INIT_39 => X"E8BFF5D2ABDF55F7AABDEAAF784154BA5D5140145007BE8B55087BEAB555D040",
INIT_3A => X"0020BAA2FFD54105D7FC21EFFFD16AA10FF80174AA557FC21EF082EBFFEF007B",
INIT_3B => X"FBC0155085540000FFAEBFFEFF7D1554BA5D7BC01FFFF8015410007FEAB45F78",
INIT_3C => X"87FC01EFA2FFD7545AAAE97555A2FBFDF455D556AA00A2803FF45AAFFC21EFAA",
INIT_3D => X"552EAAAAAFFD1400005D042AA00F7FBD5410085568A10FF80020AAFFAABFF550",
INIT_3E => X"0000000000000000000000000000000000000F7D1400BAFFD57FE005D043FE10",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(1),               -- Port A write enable input
DIA(0)   => data_write_a(13),        -- Port A data input
DOA(0)   => data_read_a_hi_512(13),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(1),               -- Port B write enable input
DIB(0)   => data_write_b(13),        -- Port B data input
DOB(0)   => data_read_b_hi_512(13),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_14_11 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10020A000180000284008280000281800000030000000033022000000580002",
INIT_01 => X"000008020000204D006800000030824840000000084000084200090008510200",
INIT_02 => X"0220043170010A600A4D008040080000041000000028009002000F333240800C",
INIT_03 => X"111813400008002400000000C400090011000000610200001104D83000F14000",
INIT_04 => X"0801800100A000000000540084000040000040000800200000C8100000000748",
INIT_05 => X"0100000000001000000000002000080008000000001000000024024001200020",
INIT_06 => X"819EB84028001010000000080400000000000004108000100000020020040081",
INIT_07 => X"92040608000440100102400A94810206844200021DA2A0002000340800062C80",
INIT_08 => X"000000000084400008800A001214040441481500040000000000A7F408002244",
INIT_09 => X"0A0040090002008420401004104444004000020400214A208001000002400120",
INIT_0A => X"0400002020000000000000000000080C8008088100004590111B480040120000",
INIT_0B => X"1000000200404800000504016000002114000008020000020080024000000000",
INIT_0C => X"0410000010000000000040001000000000000040000000000001000000000000",
INIT_0D => X"04810244825010004010000000000000000000000000000000080000B8002104",
INIT_0E => X"0002C38280001202020800000000001000004000000000401022000002040902",
INIT_0F => X"20000587050001404E8084341CBA3404800828805200008000E0E0A000080002",
INIT_10 => X"4D18178E012010C00224004091C3514072C000444A0400080001C1C140001000",
INIT_11 => X"51709A07424142084458476001003809D0104B01C5710044020C4006010500C5",
INIT_12 => X"C26EE3803180C18006519462A00005001460E4730000050A1011004001060049",
INIT_13 => X"01F9E00660318000000538318740000140000001B4600CE80001400000002B62",
INIT_14 => X"0000000AD89857B0E0684411800000003799EB764D000330C300000000E3554B",
INIT_15 => X"0000021002002C000024008284001A0902000422E3F5960080480A0216A07240",
INIT_16 => X"4090240902409024090240902409024090081021020080015134920800480010",
INIT_17 => X"0902409024090240902409024090240902409024090240902409024090240902",
INIT_18 => X"9024090240902409024090240902409024090240902409024090240902409024",
INIT_19 => X"F5579B4E5C8FF0F7BE9D5F7DF650400200000000000000000000409024090240",
INIT_1A => X"9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7BF7DDDDDFCF3CF3D",
INIT_1B => X"F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE79E7",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000003FFF03F9FCFE7F3F9FCFE7F3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"420BA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"BD54AAF7FBC01FFA2802ABEFA2FBE8B55A2AE80000F7D5555555D2AAAABAAAD1",
INIT_29 => X"AA801FFA28402000AAAE955455500155EF0804155EFAAD5554BA087FFFF55557",
INIT_2A => X"7AEA8B45080417400AA843FE0008557DFFF0800020105D557FEAA00557DE10A2",
INIT_2B => X"087FFFFEF557BEAB45552E80155AA802AB4500516AA00A2AE800BAFFFFC20BAF",
INIT_2C => X"0AA80000AA005568ABAA28402010A2843FEBAFFFBD7410A2D168BFF087BD75EF",
INIT_2D => X"005D7FFDF4555517DFEF00043FEAA082ABDF5508557DF45002ABDFFFF7803DE1",
INIT_2E => X"000AAD1420AA087BD7555FFD168AAAFFAE820AA5D5557555002E80155A280000",
INIT_2F => X"0555412AA8ABAAADB40092000000000000000000000000000000000000000000",
INIT_30 => X"50482147FFAF554971D0492E3F1C71C7BE8A2ABD7A2FFEDB55B6A080038E3DB5",
INIT_31 => X"B7AE921C517DE10A2AE851FFB68402038AAAA955554900105FF0800175D7A2DB",
INIT_32 => X"A0800BAE3F1C0092EBAAADB6D080A12410BE803AE38145B78FD7000005010495",
INIT_33 => X"2D568BC71C71D25D7007FFAFD7497BE8B5555208217DBE8A2AB451C556FA00A2",
INIT_34 => X"142ABDFC7F78E3FE28B684070AA00516DABAA28402038B6803DE82F7F5D5410A",
INIT_35 => X"D002A80155B680000105D7FF8F455D5F78FD7000E3FEAA002EBDF6D005B78F7D",
INIT_36 => X"00000000000000000000AADF47092147FD257DFFD568A82FFA4870BA555F5056",
INIT_37 => X"F55FF84000AAAAFBC0145002AA8AAAAAFFC20000000000000000000000000000",
INIT_38 => X"01EF080417555A2FFC00105D7BE8B55085142010AAD157545F7AEA8B55A2FBFF",
INIT_39 => X"EAB45080015410007FEAA0055517DE00A2AA955FFFF80020BAAAAA9754508000",
INIT_3A => X"AA8B555D557FE00A280020BAAAD140000A2AEBFFEF082A82010F7802AABA5D7F",
INIT_3B => X"803DE00FFD557400AAD56AB455D5140145007BE8B55087BEAB555D04001EFF7A",
INIT_3C => X"82EBFFEF007BE8BFF5D2ABDF55F7AABDEAAF784154BA08557FEAAA284000AAFF",
INIT_3D => X"FF80174AA557FC21EF082A80145F780020105D7BEAB45557BE8B45082EBFEBA0",
INIT_3E => X"0000000000000000000000000000000000000A2FFD54105D7FC21EFFFD16AA10",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(1),               -- Port A write enable input
DIA(0)   => data_write_a(14),        -- Port A data input
DOA(0)   => data_read_a_hi_512(14),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(1),               -- Port B write enable input
DIB(0)   => data_write_b(14),        -- Port B data input
DOB(0)   => data_read_b_hi_512(14),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_15_11 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000A000000000284000280000001800020030000000033022000000180002",
INIT_01 => X"8000080000000048000000000000026040000000080000080200000000110200",
INIT_02 => X"0020042004010E60004C0080000800000410000000020090020000300245E005",
INIT_03 => X"0000010000080400000000408400480111000000610008000000C00000E54400",
INIT_04 => X"980000010000000088C2550080000040000040000008A00028C8100000120000",
INIT_05 => X"020004012E025000000001322000000A28008000011000000220004D41000000",
INIT_06 => X"819588000800101000011008040000100001060418800510000A620000000092",
INIT_07 => X"0000000800044004010C20008440810284020002102220002000340800062480",
INIT_08 => X"0000000001140800002C0A001214050540C800400406180000002DF004000244",
INIT_09 => X"1E00400900000000000016041044400440000000000042008001000000000022",
INIT_0A => X"0000000000000220000000000000080C00000081000045901118000040000000",
INIT_0B => X"0000000200404000010500004000000114000009000000000000004200000000",
INIT_0C => X"0000000000000000000040001000040001000000000000000001000020000800",
INIT_0D => X"000000000000001001208000180800000000030200000180800C400030002000",
INIT_0E => X"0000000000002600020800000000001080004000000000000002000000000000",
INIT_0F => X"A400000000000000000008000000000000000000000014800000000000000052",
INIT_10 => X"0000000000000000000000010240000000000000000000290000000000000000",
INIT_11 => X"2001C05838120800000000000000000000010000000000000000000000001804",
INIT_12 => X"081004000000000000A010000000000000902000000000180010002020000000",
INIT_13 => X"6600000000000000000024080000000000000000280400000000000000000000",
INIT_14 => X"0000000000200801000000000000000000501001920000000000000000000A40",
INIT_15 => X"0000020000000000000000003000000000000000000A101C3614000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000080000120980000000010",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000400200000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"28BEF00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"5555555D2AAAABAAAD1420BAFF8000010082A954BA00003DFEF085155400F784",
INIT_29 => X"AE95555A2FBE8BEFA2843DE00AA8015400FF84001EFA2FBE8B55A2AE80000F7D",
INIT_2A => X"2FBEAB45F7D56AABAAAD5554BA087FFFF55557BD54AAF7FBC01FFA2802ABEFF7",
INIT_2B => X"A28402000AAAE955455500155EF0804155EFFFFBE8BFF0800174AA557BFDE10A",
INIT_2C => X"A00557DE10F7D1574AAA2D16AB55FFD568BEF087FE8A1055003FE00A2AA801FF",
INIT_2D => X"00AA802AA00AAAE800BA5D0015545AA843FE0008557DFFF0800020105D557FEA",
INIT_2E => X"00000516AA00A2AE800BAFFFFC20BAF7AEA8B45080417400FFFFC21450800154",
INIT_2F => X"8FD7005150438F78A2DBFF000000000000000000000000000000000000000000",
INIT_30 => X"EDB55B6A080038E3DB50555412AA8ABAAADB40092E38E070280024904AA1C043",
INIT_31 => X"1C71C7BE8A2ABD7E3AA9257DA2FFE8BC7BE8E38E10A28017400E38A051FFA2FF",
INIT_32 => X"00124AA557FFDE10A2FBEDB6DF7D16AABAA2DB50482147FFAF554971D0492E3F",
INIT_33 => X"10038E38A2AE851FFB68402038AAAA955554900105FF0800175D7E3FFEFBD700",
INIT_34 => X"000005010495B7AE921C517DE10FFDF50482A2DB6AB45FFD56DBD7087BEAA384",
INIT_35 => X"0FFF1C017D140410400BE8E28A10AAA085082550A1057DBE803AE38145B78FD7",
INIT_36 => X"000000000000000000001C556FA00A2A0800BAE3F1C0092EBAAADB6D080A1241",
INIT_37 => X"4AA0800020BA550028B550855400AAF7AEBDFEF0000000000000000000000000",
INIT_38 => X"7400AAAE975EFA2FBFFF55FF84000AAAAFBC0145002AA8AAAAAFFC2000AAAA97",
INIT_39 => X"E8B55085142010AAD157545F7AEA8B55AAAE821EFAAFBEAB55F7AAA8A00AA841",
INIT_3A => X"417555AAFFFDF450804020AA557BFFE10A2FFFFFEFF7D568ABAA2FFC00105D7B",
INIT_3B => X"D17DF45007FE8AAA08002AAAAA2AA955FFFF80020BAAAAA975450800001EF080",
INIT_3C => X"7802AABA5D7FEAB45080015410007FEAA0055517DE00FFFBC2000AAFBE8B55F7",
INIT_3D => X"A2AEBFFEF082A82010FFD5421EF5D0000010F7AAA8A10AA8017400552A801EFF",
INIT_3E => X"00000000000000000000000000000000000005D557FE00A280020BAAAD140000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(1),               -- Port A write enable input
DIA(0)   => data_write_a(15),        -- Port A data input
DOA(0)   => data_read_a_hi_512(15),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(1),               -- Port B write enable input
DIB(0)   => data_write_b(15),        -- Port B data input
DOB(0)   => data_read_b_hi_512(15),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_16_11 : RAMB16_S1_S1
generic map (
INIT_00 => X"DA22C618B1000482B688B186588884862A400438255FC38381441205BA803003",
INIT_01 => X"7045A80028404C211203A952A90341080B173340412000E1005D628000820484",
INIT_02 => X"428406A4000850848330118D0AAC55001349B108818005460229044001C01784",
INIT_03 => X"092C4020000500020000500986812C405000001A48202050000A214AC0650115",
INIT_04 => X"4804A55440256F504025E003A054F46415A4E62B6FE3307943965A00001A1152",
INIT_05 => X"0000001C40A5B950ADB8EA097057ECE14C86D2B7F85AAD17F4B100000B88148C",
INIT_06 => X"415401DCDCF2C0A8030140BCB0820A200342A1C641C1E8782F508F2B00003584",
INIT_07 => X"002701881A3202080AE00480A2002840BE1480FA004342AA6F12000054004867",
INIT_08 => X"08C54828091002000002B32A8C19064E486A8001510000014140C1E2A14891E0",
INIT_09 => X"015452B103020814004088B64102680B6596594800400413CAC0208944800000",
INIT_0A => X"96AA000484094C000000000000012C9000A0000D0A80000BF8028E87C1B99270",
INIT_0B => X"014808A02004200E540480212000A448C0082024AE50064B44000000000002A2",
INIT_0C => X"0004000D5846256AAEA811150445411150445411150445411150422A088A8200",
INIT_0D => X"00000004010042A204A0C5817D00005034052E40000817D00440004004AD3240",
INIT_0E => X"632B2673FA4587978A2004102800809225545155121740000004900090000000",
INIT_0F => X"00C6564CE7F4EA4B940076D296D003030800462CBD320018CAAAACFE9164C800",
INIT_10 => X"28834ADB1440A114793A4A30A40839AA14910D08DCB2640031955559FD3AC990",
INIT_11 => X"594AB0B1A025371CA0E034E8443C097A800EB090D4AAC91208ED2FA0CE5E09B1",
INIT_12 => X"7B50446083001B94BB38C540EBE61284BB304880E3E4579EDC00992980D58033",
INIT_13 => X"5511121840E7A2CD952ECC12ABC3E6ACB3DFB12ECE315000F61FF1727A85FDBC",
INIT_14 => X"75DEB07F6F2E7084517F126F8395CB2BEFBAB8BA8AF698228CC5E2F08ECA5159",
INIT_15 => X"5580A840A8009F8B108C80A1021B080AFC0DF6422C6077F4A77F20D0C0E21084",
INIT_16 => X"0000000000000000000000000000000000044000102A0001148442A110810359",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"558D11544C690DA64C1C4F68A360400000000000000000000000000000000000",
INIT_1A => X"14D14D14D14D14D14D14D14D14D14D14D14514514514514529E5F87869E79E78",
INIT_1B => X"D1E8F47A3D1E8F47A7D3E9F4FA7D3E9F4FA7D3E9F47A7D1E9F47A7D1E9F4D14D",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000007D3E9F4FA7D3E8F47A3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"C00AA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"03DFEF085155400F78428BEF087FFFFEFF7D168B55AAD17FFFF552EBFE00007F",
INIT_29 => X"2E975EFF7D568BFFFF80175EF0004000BA552A821FFFF8000010082A954BA000",
INIT_2A => X"55540000082EAABFFA2FBE8B55A2AE80000F7D5555555D2AAAABAAAD1420BA5D",
INIT_2B => X"A2FBE8BEFA2843DE00AA8015400FF84001EF0000020AA5D00154005D043FF455",
INIT_2C => X"FA2802ABEF557BEABEF5D0415410087FD74BAAAAEBFFEF557FC00AAF7AE95555",
INIT_2D => X"FFFFAABFEAAFF84001FF002A821FFAAD5554BA087FFFF55557BD54AAF7FBC01F",
INIT_2E => X"000FFFBE8BFF0800174AA557BFDE10A2FBEAB45F7D56AABA082A97545F7D16AB",
INIT_2F => X"FFEF552AB8E38087FC2092000000000000000000000000000000000000000000",
INIT_30 => X"070280024904AA1C0438FD7005150438F78A2DBFF0871F8FC7E3D56AB6DBEDB7",
INIT_31 => X"AA8ABAAADB400924920925EFF7D16ABFFE38E175EF1400000BA412E871FFE38E",
INIT_32 => X"0A1240055003FF6D5551420101C2EAFBD7A2FFEDB55B6A080038E3DB50555412",
INIT_33 => X"57FC00BAE3AA9257DA2FFE8BC7BE8E38E10A28017400E38A051FF0804050BA41",
INIT_34 => X"4971D0492E3F1C71C7BE8A2ABD74975EDBC7550E12410087FD74AAB6AABFFC75",
INIT_35 => X"A08249756DF7D168BC7F7AABAEAAF780051C70824851D7A2DB50482147FFAF55",
INIT_36 => X"00000000000000000000E3FFEFBD70000124AA557FFDE10A2FBEDB6DF7D16AAB",
INIT_37 => X"B55A2D16ABEFFFFBFDFFF552AAAAAA007BC00000000000000000000000000000",
INIT_38 => X"20AA002A955EFAAAA974AA0800020BA550028B550855400AAF7AEBDFEF08516A",
INIT_39 => X"000AAAAFBC0145002AA8AAAAAFFC20000000021EFF7D568BFFA2AA955FF5D040",
INIT_3A => X"E975EF0800174BA002E820105D003DFEF5D51420005D2ABFF45A2FBFFF55FF84",
INIT_3B => X"7BD74AAF7AEBDF455D7BC20BAAAAE821EFAAFBEAB55F7AAA8A00AA8417400AAA",
INIT_3C => X"2FFC00105D7BE8B55085142010AAD157545F7AEA8B5500557DF45552A8200000",
INIT_3D => X"A2FFFFFEFF7D568ABA0804155FFF7D568B55FFAAAAABAFF8415545000015555A",
INIT_3E => X"0000000000000000000000000000000000000AAFFFDF450804020AA557BFFE10",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(2),               -- Port A write enable input
DIA(0)   => data_write_a(16),        -- Port A data input
DOA(0)   => data_read_a_hi_512(16),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(2),               -- Port B write enable input
DIB(0)   => data_write_b(16),        -- Port B data input
DOB(0)   => data_read_b_hi_512(16),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_17_11 : RAMB16_S1_S1
generic map (
INIT_00 => X"5284CE4FB7BD2C8994A13392DBD02E14006B82AC7E800D44D3DD2FD5F9B961C0",
INIT_01 => X"2EACD01F7E03FC6793F2199B39FC233C11D93AE6F3BB92B32091DBC339B24542",
INIT_02 => X"E63CCCC00A82C08092A2AFAE667033DB50853379C10BFDC5C6F4044443C817C6",
INIT_03 => X"7FF183635AEF9E3635AEF9E18E237040404446965C0607EE6DB7854AC4DE060C",
INIT_04 => X"D78AC33FB604488B000892EF17BE6D84196482236FE100294152E294350FB697",
INIT_05 => X"081B5F9B409420D0CDB47A05403F6CE0C08A4AB7F840EDB6F48100DFC8081081",
INIT_06 => X"768465354781CBC30316367077B4BDB50646E8D87100A8201ED01C19C020F71A",
INIT_07 => X"4002A110C922480A82D0841147162C48EBB9537A0022DC67987042EE976ABEA7",
INIT_08 => X"DB931BFEF91C00002CC0E019C0C82A4E4820C15A2330E004401891181168C4D1",
INIT_09 => X"09F3A1BC11EFBC66DB65307071477FF1030C397C060B4254064302042F803A69",
INIT_0A => X"3F330802162F3B7EE3F3EC7C7DEF207000F00059D2ED56D7EED2ED3C9A867DC0",
INIT_0B => X"185C44B91BC1740B7605040BE0018CFC7429F326B9E822FFC00074D5A0AB033A",
INIT_0C => X"00367A28FC1B7F7FEFFCFBFF3EFFCFBFF3EFFCFBFF3EFFCFBFF3EFFE7DFF9E00",
INIT_0D => X"0000000008004BA78428C7AD7FC94B533F5B4FFBD2FAD7FCCA786D43FE67C218",
INIT_0E => X"BA494CEBFD4F2667ABB6F68B29760593F33FA0CF170F40006001B1A05C000000",
INIT_0F => X"7F749299D7FAEB237DFE5865B6D2BF23265CBACE542A6FEE92333AFF33E0A9BF",
INIT_10 => X"F6C24B6D18C3C9F8E2881F3F787D776B5DB94A09955054DFDD246675FE7AC153",
INIT_11 => X"BFB349E08FF9A27EDE9FA8AEFD9E7467BFCB195CFEB56A1A70D34D1706FFFA3E",
INIT_12 => X"6FE219CA80725B875EED723FF7FCB2875EDAAFEAF7FD929BFD55BBC71D79F639",
INIT_13 => X"546670D018E7A6E581D7B6AB75FDFCECA6E581D7BB5DDFC6FF0EB7D7E859FDB5",
INIT_14 => X"B978177F6D6AF5ECDB5FB76A5F5FA165B456E0FB308710C49FCFB741598B9C7E",
INIT_15 => X"CFDAAB00AC00A8BBFC8B501CF7A0FED9A540EA1952586CEB54D143ACFF9A3BA9",
INIT_16 => X"000000000000000000000000000000000026E100002F382DBD9ECFE117805F20",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"4372003009EDCC4052E917114F981800C0000000000000000000000000000000",
INIT_1A => X"BA69A69AEBA69AEBA69A69AEBA69AEBA69A69A69A69A69A68698686981D75D74",
INIT_1B => X"6A351A8D46A351A8D068341A0D068341A0D068341A0D46A341A0D46A341A69AE",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000000000046A351A8D46A351A8D4",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"7FEAA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"17FFFF552EBFE00007FC00AA087FFFFFFFFFFFFFEFF7FBEAB450804001EFAAD5",
INIT_29 => X"D168A000004020AA5D7BE8B450051401EF087FD74AA087FFFFEFF7D168B55AAD",
INIT_2A => X"D7FEAB55FF80175EFFF8000010082A954BA00003DFEF085155400F78428BEFAA",
INIT_2B => X"F7D568BFFFF80175EF0004000BA552A821FF5D00020BA552A82000552A821555",
INIT_2C => X"AAAD1420BAFFFFFDF45AAD17FFFFAAFBC01EF5D0015555557BFDEBA5D2E975EF",
INIT_2D => X"BA007FEABEF005555555A2D1554BAA2FBE8B55A2AE80000F7D5555555D2AAAAB",
INIT_2E => X"0000000020AA5D00154005D043FF45555540000082EAABFF00516AA10552E820",
INIT_2F => X"8B550000071EFB6DF7AE92000000000000000000000000000000000000000000",
INIT_30 => X"F8FC7E3D56AB6DBEDB7FFEF552AB8E38087FC2092147FFFFFFFFFBFDFC7EBF5E",
INIT_31 => X"150438F78A2DBFFBED16AA381C0A07082497FEFB6D1451471EF007BD04920871",
INIT_32 => X"2A850105D2A80155417BEFB6DEB8E175FFE38E070280024904AA1C0438FD7005",
INIT_33 => X"D7BFAEBA4920925EFF7D16ABFFE38E175EF1400000BA412E871FF550A0009249",
INIT_34 => X"E3DB50555412AA8ABAAADB40092FFF5FFF6DAADF7FFD7B6F1C71EF55001756D5",
INIT_35 => X"7145B6AA28492487082007FEDBD700515556DA2DF50492A2FFEDB55B6A080038",
INIT_36 => X"000000000000000000000804050BA410A1240055003FF6D5551420101C2EAFBD",
INIT_37 => X"FEFF7FBFFF55A2D16AB550000175EFFFFBEAA000000000000000000000000000",
INIT_38 => X"55EF087FC200008516AB55A2D16ABEFFFFBFDFFF552AAAAAA007BC0000557FFD",
INIT_39 => X"020BA550028B550855400AAF7AEBDFEFF7D568AAA5D2A97410007BFFFFF55515",
INIT_3A => X"A955EF5D2E80010002A954005D2A82155087FFFFEFAAAA975EFAAAA974AA0800",
INIT_3B => X"D1575FF5504175EF5D7FEAAAA0000021EFF7D568BFFA2AA955FF5D04020AA002",
INIT_3C => X"2FBFFF55FF84000AAAAFBC0145002AA8AAAAAFFC2000FFD57DFFFAAFFFDF55FF",
INIT_3D => X"5D51420005D2ABFF45557FE8AAA000415410007BFFF450051555EFA2FBC0000A",
INIT_3E => X"00000000000000000000000000000000000000800174BA002E820105D003DFEF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(2),               -- Port A write enable input
DIA(0)   => data_write_a(17),        -- Port A data input
DOA(0)   => data_read_a_hi_512(17),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(2),               -- Port B write enable input
DIB(0)   => data_write_b(17),        -- Port B data input
DOB(0)   => data_read_b_hi_512(17),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_18_11 : RAMB16_S1_S1
generic map (
INIT_00 => X"69844019080000A21A611406840014122A641074155FC28A2024001001801003",
INIT_01 => X"7443D920034004180005E9E3C90360C0041C0181002001602025800008440084",
INIT_02 => X"E2DCCCE61D5C008103F2000781FC0FEDEAC2161B0B8FB0008620044443006010",
INIT_03 => X"884E300802006900802006995C896D605200000856E24A040000640052141103",
INIT_04 => X"480520FC026125AC0025C9122644E3E40EC8E2001001302281841A009038A86A",
INIT_05 => X"432000040089983070019400F01010004C8DB841405A80A100B586200FAC24AE",
INIT_06 => X"09044359DC7040000000002C109B0E0A00A1104641C0803804000707284600E1",
INIT_07 => X"400D10100400481D5EB08501620000007500CE801241021FE78E404860140060",
INIT_08 => X"00880C0106A0528020019307CC082A0A4A6A01ED725021400040D028000A9729",
INIT_09 => X"00117063038000282081402E4106400B6186128040600C10C1C0200950508110",
INIT_0A => X"C0C30C2E21580C874004008080003C32A10A19090C02010E1022944061688000",
INIT_0B => X"0180A8062026000DC425C0301311324AA2373088479105D044A1022000001835",
INIT_0C => X"0D89844703649000000200000000000000000000000000000000000000000010",
INIT_0D => X"0D8306C182701404C1973010802020404084001E00010802046092B5001FB365",
INIT_0E => X"528EB314068AB8B803DB00002900800400FC503F08180050942E4200020C1B06",
INIT_0F => X"40A51D66280D6032C5F96D3C51555D5D7D5AA87285820814A3CCC501C2A60820",
INIT_10 => X"8B35A3FEBF1FEDFD9C2B30E0468AAAD5D48F37E8FC1304102947998A03984C10",
INIT_11 => X"440FE1DD772D37A0A321BC6968F32658BF2D4F2A80BF8FE3F9FE3AC362080529",
INIT_12 => X"5487910D7E5A6D961A28456A1832E5161A100DD5182BC54020EA67A189C6ED36",
INIT_13 => X"AA444CAF91EDD1B725868403BE06323551B725868A100ABD119753B70964122B",
INIT_14 => X"EDC259048ACD868EE3803D65CEDC258A8F80D55E007C3F8EBB56F4C5362C978F",
INIT_15 => X"3F240014BE84370001B6922070440556B15F7FABBC0031BCF2257C41634B14D4",
INIT_16 => X"C1B06C1B06C1B06C1B06C1B06C1B06C1B0491069068000004060300A005A0118",
INIT_17 => X"1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06",
INIT_18 => X"B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C",
INIT_19 => X"B28BBECEB80EE173C2300F7DF16000000000000000000000000041B06C1B06C1",
INIT_1A => X"8A28A28AAAAAAA28A28A28AAAAAAA28A28A28A28A28A28A2910591505C104104",
INIT_1B => X"28944A25128944A25128944A25128944A25128944A2552A954AA5128944AAAA2",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000128944A25128944A251",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"9540000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"BEAB450804001EFAAD57FEAA087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974BA082E",
INIT_29 => X"7FFFFFFFFFBFDF45AAD568B55080028B55002E82000087FFFFFFFFFFFFFEFF7F",
INIT_2A => X"0043DE10AA843DE00087FFFFEFF7D168B55AAD17FFFF552EBFE00007FC00AA08",
INIT_2B => X"0004020AA5D7BE8B450051401EF087FD74AAAAFFFDF45A2D16AB55F7FFFFFFF0",
INIT_2C => X"0F78428BEFAA80000000804154BA55042ABEF5D7FD75FFAAD540145AAD168A00",
INIT_2D => X"00082E95555085168A10557FD7545FF8000010082A954BA00003DFEF08515540",
INIT_2E => X"0005D00020BA552A82000552A821555D7FEAB55FF80175EF5D00020105D2A974",
INIT_2F => X"DFFF5D2A954AA082A92428000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFBFDFC7EBF5E8B550000071EFB6DF7AE921C7FFFFFFFFFFFFFFFF7FBF",
INIT_31 => X"AB8E38087FC2092087FFDFC7E3F1FAF55A2DF6DB7D1C002AB7D002A82028147F",
INIT_32 => X"DF6DB7DE3F5FAFC708003DE28B68E38E280871F8FC7E3D56AB6DBEDB7FFEF552",
INIT_33 => X"ADF4516DBED16AA381C0A07082497FEFB6D1451471EF007BD0492B6F1F8F55AA",
INIT_34 => X"1C0438FD7005150438F78A2DBFFA28407038140410492550A2ABC7497BD25FFA",
INIT_35 => X"F5D0E05000492097428002E9557D1C516FA28417BD5545E38E070280024904AA",
INIT_36 => X"00000000000000000000550A00092492A850105D2A80155417BEFB6DEB8E175F",
INIT_37 => X"FFFFFFFFDFEFF7FBFFFEF552E974AA082A820AA0000000000000000000000000",
INIT_38 => X"ABEF002A800AA557FFDFEFF7FBFFF55A2D16AB550000175EFFFFBEAA00557FFF",
INIT_39 => X"6ABEFFFFBFDFFF552AAAAAA007BC0000087BFDF45AAD568B55AAFBFDFEF55042",
INIT_3A => X"FC2000FFD56AB45A2FFFDFFFAAD16AB4500043DEAAFFAEAAAAA08516AB55A2D1",
INIT_3B => X"2AA8B45087FC01EFA2FFD55EFF7D568AAA5D2A97410007BFFFFF5551555EF087",
INIT_3C => X"AAA974AA0800020BA550028B550855400AAF7AEBDFEFA280154BA55040000055",
INIT_3D => X"087FFFFEFAAAA975EF5D2E974000804154BA082A975EF5D517DEAA007BD5545A",
INIT_3E => X"00000000000000000000000000000000000005D2E80010002A954005D2A82155",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(2),               -- Port A write enable input
DIA(0)   => data_write_a(18),        -- Port A data input
DOA(0)   => data_read_a_hi_512(18),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(2),               -- Port B write enable input
DIB(0)   => data_write_b(18),        -- Port B data input
DOB(0)   => data_read_b_hi_512(18),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_19_11 : RAMB16_S1_S1
generic map (
INIT_00 => X"042200000000000041088001001AA00000000000000000000000500802000003",
INIT_01 => X"040048000024000000000404000000000A22000800000800004A200000000001",
INIT_02 => X"200C8840085EB00480060000001C008002489E0F000405EA0004040404000000",
INIT_03 => X"24004000000000000000000900002C4050000000000069500208400002E14100",
INIT_04 => X"4800200C0000000044002000C80020E40000E200000130200188000000800100",
INIT_05 => X"000000000080181000000000701000004C8000000058800000B1000009880480",
INIT_06 => X"80500081081040000000002C100040400000004641C080380400070100000000",
INIT_07 => X"4020109801A4CE005C00048380142810010564C4100114012002402028044808",
INIT_08 => X"0070700000000000000083004C3902420062000020E0000100004082A140102B",
INIT_09 => X"001150200000000000000026400000016186100000000010C04002C000000000",
INIT_0A => X"007C00008082C0002000000000002C3000000004050001030102040000000000",
INIT_0B => X"0000000000000000000000000000010000800011000000000000000000000BC0",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"000000000000000000000000000000042000760000000000000000010004B200",
INIT_0E => X"0D74002280300F0002FB069040000060000C5003000800000000000000000000",
INIT_0F => X"C01AE8004500744C780687DBA828008080A5FC0D385598035D0008A00C015660",
INIT_10 => X"39D8140040201BF861F0E7D693E6170022408116DFE0AB3006BA0011401D02AC",
INIT_11 => X"5412E4997F5249FD005043B8680CC98F00D0F2DD0140100406FE053A98F6ECC7",
INIT_12 => X"7418663001858040E153888000010840E165D0000000285C246A181C03FE4662",
INIT_13 => X"8199830066F0020858385974000001260208583854E2200000660208D6B1423F",
INIT_14 => X"8235AC508FCE8811042040F008235AE04420C040CF00C031C80009B8F224978B",
INIT_15 => X"030004E00000C220010808C10D9A92A74CD7CF4A09051110AD5A3C9200B7F280",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000118",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"07208BBA3F0C7010C660C7441920000000000000000000000000000000000000",
INIT_1A => X"861869A61861861861869A61861861861861861861861861A8208C4C1534D34C",
INIT_1B => X"984C26130984C26130984C26130984C26130984D26930984C26130984C261861",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000984C26130984C26130",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"174BA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFDFEF5D2A974BA082E95400F7FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0004",
INIT_29 => X"FFFFFFFFFFFFFFFFF7FBFDFFF552E974BAA2FFFFE10087FFFFFFFFFFFFFFFFFF",
INIT_2A => X"004001EFAAAEA8ABA087FFFFFFFFFFFFFEFF7FBEAB450804001EFAAD57FEAAF7",
INIT_2B => X"FFFBFDF45AAD568B55080028B55002E82000F7FFFFFFFFFFFFDFEFA2D568B550",
INIT_2C => X"0007FC00AAF7FFFFFFFF7FBE8B55AAD16ABEF5D2ABFF55080402010087FFFFFF",
INIT_2D => X"55A2FFFDFEF5D2EBFE00AAFFFFEBA087FFFFEFF7D168B55AAD17FFFF552EBFE0",
INIT_2E => X"000AAFFFDF45A2D16AB55F7FFFFFFF00043DE10AA843DE00557FFDFEFA2D16AB",
INIT_2F => X"FFEF552A974AA0000104AA000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFF7FBFDFFF5D2A954AA082A92428E3FFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"0071EFB6DF7AE92EBFFFFFFFFFFFFDFEFF7F5FAFC7492A974AAB6F5F8E101C7F",
INIT_32 => X"F1F8FD7AAD16AB450000001FFBEA4A8AAA147FFFFFFFFFBFDFC7EBF5E8B55000",
INIT_33 => X"00000010087FFDFC7E3F1FAF55A2DF6DB7D1C002AB7D002A82028FFFFFFFEFF7",
INIT_34 => X"BEDB7FFEF552AB8E38087FC2092F7FBF8FC7E3F5EAB45B6DF6FBEF5D2AB8F7D0",
INIT_35 => X"84971F8FC7AAD56DB6DBEF5F8FD7412ABFE28B6F5F8E820871F8FC7E3D56AB6D",
INIT_36 => X"00000000000000000000B6F1F8F55AADF6DB7DE3F5FAFC708003DE28B68E38E2",
INIT_37 => X"FFFFFFFFFFFFFFFFFDFEF552E954AA0004000AA0000000000000000000000000",
INIT_38 => X"54AAF7D568A00557FFFFFFFFFFFDFEFF7FBFFFEF552E974AA082A820AAA2FFFF",
INIT_39 => X"FFF55A2D16AB550000175EFFFFBEAA00A2FFFFFFFF7FBFDFFFFFD568B55002A9",
INIT_3A => X"A800AAF7FBFDFEFF7D56AB45AAD56AB450004001EFFF842AAAA557FFDFEFF7FB",
INIT_3B => X"FFFFFFF552AA8BEF080402000087BFDF45AAD568B55AAFBFDFEF55042ABEF002",
INIT_3C => X"8516AB55A2D16ABEFFFFBFDFFF552AAAAAA007BC0000FFFBE8B55AAD168B55F7",
INIT_3D => X"00043DEAAFFAEAAAAA08556AB55A2D57FFFFF7D568B45002ABDEAAFFD16AA000",
INIT_3E => X"0000000000000000000000000000000000000FFD56AB45A2FFFDFFFAAD16AB45",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(2),               -- Port A write enable input
DIA(0)   => data_write_a(19),        -- Port A data input
DOA(0)   => data_read_a_hi_512(19),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(2),               -- Port B write enable input
DIB(0)   => data_write_b(19),        -- Port B data input
DOB(0)   => data_read_b_hi_512(19),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_20_11 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000003",
INIT_01 => X"F55FF80000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"E05022020800008400F655001FFCFF80018FA804400000000000004400000001",
INIT_03 => X"00000000000000000000000900002CC07000000000000000000000000000013F",
INIT_04 => X"68002FFE40900010000180000001FFEC0012EE0C001370F40780000000000000",
INIT_05 => X"0840000880FCBBF0100E204DF0F88311DD8005080679800000F3000029980580",
INIT_06 => X"001000030817C8E8840155FDF9001001050023F6C3C3D0F87FA19F7F011000E4",
INIT_07 => X"000000090492260800008000EE00000000000000002101FF2002C00000004018",
INIT_08 => X"2A040001071004000013FF7FCA302C0C0008214800002101554031F800000000",
INIT_09 => X"801F57F200000090000489FEC0000001EFBEF0040008023FDFC0000000004006",
INIT_0A => X"0000000008000000000000000000ADF000000200000008000008028300110230",
INIT_0B => X"0000000000000800080000000000000000000000000000000800800A40000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"000000040900005C848538000020000000800000080000020000800101FFB600",
INIT_0E => X"00800000003A010003000000000000600FFC53FF001800000002004080000000",
INIT_0F => X"0001000000007408040000004000000004E9000008020000200000000E800800",
INIT_10 => X"00200000000313100010002000008000000000129600040000400000001D0010",
INIT_11 => X"81C012060000000000218F7840000100800004000000000066C0000080080000",
INIT_12 => X"800000000017C000100000000001A800080000000001A8040000002840008185",
INIT_13 => X"0000000006F00000100200000000012600001004000000000066000000801040",
INIT_14 => X"0000200410100000000005F00000020080090A0000000085C800002000586000",
INIT_15 => X"FF00400000000000020020020001000040283024E4F2860400008000030ED080",
INIT_16 => X"00000000000000000000000000000004010201001003020200000000000127DB",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"A0700030038200010089120104D2040020000000000000000000000000000000",
INIT_1A => X"2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2C30C30C30C30C306982121A1E79E79",
INIT_1B => X"32190C86432190C86432190C86432190C86432190C86432190C86432190CB2CB",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000432190C86432190C864",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0201000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF552A974AA0004174BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA0804",
INIT_29 => X"7FFFFFFFFFFFFFFFFFFFFFFEF552E954AA000400000F7FFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E954BA007FC00BA087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974BA082E9540000",
INIT_2B => X"FFFFFFFFFF7FBFDFFF552E974BAA2FFFFE10FFFFFFFFFFFFFFFFFFFFFBFDFFF5",
INIT_2C => X"FAAD57FEAA007FFFFFFFFFFFFFEFF7FBFFF550800020BAAAD56AAAAF7FFFFFFF",
INIT_2D => X"EFF7D56AB450000021EFA2D57DE10087FFFFFFFFFFFFFEFF7FBEAB450804001E",
INIT_2E => X"000F7FFFFFFFFFFFFDFEFA2D568B550004001EFAAAEA8ABA5D7FFFFFFFFFFFDF",
INIT_2F => X"FFFF5D2E954AA080005000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFEF552A974AA0000104AAFFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"A954AA082A92428087FFFFFFFFFFFFFFFFFFBFDFEF5D2E974AA000A07000E3FF",
INIT_32 => X"FFFFFEFF7FBFFFFF552E974AA0071C50BA1C7FFFFFFFFFFFFFFFF7FBFDFFF5D2",
INIT_33 => X"EDF6FABAEBFFFFFFFFFFFFDFEFF7F5FAFC7492A974AAB6F5F8E10E3FFFFFFFFF",
INIT_34 => X"EBF5E8B550000071EFB6DF7AE921C7FFFFFFFFFBFDFEFE3F5F8F450004050AAB",
INIT_35 => X"A497FFFFFFF7FBF8FC7EBD168B450804021FFB6D57DE28147FFFFFFFFFBFDFC7",
INIT_36 => X"00000000000000000000FFFFFFFEFF7F1F8FD7AAD16AB450000001FFBEA4A8AA",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2A954AA0800174100000000000000000000000000",
INIT_38 => X"74AA002E95410A2FFFFFFFFFFFFFFFFFFFFFDFEF552E954AA0004000AAFFFFFF",
INIT_39 => X"FDFEFF7FBFFFEF552E974AA082A820AA087FFFFFFFFFFFFFEFF7FBFDFFF5D2A9",
INIT_3A => X"568A00AAFFFFFFFFFFBFDFEFFFFFFDFEF5D2E954AA0051554BA557FFFFFFFFFF",
INIT_3B => X"D16AB450804174AAFFFFFFEBAA2FFFFFFFF7FBFDFFFFFD568B55002A954AAF7D",
INIT_3C => X"57FFDFEFF7FBFFF55A2D16AB550000175EFFFFBEAA005D7FFFFEFF7FBFDFFFAA",
INIT_3D => X"0004001EFFF842AAAA087BFDFEFF7FFEAB45A2D568B550804001EFF7D57DEBA5",
INIT_3E => X"0000000000000000000000000000000000000F7FBFDFEFF7D56AB45AAD56AB45",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(2),               -- Port A write enable input
DIA(0)   => data_write_a(20),        -- Port A data input
DOA(0)   => data_read_a_hi_512(20),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(2),               -- Port B write enable input
DIB(0)   => data_write_b(20),        -- Port B data input
DOB(0)   => data_read_b_hi_512(20),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_21_11 : RAMB16_S1_S1
generic map (
INIT_00 => X"4A302428B824900A128C090A5C1800261500213C005FE812D10420054085A202",
INIT_01 => X"001FFE3440B609703B0427F801A40B8115BC4F655300340288A40D30040E4DD8",
INIT_02 => X"E00424256888D8819801000F9FFFFFFFF149FF1FCA448046C60A0D2437C517F9",
INIT_03 => X"20030640003250640003250F06002CC1740002019824E001CD357832440001FF",
INIT_04 => X"EA2C3FFD400006E04401A8837001FFFC004AEF00080B70E08FB5789421007C5C",
INIT_05 => X"00011A0C40F9FFF80920954FF0F00809DF84A0202879800000F3000029980780",
INIT_06 => X"0805984B7A1FC0A0000101FFF0480080002281F7C3C381F87C03DFFF00009004",
INIT_07 => X"B424068086A205481A60A19000908204A855B000A08A61FF20C3D004D331D340",
INIT_08 => X"1BFA0001600802000023F7FFC08D234B40C2028253000040114200000D0226C0",
INIT_09 => X"EF1F5FF054096C6ADBA169FFC202B1C1FFBEF0440021083DFFCE22DC2880E24D",
INIT_0A => X"45FF0C004041D84862A28C54518DBFF00020004C0A6044901112A0908AA0A300",
INIT_0B => X"018C241102068006C620C03882019480E63180855A492712CC01C49C20201BFE",
INIT_0C => X"08A9464116544302C02D92236488D92236488D92236488D922366446C911B210",
INIT_0D => X"08800444021048034004001890000806002804A0822189000900D80621FFBE00",
INIT_0E => X"060580261013813A2CC396506102C4053FFD5BFF00A04A00200602CA52001100",
INIT_0F => X"080C0B004C202621A85C09411500135844C196D3606941018150098404C1A304",
INIT_10 => X"B02901013416181C96C2C9C600890A2028172192C460D1820302A0130809834A",
INIT_11 => X"9C5E803408250180AC268D185DB3F4350B811068C00049A0A4AA68F05C96A001",
INIT_12 => X"002C006560138F032B1804101244C883052208209040CC849063A747512B7678",
INIT_13 => X"41401E240665750440C9488280254530314080C2C601040420352148A00501B1",
INIT_14 => X"500811204D000700114204A70422016149916011008CAA8858850B00C32591C0",
INIT_15 => X"FFC06E60AC0496022300233104663040808E991765205000070121D41D18D098",
INIT_16 => X"40100401004010040100401004010040102090010008000001C0E010020007DF",
INIT_17 => X"0100401004010040100401004010040100401004010040100401004010040100",
INIT_18 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_19 => X"FFEF9FEEFF7FFDF7FF3E3DFDF7E0000000000000000000000000401004010040",
INIT_1A => X"BEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBFFDFDFFFCF3CF3F",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFEFF7FBFDFEFF7FBFDFEFBEF",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000FFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0001000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E954AA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0004",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA0004154BAFFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"52E974BA0804000AAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0004174BAFF",
INIT_2B => X"FFFFFFFFFFFFFFFFEF552E954AA000400000007FFFFFFFFFFFFFFFFFFFFFFEF5",
INIT_2C => X"A082E95400007FFFFFFFFFFFFFFFFFFFFDFEF5D2E974BA002E97400007FFFFFF",
INIT_2D => X"FFFFFBFDFEF5D2A954AA002E974BA087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFBFDFFF5D2E954BA007FC00BA5D7FFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA000002000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080005000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"A974AA0000104AAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974BA0000174AAFFFF",
INIT_32 => X"FFFFFFFFFFFFDFEF552E954BA080A000AAE3FFFFFFFFFFFFFFFFFFFFFFFEF552",
INIT_33 => X"02A95400087FFFFFFFFFFFFFFFFFFBFDFEF5D2E974AA000A07000007FFFFFFFF",
INIT_34 => X"F7FBFDFFF5D2A954AA082A924281C7FFFFFFFFFFFFFFFFFFBFDFEF5D2A974BA0",
INIT_35 => X"A557FFFFFFFFFFFFFFFF7FBFDFFF552E974BA0020924BA1C7FFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000E3FFFFFFFFFFFFFFEFF7FBFFFFF552E974AA0071C50B",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0000020000000000000000000000000000",
INIT_38 => X"74BA0000174BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954AA080017410FFFFFF",
INIT_39 => X"FFFFFFFFFFDFEF552E954AA0004000AAF7FFFFFFFFFFFFFFFFFFFFFFFEF552A9",
INIT_3A => X"E95410087FFFFFFFFFFFFFFFF7FBFDFEF5D2A954BA082E800AAA2FFFFFFFFFFF",
INIT_3B => X"FBFFFFF552E954BA002E97410087FFFFFFFFFFFFFEFF7FBFDFFF5D2A974AA002",
INIT_3C => X"57FFFFFFFFFFFDFEFF7FBFFFEF552E974AA082A820AA557FFFFFFFFFFFFFEFF7",
INIT_3D => X"5D2E954AA0051554BA5D7FFFFFFFFFBFDFEFF7FFFFFEF5D2A974BA0000020AA5",
INIT_3E => X"0000000000000000000000000000000000000AAFFFFFFFFFFBFDFEFFFFFFDFEF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(2),               -- Port A write enable input
DIA(0)   => data_write_a(21),        -- Port A data input
DOA(0)   => data_read_a_hi_512(21),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(2),               -- Port B write enable input
DIB(0)   => data_write_b(21),        -- Port B data input
DOB(0)   => data_read_b_hi_512(21),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_22_11 : RAMB16_S1_S1
generic map (
INIT_00 => X"5290F4CDE914905A14A43D33F488243E17122300F55FEB189B343A1140548380",
INIT_01 => X"A54007B259F6A975386262000C344BA9573C6FF57B18A5FB0ABFCD3C2C5F4F0C",
INIT_02 => X"021DFF8C38B3C009D203551040030071869D0040180AA2DC53DB89BEA8204001",
INIT_03 => X"2603475A969D0475A969D0460EAA401005111011BD506954EDB40F5EF41434C0",
INIT_04 => X"922D9002100ED69E443D988B0D5400103E48003D0800011E803B06B5B9125A15",
INIT_05 => X"281B5A0C06000408F4DF9422010D8802022F2124A8022492580040440002021C",
INIT_06 => X"F780C4C052881ADA0E05440205DA50930FA182010004700083E220800440B588",
INIT_07 => X"049D028B93FB561833D8094A02F5EA92FD7247E10305C40040D136E6A023F7FC",
INIT_08 => X"00028241680A0E002A9400803A884B5B5206B7C2E53CA25144009007A64EBD64",
INIT_09 => X"41008810240240C6694008010392354010000560141801002028A83D2A08E06D",
INIT_0A => X"34000000848BCA6902A29C54539C020E11810098D4067EFF9FF284D483E2AB41",
INIT_0B => X"500001840000C80B410014088040F4A944B1AA313C0022AA0011C0DC00028001",
INIT_0C => X"80B14004D158C8CA24A1C2A870AA1C2A870AA1C2A870AA1C2A872550E1543800",
INIT_0D => X"80A14050A01509E050854498B5281A1C34E506A2C6898B52A154DAC6B6000850",
INIT_0E => X"0B03001A483A4146603050080410089180008800143D83888281A2034A850142",
INIT_0F => X"A4160600349075238473F1210006133835E92273612B3482C090068A0E84AC56",
INIT_10 => X"30060181BA1B13959DC08DA902458870201970B29602562B0581200D141D0959",
INIT_11 => X"E042021C040D0152C8058B3840F044708E7E1C20A0106EA166C13AFC14AA3804",
INIT_12 => X"080E004B0C17C1439A9838301DC1A8438EA32C009DC1A8255300650458A1D588",
INIT_13 => X"018010E186F110A908E3A8CB0026C9A610A908E6A60F0807626610E160589C4C",
INIT_14 => X"2A701667334005800B1605F043858125E0D04110408D2485CA034681E43A1E40",
INIT_15 => X"00646002304244A91102C93A2D608D2A258DF8034188200C050171A41108F084",
INIT_16 => X"110441104411044110441104411044110466C440446CA06951D4EA8010009804",
INIT_17 => X"0040100401004411044110441104411044110441104411044110441104411044",
INIT_18 => X"0401004010040100401004010040100401004010040100401004010040100401",
INIT_19 => X"F7DFBFDEFE8FF1F7DEBDDF7DF7D05122890000000003FFFFFFFF900401004010",
INIT_1A => X"9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7BFFDFD7DDDF7DF7D",
INIT_1B => X"F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE79E7",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000003F9FCFE7F3F9FCFE7F3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA000400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0800",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000002000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2A954BA000015400FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080402010FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2A954BA0004154BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A0004174BAFFFFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0800154AAFFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF552A974AA0000174BAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974A",
INIT_2E => X"000007FFFFFFFFFFFFFFFFFFFFFFEF552E974BA0804000AAA2FFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080400010000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E954AA080005000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000402010FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2A954BA000417410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"804154BAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974BA0000174AAFFFFFFFFFFF",
INIT_34 => X"FFFFFFFEF552A974AA0000104AAE3FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0",
INIT_35 => X"AA2FFFFFFFFFFFFFFFFFFFFFFFEF552E954BA000E124BAE3FFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000007FFFFFFFFFFFFFFFFFFFFDFEF552E954BA080A000A",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804000100000000000000000000000000",
INIT_38 => X"54AA000400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2A954AA080017410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"0174BAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A954BA000415400FFFFFFFFFFFFF",
INIT_3B => X"FFFDFEF552E974AA0804174AAF7FFFFFFFFFFFFFFFFFFFFFFFEF552A974BA000",
INIT_3C => X"2FFFFFFFFFFFFFFFFFFFFFDFEF552E954AA0004000AAA2FFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2A954BA082E800AAAAFFFFFFFFFFFFFFFFFFFBFDFEF5D2E954BA002A820BAA",
INIT_3E => X"0000000000000000000000000000000000000087FFFFFFFFFFFFFFFF7FBFDFEF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(2),               -- Port A write enable input
DIA(0)   => data_write_a(22),        -- Port A data input
DOA(0)   => data_read_a_hi_512(22),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(2),               -- Port B write enable input
DIB(0)   => data_write_b(22),        -- Port B data input
DOB(0)   => data_read_b_hi_512(22),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_23_11 : RAMB16_S1_S1
generic map (
INIT_00 => X"EF20906D902424807BC8241BC81801B97D38AD3C0800103362A6741C80A12A02",
INIT_01 => X"001FFF8409F089003B4422000D80C80106804A7951C5B9D1C828043EA28838F9",
INIT_02 => X"E01CEE21649C82C40800000F9FFEFF8E72CA7F5FC2E22809925A0D3611C877F8",
INIT_03 => X"24000400402670400402670D48222DC1764446838624000080007460C40001BF",
INIT_04 => X"68403FFC020560E0443E21037C01FFFC0002EE00628BF0E02FAD781014085014",
INIT_05 => X"0112000202FBFFF00920017FF0F0628BFF8488890979800002F702002BB807A0",
INIT_06 => X"EF85788B681FC000000001FFF0010000000001F7CBC385F87C0BFFFF20040001",
INIT_07 => X"F6E200000000C1440E3AE408009120071070FA07A1CB23FFA403F0C4D23BF7C0",
INIT_08 => X"0BF87CA400804000003FF7FFD8880A034AC09662305AB10555421006891A1089",
INIT_09 => X"BE1F5FEA10092C0896A243FFC0008087FFBEF2000000001DFFC612C0C0400100",
INIT_0A => X"41FF0C2060501000600000000001BFFA800808189A657EF81DD0C00079CC8001",
INIT_0B => X"018C24110A860006C620C0312241C482B20400CC52492710CC80060020A81BFE",
INIT_0C => X"0C08866907048320C20C10030400C10030400C10030400C10030400608018210",
INIT_0D => X"040002000041500300100040000500C000801000C02400000952800001FFBF04",
INIT_0E => X"FC850015385380380CDB86106502C5043FFD5FFF00A04BC010A7724B10000800",
INIT_0F => X"89F90A002A70A710A51C01C05904014861433602A1CAF13F2110055614C72FC0",
INIT_10 => X"E02D02001C1E14981B43253EE50C8220180F1082E06397E07E42200AAC298E57",
INIT_11 => X"8421802400A90022B0070FAE18019214A380344920080B21A58B02AC60BACDF0",
INIT_12 => X"0A2A000C480B0704B54028101AC49C84BB4100009AC49C80857A82D20CE8CB22",
INIT_13 => X"01E00C8103416445C12ED0400027C5292445C12D500B0005A62D344CB241D095",
INIT_14 => X"132C907425604680038706A35132C94BDD011010404428886AC91B11311C8280",
INIT_15 => X"FF000470BE0692020328CA0028042054A92771C50FC070110001C1680809591D",
INIT_16 => X"00802008020080200802008020080200800800200200000000000008004807DF",
INIT_17 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_18 => X"8020080200802008020080200802008020080200802008020080200802008020",
INIT_19 => X"0000000000000000000000000000000000000000000000000000008020080200",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080002010FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974AA000400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000400010FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974AA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080000010FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E954AA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954A",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA000015400FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080002010FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974AA000400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000402010FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E954AA080005000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA080407000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA00041741",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080000010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000402010FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2A954AA080002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954AA080017410FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"552A954BA000415400F7FFFFFFFFFFFFFFFFFFFFFFFFF552A954BA080015410F",
INIT_3E => X"0000000000000000000000000000000000000F7FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(2),               -- Port A write enable input
DIA(0)   => data_write_a(23),        -- Port A data input
DOA(0)   => data_read_a_hi_512(23),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(2),               -- Port B write enable input
DIB(0)   => data_write_b(23),        -- Port B data input
DOB(0)   => data_read_b_hi_512(23),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_24_11 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100600007FFF000080108004000800020000840041000080808",
INIT_02 => X"FC5CA803400EB8209000000F9FFEFF8E7240FF1FC22409EA04018E50074017F0",
INIT_03 => X"11100400000000400000000D00002CC07400000090C080019001010A000001BF",
INIT_04 => X"68003FFC00040000000000008001FFFC0002EE00000370E007A100000000E468",
INIT_05 => X"0000000000F8BFF00920004DF0F00001DF8000000079800000F3000029980780",
INIT_06 => X"6E461803081FC000000001FFF0000000000001F7C3C380F87C019FFF00000000",
INIT_07 => X"600C2400013649609C8000980040814210254000A00B21FF2003F2A80D500000",
INIT_08 => X"0BF80000000000000003F7FFD88D2B4A02C0940062EC2804001610020408178B",
INIT_09 => X"8E1F5FE010092C0892A041FFC0000001FFBEF0000000001DFFC002C000000000",
INIT_0A => X"41FF0C0000000000600000000001BFFA0000005501AA00000CE2000009400000",
INIT_0B => X"018C0411020600048620C030020502000200000400490510CC00040020201BF4",
INIT_0C => X"0808064106040300C00C10030400C10030400C10030400C10030400608018210",
INIT_0D => X"0000000000004003000000000000001200580000000000000000000001FFBE00",
INIT_0E => X"0086C022005381380FDB96516140C6043FFD5BFF000041000000004110000000",
INIT_0F => X"80010D804400A7240C840C201D0210840043B4804012500021E0088014C04940",
INIT_10 => X"4109038041021C980200D06410C1924030008142E06024A00043C01100298092",
INIT_11 => X"587CC200002100C14428090A1D02348190814C09C010104025AA40041A0D8005",
INIT_12 => X"022E0030300B0E46177004208000D8C61D7004300000D884817B00011306B2D9",
INIT_13 => X"01E003060344710009875C018100013831000985DC000C20003C310006143B70",
INIT_14 => X"4001850EDC004780144806A64400186CBF8961104000C3807884000846EB9500",
INIT_15 => X"FF0006E08C063C0220002201490418082010A57263E0100008000290161E711C",
INIT_16 => X"00000000000000000000000000000000000000000000000000000000000007DF",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"F2D0AEEAF6E7CC1132CDB4441990000000000000000000000000000000000000",
INIT_1A => X"BEFBE79E79E79E79E79EFBEFBEFBEFBEFBEF9EF9EF9EF9EFA69861219575D75F",
INIT_1B => X"783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1EFBEF",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000783C1E0F0783C1E0F0",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0201000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A000400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA000400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000400000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402010000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"00002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080002010FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000400010FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA00040000",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020100000000000000000000000000",
INIT_38 => X"74BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"000010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA000002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974AA000402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000002010F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(3),               -- Port A write enable input
DIA(0)   => data_write_a(24),        -- Port A data input
DOA(0)   => data_read_a_hi_512(24),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(3),               -- Port B write enable input
DIB(0)   => data_write_b(24),        -- Port B data input
DOB(0)   => data_read_b_hi_512(24),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_25_11 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100200002000000080100004000000020000800041000080808",
INIT_02 => X"FC400086000000800000000F9FFEFF8E738FFF1FC204010000000111568DD7F8",
INIT_03 => X"00000400000000400000000D00002CC4740000008000000080000000000001BF",
INIT_04 => X"68003FFF64A564AC000000000001FFFE0082EF00010370E007A1000000004000",
INIT_05 => X"0A00040148F8BFF80920804DF0F00101DFC040000079C92484F30499299837C1",
INIT_06 => X"66041803081FC0E0801101FFFD000E41002299F7E3C380F87C019FFF81200096",
INIT_07 => X"000000080480AE00000080000000000000000000A00B21FF2003E00000000000",
INIT_08 => X"1BF80000400A02000003F7FFFA0008000200A0400008A0000014100200081000",
INIT_09 => X"8E1F5FFA53EFBCACB2E369FFE0010001FFBEF80C40630C7DFFEEBAF000800202",
INIT_0A => X"41FF0C0600000000600000000001BFFE00301000000000000CC020000140000C",
INIT_0B => X"01DCCC31222730A49620C030020100000200000400490D10EC00040220201BF4",
INIT_0C => X"0808064106240300C00C10030400C10030400C10030400C10030400608018210",
INIT_0D => X"0883044582114013412080000000000000000000000000000012800001FFBE00",
INIT_0E => X"00040020000180380FC386106140C6043FFD5BFF00A04B80608003CB120C1106",
INIT_0F => X"0000080040000200040400000100000000009480000240000100080000400900",
INIT_10 => X"0001000000000808000000240000020000000100006004800002001000008012",
INIT_11 => X"0001001808220000002004001900000080800008000000000022400000088000",
INIT_12 => X"0010000000000E00110000000000408009000000000040808063004000008200",
INIT_13 => X"6000000000046100000240000000001021000004400000000010210000001010",
INIT_14 => X"4000000404000800000000060400000088000001800000001084000000088000",
INIT_15 => X"FF800C608C041002000002000006100000002100000000180600000000100018",
INIT_16 => X"4110441104411044110441104411044510629041040D180400000010028047DF",
INIT_17 => X"1104411044110441104411044110441104411044110441104411044110441104",
INIT_18 => X"1044110441104411044110441104411044110441104411044110441104411044",
INIT_19 => X"FBA2894A196A8C5A2932EC15DA080800002FFFFFFFFFFFFFFFFFC11044110441",
INIT_1A => X"2492492492492492492410410410410410410492410492412000531215A69A6B",
INIT_1B => X"158AC562B158AC562B158AC562B158AC562B1588C46231188C46231188C49249",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000B158AC562B158AC562B",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080000010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000010FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08000000",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(3),               -- Port A write enable input
DIA(0)   => data_write_a(25),        -- Port A data input
DOA(0)   => data_read_a_hi_512(25),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(3),               -- Port B write enable input
DIB(0)   => data_write_b(25),        -- Port B data input
DOB(0)   => data_read_b_hi_512(25),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_26_11 : RAMB16_S1_S1
generic map (
INIT_00 => X"E9264EAB20190CA3BA4997AA9002AE9C001006B0778015CFA17E0811039879C7",
INIT_01 => X"2FFFF9BB1F773C7F9BB07DFFFDD863FC5FFF3FEFFBBF9FFB22FFFBC7B9F30686",
INIT_02 => X"E06CCC62052E708180F6FFBFFFFCFFFFF9C7FF7FC24332E642090000074037F6",
INIT_03 => X"428003739CD9863739CD9869FE2B7DEAF300029E4E300DFE69A6E644E6FF473F",
INIT_04 => X"7C2FEFFFF5BA124F003DD31EAFFFFFEE9FF7EE6F4C0770FFD7DC7CA53997B2B1",
INIT_05 => X"DFFB5421C1F8BBFAFDBFFACDF0FFCC05DDDBFF3690F9EDB7F5F7AFF639BD7DE3",
INIT_06 => X"EFD044ABC817C3E3A74667FDFFB6FF5727CC3BFEF7C3FAF87FF59F7FFBFEF69F",
INIT_07 => X"00003002132462052E708180EF060C18E5BEFB051225CDFF7002C4EEDE77F6E0",
INIT_08 => X"3FFF7D5000EC75088ED3FF7FC8790E46426CE06CB1F8E041051831FA3068D77E",
INIT_09 => X"C05FD7FF9BEFBDCEFBEE59FEF44F6603EFBEFAFCC2E35E7FDFD147CCF3F583FA",
INIT_0A => X"67FF1C7FBFADEB31E35768E8ED6BFDF3EB3EBF9DDBCE7FDC1DF8A760F3EACC02",
INIT_0B => X"5BDDCC3B336F7C548667D47B7737AF3FD62601EDC25B3533DCEB07F262213FFC",
INIT_0C => X"5F9A06E19F4D93A0EA0F78C35E30D78C35E30D78C35E30D78C35E986BC61AE31",
INIT_0D => X"5FD7AFEFDFFAF59B6FF28FE1D80D73D840607307DCFE1D80EF69A004DFFFF7FF",
INIT_0E => X"0004001F8041897B2FFFC6D86D70CE04FFFFF3FF1F5F5475BD7F72E4D75EBFAF",
INIT_0F => X"F60008003F008237B0040A00010003E020023E0201F45EC0010007E01047D17B",
INIT_10 => X"00010001DC0004C81003DE050A700200001DC0006863E8BD8002000FC0208FA2",
INIT_11 => X"2200E400002801E1A00004C21C0206F60081800800007B00010F02007EC09A0E",
INIT_12 => X"0880007E000807C7C1A612001E0015C7C19C22001E0015C59DFE82011A311AA0",
INIT_13 => X"00001BC00101F60409F0670840070809760409F06984800780097604067D0010",
INIT_14 => X"81019F40042100001F800203D81019EC085614000085C80023D81009CF008A74",
INIT_15 => X"FF802FFDFFAFD082003B032FB987E04021D481D4000819060801E0D00001231D",
INIT_16 => X"EBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEFFBFBFBFBBFCFBB0FFDFEFFEF2DFFFFFB",
INIT_17 => X"BFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAF",
INIT_18 => X"FAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFE",
INIT_19 => X"475B15BCF491E166CC8553F86EDB5C88646FFFFFFFFFFFFFFFFFEBFAFEBFAFEB",
INIT_1A => X"861861861861861861861861861861861861869A69A61861AFBD54D5F871C71D",
INIT_1B => X"984C26130984C26130984C26130984C26130984C26130984C26130984C261861",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000984C26130984C26130",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040201",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(3),               -- Port A write enable input
DIA(0)   => data_write_a(26),        -- Port A data input
DOA(0)   => data_read_a_hi_512(26),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(3),               -- Port B write enable input
DIB(0)   => data_write_b(26),        -- Port B data input
DOB(0)   => data_read_b_hi_512(26),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_27_11 : RAMB16_S1_S1
generic map (
INIT_00 => X"00080A40000A41248002029000050A088000008242A0004404480002000A1155",
INIT_01 => X"2FFFF1C11F781C129C107DFFFE0860941E81258CA2B71C2220EC1B86E1A00002",
INIT_02 => X"E1000000810000014400FF6FFFF0FFFFF8007F1FC21110005080200000221FF0",
INIT_03 => X"4080026318C18226318C1821302232EAE00002BE001115FE48620040840A863F",
INIT_04 => X"643D4FFC2530000F003D821C0BFFFF8E9EF79E6D440748FED70060842105B0B0",
INIT_05 => X"D6F39020D1F8A3FAFDBFBACDC8FDC405D1DB7F1490E5EDB7D5CBADB2385D79C3",
INIT_06 => X"6FE000A38007C3032646EFF1F0B6FF46A78C39F8E723F2E47FE59C7F9ADA2612",
INIT_07 => X"00002820000000810000014401060C180190310540118DFF1000C0849673F6C0",
INIT_08 => X"3FF779100062B12A8EC3F47FC80208808210880C00082050000110023068D030",
INIT_09 => X"005F07E09BFFBD07FBAC09F8E42922038F7DF8BEC2E39C5F1FD047CEF1B582D8",
INIT_0A => X"63FF5D5F9FADE911E81C09818109E1F16B16B71092CE7ED81CF403601228C402",
INIT_0B => X"1BFDCC39732F3554866AD57C37BEAF1C152201A4C05B7531D56B05B06A213FF8",
INIT_0C => X"5BCA06F18FC59380F00E34430D10C34430D10C34430D10C34430F0861A2186B5",
INIT_0D => X"5B56ADAB5FAAE58B2F628EA0C80FA3F04040510768EA0C80CC61A0044DFFC6EB",
INIT_0E => X"0004001D800188792CE79715710AE4047FFD23FF315D54358D593474955AB6AD",
INIT_0F => X"520008003B000297B0040200010003E020001F0201E44A400100076000579129",
INIT_10 => X"00010001DC00004A10035E0408300200001DC000086BC8948002000EC000AF22",
INIT_11 => X"02002400002801E1A00000C01E0202F60080800800007B00000782006EC0820A",
INIT_12 => X"0080007E000006A7C10602001E0001A7C10C02001E0001C18DE282010A311AA0",
INIT_13 => X"00001BC00000FE0401F04300400708007E0401F04180800780007E04047D0010",
INIT_14 => X"81011F40040100001F800002F81011EC080604000085C80001F810094F008034",
INIT_15 => X"FF800C6DDDAFD082001B03249887E04001D481D4000009020801E0D00001021F",
INIT_16 => X"AB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6BF1EBDABD8E270BF84A25C6ACB777E3",
INIT_17 => X"B6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6AD",
INIT_18 => X"6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADA",
INIT_19 => X"490E2168100481CA860402104A471688747FFFFFFFFFFFFFFFFFAB6ADAB6ADAB",
INIT_1A => X"000000000000000000000000000000000008200000000000200072F210000001",
INIT_1B => X"05028140A05028140A05028140A05028140A0500804020100804020100800000",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000A05028140A05028140A",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040201",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(3),               -- Port A write enable input
DIA(0)   => data_write_a(27),        -- Port A data input
DOA(0)   => data_read_a_hi_512(27),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(3),               -- Port B write enable input
DIB(0)   => data_write_b(27),        -- Port B data input
DOB(0)   => data_read_b_hi_512(27),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_28_11 : RAMB16_S1_S1
generic map (
INIT_00 => X"02200AA400180030808802A900002A08001280A08A801044104A1000001818C3",
INIT_01 => X"0AA00011460214428114180000882214413D0A71592A01D92213D28005210202",
INIT_02 => X"0451110A012100884000AA30200000000C100040104112101100008888200000",
INIT_03 => X"448000318C52A20318C52A20148810200111100C211004AA00034204200A2200",
INIT_04 => X"04004001001A90110000121402AA0000003C00000500000040080421080D0080",
INIT_05 => X"4060000C8001000000002E000000050000001610300000010000802202040012",
INIT_06 => X"1000002080001111001222000425A1040026A008000000000000000009328280",
INIT_07 => X"2491008A00491201210088400122448908A20402000408001000040820000000",
INIT_08 => X"20058310402A160026500000028040101004200C840082115554000112244814",
INIT_09 => X"4140000800000060000720000102028000000490160801020002200011100010",
INIT_0A => X"020000081B34211082B694D4D294000020020381040000000200032040004400",
INIT_0B => X"4800210C19808400500010009110091500020B408810000100200020408B0000",
INIT_0C => X"01028000080118020023604858121604858121604858121604858090B0242C00",
INIT_0D => X"010000800920040804020A6058003108402043058C460580653020005A004039",
INIT_0E => X"00000002800008014004104104420A00C000200005000010040A0020CC000200",
INIT_0F => X"520000000500000010000200000000000000280000040A40000000A000001029",
INIT_10 => X"00000000000000C0000002000830000000000000480008148000000140000020",
INIT_11 => X"020024000000000000000440000000020000800000000000000C00000040020A",
INIT_12 => X"00800000000001804006020000000500400C0200000005400A90000000100000",
INIT_13 => X"0000000000018200001003004000000142000010018080000001420000200000",
INIT_14 => X"8000080000010000000000018800008000060400000000000310000008000034",
INIT_15 => X"000002040080000000110006B081400000400000000009020000000000002200",
INIT_16 => X"802008020080200802008020080200802101210810C39A66A90A85420413A820",
INIT_17 => X"0200802008020080200802008020080200802008020080200802008020080200",
INIT_18 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_19 => X"DE21102C110A00246972BD89A40A0C22E1000000000000000000002008020080",
INIT_1A => X"2082082082082082082082082082082082082082082082080D35050758C30C31",
INIT_1B => X"0582C160B0582C160B0582C160B0582C160B0580C06030180C06030180C08208",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000B0582C160B0582C160B",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(3),               -- Port A write enable input
DIA(0)   => data_write_a(28),        -- Port A data input
DOA(0)   => data_read_a_hi_512(28),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(3),               -- Port B write enable input
DIB(0)   => data_write_b(28),        -- Port B data input
DOB(0)   => data_read_b_hi_512(28),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_29_11 : RAMB16_S1_S1
generic map (
INIT_00 => X"79964E4BA01DACAB9E659792D00AAE160002829C7FDFEFCEE97C2815039D70C3",
INIT_01 => X"0ABFF9AB0775343F9AB01DF80D5821FC0FFF3FEFD1AF9FF1207FFBC7B9720586",
INIT_02 => X"002CCC60050E700080F6AAA7BFFC007189C7FF2FC00330E602800000074037F6",
INIT_03 => X"468003210868A63210868A68DA017D207200021C4E200CAA6186A40042FF4300",
INIT_04 => X"7C2FE002F0900001003C5316A6ABFFE21F36E02F0D03701F47D41800109FB281",
INIT_05 => X"4979440580F9B808F49F6A4DF00F8D01DC4B97369078249370F482E62BA41462",
INIT_06 => X"B250442BC81001E1870223FC0BF7F11507C423FE33C078F803F19F00E936721D",
INIT_07 => X"00011080012460050E700080EF020408EC8CFA01122149FF700200665A35D260",
INIT_08 => X"2BFD055040A452000443FF00007906464068406C31F84000000831FA1028575A",
INIT_09 => X"805FD017102690AA694551FE30444681E0820AD40201423FC00122C493500172",
INIT_0A => X"0600002AFFBE2330815568A8AD6ABC02A02A0B0CCB463B4C0748A720B1EA4C00",
INIT_0B => X"0850400A11414C005005000B51158936D20601A98A10200308A002E240010BFC",
INIT_0C => X"05928020194918A22A2268C81A32068C81A32068C81A32068C81A99034640C00",
INIT_0D => X"058102C48970541944B20FA1580561D040406305587A158046282000DBFFF13D",
INIT_0E => X"000000028040890327DCD28928324400DFFFF0001F1F0050342D42A086040B02",
INIT_0F => X"F60000000500802010000A000000000000022A0000141EC0000000A01000507B",
INIT_10 => X"00000000000004C0000082010A700000000000006800283D80000001402000A0",
INIT_11 => X"2200E4000000000000000442040004020001800000000000010D000010401A0E",
INIT_12 => X"08800000000801C040A6120000001540409C2200000015441DAC800010100000",
INIT_13 => X"0000000001019600081027084000000956000810298480000009560002200000",
INIT_14 => X"800088000021000000000201D800088000561400000000002358000088000A74",
INIT_15 => X"00802594A282C0000033010FB181E00020400000000819060000000000002305",
INIT_16 => X"C0B02C0B02C0B02C0B02C0B02C0B02C4B12B312912831A27FCFE7FFB175B6FF8",
INIT_17 => X"0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02",
INIT_18 => X"B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C",
INIT_19 => X"BBCF9F96EE7FFDF7FE783FFDFFEA0C00602FFFFFFFFFFFFFFFFFC0B02C0B02C0",
INIT_1A => X"EFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEEBAEBAEBAEBAEBBFFDF9FBEFFFFFFE",
INIT_1B => X"BFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFBEFB",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000FBFDFEFF7FBFDFEFF7F",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(3),               -- Port A write enable input
DIA(0)   => data_write_a(29),        -- Port A data input
DOA(0)   => data_read_a_hi_512(29),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(3),               -- Port B write enable input
DIB(0)   => data_write_b(29),        -- Port B data input
DOB(0)   => data_read_b_hi_512(29),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_30_11 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"F7FFBFFEFF9FE1F7FFBFFFFDFFD0000000000000000000000000000000000000",
INIT_1A => X"9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7AFBD75F5FDF7DF7F",
INIT_1B => X"F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE79E7",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000003F9FCFE7F3F9FCFE7F3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(3),               -- Port A write enable input
DIA(0)   => data_write_a(30),        -- Port A data input
DOA(0)   => data_read_a_hi_512(30),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(3),               -- Port B write enable input
DIB(0)   => data_write_b(30),        -- Port B data input
DOB(0)   => data_read_b_hi_512(30),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_31_11 : RAMB16_S1_S1
generic map (
INIT_00 => X"129000008004A00804A40000400800020000000C005FEA005800200400050100",
INIT_01 => X"255FF18019700810180065FFFC0040801E80258CA2951C2200EC0906A0804140",
INIT_02 => X"E0000000000000011000550FDFF0FFFFF0007F1FC200000044000000000817F0",
INIT_03 => X"0000024210A30024210A3001002220C06044469200040154482000408400043F",
INIT_04 => X"602D0FFC2420000E003D80080955FF8E1ECA8E2D400340FE870060842100B030",
INIT_05 => X"0213100040F8A3F8FDBF944DC0FDC001D1CB6904A061EDB6D4C30490281831C1",
INIT_06 => X"6FC000830007C202060445F1F0D25E4207A099F0E303F0E07FE19C7F80402412",
INIT_07 => X"0000200000000000000001100004081001103107000185FF0000C0849673F6C0",
INIT_08 => X"1BF27A00000000000883F47FC800080002008000000820440000100220489020",
INIT_09 => X"011F07E013EFBC06FBA009F8E00120038F3CF82C44630C5D1FC002CCE0808248",
INIT_0A => X"61FF0C06C48BC801600000000001A1F00110101092CE7ED81CF0004012288000",
INIT_0B => X"11DCCC31222730048620C4382204A608142002A440492530C401049020221BF8",
INIT_0C => X"0888066187448380E00C10030400C10030400C10030400C10030600608018210",
INIT_0D => X"080204010200418301208480800D02D00040100240A808008840800405FF8640",
INIT_0E => X"0004001D000180780CE386106100C4043FFD03FF101D40008001304018081004",
INIT_0F => X"000008003A000217A0040000010003E02000160201E040000100074000478100",
INIT_10 => X"00010001DC00000810035C0400000200001DC0000063C0800002000E80008F02",
INIT_11 => X"00000000002801E1A00000801C0202F40080000800007B00000302006E808000",
INIT_12 => X"0000007E00000607810000001E000087810000001E000081846282010A211AA0",
INIT_13 => X"00001BC00000740401E0400000070800340401E04000000780003404045D0010",
INIT_14 => X"01011740040000001F8000025010116C080000000085C80000C8100947008000",
INIT_15 => X"FF800C609C06D082000A03200806A040019481D4000000000801E0D00001001D",
INIT_16 => X"010040100401004010040100401004010060C040040C200950402090128057C3",
INIT_17 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_18 => X"0040100401004010040100401004010040100401004010040100401004010040",
INIT_19 => X"00000000000000000000000000001000802FFFFFFFFFFFFFFFFF810040100401",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(3),               -- Port A write enable input
DIA(0)   => data_write_a(31),        -- Port A data input
DOA(0)   => data_read_a_hi_512(31),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(3),               -- Port B write enable input
DIB(0)   => data_write_b(31),        -- Port B data input
DOB(0)   => data_read_b_hi_512(31),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_0_10 : RAMB16_S1_S1
generic map (
INIT_00 => X"ED39BA795990D275FB4A6E96ACC4731DEA4598B0AFB54867F6EE4618C3749803",
INIT_01 => X"8AA0047D8607944AC7DA180001ECA2444042106208408208C20022E9173734B3",
INIT_02 => X"1A7DDD79F9A73E6CCA7DAAF00001000008478020113D98E382FEDF333027C80F",
INIT_03 => X"75D341110C58F31110C58F32A208921F8051500147A0E4AB3493FB3A01EBE240",
INIT_04 => X"86424001531009B100425A97B2AA0001E03501D0A39C8F0078420001106D0C4C",
INIT_05 => X"BCC8CA2EBF03400700402BB20F00239E20341699198600000B08694B16434804",
INIT_06 => X"103FB860B2800161F8432200012DA185F80F24081C3C0707800E600056881308",
INIT_07 => X"B24197ABCDA467F9A73E6CCAFDC3870EEEEC44E2BDFE220094D03022210C011C",
INIT_08 => X"240581B5695EAA80262C080032BF07C7C1FC3F8E94F65B11555EAFFC1C306758",
INIT_09 => X"7E40000BEC004170040DB60017FED1CC0001045002984202003DB931192D60A5",
INIT_0A => X"120071411A74315881A28C141118000C5A85A60444210123820B43B40804674D",
INIT_0B => X"0820008E514045BB514F0106D1D8599581D3A958BC104A89215AC14C48898403",
INIT_0C => X"C261C01C48B1584A0CA3E2687A9A1E2687A9A1E2687A9A1E26870CD061343885",
INIT_0D => X"D274E93A758FA8683AC54B287522E10A74AF4AA59C568752662F5AC218000002",
INIT_0E => X"FF83C002783A0904231C70470C7E0B92800224008AE09FAD4BD48D1FC5D3A4E9",
INIT_0F => X"5BFF078004F075885DFBF7E15C06101C55E921F1F80FAB7FE0F0009E0E903EAD",
INIT_10 => X"F12E0380231F13978FF023FAFDBD9870380230F2D6081F56FFC1E0013C1D207D",
INIT_11 => X"DE7F263C0C8700125C0F8F3C43F1F10BBF7EFC61E01804E1E6C8F8FE807F67FB",
INIT_12 => X"02BE00017C17C1007E5E2E3081C5AC007E6F0E3081C5AC44418D65FE45DEE55B",
INIT_13 => X"61E0042786F103E9F01F9BC3C120C5A703E9F01F978B8C20666703E9F8A0FFED",
INIT_14 => X"FA7E283FFB414F80005F05F10FA7E283F78F6511C048278DCA174FF038FF15B4",
INIT_15 => X"0066A20B61692F293185D8D724E15D3FCC6B7C236FE0691B0700132C1F0EF880",
INIT_16 => X"3A4E93A4E93A4E93A4E93A4E93A4E93A4F942F92E9628540AD2A91442525A000",
INIT_17 => X"A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E9",
INIT_18 => X"4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93",
INIT_19 => X"55F3898E09B56C74DAB15D1CF13501AA495000000000000000003A4E93A4E93A",
INIT_1A => X"082082082082082082082082082082082082082082082082082084E41DC71C71",
INIT_1B => X"E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F82082",
INIT_1C => X"FFFFFFFFFFFFFFF94A5294A5294A5294A5294A52800003E1F0F87C3E1F0F87C3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"3060C183060C187FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"BDEBA0000000000000000000000000000000000000000000003060C183060C18",
INIT_28 => X"168ABA002E82145085155545F7AA975EFFFAABDE00FFAEBDFFF5D2EAAAAAF7AE",
INIT_29 => X"7FFFE10005542145557FD5545FF8000155087FC0155F7D168B55007BFDF45085",
INIT_2A => X"7FFC0010080017555555568AAAFFFFD7545AA8028A00A2802AABAFF8028BEF5D",
INIT_2B => X"FF842AABAA2AE95545FFD168ABAF7AEAAAAAA2FFFDF4500043FE105D2E954BAF",
INIT_2C => X"5007FD7400550415410002E974BA5D5168A00A2D142155005142010FFAE820AA",
INIT_2D => X"FFF780000BA007FE8AAAFF803FFFF5D2A821550000000BA007FD55FF5D7FC014",
INIT_2E => X"000AAFBEAA00007BFDFFF082EBDF455D5142000082E82145FFD17DFEFFFD168B",
INIT_2F => X"DFD75D2AA8A80EA8E2FE3F000000000000000000000000000000000000000000",
INIT_30 => X"68B551475FAF6D1C556F0AA1C24AABEA495FC716F002A975FFE3AA95E00EBAEB",
INIT_31 => X"42A0070071C50BAFEF1FAE0016D56A16D557BC257D415E0216FA3F1E8FC0145B",
INIT_32 => X"8010E004924874825D7FEAA85487FD24AFE3D02DAAAE12BD5545A2803AA00005",
INIT_33 => X"120155EA568E870BAEB8A05A2AEA8B50F55A2F150005A3A438BD04AFAB8F550A",
INIT_34 => X"545E055FFBE81D0BE8EA8A3AA05A2A5504001C74BA42A1571E8028E3DB7816D0",
INIT_35 => X"A5C7E3DFFFE90B45B47ABA497A82FFAFD2A82485FD2415A105C21451ED42A002",
INIT_36 => X"00000000000000000000B55EAAA100AA1D0F6F480B6A555A2A57A002A3D5FDB6",
INIT_37 => X"5EFAAAAB5E1AF3AABFF45592E88A0AFE80A8B0A0000000000000000000000000",
INIT_38 => X"65F520EBE9EF67D7BEA1FD5D556ABEF5D557FEBA55022A3F70C6B405F4D2AE97",
INIT_39 => X"C114728007521170821CE0FDE69411A8DED57CE1055555E5F58EFFC01FE2CACB",
INIT_3A => X"42341D5DEEBEF55080034E0A592A4AD0079C75D6070CC5CBB0280C029ABAA3EB",
INIT_3B => X"7F353AAF6C77F7F20D968BF57812A95E02A2AAB5EB0F280800EFAEE9F5D18F31",
INIT_3C => X"C91565455C141E41887D58AC448B69C30E02116220415A9540AA854140A0A204",
INIT_3D => X"DE6BE93172D7D625B556EEAB157ABEBE1B4D792A4AD1183454180DD3FDCAAAB7",
INIT_3E => X"F0000001FF0000001FF0000001FF0000001FF01EABC4B8014174FF7DA80F52FE",
INIT_3F => X"FF0000001FF0000001FF0000001FF0000001FF0000001FF0000001FF0000001F")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(0),               -- Port A write enable input
DIA(0)   => data_write_a(0),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(0),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(0),               -- Port B write enable input
DIB(0)   => data_write_b(0),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(0),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_1_10 : RAMB16_S1_S1
generic map (
INIT_00 => X"212C001411984004084D000508C53810A03D1450E839B003342114428A000803",
INIT_01 => X"00000019400B100A8196000000CC004400400002000000000000028001340000",
INIT_02 => X"052137AE8031800C0044009000000000061800001CD4019802AD04CCCFC20004",
INIT_03 => X"04514108C60C21008C6042108400000201440020505100000043C30E10E9F000",
INIT_04 => X"02104001011DEFE088805681920000008000004001900800004002108C280008",
INIT_05 => X"040002340105000200000000080001900010000108040000000008411600401C",
INIT_06 => X"1034001042800808201000000001000820020000102000040000000000800180",
INIT_07 => X"64BF81A15EDFDE8031800C00843060C19E030022103600000450020800040004",
INIT_08 => X"00008004691687AA840008000090248CC84E000046000311555521F183060AC5",
INIT_09 => X"0820800D08100171000DB000154440C800400500000852020011200201012021",
INIT_0A => X"02000040001000880A2A04445004000102002041000001008208001440004140",
INIT_0B => X"4820018A1140440078050040511000102000A008183000010002404400000000",
INIT_0C => X"1000C80008000C030030880C2A030A00C28030A80C2A030A00C28018D4061401",
INIT_0D => X"10040802050080200284401C0022880F009E08008205C0020118088018000000",
INIT_0E => X"0F03C00280000000420860C60C0C0B92C0000000004000010042000040102008",
INIT_0F => X"001E078005000108400005E11C0610000000288058000003C0F000A000100000",
INIT_10 => X"F10E0380000000C202300000008D187038000000480800000781E00140002000",
INIT_11 => X"806302380C870010000004400100110800007861E0180000000C400680000001",
INIT_12 => X"023E00000000018000580C308000050000610C30800005000215006800000101",
INIT_13 => X"61E0000000018100B0001843812000014100B00016030C20000141002880026D",
INIT_14 => X"400A20009B404F80000000018400A20044096111C04000000304026000501580",
INIT_15 => X"0046820040082300218450C2800010094000482141E060190700100000002200",
INIT_16 => X"020080200802008020080200802008020080008008600500A82A1100A8000000",
INIT_17 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_18 => X"0080200802008020080200802008020080200802008020080200802008020080",
INIT_19 => X"81328A46BABEFC54A0810C7452B4428A14000000000000000000020080200802",
INIT_1A => X"AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA28A28A28A28A2A8218D2C0C924925",
INIT_1B => X"E974BA5D2E974BA5D2E974BA5D2E974BA5D2E975BADD6EB75BADD6EB75BAAAAA",
INIT_1C => X"FFFFFFFFFFFFFFFD8C6318C6318C6318C6318C63000002E974BA5D2E974BA5D2",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"70E1C3870E1C387FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"5555500000000000000000000000000000000000000000000070E1C3870E1C38",
INIT_28 => X"EBDF455D2EAABEFF7FFE8BFF5D0002155557FFFFFF007FC21EFA2FFD74AAAAD5",
INIT_29 => X"AA95400552AAAABAFFD1574105D7FD75FFAAAA800AAF7AA974BAFFFBE8B45F7A",
INIT_2A => X"0517DF555D2EAAA1055000015500557DF45AAD1400BAA2AE801550051555EFF7",
INIT_2B => X"FFD540155557FD5400F78028BFFFFFBEAB55F780020AAAA80020AA082EAAB550",
INIT_2C => X"AFF842ABEF5D517DF55552A974AAF7AE820AA0851574BAA2D1574AA5D7BFDEBA",
INIT_2D => X"EFAAD1575EF557FFFE10557FFFFFFFFD56AAAAFFFFD7555AAD168B45AAAEAAAB",
INIT_2E => X"0005D7FFDF4500043FE105D2E954BAF7AE80010082A97410557FEABFFAAFBE8B",
INIT_2F => X"51C7A2FBD5490BFD1C056A000000000000000000000000000000000000000000",
INIT_30 => X"974BAF7FFEFB45FFAABDF55492AA8BC2EBDFEAF7F1F840017D4975D2FEF147FC",
INIT_31 => X"080BEF495FC71D54124924385FAAA8AAAE3D145410F7F1D55D71C002DABAEBAA",
INIT_32 => X"002D082082AB8B6DBEDB7DF7F540E2AE85028B40155145F7AF6DBED5450AA1C2",
INIT_33 => X"78E021FF1471FDEAAFFD56F16D5571D2E28E38E0216FA2D1E8E80140F45082B4",
INIT_34 => X"A2DA3FB7DAAD4AAAAF487BC70BFA97F7AF6D417E92482BF84020BA495557E3FF",
INIT_35 => X"55554ADBD7A2FFC7BEFF6FFD7FC7002FD74951D71EDFFABFD16FAAAE92BD5545",
INIT_36 => X"00000000000000000000547AB8F550A8010E00492487482FFFE82A85EBAE2FFC",
INIT_37 => X"1EF005162BEF047FD5545AAFBF7400FBF9424F70000000000000000000000000",
INIT_38 => X"714F8338AAAA1D0AE974AAF7FFFDF55F7AABFF55082CA8B4DF6C1E8F5E540002",
INIT_39 => X"EABEF75550ACBB7582225FF5843404547184164AA5D2EBEEB0A2D555410D3555",
INIT_3A => X"FEAAEB083BC1000FF8409000512AEABFFDF79DCBF755962010BDCBBC21455D7F",
INIT_3B => X"801F8BA0C57740BDAA0688E5405D57D412F7D55F5E50C7F401BAAE8403CF5A3F",
INIT_3C => X"5D16BABAA3EBC3157ABD5FFE55F2AA9FEAFDF7F431A9F7FFE81FF013A8001AFF",
INIT_3D => X"FB863550229BCABEB7DA403FFFDA2FBF7FED2C7F955445079E280A00C56145EF",
INIT_3E => X"0000000000000000000000000000000000000596EBEF55080034E0A592A4AD00",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(0),               -- Port A write enable input
DIA(0)   => data_write_a(1),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(1),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(0),               -- Port B write enable input
DIB(0)   => data_write_b(1),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(1),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_2_10 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10E006600180111284380310006289800480032283E000A34301002001A0817",
INIT_01 => X"0005A00810790848048044A54E404350404000720885800802000906E4910200",
INIT_02 => X"407004208400408044C600C50AA055254010541A110222841200000002402544",
INIT_03 => X"0600011004182401004102408C28414043101000408118000145840440F5C415",
INIT_04 => X"5035855703A2900A000CD3088400F40688C9844409060850925E58A4081A0221",
INIT_05 => X"0200840D1021A15AC50494894850890540D1E12020C6E510818500440A280090",
INIT_06 => X"113044094002801020440090A8011A1224AB9380552102442884882A20004097",
INIT_07 => X"000100880004428400408044860000008C022402102100AA40004404B5075460",
INIT_08 => X"15C23440408C862A2A12382A8A5244145048C06085008010141521F000001240",
INIT_09 => X"400582B9033AA0E7AA4110B0506744810554542450694E710A836188C2C00222",
INIT_0A => X"443518360012C2210B020414109130A28038188096A06B8C120CA440A9C00802",
INIT_0B => X"1345E53300EC68005605002964AF222A5704004D080211121C80024200821780",
INIT_0C => X"181080C1110C882202211488452213C88472213C88472213488441109A442231",
INIT_0D => X"008204440210091341208041000810C00000300220201800A908000038AD0284",
INIT_0E => X"00040002804180300E88D28D206A40000554815500481440300000C44A081100",
INIT_0F => X"000008000500828700000000010000000002380000A00000010000A010050000",
INIT_10 => X"00010000000004CA000214000000020000000000684280000002000140200500",
INIT_11 => X"000000000020000000000442100002840000000800000000010C000026000000",
INIT_12 => X"00000000000805A4800000000000152300000000000015801272000100210020",
INIT_13 => X"000000000101C00000C000000000000940000120000000000009600004050000",
INIT_14 => X"0000130000000000000002018000106000000000000000002380000141000000",
INIT_15 => X"55000190000000000002000280000000011080C0000000000000000000002310",
INIT_16 => X"40902409064190641906419024090244902A9003004800415120D4A190804241",
INIT_17 => X"0900409004090641906419064190240902409024090641906419064190240902",
INIT_18 => X"9044090040900409004190441904419044090040900409004190441904419044",
INIT_19 => X"75960040138D70C030B51C50C7D100A2052F81F81F83F03F03F0419044190441",
INIT_1A => X"0410410410410410410410410410410410410410410410410248602081659659",
INIT_1B => X"5128944A25128944A25128944A25128944A25128944A25128944A25128941041",
INIT_1C => X"FFFFFFFFFFFFFFFE1084210842108421084210843FFF825128944A25128944A2",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"7FD5FF555815607FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"2AA000000000000000000000000000000000000000000000007FD5FF55581560",
INIT_28 => X"FC21EFA2FFD75EFAA8415410AA8415555087BFFF55A2AA800BAFFAE954000800",
INIT_29 => X"84155EFA2AEBDEAAA2FBEAABA5D7FE8B555551421455D0002145552EBFEBA007",
INIT_2A => X"2AEBDF555D2E954BAA2AA974BAFFFFE8B45552EBDF45FFAEAABFFF7FFE8B55F7",
INIT_2B => X"AAAAAAAAAFFD1574105D7FFFF555D2AAAAAA5D2E820BAA2FBEAB5555557DF55A",
INIT_2C => X"50055575EFFF84021555D043DEAA5D04021EF557FC21FFAA8428BFFAAAA954AA",
INIT_2D => X"10085568A00FF80175FFA2D17DFEFF7800215500557DF55AA80001FFAA800015",
INIT_2E => X"0005D00020AAAA80020AA082EAAB5500517DF555D042AA10A284154005D00154",
INIT_2F => X"00AAFFAA9543A080038A2A000000000000000000000000000000000000000000",
INIT_30 => X"0017D5D20B8EAA007FC51C7A2FBD55D2BE800042AFE8E1557D0075D2F45BEAA8",
INIT_31 => X"AA8BC7EBDFEAFEFFD00105FFBC20BDEAAA2FBF8AAA557BE8B6D5D5FFABEF4904",
INIT_32 => X"FFEFB6D555578F7DB6A0BDF7D480E174BFA02A974BAF7F5EFB455D2ABDF55492",
INIT_33 => X"ED1FDE90E3A497492B6AAADAAAE3D155E105571D55D71C002DABA5524820BAB6",
INIT_34 => X"BE8F401D7B6A0001470155C51D0092A071555D5E3AE821D00001FF0871C016DB",
INIT_35 => X"5BE8555400550A38428007FED000E3DA3DFD5E3DFFFBD5A38A021551C5F7AF6D",
INIT_36 => X"00000000000000000000410F45082B4002D082082AB8B6D1C5B7DF7FF78E075C",
INIT_37 => X"5EF005560B55F7AA800AAF7AA954AA00042AAA20000000000000000000000000",
INIT_38 => X"ABEF057D68F5F5A00021EF55042AAAA007FD5555AAFBD7545FBB8020A3F7AE97",
INIT_39 => X"7DF55D7AABFF5428ACA8F45A6C1E8F5EFF84165EFF7802BAB0A2FFEAABA557BE",
INIT_3A => X"CA8AA80800020AAF7FBFFFEF04552ABFFFF841FFE75CA882108202E974AAF7D5",
INIT_3B => X"00151FF0C57401E5F3D1E00A1A884174A8FFAEBFEB0A2D55541051555694F002",
INIT_3C => X"2AA801455D7FE8BFFF680800FFF7AAA155F595542455512A975455D3AA8A0055",
INIT_3D => X"5D79FCAF774AE005BE7895554005D2A8A0B882FFFFE10AAAAAB755A66B6AF56A",
INIT_3E => X"00000000000000000000000000000000000000C3BC1000FF8409000512AEABFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(0),               -- Port A write enable input
DIA(0)   => data_write_a(2),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(2),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(0),               -- Port B write enable input
DIB(0)   => data_write_b(2),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(2),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_3_10 : RAMB16_S1_S1
generic map (
INIT_00 => X"210C00A20020000108430020001600B8156021104940741B3530400E02B92203",
INIT_01 => X"014C9BCA58B1296D24A402C992500B69404040028804A0080A000416A8D90A08",
INIT_02 => X"C12026A484318004404405C9C66E331352180D468B8203980300204442E02B34",
INIT_03 => X"04000748D60D24648D60524C88804D0215011020D15018148040C10A70E1D58C",
INIT_04 => X"18283333240FE41244187308C9104D70944852640901083801750EB0A418C220",
INIT_05 => X"0613142D01912CC2A1B4140528348900C612A104201C689044340ED413A07649",
INIT_06 => X"119000034019881822104C5E68035250A222829710A0A02C18C01A9920842413",
INIT_07 => X"402F00AB0016CA0431800444841020509D038B021230C1990001C644C8273200",
INIT_08 => X"16905000408482088290E8E64010248C4A5AA840C2000110001521F0810A92E7",
INIT_09 => X"0003CE6581BD016342A951AB146C4480530C3B2A8088D3542651670200C1826A",
INIT_0A => X"00735D36209A8A20020894004284B660821030C8990467401218004041020002",
INIT_0B => X"512445B740457154562F957CC08B00093700080D0A4851001D8302D20A0A1530",
INIT_0C => X"00508650008008021021A40861021840869021A408610218C0869810D6043095",
INIT_0D => X"1C8508438450801043A08090380A8834207007022209038080190000999C8F84",
INIT_0E => X"000400200000C0002A48A206204C4205F3304B33004C0041006240140A1C310A",
INIT_0F => X"0000080040000083800400000100000000008400018040000100080000510100",
INIT_10 => X"0001000000000800000244040000020000000100002A0080000200100000A702",
INIT_11 => X"000000000020000000200000080002C000800008000000000022000006808000",
INIT_12 => X"0000000000000A2281000000000040A3810000000000402001400000022002A0",
INIT_13 => X"000000000004200001C0400000000010200001C0400000000010000004490010",
INIT_14 => X"0001070004000000000000060000104C08000000000000001000000903008000",
INIT_15 => X"CC004050CA0C00020220200070040000010401C4000000000000000000100008",
INIT_16 => X"4310E4310A4210A4210A4210A4210A4210A8D0830A68010001B4DA881048061C",
INIT_17 => X"21084290A4210A4210A4210A4210A4210A4210A4210E4310E4310E4310E4310E",
INIT_18 => X"90A421084290A421084390E4310C4390E4310C4390E4310C4290A421084290A4",
INIT_19 => X"015303C0C78C706428A14C586291000A044001FFE000003FFC004290A4210842",
INIT_1A => X"2492492492492492492492492492492492410410410410412821600001249249",
INIT_1B => X"51A8D46A351A8D46A351A8D46A351A8D46A351A9D4EA753A9D4EA753A9D49249",
INIT_1C => X"FFFFFFFFFFFFFFFC00000000000000000000000038F56351A8D46A351A8D46A3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"55AB02055AB0207FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"420000000000000000000000000000000000000000000000007FFFAB57FFFAB5",
INIT_28 => X"A800BAFFAE9554508002AA00AA843DF55FFAA955EFA2D168B55557BEAA000055",
INIT_29 => X"002AB55AAAA955EF005568A00087BE8BFFA2D155410AA8415555087BFFF55A2A",
INIT_2A => X"AAABFF5508003FF555D0002145552ABFEBA007FC21EF007FD75FFAA841541008",
INIT_2B => X"082EBDEAAA2FBEAABA5D7FC0155005168B455D042AB45F7FFD741000042AA10A",
INIT_2C => X"FF7FBEAB55F7AABDEBA5D7FC2010A2D1575FFF7AA975555D2E80145F78415545",
INIT_2D => X"EF5555554AA087BC01FFFFAAAAB55552A954BAFFFFE8B55552EBDE00F7AEAABF",
INIT_2E => X"000082E820BAA2FBEAB5555557DF55A2AEBDF555D2E954BA002EAAABA002A821",
INIT_2F => X"FB7D5D7FEAA3808554203A000000000000000000000000000000000000000000",
INIT_30 => X"1557D1475FAF45BEAA800AAFFAA95578080038A2AA28E3AF55E3A0BA5D7AADB6",
INIT_31 => X"BD55D7BE80004AA1E8E2AB55B6A0925D7085F6AA10087FEABD7AAD57AEBAB68E",
INIT_32 => X"F5D0438140E2FA38B6AEBFF6D1D04AAFFA41040017D5D20B8EAA007FC51C7A2F",
INIT_33 => X"D0A901FFFF801557D1C20B8EAAA2FBE80AA557BE8B6D5D5FFABEF49002FB55FF",
INIT_34 => X"5D20BDE00EBAAA8BC7EBDFEAFEFAB8ABAE925D21C7010EADB525D7FFAE975C75",
INIT_35 => X"F002EADA921420871D74971D24820875C21D5EB8AA8FFF012A954BAFFF5EFB45",
INIT_36 => X"000000000000000000001C24820BAB6FFEFB6D555578F7DB6A0BDF7DEB8E125F",
INIT_37 => X"B55A28408145AAFFFFFFF5D7FEAABA0051400A20000000000000000000000000",
INIT_38 => X"AB55FAD568AA2AFAE975EF555168B55F7AA800BAF7AA955EF00042AAA2A2AEAA",
INIT_39 => X"2AAAA007FD55558A7BD7145FBB8020A35D2ABEF55F7800015F087FEAA00007FE",
INIT_3A => X"968F575D003FF55F7D5420BA5D2ABFEAAF7AE9DFF759A82AEF70800021EF5504",
INIT_3B => X"FFD5145FBAC9755F05040255FFD84175EF55002AAB0A2FFEAABA557BEA3EF057",
INIT_3C => X"82E974AAF7D57DF45552A3FF10AA8429F45A7D5EAF5FFBAEAAA10554155400AA",
INIT_3D => X"FF843FFE77C80825BC052ABFE10550415557085540000005156155FE90A8F5C0",
INIT_3E => X"00000000000000000000000000000000000005500020AAF7FBFFFEF04552ABFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(0),               -- Port A write enable input
DIA(0)   => data_write_a(3),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(3),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(0),               -- Port B write enable input
DIB(0)   => data_write_b(3),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(3),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_4_10 : RAMB16_S1_S1
generic map (
INIT_00 => X"A108400020612C80284210081034849800A00030300004833522C82D04A16002",
INIT_01 => X"2043998A1839284D1CA0650E1E504368403008418984014902030806A0D10200",
INIT_02 => X"C120042200000000044441CE01E80F00A49043118680008002000000026208E4",
INIT_03 => X"040001020019200020011209CC0164C060000000690111040144800042F5C403",
INIT_04 => X"7029AF0F81A00010CCA47700CC513CAC0D0B8E02010740E19754080108988021",
INIT_05 => X"02139405007133C0712244CD20F20105D583000020E9892201D304D42A9835E1",
INIT_06 => X"9190440300078002014405D9EE814C0284A883B6D7038AE079059B7800048092",
INIT_07 => X"000100AA0004408000000004840400008D200102503000782000C00C8025C000",
INIT_08 => X"00728A00408403220811991E02120C044058080004000001101121F220000260",
INIT_09 => X"811001E1185B38AD23C3707AD46440818F3CF80EC423CA7D01D123C80200816A",
INIT_0A => X"45810810A01B40216361056D6150F41200280001900439001FD8A00041400000",
INIT_0B => X"11FC88076266E800D605402962A820211500024808010512C40106D222223B14",
INIT_0C => X"0408804116040B02C02C500B0C02C100B0C02C100B0402C300B0401618058611",
INIT_0D => X"040200050200501301208482200D00D0A0408402C4282200A84800009B878680",
INIT_0E => X"00000020000100024AC88300300060090F0D830F00025400300204D018000804",
INIT_0F => X"8000000040000206A2000800000000000000950002E010000000080000588040",
INIT_10 => X"0000000000000808000554000200000000000100006D0020000000100000BB00",
INIT_11 => X"0000400000000000002000001A0002504001000000000000002280000D800800",
INIT_12 => X"0800000000000E2C802000000000408D801000000000408012440000200110A0",
INIT_13 => X"000000000004680003A0040000000010280003800800000000102800000B0000",
INIT_14 => X"000005C0002000000000000620000158000010000000000010A0000B00000200",
INIT_15 => X"C30146200400104002602600400000000294004000000004000000000010001A",
INIT_16 => X"0080200000008020000000802000000080080000004090014134DA101288C6DB",
INIT_17 => X"0802000000000401806010040180601004018060100000802000000080200000",
INIT_18 => X"8060180601004010040080200802000000000000802008020000000000008020",
INIT_19 => X"C0A28A063807E0500014063450404882846FFE000003FFC00000010040100401",
INIT_1A => X"AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA28A28A28A28A2934C8D0CCD145144",
INIT_1B => X"68341A0D068341A0D068341A0D068341A0D068351A8D46A351A8D46A351AAAAA",
INIT_1C => X"FFFFFFFFFFFFFFFC0000000000000000000000001FE32068341A0D068341A0D0",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"408102040810207FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"800AA00000000000000000000000000000000000000000000040810204081020",
INIT_28 => X"168B55557BEAB4500554200000557FE10FFFBEAA10007FD7410FFAA97555082A",
INIT_29 => X"55574105D2A800AA00043FEBA5D7FEAA00007BE8AAAAA843DF55FFAA955EFA2D",
INIT_2A => X"57BC00AAA2FFEAAAAAA8415555087BFFF55A2AA800BAFFAE9555508002AA0000",
INIT_2B => X"A2AA955EF005568A00087BE8BFFA2D17DE1000517FE10AAAAA8AAA002E975455",
INIT_2C => X"FAA8417410A2D140000F7FBC2010A2D157400AAAE974AAAAAA974BA08002AB55",
INIT_2D => X"EFA2AABDEAA087BEAAAAA2FBD54BA080002145552ABFEAA007FC21EF007FD75F",
INIT_2E => X"00055042AB45F7FFD741000042AA10AAAABFF5508003FF55F7D568A00552EA8B",
INIT_2F => X"5400F7A49057D0824850B8000000000000000000000000000000000000000000",
INIT_30 => X"3AF55F7A0925D7AADB6FB7D5D7FEAB7808554203A145178E00FFFBE8A101475D",
INIT_31 => X"A9557D080038AAA145157428492E8008200043FE925571EFA380871C7028A28E",
INIT_32 => X"AEA8A9200249056D4175C5092AAF5FDA38BE8E1557D1475FAF45BEAA800AAFFA",
INIT_33 => X"AA4954281C0E2FB55B6A0925D7085F6AA10087FEABD7AAD57AEBA08517DE00AA",
INIT_34 => X"007FC51C7007BD55D7BE80004AAFEDB42028EBFBC2028BED152438AAA092492A",
INIT_35 => X"AF7DF6AA00412EAABFFAA803DEBA0875EDA80BEF1C743840040017D5520B8EAA",
INIT_36 => X"0000000000000000000041002FB55FFF5D0438140E2FA38B6AEBFF6DBE84AAEB",
INIT_37 => X"A00FFFFEAA105D5155410FF84021EF0800154B20000000000000000000000000",
INIT_38 => X"DEBA0851574B2AAAEAAB55F78400145AAFFFFFEF5D7FEABFF0051400A25D5568",
INIT_39 => X"68B55F7AA800BAF7AA955EF00042AAA25555410BA082E8201000043FE005D517",
INIT_3A => X"568AA200557DE00AAAAAAA000804001FF005575408AA557FEB2FFAE975EF5551",
INIT_3B => X"D1550AAAA8002010F2AC154B25F2ABFF55F7800015F087FEAA00007FEAB55FAD",
INIT_3C => X"800021EF55042AAAA007FD5555087BD6145FAAC000A2A6FBC00BAAAFBC00BAF7",
INIT_3D => X"F7AEBDFF779A82AA43F7FBE8A00082EA8BFFAA843FEBA08517DE00F3F9574B30",
INIT_3E => X"000000000000000000000000000000000000008003FF55F7D5420BA5D2ABFEAA",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(0),               -- Port A write enable input
DIA(0)   => data_write_a(4),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(4),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(0),               -- Port B write enable input
DIB(0)   => data_write_b(4),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(4),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_5_10 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50DF4A0791B3FCB694379283C81FD996A091832102004A336A20E03C040C002",
INIT_01 => X"805FBDC69830A84D5C6A60000C34C26841280A00084000C8C212892EEAD53235",
INIT_02 => X"3B2026B578918E640A4F01CF8011FF0002080000082CA9998276DF7772C7C80D",
INIT_03 => X"37134108420D700084205702A4008A1D9100002171C0E0051554D93A11F5D140",
INIT_04 => X"8A41A0FC03A56DA000425A819410E3816C086198A388B702A8CA1210844A0C4C",
INIT_05 => X"B1808A062E8BC835F5E84532D708238A282F00A9291224800A2861490343082C",
INIT_06 => X"903FB8483A90581859050424100940825C6184401CDC451B860A6507160C4100",
INIT_07 => X"D26F068BCC96CDF8918E640E96D1A3469D6300E2FFEA27F8E4D23248130E259C",
INIT_08 => X"0BFA82E568442B2A082C0A7E3014250D49DA37A2420619000002AFF48D1222E5",
INIT_09 => X"3F005001E40969289429360416DCD1C46083030604B1CA20C03DF83B0A2C60A5",
INIT_0A => X"14613C71005A10492B888120288F480D58858449026145B3830F449449062B4F",
INIT_0B => X"11AC04934AC648BFD727C031E64170A137D5AA5C3E4B0F8A3C58C34C002290E3",
INIT_0C => X"CA29C6CC50384B6AC6AC86AB31AACA6AB39AAC86AB39AACA6AB3055643559C31",
INIT_0D => X"C673E33CF28F38603855401985228A0614BD30A0A2819852011E5AC2B87F9182",
INIT_0E => X"FF87C002F87A803E460B2516510CA594FF0044FFA4B08BAC4BB2CD0F09CF84E3",
INIT_0F => X"0DFF0F8005F0F5100DFFF5E15D06101C55EB29F1E00BE53FE1F000BE1E802F94",
INIT_10 => X"F12F0380231F17D78FC029FFF58D9A70380230F2FE0017C37FC3E0017C3D005F",
INIT_11 => X"FC7F023C0CA700125C0F8F7E43F1F001BFFE7C69E01804E1E7CCF8FC003FF5F1",
INIT_12 => X"023E00017C1FC1A4BFD82C3081C5BD27BFE30C3081C5BD00C02365D645CEEF5B",
INIT_13 => X"61E0042787F181E9C1EFD8CB8120C5AF41E9C18FD60F0C20666F41E9F009FFFD",
INIT_14 => X"7A7C077FFF404F80005F07F187A7D14BFFC96111C048278DEB074F9930FF9D80",
INIT_15 => X"C064014B8B652E2B3120C81284641D3E8DBF7D636FE860190700132C1F0EFB80",
INIT_16 => X"38CE1384E3384E338CE138CE1384E33C4E3ECE32E128882551349A1CBAA44103",
INIT_17 => X"84E3384E3384E3384E338CE138CE1384E3384E338CE138CE1384E3384E338CE1",
INIT_18 => X"CE138CE138CE138CE1384E3384E3384E3384E338CE138CE138CE138CE1384E33",
INIT_19 => X"F5E5BB4E7F7B9DB7FF3A1B6DB7E8410A8C000000000000000000384E3384E338",
INIT_1A => X"BEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEF9F7CFDFDDCF3CF3D",
INIT_1B => X"BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEFBEF",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000001711C7BBDDEEF77BBDDEEF77",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"FDFFF00000000000000000000000000000000000000000000080000000000000",
INIT_28 => X"FD7410FFAA97410082A800AAAAAE955450055421FFFFFBC0010AAD5574BA557F",
INIT_29 => X"7FD74000055574BA5D7FD7555A2D5575EF55517FF5500557FE10FFFBEAA10007",
INIT_2A => X"0002AABA5D2ABFFFFAA843DF55FFAA955EFA2D168B55557BEAB5500554200000",
INIT_2B => X"5D2A800AA00043FEBA5D7FEAA00007BC00AAAAAEBDF45A28428B45FFD168BFF0",
INIT_2C => X"5080028A00A2FFFDE00F7D57FEBAFF80174BAAAD1555EF555555555005557410",
INIT_2D => X"BA5D2E821FFA2D5554BA557BD75FFAA8415555087BFFF55A2AA800BAFFAE9555",
INIT_2E => X"00000517FE10AAAAA8AAA002E97545557BC00AAA2FFEAAAA082A97545F7D5420",
INIT_2F => X"7010BEDF524AA5571FDFEF000000000000000000000000000000000000000000",
INIT_30 => X"78E00EBFBE8A101475D5400F7A49043D0824850B8A2AE9756D145B401FFFFFFC",
INIT_31 => X"FEAB7D0855420BA1471D74380851524BA5571D757DB6D5525EF555178F6D1451",
INIT_32 => X"8A28B6DEBDF6DBEF1C0A28AAA5524BFFFFA28E3AF55F7A0925D7AADB6FB7D5D7",
INIT_33 => X"5555057D145152428492E8008200043FE925571EFA380871C7028B6AEBDF45B6",
INIT_34 => X"BEAA800AAFFAA9557D080038AAAA2FBF8E10EBD578EAAFF8415482BED1555EF5",
INIT_35 => X"81C209256DFFDF420BA552A821FFB6DF574A85575C55EFBE8E1557D1475FAF45",
INIT_36 => X"0000000000000000000008517DE00AAAEA8A9200249056D4175C50920875FDA3",
INIT_37 => X"5FF5D7BC21EFF7FBD7400F7FBC00BA55557DFF70000000000000000000000000",
INIT_38 => X"01FF5D5568BE7555568A00AAFFEAA105D5155410FF84020AA0800154B2AAAA97",
INIT_39 => X"00145AAFFFFFEF5D7FEABFF0051400A25551554BA0051400BA5551575EFF7D14",
INIT_3A => X"1574B2FFAABFF45FFAAAABFFAAFFFDFFF552EA8AAA55043DFF7AAAEAAB55F784",
INIT_3B => X"8002410FFD5575EF5555421E75555400BA082E8201000043FE005D517DEBA085",
INIT_3C => X"FAE975EF555168B55F7AA800BAF7AA955EF00002AAA2A2FBE8A00A2D16AAAAFF",
INIT_3D => X"0055554088A557FEB25D00021FFFFFFC00BA552A821EFFFFFD74BA5D51575F7F",
INIT_3E => X"000000000000000000000000000000000000000557DE00AAAAAAA000804001FF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(0),               -- Port A write enable input
DIA(0)   => data_write_a(5),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(5),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(0),               -- Port B write enable input
DIB(0)   => data_write_b(5),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(5),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_6_10 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10800B0061A01002840002C03002818000402322520070B313301C4389B2082",
INIT_01 => X"250041CA3839684D18A160000C52426841000000090800090210080008110200",
INIT_02 => X"0020042080010000044654C0000C008010000000001020900200200002620814",
INIT_03 => X"060881021088200021080200E4000A0891000020610111500104C00000F14400",
INIT_04 => X"0880000100000002000052288144004281C050400100280000C8100000080001",
INIT_05 => X"928080840001100A08009000280201000850E022401400002028214043410820",
INIT_06 => X"10100518090012122100C808049310002040000410A0001400000200120840D2",
INIT_07 => X"000100800004400001000000860408108C22000A502010074120044800040001",
INIT_08 => X"50000040D0C4E2088003FD01C01004044058082004000000000121F020408244",
INIT_09 => X"00BF17E9001205A5204911F814444080400100020000D200DFD16400C2A40AA0",
INIT_0A => X"04611C17849000022862A1596C8B5DF04834948900000100220C244840000880",
INIT_0B => X"03AD0413424E4044D665C070C22602291504400D084915020448114080201000",
INIT_0C => X"5E08864011088B22D22C008B0022C408B1022C208B0822C608B1111600458010",
INIT_0D => X"4251A12CD28A300429688001000800000020280204001000A00804309A002182",
INIT_0E => X"0000000280402400420800000000006200FC10002442042429324294014E8CA7",
INIT_0F => X"A40000000500800840000800000000000002280018001480000000A010100052",
INIT_10 => X"00000000000004C2003000010240000000000000680800290000000140202000",
INIT_11 => X"2000C0000000000000000442000001080001000000000000010C000280001804",
INIT_12 => X"08000000000801C300A010000000156000902000000015101200002800000000",
INIT_13 => X"000000000101800038002408000000094000386028040000000940000ED40000",
INIT_14 => X"0003B000002000000000020180002A24005010000000000023000060C7000A40",
INIT_15 => X"3F0280090321000040A410C28108000160008094000810040000000000002300",
INIT_16 => X"284A5284A728CA5284A528CA728CA52C4A5A0A32A300940101349A0408240818",
INIT_17 => X"9CA1294A329CA5284A728CA7284A5284A728CA5284A528CA728CA5284A728CA7",
INIT_18 => X"CA3294A129CA3294A129CA1294A329CA1294A3294A129CA3294A129CA3294A32",
INIT_19 => X"F5F78BCE7F8FF0F4FA955F7CF7F40A80145D55555556AAAAAAAAA94A329CA129",
INIT_1A => X"8E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E39B6CEDECDDF7DF7D",
INIT_1B => X"F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE38E3",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000001A1A33F9FCFE7F3F9FCFE7F3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"555FF00000000000000000000000000000000000000000000080000000000000",
INIT_28 => X"BC0010AAD5574BA557FFDFFF087BFDF45F7AA974AAAAAA97555F784174BAF7D5",
INIT_29 => X"515555508043FE00F7AA97555A2FBD7410AA8428AAAAAAE955450055421FFFFF",
INIT_2A => X"7D1575EFFFAA9555500557FE10FFFBEAA10007FD7410FFAA97400082A800AA08",
INIT_2B => X"0055574BA5D7FD7555A2D5575EF55517FF55A2AA97400552AAAB45082E80155F",
INIT_2C => X"500554200000003DE10FFD5401FFF7AAA8A10082EAAB45A2FFC2000007FD7400",
INIT_2D => X"10AA803FE105D516AABAFF843FFFFAA843DF55FFAA955EFA2D168B55557BEAB5",
INIT_2E => X"000AAAEBDF45A28428B45FFD168BFF00002AABA5D2ABFFFF087BD5545007BFDE",
INIT_2F => X"256DEB84104BAFFD1525FF000000000000000000000000000000000000000000",
INIT_30 => X"9756D145B401FFFFFFC7010BEDF524AA5571FDFEF1C7BFFF55FFA095482B6A49",
INIT_31 => X"4904380824850381C5B5057D1C003DE28F7A49057DAAF5D2428A2842AAAAA2AE",
INIT_32 => X"2AAFB451C2A8017DE3DF525FFFFA49756D145178E00EBFBE8A101475D5400F7A",
INIT_33 => X"2F1C50381471D74380851524BA5571D757DB6D5525EF555178F6DAAA49542841",
INIT_34 => X"AADB6FB7D5D7FEAB7D0855420BA1C0E3FE00E3DB471EFE3AAAAA00082EA8B6DA",
INIT_35 => X"F1C7BD057D1C71FFE10A28038E1049516AAB8FF8428FEFA28E3AF55F7A0925D7",
INIT_36 => X"00000000000000000000B6AEBDF45B68A28B6DEBDF6DBEF1C0A28AAA5524BFFF",
INIT_37 => X"F55F78017400F780001FFAA84000AAFFD1401E70000000000000000000000000",
INIT_38 => X"20BAAA8428AA2AAAA975FF5D7BC21EFF7FBD7400F7FBC00BA55557DFF7557BFD",
INIT_39 => X"EAA105D5155410FF84020AA0800154B2557FC01EF55043FEAAFF80021EFA2D14",
INIT_3A => X"568BE7AA80174AA082ABDF555D2A821EFAAFBC01FFF780155F7555568A00AAFF",
INIT_3B => X"AEA8A10082EA8BEFAAD5554B25551554BA0051400BA5551575EFF7D1401FF5D5",
INIT_3C => X"AAEAAB55F78400145AAFFFFFEF5D7FEABFF0051400A25D2EBFE10AAFFD55EFA2",
INIT_3D => X"552EA8AAA55043DFF7557BC01EF55557DE00AA842AA0000516AABAFF8428BE7A",
INIT_3E => X"0000000000000000000000000000000000000FFAABFF45FFAAAABFFAAFFFDFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(0),               -- Port A write enable input
DIA(0)   => data_write_a(6),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(6),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(0),               -- Port B write enable input
DIB(0)   => data_write_b(6),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(6),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_7_10 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10844B00482258A2842112C02450418800002300500030B313300C418992002",
INIT_01 => X"000009CA3839684D1CA0E0000E51424840000000080000080200080008510204",
INIT_02 => X"0120042086010000044600C00008000004100000000260900200000002402004",
INIT_03 => X"8628A10000082400000002408400080011000000610008000208C00000E14400",
INIT_04 => X"0911800100A000000000524084000040000050001140200100C8100000080102",
INIT_05 => X"0300812401011000000000002000114008008060441000000020024093000000",
INIT_06 => X"9190431C0D4010100000880804010010800000041080081000000200010424B2",
INIT_07 => X"000100AA0004408601000004860000008C02000A103010006928040800062481",
INIT_08 => X"84000048D484C20888000A0002120484C048007004000000000021F000000244",
INIT_09 => X"00A06009881201A520491004106C48A04040002400A15A208001650004001020",
INIT_0A => X"C99E1060201002044809C1040140A001004808810000459033189C0A400118A0",
INIT_0B => X"102000024040484050050041648A0041140C500B08821054C000264120000400",
INIT_0C => X"0404A083260E0832132011880462011880462051881462051881D31018C40620",
INIT_0D => X"0001000080001000813094801A8F80F00A600B52602801A88848011118003700",
INIT_0E => X"000003C007C002808228010410082042C000C000000004001002000400040002",
INIT_0F => X"A4000007800F80C840000800009864038A1200081C0014800000F001F0200052",
INIT_10 => X"00002C0E00E0E4004038000102400002C0E00E0D20100029000001E003E04000",
INIT_11 => X"2000C04031100E0403D0700300080908000100000661801E1900040380001804",
INIT_12 => X"0840878083E8003780A01043203A101780902043203A10082410082880000000",
INIT_13 => X"0601E0187900181035E0240806483248181035E0280410C8198818100DDD0000",
INIT_14 => X"0403774000201021E020FA006040376C00501022131210722060806D47000A40",
INIT_15 => X"00928A0002000110888600C032128201519480D40009902430160403E0E00506",
INIT_16 => X"01000000020080601802000000000405000A0020020081014134928820480010",
INIT_17 => X"0802018040000000006018020080200804010000000000806018020080000004",
INIT_18 => X"0000000001806008020000001006008020080001004008020080201004000020",
INIT_19 => X"0000000000000000000000000000400A004618618618C30C30C3000020180600",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000000B0840000000000000000000",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"1555500000000000000000000000000000000000000000000080000000000000",
INIT_28 => X"A97555F784174BAF7D5555FFF780155EFAAAEA8ABAAAFBFDE0055556AA005D04",
INIT_29 => X"55555EFAAFFFDFEFAAAAAAB455D556AA00FFAE95555087BFDF45F7AA974AAAAA",
INIT_2A => X"02EAAAAA082EA8A00AAAE955450055421FFFFFBC0010AAD5574BA557FFDFFF55",
INIT_2B => X"08043FE00F7AA97555A2FBD7410AA8428AAA557BFDFFF55003DFFFF7FBEAA000",
INIT_2C => X"0082A800AAF7AE975FFA28000010552EBDE00007BEAAAAA2D140000085155555",
INIT_2D => X"45087FEAB455D516AB55557BD55FF00557FE10FFFBEAA10007FD7410FFAA9740",
INIT_2E => X"000A2AA97400552AAAB45082E80155F7D1575EFFFAA955555D51574AAAAFFD55",
INIT_2F => X"AE105D556AA10410E17555000000000000000000000000000000000000000000",
INIT_30 => X"FFF55FFA095482B6A49256DEB84104BAFFD1525FFFF8E175C7A2AAAAA82A2F1F",
INIT_31 => X"F524AA5571FDFEF415B575D7AAF1FFFD7AAAAAFB7D495F6AA10E3AE905551C7B",
INIT_32 => X"003AFEFEBFBEAA001C2EA8A821C2EAAA00A2AE9756D145B401FFFFFFC7010BED",
INIT_33 => X"EDB470101C5B5057D1C003DE28F7A49057DAAF5D2428A2842AAAA497BFAFFF49",
INIT_34 => X"1475D5400F7A490438082485038F7A4905C7A28A070384120BDE100075EAA82B",
INIT_35 => X"D495150492BEF1D2555087BE8B7D555F6AB57417BC05D7145178E00EBFBE8A10",
INIT_36 => X"00000000000000000000AAA495428412AAFB451C2A8017DE3DF525FFFFA49756",
INIT_37 => X"555A2AEA8A10AAD568A00555168A10002E9754D0000000000000000000000000",
INIT_38 => X"8A10AAAE8215D557BFDF55F78017400F780001FFAA84000AAFFD1401E7FFAA97",
INIT_39 => X"C21EFF7FBD7400F7FBC00BA55557DFF7007BD5555AAD57DF55AAAEBDFEF007BE",
INIT_3A => X"428AA2007FE8BFF080028BFFAAFFEAA105D2EAAA005D2AAAA18AAAA975FF5D7B",
INIT_3B => X"043DE0000516AA10F7FBD7408557FC01EF55043FEAAFF80021EFA2D1420BAAA8",
INIT_3C => X"55568A00AAFFEAA105D5155410FF84020AA0800154B2FF8402145A2AA954AA00",
INIT_3D => X"AAFBC01FFF780155F7005140000FFD140145007FE8BEF557BEAB55087FC215D5",
INIT_3E => X"0000000000000000000000000000000000000AA80174AA082ABDF555D2A821EF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(0),               -- Port A write enable input
DIA(0)   => data_write_a(7),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(7),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(0),               -- Port B write enable input
DIB(0)   => data_write_b(7),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(7),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_8_10 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00000648E2840112C00000418000002700500030B3132000400812082",
INIT_01 => X"100008480009004C04A100000252024840000000180800080200010040110204",
INIT_02 => X"0020042000490000004600804008000005100000000024900200000002400004",
INIT_03 => X"0A0C33400008082400000080A4004B0891000020610112000040C00000E5C000",
INIT_04 => X"18800001000000000000512080000040800150400824280110C8100000120200",
INIT_05 => X"908084A10100100200004080280008240810802206940000012C214451610800",
INIT_06 => X"81B000080860109021400008040000202048020414A0021400040200322824C1",
INIT_07 => X"000000080004408049000004860000008402001A50208000630C040800062483",
INIT_08 => X"440000428644212280800A00021004044048002124000000000021F000000244",
INIT_09 => X"00004009001001010008100414644410400102228000D20080114502006409A2",
INIT_0A => X"000051312000042200294429148A4801C80C8C81000045907118040340020832",
INIT_0B => X"4020000240404140004D0544C4AA0001150410090302500011C813428A000400",
INIT_0C => X"46501090008820240240409000240009000240009000240009000120204808A5",
INIT_0D => X"42D1A168D09A301468402480004780F00140080860280004085904309A002196",
INIT_0E => X"00783FC00044340242280000000000020000C0000442106419120004034685A3",
INIT_0F => X"8000F07F800088A80000081EA2F9EC0000064004081010001E0FF00011104040",
INIT_10 => X"0ED0FC7E00000422201080000202658FC7E0000021882020003C1FE000222080",
INIT_11 => X"018059C3F350FE0C00000002A0040500000103961FE780000110010090000800",
INIT_12 => X"FD41FF80000830200021C1CF600012200010D1CF600012121600100810000004",
INIT_13 => X"9E1FE000010A1802100004343ED8000898021000087073D80008980200800002",
INIT_14 => X"0080200000BEB07FE00002086008020000209AEE3F300000246020200000620B",
INIT_15 => X"0088881903210000440610C8000A808040000208901786E4F0FE0C0000000166",
INIT_16 => X"685A1685A769DA368DA368DA769DA36CDA121A11A141800011309284002C0810",
INIT_17 => X"95A5685A1685A5695A368DA368DA769DA368DA368DA7695A1685A1685A5695A1",
INIT_18 => X"5A1695A568DA368DA369DA768DA1685A1695A5685A168DA369DA768DA368DA16",
INIT_19 => X"A4028A0A543EBC57A10A1E75D64108080468618618630C30C30C69DA5685A168",
INIT_1A => X"9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7BF3CCD8DF5B2DB2C",
INIT_1B => X"F87D3E1F4F87D3E1F4F87D3E1F4F87D3E1F4F87C3E1F0F87C3E1F0F87C3E79E7",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000006A6D4F87D3E1F4F87D3E1F4",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"155FF00000000000000000000000000000000000000000000080000000000000",
INIT_28 => X"BFDE0055556AA005D0415555080000000087BEAA10F7803DE00FFAEBFFFF0800",
INIT_29 => X"2AA8AAA557FC0010F780154105D7FC2145005155555F780155EFAAAEA8ABAAAF",
INIT_2A => X"7FFFFF55AA80155FF087BFDF45F7AA974AAAAAA97555F784174BAF7D5555FF55",
INIT_2B => X"AAFFFDFEFAAAAAAB455D556AA00FFAE95555AAFFE8A00552EBFE00F7D17FF45F",
INIT_2C => X"A557FFDFFF5504000AAAAAAA8B55F7D140010552E821EFAAAABDF555555555EF",
INIT_2D => X"55AA8028A00A2D57FF45557BE8A00AAAE955450055421FFFFFBC0010AAD5574B",
INIT_2E => X"000557BFDFFF55003DFFFF7FBEAA00002EAAAAA082EA8A00002AA8A10F784021",
INIT_2F => X"FE10F7AEBAFFF080A175D7000000000000000000000000000000000000000000",
INIT_30 => X"175C7A2AAAAA82A2F1FAE105D556AA10410E17555080E000280071E8A00EB8E3",
INIT_31 => X"4104BAFFD1525FF492EA8AAA5571C2000FF8A17400557FC015514555757DFF8E",
INIT_32 => X"2ABDE10EBDF7AF6DE3FFF8F7DB68A105D71C7BFFF55FFA095482B6A49256DEB8",
INIT_33 => X"AA0BDF6D415B575D7AAF1FFFD7AAAAAFB7D495F6AA10E3AE90555A2FBE8A3849",
INIT_34 => X"FFFFC7010BEDF524AA5571FDFEF550E00082B6A0AFB55F7D1420104124821D7A",
INIT_35 => X"01C2EA8A00F7800017DA2842FA00B6D578F6D557FFDA00A2AE9756D145B401FF",
INIT_36 => X"00000000000000000000497BFAFFF49003AFEFEBFBEAA001C2EA8A821C2EAAA0",
INIT_37 => X"0BA08556AA00AAAABFE00F7AEAABEF082E955450000000000000000000000000",
INIT_38 => X"21555D51575EFFFAA97555A2AEA8A10AAD568A00555168A10002E9754D082E82",
INIT_39 => X"17400F780001FFAA84000AAFFD1401E7082EAAABA5D5140010F7AE974105D7BC",
INIT_3A => X"E8215DA2FFE8ABA082ABFE00AAFBEABFFAAFBEABFFF7AA80145557BFDF55F780",
INIT_3B => X"D540000000402145AA843FFFF007BD5555AAD57DF55AAAEBDFEF007BE8A10AAA",
INIT_3C => X"AAA975FF5D7BC21EFF7FBD7400F7FBC00BA55557DFF75D2E82010F7843DF45FF",
INIT_3D => X"5D2EAAA005D2AAAA185D2AAAA10F780021FFA2803DE10FFD16ABFF5D7BFDE10A",
INIT_3E => X"0000000000000000000000000000000000000007FE8BFF080028BFFAAFFEAA10",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(1),               -- Port A write enable input
DIA(0)   => data_write_a(8),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(8),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(1),               -- Port B write enable input
DIB(0)   => data_write_b(8),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(8),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_9_10 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00018248A2840112C00002C18000002300500030B3132000400812006",
INIT_01 => X"400008000000004C0020000000100248413C0A61590001D90213C10008110204",
INIT_02 => X"01A0042080010000054600C04008000004100000001020900200200002420804",
INIT_03 => X"024003400008012400000010E4004B0891000020610310000144C00000F5C000",
INIT_04 => X"1801800100E000000000510084000040010050020810200000C8900000320200",
INIT_05 => X"918004311104100000000000200008100800002000100000002C234415610820",
INIT_06 => X"81B00008080010100000980804000008800042041080001000100200322C2481",
INIT_07 => X"0000811800044080010000058600000086020002502080006000040800062C80",
INIT_08 => X"0000004001D4618008800A00061004044048002004000000000061F000000244",
INIT_09 => X"000040090802009420409004104444084001022400214A2080014400026401A2",
INIT_0A => X"04000071200000A003CA294140200800C80C8C8100004590111C040040120800",
INIT_0B => X"12210002404848502847040164880021150400080222000200C8034200000000",
INIT_0C => X"4610088010080421021040841021000841021000841021000841010800420820",
INIT_0D => X"42D0A16C529A321068500484000500D10042080040284000084900001A002196",
INIT_0E => X"00000002804000004228010410082002C000C0002400046419120410034285A1",
INIT_0F => X"A00000000500800800000800000000000002290008001080000000A010100042",
INIT_10 => X"00000000000004C2001000000240000000000000680800280000000140202000",
INIT_11 => X"0000C0000000000000000442020001000001000000000000010C800080000804",
INIT_12 => X"08000000000801A7802010000000152780102000000015000600000800000000",
INIT_13 => X"000000000101900011E0240000000009500011E0280000000009500004DD0000",
INIT_14 => X"000137400020000000000201C000136C00101000000000002340002947000240",
INIT_15 => X"0080881901210000000600C280028000419480D4000010040000000000002304",
INIT_16 => X"68DA368DA1685A1685A1685A1685A16C5A121A13A141950051309284A82C0010",
INIT_17 => X"85A1685A1685A1685A368DA368DA368DA368DA368DA368DA368DA368DA368DA3",
INIT_18 => X"5A1685A168DA368DA368DA368DA368DA368DA368DA3685A1685A1685A1685A16",
INIT_19 => X"0157344CCCF48DE68A895C38E2540A8010100000000000000000685A1685A168",
INIT_1A => X"14514514514514514514514514514514514D34D34D34D34D28E1004039248209",
INIT_1B => X"D268341A4D268341A0D069349A0D069349A0D068341A0D068341A0D068345145",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000014D490D069349A0D068341A4",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"EAABA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"03DE00FFAEBFFFF0800155FFAAFBE8B45002A974AAAA803DFFFAA843DF45FFFF",
INIT_29 => X"7BFDE00A2FBD7400F7FBFDFFFA2AEBDE00AAFBEAABA080000000087BEAA10F78",
INIT_2A => X"055401FFF7AEAAA10F780155EFAAAEA8ABAAAFBFDE0055556AA005D041555508",
INIT_2B => X"557FC0010F780154105D7FC2145005155555557BE8BEF007FFDEAAAAD1555EF0",
INIT_2C => X"AF7D5555FFF780154AA5D2AA8A10F7AA974AA082E80010A2AAAAA10552AA8AAA",
INIT_2D => X"BAF7D17FEBAA2AEBDF45002EAAABA087BFDF45F7AA974AAAAAA97555F784174B",
INIT_2E => X"000AAFFE8A00552EBFE00F7D17FF45F7FFFFF55AA80155FF080400145FFFBEAA",
INIT_2F => X"8FC7BE8A3DF7DF7F5E8A92000000000000000000000000000000000000000000",
INIT_30 => X"000280071E8A00EB8E3FE10F7AEBAFFF080A175D7BEF1E8B6D002090482B68E3",
INIT_31 => X"56AA10410E175550871FFE00A2FBD0400FFF5FDFC7B6A0BDE38B6F5E8A92080E",
INIT_32 => X"7BFAE82A2DB555C71C5B451D7FFAAA8A38FF8E175C7A2AAAAA82A2F1FAE105D5",
INIT_33 => X"2AEADA38492EA8AAA5571C2000FF8A17400557FC015514555757D5D71E8BEF14",
INIT_34 => X"B6A49256DEB84104BAFFD1525FFFF84174BA5D20AAA00E3AA904BA142A87010A",
INIT_35 => X"7000400155FFFBEDA82FFD57DEBAAAA0BFF7D0024ADA921C7BFFF55FFA095482",
INIT_36 => X"00000000000000000000A2FBE8A38492ABDE10EBDF7AF6DE3FFF8F7DB68A105D",
INIT_37 => X"BEF080402000F7AAA8B55FFAABDFEFF7D16AA000000000000000000000000000",
INIT_38 => X"FEAAFFD16AA00082E820BA08556AA00AAAABFE00F7AEAABEF082E95545F7D568",
INIT_39 => X"A8A10AAD568A00555168A10002E9754D00517DE00A2FFC2000F7D17FF55FF803",
INIT_3A => X"1575EF555568BEF5D7FE8A10AAFFD55555D7FD5555FFAAA8AAAFFAA97555A2AE",
INIT_3B => X"AE800AA552A97400A2AEBDEAA082EAAABA5D5140010F7AE974105D7BC21555D5",
INIT_3C => X"57BFDF55F78017400F780001FFAA84000AAFFD1401E7FF80174AA5D0028A00AA",
INIT_3D => X"AAFBEABFFF7AA80145080002145F7FBFFE00FFD17FEAAA2803DFEF08043FE005",
INIT_3E => X"0000000000000000000000000000000000000A2FFE8ABA082ABFE00AAFBEABFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(1),               -- Port A write enable input
DIA(0)   => data_write_a(9),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(9),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(1),               -- Port B write enable input
DIB(0)   => data_write_b(9),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(9),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_10_10 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00018248A2840112C00002C18000202300500030B3132000400992006",
INIT_01 => X"254008000000004C002000000010026840000000080000080200010008110204",
INIT_02 => X"0020042000010000004455800008000004100000000000900200000002400004",
INIT_03 => X"020001021089000021081000C400090011000000610001540104C00000F14400",
INIT_04 => X"0811800101A00002000050088554004200C840000000200080C8100000000001",
INIT_05 => X"030080001000100800009400200000000840E020201000000024024001200020",
INIT_06 => X"81B00008080012120004CC080492500280208004148000100000020020042493",
INIT_07 => X"0000000800044080010000048404081085020002502000006000040800062480",
INIT_08 => X"100202400084410808000A00021004044048000004000000000021F020408264",
INIT_09 => X"010040090002008420401004144440004040022484214A2080110108C2C00320",
INIT_0A => X"04004166A48A0001080000000000080080181881000045901118044040020800",
INIT_0B => X"1201000200484910000F0105602622291404020902005002018002400A022000",
INIT_0C => X"0440001011808020120004801120044800120004801120044800110002400884",
INIT_0D => X"008000440210100041308480800F82F00040180260A808008848000018002104",
INIT_0E => X"000000028040000002280104100820020000400020000440100204100A000100",
INIT_0F => X"040000000500800800000000000000000002280008000400000000A010100010",
INIT_10 => X"00000000000004C2001000010000000000000000680800010000000140202000",
INIT_11 => X"200000000000000000000442000001000000000000000000010C000080001000",
INIT_12 => X"00000000000801C0008000000000154000800000000015000410000800000000",
INIT_13 => X"0000000001019800180000080000000958001800000400000009580002800000",
INIT_14 => X"0000A0000000000000000201E0000A0000400000000000002360002080000800",
INIT_15 => X"0080881000000000000600C28102800060000000000800000000000000002306",
INIT_16 => X"401004010040100401004010040100441020D0030008840051309A90BA884010",
INIT_17 => X"0902409024090240900401004010040100401004010040100401004010040100",
INIT_18 => X"1004010040902409024090240902409024090240902409024090240902409024",
INIT_19 => X"F546890A940FE0D3971243555205428290100000000000000000401004010040",
INIT_1A => X"8A28A28A28A28A28A28A28A28A28A28A28A28A28A28A28A29554199854514514",
INIT_1B => X"2B95CAE532994CA6532995CAE572B94CA6532994CA6532994CA6532994CA28A2",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000002718E72B94CA6532994CA657",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"FDE1000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"03DFFFAA843DF45FFFFEAABA007FC2155F7D155545AA80001EFAAFBEAB45557F",
INIT_29 => X"042AB55FFD168B55AA8000010FFFBE8BFFF78402155AAFBE8B45002A974AAAA8",
INIT_2A => X"AD16AABA002ABDE10080000000087BEAA10F7803DE00FFAEBFFFF0800155FF00",
INIT_2B => X"A2FBD7400F7FBFDFFFA2AEBDE00AAFBEAABAA2FFD741055003DFEFF7AA801FFA",
INIT_2C => X"05D0415555007FD74105555555EFF7FBC0145F78028A00A2D142155087BFDE00",
INIT_2D => X"55AAD168ABA002A975FFF7AEBDEBAF780155EFAAAEA8ABAAAFBFDE0055556AA0",
INIT_2E => X"000557BE8BEF007FFDEAAAAD1555EF0055401FFF7AEAAA105D042ABFF5D556AB",
INIT_2F => X"71D7AAFBEFB455D71F8E00000000000000000000000000000000000000000000",
INIT_30 => X"E8B6D002090482B68E38FC7BE8A3DF7DF7F5E8A92007BC217DEBDB55555AA8E0",
INIT_31 => X"EBAFFF080A175D700042AB7DEBDB6DB55BE8E05000EBFFE8BC7E38E07145BEF1",
INIT_32 => X"0A3DFD7F7A4821D7A2D16FA82142EB8E00080E000280071E8A00EB8E3FE10F7A",
INIT_33 => X"ED1421450871FFE00A2FBD0400FFF5FDFC7B6A0BDE38B6F5E8A92B6FBD541049",
INIT_34 => X"A2F1FAE105D556AA10410E175550071D54104951555D7EBF5C5155E3842AA00B",
INIT_35 => X"8410E2ABD749516FB55BED16FA820820955EFE3AEBDEAAFF8E175C7A2AAAAA82",
INIT_36 => X"000000000000000000005D71E8BEF147BFAE82A2DB555C71C5B451D7FFAAA8A3",
INIT_37 => X"1EFA2FFD7545AAAE97555A2FBFDF455D556AA000000000000000000000000000",
INIT_38 => X"8B45AAAA95545F7D568BEF080402000F7AAA8B55FFAABDFEFF7D16AA00087FC0",
INIT_39 => X"6AA00AAAABFE00F7AEAABEF082E9554500042ABFFA2FFFFF45F7AE97400AAFFE",
INIT_3A => X"16AA00FFFBD5400082EBFF45F78400155A2D57FE00552EA8A00082E820BA0855",
INIT_3B => X"D557555A2802AA10FFD54214500517DE00A2FFC2000F7D17FF55FF803FEAAFFD",
INIT_3C => X"FAA97555A2AEA8A10AAD568A00555168A10002E9754D085155410085557555AA",
INIT_3D => X"5D7FD5555FFAAA8AAA002AAAB4508557DF55F7D17FE000804155FFAAAABDEAAF",
INIT_3E => X"0000000000000000000000000000000000000555568BEF5D7FE8A10AAFFD5555",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(1),               -- Port A write enable input
DIA(0)   => data_write_a(10),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(10),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(1),               -- Port B write enable input
DIB(0)   => data_write_b(10),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(10),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_11_10 : RAMB16_S1_S1
generic map (
INIT_00 => X"A101C4B05A0034CA2840712C2D001419000002300500030B31B20084EC992002",
INIT_01 => X"90000986B83028491800E0000C26426040000000080000088200080802512224",
INIT_02 => X"1A2004205E010640024D00800008000004100000040EC090820018003241A00C",
INIT_03 => X"28639100000C5C00000045C08400C8001100000061806A001618C03001E54400",
INIT_04 => X"1A800001000009A0804059A190000040400040008058220008C8100000120D4E",
INIT_05 => X"02000E81080250010000002022000058080400000E1200000020004401000004",
INIT_06 => X"819435143F20101010001008040800B8100102041088011100022200000024B2",
INIT_07 => X"90640D280884453E01064002944180008402001295BA100022E4340800062D82",
INIT_08 => X"400000093204802200280A0012160585C1D808D004000000000323F40C102244",
INIT_09 => X"380040098010001100009204107C5950400000220080C200800900020C006827",
INIT_0A => X"80007100004016EA080801010000080D00200081000045B0511D289940103399",
INIT_0B => X"002000024040410A000D0104408810C115D9C008050042400100D04E88000002",
INIT_0C => X"00655010009264201200C7B421ED0C7B421ED0C7B431ED087B43176843DA1085",
INIT_0D => X"0401020080400A10012494881A4F80F209500BB2602881A488485C1318002000",
INIT_0E => X"6619A540124814800228010410082022C00040002020090020220C9600040802",
INIT_0F => X"ACCC334A802491600C587949B6D0141B4CC600D5761B1599865A500490B86A56",
INIT_10 => X"BAC845542056A61686EC81E3A6CB68AA2C622C9A251C352B330CB4A0092170D8",
INIT_11 => X"BCCAD0B5A81536080CC6B21A21B1FC09CB0F1076D4A200B2AD4068F4101639B5",
INIT_12 => X"4D2CC281E31AA0103AB8D5514066380804B268A2E060901204112566F10AC418",
INIT_13 => X"D551443C47281002540B2C9AAAA8662A1152B202AE3554403028115AA88201A1",
INIT_14 => X"548A20A0492A2724A0621620402A020141F172FB182A32AB6845AB6200251BC9",
INIT_15 => X"00C00A000200074044E6801832728080D00A380B753952C4877E0104DDE4D124",
INIT_16 => X"0080200802008020080200802008020480080022020081010124988800400010",
INIT_17 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_18 => X"0000000000802008020080200802008020080200802008020080200802008020",
INIT_19 => X"55062608804180C0B10A42104201400204000000000000000000000000000000",
INIT_1A => X"00000000000000000000000000000000000820820820820801C4149470000000",
INIT_1B => X"0000000000000000040200000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000007E0F0000000000000100800",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"000AA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0001EFAAFBEAB45557FFDE10082ABDF5508557DF45002ABDFFFF7803DE10AA80",
INIT_29 => X"AEBFF45FFAEBFEAA002A801FFF7FFE8A10A28000000007FC2155F7D155545AA8",
INIT_2A => X"2AABFE10082ABFFEFAAFBE8B45002A974AAAA803DFFFAA843DF45FFFFEAABAA2",
INIT_2B => X"FFD168B55AA8000010FFFBE8BFFF78402155AAD155555A28428BFF002ABDE00A",
INIT_2C => X"F0800155FF00557FF45557FC2010002A80010A2842AAAA007BFFF4500042AB55",
INIT_2D => X"FF5D00154BAF7FBE8BEFFFD540000080000000087BEAA10F7803DE00FFAEBFFF",
INIT_2E => X"000A2FFD741055003DFEFF7AA801FFAAD16AABA002ABDE10A2D168A10A284021",
INIT_2F => X"DFC7F78E3FE28B684070AA000000000000000000000000000000000000000000",
INIT_30 => X"C217DEBDB55555AA8E071D7AAFBEFB455D71F8E00002EBDF6D005B78F7D142AB",
INIT_31 => X"A3DF7DF7F5E8A92BEAEBFF7DEBA0BDEAA1C2A801C7E3FFEFA10B68407038007B",
INIT_32 => X"8A28BFF082ABAE10B6AAB8E280820B8FEFBEF1E8B6D002090482B68E38FC7BE8",
INIT_33 => X"07FF8F7D00042AB7DEBDB6DB55BE8E05000EBFFE8BC7E38E07145B6D15756DA2",
INIT_34 => X"EB8E3FE10F7AEBAFFF080A175D708517DF7D497BC5028142A87000A28A2AA920",
INIT_35 => X"0B6DB6AA28A280001FF5D0A10482FFFFEFBC7E3DF42028080E000280071E8A00",
INIT_36 => X"00000000000000000000B6FBD5410490A3DFD7F7A4821D7A2D16FA82142EB8E0",
INIT_37 => X"FEF007BE8BFF5D2ABDF55F7AABDEAAF784154BA0000000000000000000000000",
INIT_38 => X"DE00FF84154BA087FC01EFA2FFD7545AAAE97555A2FBFDF455D556AA00082EBF",
INIT_39 => X"02000F7AAA8B55FFAABDFEFF7D16AA00FFAEBFFEFAA803DEBA5D2E82155A2FBF",
INIT_3A => X"A95545F7D5555FFAAAAA8BFF002AAAA00FFAAA8AAA080028BFFF7D568BEF0804",
INIT_3B => X"2E95400A2AEA8A00007FEABFF00042ABFFA2FFFFF45F7AE97400AAFFE8B45AAA",
INIT_3C => X"82E820BA08556AA00AAAABFE00F7AEAABEF082E9554508557DFFF007BD54BA5D",
INIT_3D => X"A2D57FE00552EA8A00FFFFE8AAAAA80001FF5D2E82000F7FFFFF45AAFFC20BA0",
INIT_3E => X"0000000000000000000000000000000000000FFFBD5400082EBFF45F78400155",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(1),               -- Port A write enable input
DIA(0)   => data_write_a(11),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(11),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(1),               -- Port B write enable input
DIB(0)   => data_write_b(11),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(11),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_12_10 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50080B01BC002006940202C0DE041196A83183000000023322287E0FC000006",
INIT_01 => X"75400D849830C84C5823E0000C17424840000000080000088200002802153231",
INIT_02 => X"18A026B43ED180040147558040090000061800000C06ED9802768F4472C52005",
INIT_03 => X"2A67E34A528D0524A52850528400C8001100000171C02B550618C91A10E55440",
INIT_04 => X"1BC0000100056C8280825DE98154004300C840800850240080CA921084520A07",
INIT_05 => X"02000F832000500C0000941024000852084060202E100001002000448100000C",
INIT_06 => X"819A1D1C3FE01A1A40045408049A50BA4020C6041090001200006200000000F2",
INIT_07 => X"C26A0719CC96CC6ED18A64019695A854870300FA3968B20068FC06080106249F",
INIT_08 => X"D002024B3E040800008C0A002610240D494A06F3460409000000E3F0AD5282E5",
INIT_09 => X"27A06009200040000400120412445D78400001000410420080218029CC807A27",
INIT_0A => X"18000006848A026F000000000000080000F010C100204593F11A6CDF48003BF8",
INIT_0B => X"000000820040402B28050400400432C9349DF21A31A00ACC0000F04F80020001",
INIT_0C => X"00357804611AE45D05D0833430CD0833420CD0C33420CD0833430668619A1000",
INIT_0D => X"0000000000000A74812DF00E87E80A079F9F90FA0280E87E800C7FF3B8002000",
INIT_0E => X"3B6B0E404D26160682082002000401EA0000C40000800A006002818808000000",
INIT_0F => X"A476D61C809A4DA84272592D6246FC1B17B541F97E1B348EDA93900B2B286C56",
INIT_10 => X"30C669E622DBC325CFD881A962454CFBE5403AB99594362B1DB52720165650D9",
INIT_11 => X"F8D2D39A3745261E4A95A110A3F855000E4B1D32BAB504BB7490FCFF912A3834",
INIT_12 => X"B90E9B018C7530200AB8F8BF41F9A22006B37DC8E1F9A21A70116D4C5080651C",
INIT_13 => X"118780319CCA08AB1001ACDF34B8F1C688AB1002AE3F7B807B6289F368828C4C",
INIT_14 => X"2AF020233376A5ECC016B1A827CDA21160F051DE610A34C50427E6E220323E4A",
INIT_15 => X"0077020000000439FDC05C5806781FAB46095A0B5199B0AC55521524F1864022",
INIT_16 => X"000000000000000000000000000000000026C000002884000130921092804010",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"8020080200000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0051B946088881360A95090CB054420290100000000000000000008020080200",
INIT_1A => X"041041041041041041041041041041041049249249249249200100002D451451",
INIT_1B => X"92C964B2592C964B2592C964B2592C964B2592C86432190C86432190C8641041",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000003800F592C964B2592C964B25",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"7DE1000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"ABDFFFF7803DE10AA80000AAAA843FE0008557DFFF0800020105D557FEAA0055",
INIT_29 => X"D5420000051555FFA2AA8200000557DFFFF7AA80000082ABDF5508557DF45002",
INIT_2A => X"82AA8AAAAAFFC00BA007FC2155F7D155545AA80001EFAAFBEAB45557FFDE10AA",
INIT_2B => X"FFAEBFEAA002A801FFF7FFE8A10A28000000A2D155410F7FFFFEBA08003FE000",
INIT_2C => X"5FFFFEAABA000028A105D2ABFE10A2AABFE1055516ABEF5D517DEAAA2AEBFF45",
INIT_2D => X"55002A820AA08557DFFFF7AA82155AAFBE8B45002A974AAAA803DFFFAA843DF4",
INIT_2E => X"000AAD155555A28428BFF002ABDE00A2AABFE10082ABFFEF0855420000004175",
INIT_2F => X"5010495B7AE921C517DE10000000000000000000000000000000000000000000",
INIT_30 => X"BDF6D005B78F7D142ABDFC7F78E3FE28B684070AABE803AE38145B78FD700000",
INIT_31 => X"BEFB455D71F8E00BED547038145B505FFB6A487000005F7AFD7F7A482038002E",
INIT_32 => X"F1FDE821C003FE001C2EAAAAAB6F5C2082007BC217DEBDB55555AA8E071D7AAF",
INIT_33 => X"D517DEAABEAEBFF7DEBA0BDEAA1C2A801C7E3FFEFA10B68407038B6D550428FF",
INIT_34 => X"B68E38FC7BE8A3DF7DF7F5E8A9200002FA285D20BDE28A2A4B8E10555B68BEF5",
INIT_35 => X"F085F47038140010555142082082005F7DFD7F7A482155BEF1E8B6D002090482",
INIT_36 => X"00000000000000000000B6D15756DA28A28BFF082ABAE10B6AAB8E280820B8FE",
INIT_37 => X"ABA5D7FEAB45080015410007FEAA0055517DE000000000000000000000000000",
INIT_38 => X"AB45F780020BA082EBFFEF007BE8BFF5D2ABDF55F7AABDEAAF784154BAF7802A",
INIT_39 => X"D7545AAAE97555A2FBFDF455D556AA00F7D1554BA5D7BC01FFFF8015410007FE",
INIT_3A => X"4154BAF7D1400BAFFD57FE005D043FE10552EAAAAAFFD140000087FC01EFA2FF",
INIT_3B => X"8428A105D7FEABEF55557DEBAFFAEBFFEFAA803DEBA5D2E82155A2FBFDE00FF8",
INIT_3C => X"7D568BEF080402000F7AAA8B55FFAABDFEFF7D16AA0008003FEBA55003DEBAA2",
INIT_3D => X"FFAAA8AAA080028BFF087BD54AA550402145550000010087FFFF45F78402145F",
INIT_3E => X"0000000000000000000000000000000000000F7D5555FFAAAAA8BFF002AAAA00",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(1),               -- Port A write enable input
DIA(0)   => data_write_a(12),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(12),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(1),               -- Port B write enable input
DIB(0)   => data_write_b(12),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(12),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_13_10 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10154A0441836CA2840512822007C18000E02700500030B31B300040081A042",
INIT_01 => X"00000804A000C04800020000000002404001000008220008A200100802110204",
INIT_02 => X"02200430000104000A4700804008000004100000000420918204D3033240400D",
INIT_03 => X"AA4003400008592400000590C40009141100000C6180C0000000C00001E14000",
INIT_04 => X"0800000102400120088054019000004160004190BAA0270000C8100000600206",
INIT_05 => X"21000012040610050040000227003AA0082400E94C1200000824424005220020",
INIT_06 => X"81963B180C001010580000080400000058000004109C00138000020024142581",
INIT_07 => X"002C8008000441600106400A9600010494020002B8AAA000EF003408000E2580",
INIT_08 => X"000000E48194408000A00A001210040441C80320040210000002ABF004102244",
INIT_09 => X"2A004009640040100400940412D4C4004000022000104200802D983000480120",
INIT_0A => X"8000202020401480000000000000080C90090881000145B0111A14004015080D",
INIT_0B => X"00000002004040AA08050400404040C11444000805200A402090024000008002",
INIT_0C => X"8410000A00280020020040800020040800020000801020000800010020400000",
INIT_0D => X"84A14250A055100050100490000500D00040080040290000084E4000B800610C",
INIT_0E => X"DCD13042BEDA36820228000000000000C000400081A08BC812A2092B02850942",
INIT_0F => X"89B9A260857DB400431969CA985D480949D32804A40AB137341C10B7D6A02EC0",
INIT_10 => X"E6ACA678001CE7D0296C213A460CA4271CA2168AEC1017606E6838216FAD4055",
INIT_11 => X"84AD4961C281B20213073C5FC0058008632D30D522CE80239DCC01AB013A4D20",
INIT_12 => X"2E6B13804A4B01D83461299900F6BD583A519104A0EEBD1A141010B2A4C8E116",
INIT_13 => X"89E5E40913419151EE0E94641828F72B5151EE0D184B321037AF5158BB02D085",
INIT_14 => X"562EC0B42162D68EE0073AE1C562EC13D521921A4170300B2B458B56B01C2280",
INIT_15 => X"00888A120240034000E6DC8285028014B82372011FC1E4F5E0A00929684EAF84",
INIT_16 => X"50942509425094250942509425094254940A1421420082020120908800480030",
INIT_17 => X"0942509425094250942509425094250942509425094250942509425094250942",
INIT_18 => X"9425094250942509425094250942509425094250942509425094250942509425",
INIT_19 => X"F7EFBBEEFF3F7DF7FF3E9F7DF7E2450228000000000000000000509425094250",
INIT_1A => X"BAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBF7DFDFDDD555555",
INIT_1B => X"EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAEBAE",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000000000F7EBF5FAFD7EBF5FAFD7",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"2ABEF00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0020105D557FEAA00557DE10AAD5554BA087FFFF55557BD54AAF7FBC01FFA280",
INIT_29 => X"7BD75EF087FFFFEF557BEAB45552E80155AA802AB45AA843FE0008557DFFF080",
INIT_2A => X"FAE820AA5D5557555082ABDF5508557DF45002ABDFFFF7803DE10AA80000AA08",
INIT_2B => X"0051555FFA2AA8200000557DFFFF7AA80000AAD1420AA087BD7555FFD168AAAF",
INIT_2C => X"5557FFDE10AAAEA8BFFA2FBD7545FFD157555085140010F7AEAABFFAAD542000",
INIT_2D => X"BA557BE8A10A284154BAFFAAAAB45007FC2155F7D155545AA80001EFAAFBEAB4",
INIT_2E => X"000A2D155410F7FFFFEBA08003FE00082AA8AAAAAFFC00BA00002AAAAF7D5574",
INIT_2F => X"0492E3F1C71C7BE8A2ABD7000000000000000000000000000000000000000000",
INIT_30 => X"3AE38145B78FD7000005010495B7AE921C517DE10A2DB50482147FFAF554971D",
INIT_31 => X"E3FE28B684070AA1C71D25D7007FFAFD7497BE8B5555208217DBE8A2AB45BE80",
INIT_32 => X"7FD257DFFD568A82FFA4870BA555F5056D002EBDF6D005B78F7D142ABDFC7F78",
INIT_33 => X"FAAAFBFFBED547038145B505FFB6A487000005F7AFD7F7A482038AADF4709214",
INIT_34 => X"AA8E071D7AAFBEFB455D71F8E00A2A0ADBC7A2FFD257DE3DF52555085142000F",
INIT_35 => X"21C002AA92FFDF574824171EAA10B680124BAFFAAAFB45007BC217DEBDB55555",
INIT_36 => X"00000000000000000000B6D550428FFF1FDE821C003FE001C2EAAAAAB6F5C208",
INIT_37 => X"0105D7BE8B55085142010AAD157545F7AEA8B550000000000000000000000000",
INIT_38 => X"01EFF7AAA8B55F7802AABA5D7FEAB45080015410007FEAA0055517DE00A2FFC0",
INIT_39 => X"E8BFF5D2ABDF55F7AABDEAAF784154BA5D5140145007BE8B55087BEAB555D040",
INIT_3A => X"0020BAA2FFD54105D7FC21EFFFD16AA10FF80174AA557FC21EF082EBFFEF007B",
INIT_3B => X"FBC0155085540000FFAEBFFEFF7D1554BA5D7BC01FFFF8015410007FEAB45F78",
INIT_3C => X"87FC01EFA2FFD7545AAAE97555A2FBFDF455D556AA00A2803FF45AAFFC21EFAA",
INIT_3D => X"552EAAAAAFFD1400005D042AA00F7FBD5410085568A10FF80020AAFFAABFF550",
INIT_3E => X"0000000000000000000000000000000000000F7D1400BAFFD57FE005D043FE10",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(1),               -- Port A write enable input
DIA(0)   => data_write_a(13),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(13),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(1),               -- Port B write enable input
DIB(0)   => data_write_b(13),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(13),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_14_10 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10020A000180000284008280000281800000030000000033022000000580002",
INIT_01 => X"000008020000204D006800000030824840000000084000084200090008510200",
INIT_02 => X"0220043170010A600A4D008040080000041000000028009002000F333240800C",
INIT_03 => X"111813400008002400000000C400090011000000610200001104D83000F14000",
INIT_04 => X"0801800100A000000000540084000040000040000800200000C8100000000748",
INIT_05 => X"0100000000001000000000002000080008000000001000000024024001200020",
INIT_06 => X"819EB84028001010000000080400000000000004108000100000020020040081",
INIT_07 => X"92040608000440100102400A94810206844200021DA2A0002000340800062C80",
INIT_08 => X"000000000084400008800A001214040441481500040000000000A7F408002244",
INIT_09 => X"0A0040090002008420401004104444004000020400214A208001000002400120",
INIT_0A => X"0400002020000000000000000000080C8008088100004590111B480040120000",
INIT_0B => X"1000000200404800000504016000002114000008020000020080024000000000",
INIT_0C => X"0410000010000000000040001000000000000040000000000001000000000000",
INIT_0D => X"04810244825010004010000000000000000000000000000000080000B8002104",
INIT_0E => X"0002C38280001202020800000000001000004000000000401022000002040902",
INIT_0F => X"20000587050001404E8084341CBA3404800828805200008000E0E0A000080002",
INIT_10 => X"4D18178E012010C00224004091C3514072C000444A0400080001C1C140001000",
INIT_11 => X"51709A07424142084458476001003809D0104B01C5710044020C4006010500C5",
INIT_12 => X"C26EE3803180C18006519462A00005001460E4730000050A1011004001060049",
INIT_13 => X"01F9E00660318000000538318740000140000001B4600CE80001400000002B62",
INIT_14 => X"0000000AD89857B0E0684411800000003799EB764D000330C300000000E3554B",
INIT_15 => X"0000021002002C000024008284001A0902000422E3F5960080480A0216A07240",
INIT_16 => X"4090240902409024090240902409024090081021020080015134920800480010",
INIT_17 => X"0902409024090240902409024090240902409024090240902409024090240902",
INIT_18 => X"9024090240902409024090240902409024090240902409024090240902409024",
INIT_19 => X"F5579B4E5C8FF0F7BE9D5F7DF650400200000000000000000000409024090240",
INIT_1A => X"9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7BF7DDDDDFCF3CF3D",
INIT_1B => X"F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE79E7",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000003FFF03F9FCFE7F3F9FCFE7F3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"420BA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"BD54AAF7FBC01FFA2802ABEFA2FBE8B55A2AE80000F7D5555555D2AAAABAAAD1",
INIT_29 => X"AA801FFA28402000AAAE955455500155EF0804155EFAAD5554BA087FFFF55557",
INIT_2A => X"7AEA8B45080417400AA843FE0008557DFFF0800020105D557FEAA00557DE10A2",
INIT_2B => X"087FFFFEF557BEAB45552E80155AA802AB4500516AA00A2AE800BAFFFFC20BAF",
INIT_2C => X"0AA80000AA005568ABAA28402010A2843FEBAFFFBD7410A2D168BFF087BD75EF",
INIT_2D => X"005D7FFDF4555517DFEF00043FEAA082ABDF5508557DF45002ABDFFFF7803DE1",
INIT_2E => X"000AAD1420AA087BD7555FFD168AAAFFAE820AA5D5557555002E80155A280000",
INIT_2F => X"0555412AA8ABAAADB40092000000000000000000000000000000000000000000",
INIT_30 => X"50482147FFAF554971D0492E3F1C71C7BE8A2ABD7A2FFEDB55B6A080038E3DB5",
INIT_31 => X"B7AE921C517DE10A2AE851FFB68402038AAAA955554900105FF0800175D7A2DB",
INIT_32 => X"A0800BAE3F1C0092EBAAADB6D080A12410BE803AE38145B78FD7000005010495",
INIT_33 => X"2D568BC71C71D25D7007FFAFD7497BE8B5555208217DBE8A2AB451C556FA00A2",
INIT_34 => X"142ABDFC7F78E3FE28B684070AA00516DABAA28402038B6803DE82F7F5D5410A",
INIT_35 => X"D002A80155B680000105D7FF8F455D5F78FD7000E3FEAA002EBDF6D005B78F7D",
INIT_36 => X"00000000000000000000AADF47092147FD257DFFD568A82FFA4870BA555F5056",
INIT_37 => X"F55FF84000AAAAFBC0145002AA8AAAAAFFC20000000000000000000000000000",
INIT_38 => X"01EF080417555A2FFC00105D7BE8B55085142010AAD157545F7AEA8B55A2FBFF",
INIT_39 => X"EAB45080015410007FEAA0055517DE00A2AA955FFFF80020BAAAAA9754508000",
INIT_3A => X"AA8B555D557FE00A280020BAAAD140000A2AEBFFEF082A82010F7802AABA5D7F",
INIT_3B => X"803DE00FFD557400AAD56AB455D5140145007BE8B55087BEAB555D04001EFF7A",
INIT_3C => X"82EBFFEF007BE8BFF5D2ABDF55F7AABDEAAF784154BA08557FEAAA284000AAFF",
INIT_3D => X"FF80174AA557FC21EF082A80145F780020105D7BEAB45557BE8B45082EBFEBA0",
INIT_3E => X"0000000000000000000000000000000000000A2FFD54105D7FC21EFFFD16AA10",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(1),               -- Port A write enable input
DIA(0)   => data_write_a(14),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(14),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(1),               -- Port B write enable input
DIB(0)   => data_write_b(14),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(14),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_15_10 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000A000000000284000280000001800020030000000033022000000180002",
INIT_01 => X"8000080000000048000000000000026040000000080000080200000000110200",
INIT_02 => X"0020042004010E60004C0080000800000410000000020090020000300245E005",
INIT_03 => X"0000010000080400000000408400480111000000610008000000C00000E54400",
INIT_04 => X"980000010000000088C2550080000040000040000008A00028C8100000120000",
INIT_05 => X"020004012E025000000001322000000A28008000011000000220004D41000000",
INIT_06 => X"819588000800101000011008040000100001060418800510000A620000000092",
INIT_07 => X"0000000800044004010C20008440810284020002102220002000340800062480",
INIT_08 => X"0000000001140800002C0A001214050540C800400406180000002DF004000244",
INIT_09 => X"1E00400900000000000016041044400440000000000042008001000000000022",
INIT_0A => X"0000000000000220000000000000080C00000081000045901118000040000000",
INIT_0B => X"0000000200404000010500004000000114000009000000000000004200000000",
INIT_0C => X"0000000000000000000040001000040001000000000000000001000020000800",
INIT_0D => X"000000000000001001208000180800000000030200000180800C400030002000",
INIT_0E => X"0000000000002600020800000000001080004000000000000002000000000000",
INIT_0F => X"A400000000000000000008000000000000000000000014800000000000000052",
INIT_10 => X"0000000000000000000000010240000000000000000000290000000000000000",
INIT_11 => X"2001C05838120800000000000000000000010000000000000000000000001804",
INIT_12 => X"081004000000000000A010000000000000902000000000180010002020000000",
INIT_13 => X"6600000000000000000024080000000000000000280400000000000000000000",
INIT_14 => X"0000000000200801000000000000000000501001920000000000000000000A40",
INIT_15 => X"0000020000000000000000003000000000000000000A101C3614000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000080000120980000000010",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000400200000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"28BEF00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"5555555D2AAAABAAAD1420BAFF8000010082A954BA00003DFEF085155400F784",
INIT_29 => X"AE95555A2FBE8BEFA2843DE00AA8015400FF84001EFA2FBE8B55A2AE80000F7D",
INIT_2A => X"2FBEAB45F7D56AABAAAD5554BA087FFFF55557BD54AAF7FBC01FFA2802ABEFF7",
INIT_2B => X"A28402000AAAE955455500155EF0804155EFFFFBE8BFF0800174AA557BFDE10A",
INIT_2C => X"A00557DE10F7D1574AAA2D16AB55FFD568BEF087FE8A1055003FE00A2AA801FF",
INIT_2D => X"00AA802AA00AAAE800BA5D0015545AA843FE0008557DFFF0800020105D557FEA",
INIT_2E => X"00000516AA00A2AE800BAFFFFC20BAF7AEA8B45080417400FFFFC21450800154",
INIT_2F => X"8FD7005150438F78A2DBFF000000000000000000000000000000000000000000",
INIT_30 => X"EDB55B6A080038E3DB50555412AA8ABAAADB40092E38E070280024904AA1C043",
INIT_31 => X"1C71C7BE8A2ABD7E3AA9257DA2FFE8BC7BE8E38E10A28017400E38A051FFA2FF",
INIT_32 => X"00124AA557FFDE10A2FBEDB6DF7D16AABAA2DB50482147FFAF554971D0492E3F",
INIT_33 => X"10038E38A2AE851FFB68402038AAAA955554900105FF0800175D7E3FFEFBD700",
INIT_34 => X"000005010495B7AE921C517DE10FFDF50482A2DB6AB45FFD56DBD7087BEAA384",
INIT_35 => X"0FFF1C017D140410400BE8E28A10AAA085082550A1057DBE803AE38145B78FD7",
INIT_36 => X"000000000000000000001C556FA00A2A0800BAE3F1C0092EBAAADB6D080A1241",
INIT_37 => X"4AA0800020BA550028B550855400AAF7AEBDFEF0000000000000000000000000",
INIT_38 => X"7400AAAE975EFA2FBFFF55FF84000AAAAFBC0145002AA8AAAAAFFC2000AAAA97",
INIT_39 => X"E8B55085142010AAD157545F7AEA8B55AAAE821EFAAFBEAB55F7AAA8A00AA841",
INIT_3A => X"417555AAFFFDF450804020AA557BFFE10A2FFFFFEFF7D568ABAA2FFC00105D7B",
INIT_3B => X"D17DF45007FE8AAA08002AAAAA2AA955FFFF80020BAAAAA975450800001EF080",
INIT_3C => X"7802AABA5D7FEAB45080015410007FEAA0055517DE00FFFBC2000AAFBE8B55F7",
INIT_3D => X"A2AEBFFEF082A82010FFD5421EF5D0000010F7AAA8A10AA8017400552A801EFF",
INIT_3E => X"00000000000000000000000000000000000005D557FE00A280020BAAAD140000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(1),               -- Port A write enable input
DIA(0)   => data_write_a(15),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(15),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(1),               -- Port B write enable input
DIB(0)   => data_write_b(15),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(15),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_16_10 : RAMB16_S1_S1
generic map (
INIT_00 => X"DA22C618B1000482B688B186588884862A400438255FC38381441205BA803003",
INIT_01 => X"7045A80028404C211203A952A90341080B173340412000E1005D628000820484",
INIT_02 => X"428406A4000850848330118D0AAC55001349B108818005460229044001C01784",
INIT_03 => X"092C4020000500020000500986812C405000001A48202050000A214AC0650115",
INIT_04 => X"4804A55440256F504025E003A054F46415A4E62B6FE3307943965A00001A1152",
INIT_05 => X"0000001C40A5B950ADB8EA097057ECE14C86D2B7F85AAD17F4B100000B88148C",
INIT_06 => X"415401DCDCF2C0A8030140BCB0820A200342A1C641C1E8782F508F2B00003584",
INIT_07 => X"002701881A3202080AE00480A2002840BE1480FA004342AA6F12000054004867",
INIT_08 => X"08C54828091002000002B32A8C19064E486A8001510000014140C1E2A14891E0",
INIT_09 => X"015452B103020814004088B64102680B6596594800400413CAC0208944800000",
INIT_0A => X"96AA000484094C000000000000012C9000A0000D0A80000BF8028E87C1B99270",
INIT_0B => X"014808A02004200E540480212000A448C0082024AE50064B44000000000002A2",
INIT_0C => X"0004000D5846256AAEA811150445411150445411150445411150422A088A8200",
INIT_0D => X"00000004010042A204A0C5817D00005034052E40000817D00440004004AD3240",
INIT_0E => X"632B2673FA4587978A2004102800809225545155121740000004900090000000",
INIT_0F => X"00C6564CE7F4EA4B940076D296D003030800462CBD320018CAAAACFE9164C800",
INIT_10 => X"28834ADB1440A114793A4A30A40839AA14910D08DCB2640031955559FD3AC990",
INIT_11 => X"594AB0B1A025371CA0E034E8443C097A800EB090D4AAC91208ED2FA0CE5E09B1",
INIT_12 => X"7B50446083001B94BB38C540EBE61284BB304880E3E4579EDC00992980D58033",
INIT_13 => X"5511121840E7A2CD952ECC12ABC3E6ACB3DFB12ECE315000F61FF1727A85FDBC",
INIT_14 => X"75DEB07F6F2E7084517F126F8395CB2BEFBAB8BA8AF698228CC5E2F08ECA5159",
INIT_15 => X"5580A840A8009F8B108C80A1021B080AFC0DF6422C6077F4A77F20D0C0E21084",
INIT_16 => X"0000000000000000000000000000000000044000102A0001148442A110810359",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"558D11544C690DA64C1C4F68A360400000000000000000000000000000000000",
INIT_1A => X"14D14D14D14D14D14D14D14D14D14D14D14514514514514529E5F87869E79E78",
INIT_1B => X"D1E8F47A3D1E8F47A7D3E9F4FA7D3E9F4FA7D3E9F47A7D1E9F47A7D1E9F4D14D",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000007D3E9F4FA7D3E8F47A3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"C00AA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"03DFEF085155400F78428BEF087FFFFEFF7D168B55AAD17FFFF552EBFE00007F",
INIT_29 => X"2E975EFF7D568BFFFF80175EF0004000BA552A821FFFF8000010082A954BA000",
INIT_2A => X"55540000082EAABFFA2FBE8B55A2AE80000F7D5555555D2AAAABAAAD1420BA5D",
INIT_2B => X"A2FBE8BEFA2843DE00AA8015400FF84001EF0000020AA5D00154005D043FF455",
INIT_2C => X"FA2802ABEF557BEABEF5D0415410087FD74BAAAAEBFFEF557FC00AAF7AE95555",
INIT_2D => X"FFFFAABFEAAFF84001FF002A821FFAAD5554BA087FFFF55557BD54AAF7FBC01F",
INIT_2E => X"000FFFBE8BFF0800174AA557BFDE10A2FBEAB45F7D56AABA082A97545F7D16AB",
INIT_2F => X"FFEF552AB8E38087FC2092000000000000000000000000000000000000000000",
INIT_30 => X"070280024904AA1C0438FD7005150438F78A2DBFF0871F8FC7E3D56AB6DBEDB7",
INIT_31 => X"AA8ABAAADB400924920925EFF7D16ABFFE38E175EF1400000BA412E871FFE38E",
INIT_32 => X"0A1240055003FF6D5551420101C2EAFBD7A2FFEDB55B6A080038E3DB50555412",
INIT_33 => X"57FC00BAE3AA9257DA2FFE8BC7BE8E38E10A28017400E38A051FF0804050BA41",
INIT_34 => X"4971D0492E3F1C71C7BE8A2ABD74975EDBC7550E12410087FD74AAB6AABFFC75",
INIT_35 => X"A08249756DF7D168BC7F7AABAEAAF780051C70824851D7A2DB50482147FFAF55",
INIT_36 => X"00000000000000000000E3FFEFBD70000124AA557FFDE10A2FBEDB6DF7D16AAB",
INIT_37 => X"B55A2D16ABEFFFFBFDFFF552AAAAAA007BC00000000000000000000000000000",
INIT_38 => X"20AA002A955EFAAAA974AA0800020BA550028B550855400AAF7AEBDFEF08516A",
INIT_39 => X"000AAAAFBC0145002AA8AAAAAFFC20000000021EFF7D568BFFA2AA955FF5D040",
INIT_3A => X"E975EF0800174BA002E820105D003DFEF5D51420005D2ABFF45A2FBFFF55FF84",
INIT_3B => X"7BD74AAF7AEBDF455D7BC20BAAAAE821EFAAFBEAB55F7AAA8A00AA8417400AAA",
INIT_3C => X"2FFC00105D7BE8B55085142010AAD157545F7AEA8B5500557DF45552A8200000",
INIT_3D => X"A2FFFFFEFF7D568ABA0804155FFF7D568B55FFAAAAABAFF8415545000015555A",
INIT_3E => X"0000000000000000000000000000000000000AAFFFDF450804020AA557BFFE10",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(2),               -- Port A write enable input
DIA(0)   => data_write_a(16),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(16),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(2),               -- Port B write enable input
DIB(0)   => data_write_b(16),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(16),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_17_10 : RAMB16_S1_S1
generic map (
INIT_00 => X"5284CE4FB7BD2C8994A13392DBD02E14006B82AC7E800D44D3DD2FD5F9B961C0",
INIT_01 => X"2EACD01F7E03FC6793F2199B39FC233C11D93AE6F3BB92B32091DBC339B24542",
INIT_02 => X"E63CCCC00A82C08092A2AFAE667033DB50853379C10BFDC5C6F4044443C817C6",
INIT_03 => X"7FF183635AEF9E3635AEF9E18E237040404446965C0607EE6DB7854AC4DE060C",
INIT_04 => X"D78AC33FB604488B000892EF17BE6D84196482236FE100294152E294350FB697",
INIT_05 => X"081B5F9B409420D0CDB47A05403F6CE0C08A4AB7F840EDB6F48100DFC8081081",
INIT_06 => X"768465354781CBC30316367077B4BDB50646E8D87100A8201ED01C19C020F71A",
INIT_07 => X"4002A110C922480A82D0841147162C48EBB9537A0022DC67987042EE976ABEA7",
INIT_08 => X"DB931BFEF91C00002CC0E019C0C82A4E4820C15A2330E004401891181168C4D1",
INIT_09 => X"09F3A1BC11EFBC66DB65307071477FF1030C397C060B4254064302042F803A69",
INIT_0A => X"3F330802162F3B7EE3F3EC7C7DEF207000F00059D2ED56D7EED2ED3C9A867DC0",
INIT_0B => X"185C44B91BC1740B7605040BE0018CFC7429F326B9E822FFC00074D5A0AB033A",
INIT_0C => X"00367A28FC1B7F7FEFFCFBFF3EFFCFBFF3EFFCFBFF3EFFCFBFF3EFFE7DFF9E00",
INIT_0D => X"0000000008004BA78428C7AD7FC94B533F5B4FFBD2FAD7FCCA786D43FE67C218",
INIT_0E => X"BA494CEBFD4F2667ABB6F68B29760593F33FA0CF170F40006001B1A05C000000",
INIT_0F => X"7F749299D7FAEB237DFE5865B6D2BF23265CBACE542A6FEE92333AFF33E0A9BF",
INIT_10 => X"F6C24B6D18C3C9F8E2881F3F787D776B5DB94A09955054DFDD246675FE7AC153",
INIT_11 => X"BFB349E08FF9A27EDE9FA8AEFD9E7467BFCB195CFEB56A1A70D34D1706FFFA3E",
INIT_12 => X"6FE219CA80725B875EED723FF7FCB2875EDAAFEAF7FD929BFD55BBC71D79F639",
INIT_13 => X"546670D018E7A6E581D7B6AB75FDFCECA6E581D7BB5DDFC6FF0EB7D7E859FDB5",
INIT_14 => X"B978177F6D6AF5ECDB5FB76A5F5FA165B456E0FB308710C49FCFB741598B9C7E",
INIT_15 => X"CFDAAB00AC00A8BBFC8B501CF7A0FED9A540EA1952586CEB54D143ACFF9A3BA9",
INIT_16 => X"000000000000000000000000000000000026E100002F382DBD9ECFE117805F20",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"4372003009EDCC4052E917114F981800C0000000000000000000000000000000",
INIT_1A => X"BA69A69AEBA69AEBA69A69AEBA69AEBA69A69A69A69A69A68698686981D75D74",
INIT_1B => X"6A351A8D46A351A8D068341A0D068341A0D068341A0D46A341A0D46A341A69AE",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000000000046A351A8D46A351A8D4",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"7FEAA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"17FFFF552EBFE00007FC00AA087FFFFFFFFFFFFFEFF7FBEAB450804001EFAAD5",
INIT_29 => X"D168A000004020AA5D7BE8B450051401EF087FD74AA087FFFFEFF7D168B55AAD",
INIT_2A => X"D7FEAB55FF80175EFFF8000010082A954BA00003DFEF085155400F78428BEFAA",
INIT_2B => X"F7D568BFFFF80175EF0004000BA552A821FF5D00020BA552A82000552A821555",
INIT_2C => X"AAAD1420BAFFFFFDF45AAD17FFFFAAFBC01EF5D0015555557BFDEBA5D2E975EF",
INIT_2D => X"BA007FEABEF005555555A2D1554BAA2FBE8B55A2AE80000F7D5555555D2AAAAB",
INIT_2E => X"0000000020AA5D00154005D043FF45555540000082EAABFF00516AA10552E820",
INIT_2F => X"8B550000071EFB6DF7AE92000000000000000000000000000000000000000000",
INIT_30 => X"F8FC7E3D56AB6DBEDB7FFEF552AB8E38087FC2092147FFFFFFFFFBFDFC7EBF5E",
INIT_31 => X"150438F78A2DBFFBED16AA381C0A07082497FEFB6D1451471EF007BD04920871",
INIT_32 => X"2A850105D2A80155417BEFB6DEB8E175FFE38E070280024904AA1C0438FD7005",
INIT_33 => X"D7BFAEBA4920925EFF7D16ABFFE38E175EF1400000BA412E871FF550A0009249",
INIT_34 => X"E3DB50555412AA8ABAAADB40092FFF5FFF6DAADF7FFD7B6F1C71EF55001756D5",
INIT_35 => X"7145B6AA28492487082007FEDBD700515556DA2DF50492A2FFEDB55B6A080038",
INIT_36 => X"000000000000000000000804050BA410A1240055003FF6D5551420101C2EAFBD",
INIT_37 => X"FEFF7FBFFF55A2D16AB550000175EFFFFBEAA000000000000000000000000000",
INIT_38 => X"55EF087FC200008516AB55A2D16ABEFFFFBFDFFF552AAAAAA007BC0000557FFD",
INIT_39 => X"020BA550028B550855400AAF7AEBDFEFF7D568AAA5D2A97410007BFFFFF55515",
INIT_3A => X"A955EF5D2E80010002A954005D2A82155087FFFFEFAAAA975EFAAAA974AA0800",
INIT_3B => X"D1575FF5504175EF5D7FEAAAA0000021EFF7D568BFFA2AA955FF5D04020AA002",
INIT_3C => X"2FBFFF55FF84000AAAAFBC0145002AA8AAAAAFFC2000FFD57DFFFAAFFFDF55FF",
INIT_3D => X"5D51420005D2ABFF45557FE8AAA000415410007BFFF450051555EFA2FBC0000A",
INIT_3E => X"00000000000000000000000000000000000000800174BA002E820105D003DFEF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(2),               -- Port A write enable input
DIA(0)   => data_write_a(17),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(17),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(2),               -- Port B write enable input
DIB(0)   => data_write_b(17),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(17),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_18_10 : RAMB16_S1_S1
generic map (
INIT_00 => X"69844019080000A21A611406840014122A641074155FC28A2024001001801003",
INIT_01 => X"7443D920034004180005E9E3C90360C0041C0181002001602025800008440084",
INIT_02 => X"E2DCCCE61D5C008103F2000781FC0FEDEAC2161B0B8FB0008620044443006010",
INIT_03 => X"884E300802006900802006995C896D605200000856E24A040000640052141103",
INIT_04 => X"480520FC026125AC0025C9122644E3E40EC8E2001001302281841A009038A86A",
INIT_05 => X"432000040089983070019400F01010004C8DB841405A80A100B586200FAC24AE",
INIT_06 => X"09044359DC7040000000002C109B0E0A00A1104641C0803804000707284600E1",
INIT_07 => X"400D10100400481D5EB08501620000007500CE801241021FE78E404860140060",
INIT_08 => X"00880C0106A0528020019307CC082A0A4A6A01ED725021400040D028000A9729",
INIT_09 => X"00117063038000282081402E4106400B6186128040600C10C1C0200950508110",
INIT_0A => X"C0C30C2E21580C874004008080003C32A10A19090C02010E1022944061688000",
INIT_0B => X"0180A8062026000DC425C0301311324AA2373088479105D044A1022000001835",
INIT_0C => X"0D89844703649000000200000000000000000000000000000000000000000010",
INIT_0D => X"0D8306C182701404C1973010802020404084001E00010802046092B5001FB365",
INIT_0E => X"528EB314068AB8B803DB00002900800400FC503F08180050942E4200020C1B06",
INIT_0F => X"40A51D66280D6032C5F96D3C51555D5D7D5AA87285820814A3CCC501C2A60820",
INIT_10 => X"8B35A3FEBF1FEDFD9C2B30E0468AAAD5D48F37E8FC1304102947998A03984C10",
INIT_11 => X"440FE1DD772D37A0A321BC6968F32658BF2D4F2A80BF8FE3F9FE3AC362080529",
INIT_12 => X"5487910D7E5A6D961A28456A1832E5161A100DD5182BC54020EA67A189C6ED36",
INIT_13 => X"AA444CAF91EDD1B725868403BE06323551B725868A100ABD119753B70964122B",
INIT_14 => X"EDC259048ACD868EE3803D65CEDC258A8F80D55E007C3F8EBB56F4C5362C978F",
INIT_15 => X"3F240014BE84370001B6922070440556B15F7FABBC0031BCF2257C41634B14D4",
INIT_16 => X"C1B06C1B06C1B06C1B06C1B06C1B06C1B0491069068000004060300A005A0118",
INIT_17 => X"1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06",
INIT_18 => X"B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C",
INIT_19 => X"B28BBECEB80EE173C2300F7DF16000000000000000000000000041B06C1B06C1",
INIT_1A => X"8A28A28AAAAAAA28A28A28AAAAAAA28A28A28A28A28A28A2910591505C104104",
INIT_1B => X"28944A25128944A25128944A25128944A25128944A2552A954AA5128944AAAA2",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000128944A25128944A251",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"9540000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"BEAB450804001EFAAD57FEAA087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974BA082E",
INIT_29 => X"7FFFFFFFFFBFDF45AAD568B55080028B55002E82000087FFFFFFFFFFFFFEFF7F",
INIT_2A => X"0043DE10AA843DE00087FFFFEFF7D168B55AAD17FFFF552EBFE00007FC00AA08",
INIT_2B => X"0004020AA5D7BE8B450051401EF087FD74AAAAFFFDF45A2D16AB55F7FFFFFFF0",
INIT_2C => X"0F78428BEFAA80000000804154BA55042ABEF5D7FD75FFAAD540145AAD168A00",
INIT_2D => X"00082E95555085168A10557FD7545FF8000010082A954BA00003DFEF08515540",
INIT_2E => X"0005D00020BA552A82000552A821555D7FEAB55FF80175EF5D00020105D2A974",
INIT_2F => X"DFFF5D2A954AA082A92428000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFBFDFC7EBF5E8B550000071EFB6DF7AE921C7FFFFFFFFFFFFFFFF7FBF",
INIT_31 => X"AB8E38087FC2092087FFDFC7E3F1FAF55A2DF6DB7D1C002AB7D002A82028147F",
INIT_32 => X"DF6DB7DE3F5FAFC708003DE28B68E38E280871F8FC7E3D56AB6DBEDB7FFEF552",
INIT_33 => X"ADF4516DBED16AA381C0A07082497FEFB6D1451471EF007BD0492B6F1F8F55AA",
INIT_34 => X"1C0438FD7005150438F78A2DBFFA28407038140410492550A2ABC7497BD25FFA",
INIT_35 => X"F5D0E05000492097428002E9557D1C516FA28417BD5545E38E070280024904AA",
INIT_36 => X"00000000000000000000550A00092492A850105D2A80155417BEFB6DEB8E175F",
INIT_37 => X"FFFFFFFFDFEFF7FBFFFEF552E974AA082A820AA0000000000000000000000000",
INIT_38 => X"ABEF002A800AA557FFDFEFF7FBFFF55A2D16AB550000175EFFFFBEAA00557FFF",
INIT_39 => X"6ABEFFFFBFDFFF552AAAAAA007BC0000087BFDF45AAD568B55AAFBFDFEF55042",
INIT_3A => X"FC2000FFD56AB45A2FFFDFFFAAD16AB4500043DEAAFFAEAAAAA08516AB55A2D1",
INIT_3B => X"2AA8B45087FC01EFA2FFD55EFF7D568AAA5D2A97410007BFFFFF5551555EF087",
INIT_3C => X"AAA974AA0800020BA550028B550855400AAF7AEBDFEFA280154BA55040000055",
INIT_3D => X"087FFFFEFAAAA975EF5D2E974000804154BA082A975EF5D517DEAA007BD5545A",
INIT_3E => X"00000000000000000000000000000000000005D2E80010002A954005D2A82155",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(2),               -- Port A write enable input
DIA(0)   => data_write_a(18),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(18),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(2),               -- Port B write enable input
DIB(0)   => data_write_b(18),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(18),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_19_10 : RAMB16_S1_S1
generic map (
INIT_00 => X"042200000000000041088001001AA00000000000000000000000500802000003",
INIT_01 => X"040048000024000000000404000000000A22000800000800004A200000000001",
INIT_02 => X"200C8840085EB00480060000001C008002489E0F000405EA0004040404000000",
INIT_03 => X"24004000000000000000000900002C4050000000000069500208400002E14100",
INIT_04 => X"4800200C0000000044002000C80020E40000E200000130200188000000800100",
INIT_05 => X"000000000080181000000000701000004C8000000058800000B1000009880480",
INIT_06 => X"80500081081040000000002C100040400000004641C080380400070100000000",
INIT_07 => X"4020109801A4CE005C00048380142810010564C4100114012002402028044808",
INIT_08 => X"0070700000000000000083004C3902420062000020E0000100004082A140102B",
INIT_09 => X"001150200000000000000026400000016186100000000010C04002C000000000",
INIT_0A => X"007C00008082C0002000000000002C3000000004050001030102040000000000",
INIT_0B => X"0000000000000000000000000000010000800011000000000000000000000BC0",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"000000000000000000000000000000042000760000000000000000010004B200",
INIT_0E => X"0D74002280300F0002FB069040000060000C5003000800000000000000000000",
INIT_0F => X"C01AE8004500744C780687DBA828008080A5FC0D385598035D0008A00C015660",
INIT_10 => X"39D8140040201BF861F0E7D693E6170022408116DFE0AB3006BA0011401D02AC",
INIT_11 => X"5412E4997F5249FD005043B8680CC98F00D0F2DD0140100406FE053A98F6ECC7",
INIT_12 => X"7418663001858040E153888000010840E165D0000000285C246A181C03FE4662",
INIT_13 => X"8199830066F0020858385974000001260208583854E2200000660208D6B1423F",
INIT_14 => X"8235AC508FCE8811042040F008235AE04420C040CF00C031C80009B8F224978B",
INIT_15 => X"030004E00000C220010808C10D9A92A74CD7CF4A09051110AD5A3C9200B7F280",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000118",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"07208BBA3F0C7010C660C7441920000000000000000000000000000000000000",
INIT_1A => X"861869A61861861861869A61861861861861861861861861A8208C4C1534D34C",
INIT_1B => X"984C26130984C26130984C26130984C26130984D26930984C26130984C261861",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000984C26130984C26130",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"174BA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFDFEF5D2A974BA082E95400F7FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0004",
INIT_29 => X"FFFFFFFFFFFFFFFFF7FBFDFFF552E974BAA2FFFFE10087FFFFFFFFFFFFFFFFFF",
INIT_2A => X"004001EFAAAEA8ABA087FFFFFFFFFFFFFEFF7FBEAB450804001EFAAD57FEAAF7",
INIT_2B => X"FFFBFDF45AAD568B55080028B55002E82000F7FFFFFFFFFFFFDFEFA2D568B550",
INIT_2C => X"0007FC00AAF7FFFFFFFF7FBE8B55AAD16ABEF5D2ABFF55080402010087FFFFFF",
INIT_2D => X"55A2FFFDFEF5D2EBFE00AAFFFFEBA087FFFFEFF7D168B55AAD17FFFF552EBFE0",
INIT_2E => X"000AAFFFDF45A2D16AB55F7FFFFFFF00043DE10AA843DE00557FFDFEFA2D16AB",
INIT_2F => X"FFEF552A974AA0000104AA000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFF7FBFDFFF5D2A954AA082A92428E3FFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"0071EFB6DF7AE92EBFFFFFFFFFFFFDFEFF7F5FAFC7492A974AAB6F5F8E101C7F",
INIT_32 => X"F1F8FD7AAD16AB450000001FFBEA4A8AAA147FFFFFFFFFBFDFC7EBF5E8B55000",
INIT_33 => X"00000010087FFDFC7E3F1FAF55A2DF6DB7D1C002AB7D002A82028FFFFFFFEFF7",
INIT_34 => X"BEDB7FFEF552AB8E38087FC2092F7FBF8FC7E3F5EAB45B6DF6FBEF5D2AB8F7D0",
INIT_35 => X"84971F8FC7AAD56DB6DBEF5F8FD7412ABFE28B6F5F8E820871F8FC7E3D56AB6D",
INIT_36 => X"00000000000000000000B6F1F8F55AADF6DB7DE3F5FAFC708003DE28B68E38E2",
INIT_37 => X"FFFFFFFFFFFFFFFFFDFEF552E954AA0004000AA0000000000000000000000000",
INIT_38 => X"54AAF7D568A00557FFFFFFFFFFFDFEFF7FBFFFEF552E974AA082A820AAA2FFFF",
INIT_39 => X"FFF55A2D16AB550000175EFFFFBEAA00A2FFFFFFFF7FBFDFFFFFD568B55002A9",
INIT_3A => X"A800AAF7FBFDFEFF7D56AB45AAD56AB450004001EFFF842AAAA557FFDFEFF7FB",
INIT_3B => X"FFFFFFF552AA8BEF080402000087BFDF45AAD568B55AAFBFDFEF55042ABEF002",
INIT_3C => X"8516AB55A2D16ABEFFFFBFDFFF552AAAAAA007BC0000FFFBE8B55AAD168B55F7",
INIT_3D => X"00043DEAAFFAEAAAAA08556AB55A2D57FFFFF7D568B45002ABDEAAFFD16AA000",
INIT_3E => X"0000000000000000000000000000000000000FFD56AB45A2FFFDFFFAAD16AB45",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(2),               -- Port A write enable input
DIA(0)   => data_write_a(19),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(19),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(2),               -- Port B write enable input
DIB(0)   => data_write_b(19),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(19),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_20_10 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000003",
INIT_01 => X"F55FF80000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"E05022020800008400F655001FFCFF80018FA804400000000000004400000001",
INIT_03 => X"00000000000000000000000900002CC07000000000000000000000000000013F",
INIT_04 => X"68002FFE40900010000180000001FFEC0012EE0C001370F40780000000000000",
INIT_05 => X"0840000880FCBBF0100E204DF0F88311DD8005080679800000F3000029980580",
INIT_06 => X"001000030817C8E8840155FDF9001001050023F6C3C3D0F87FA19F7F011000E4",
INIT_07 => X"000000090492260800008000EE00000000000000002101FF2002C00000004018",
INIT_08 => X"2A040001071004000013FF7FCA302C0C0008214800002101554031F800000000",
INIT_09 => X"801F57F200000090000489FEC0000001EFBEF0040008023FDFC0000000004006",
INIT_0A => X"0000000008000000000000000000ADF000000200000008000008028300110230",
INIT_0B => X"0000000000000800080000000000000000000000000000000800800A40000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"000000040900005C848538000020000000800000080000020000800101FFB600",
INIT_0E => X"00800000003A010003000000000000600FFC53FF001800000002004080000000",
INIT_0F => X"0001000000007408040000004000000004E9000008020000200000000E800800",
INIT_10 => X"00200000000313100010002000008000000000129600040000400000001D0010",
INIT_11 => X"81C012060000000000218F7840000100800004000000000066C0000080080000",
INIT_12 => X"800000000017C000100000000001A800080000000001A8040000002840008185",
INIT_13 => X"0000000006F00000100200000000012600001004000000000066000000801040",
INIT_14 => X"0000200410100000000005F00000020080090A0000000085C800002000586000",
INIT_15 => X"FF00400000000000020020020001000040283024E4F2860400008000030ED080",
INIT_16 => X"00000000000000000000000000000004010201001003020200000000000127DB",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"A0700030038200010089120104D2040020000000000000000000000000000000",
INIT_1A => X"2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2C30C30C30C30C306982121A1E79E79",
INIT_1B => X"32190C86432190C86432190C86432190C86432190C86432190C86432190CB2CB",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000432190C86432190C864",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0201000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF552A974AA0004174BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA0804",
INIT_29 => X"7FFFFFFFFFFFFFFFFFFFFFFEF552E954AA000400000F7FFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E954BA007FC00BA087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974BA082E9540000",
INIT_2B => X"FFFFFFFFFF7FBFDFFF552E974BAA2FFFFE10FFFFFFFFFFFFFFFFFFFFFBFDFFF5",
INIT_2C => X"FAAD57FEAA007FFFFFFFFFFFFFEFF7FBFFF550800020BAAAD56AAAAF7FFFFFFF",
INIT_2D => X"EFF7D56AB450000021EFA2D57DE10087FFFFFFFFFFFFFEFF7FBEAB450804001E",
INIT_2E => X"000F7FFFFFFFFFFFFDFEFA2D568B550004001EFAAAEA8ABA5D7FFFFFFFFFFFDF",
INIT_2F => X"FFFF5D2E954AA080005000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFEF552A974AA0000104AAFFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"A954AA082A92428087FFFFFFFFFFFFFFFFFFBFDFEF5D2E974AA000A07000E3FF",
INIT_32 => X"FFFFFEFF7FBFFFFF552E974AA0071C50BA1C7FFFFFFFFFFFFFFFF7FBFDFFF5D2",
INIT_33 => X"EDF6FABAEBFFFFFFFFFFFFDFEFF7F5FAFC7492A974AAB6F5F8E10E3FFFFFFFFF",
INIT_34 => X"EBF5E8B550000071EFB6DF7AE921C7FFFFFFFFFBFDFEFE3F5F8F450004050AAB",
INIT_35 => X"A497FFFFFFF7FBF8FC7EBD168B450804021FFB6D57DE28147FFFFFFFFFBFDFC7",
INIT_36 => X"00000000000000000000FFFFFFFEFF7F1F8FD7AAD16AB450000001FFBEA4A8AA",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2A954AA0800174100000000000000000000000000",
INIT_38 => X"74AA002E95410A2FFFFFFFFFFFFFFFFFFFFFDFEF552E954AA0004000AAFFFFFF",
INIT_39 => X"FDFEFF7FBFFFEF552E974AA082A820AA087FFFFFFFFFFFFFEFF7FBFDFFF5D2A9",
INIT_3A => X"568A00AAFFFFFFFFFFBFDFEFFFFFFDFEF5D2E954AA0051554BA557FFFFFFFFFF",
INIT_3B => X"D16AB450804174AAFFFFFFEBAA2FFFFFFFF7FBFDFFFFFD568B55002A954AAF7D",
INIT_3C => X"57FFDFEFF7FBFFF55A2D16AB550000175EFFFFBEAA005D7FFFFEFF7FBFDFFFAA",
INIT_3D => X"0004001EFFF842AAAA087BFDFEFF7FFEAB45A2D568B550804001EFF7D57DEBA5",
INIT_3E => X"0000000000000000000000000000000000000F7FBFDFEFF7D56AB45AAD56AB45",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(2),               -- Port A write enable input
DIA(0)   => data_write_a(20),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(20),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(2),               -- Port B write enable input
DIB(0)   => data_write_b(20),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(20),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_21_10 : RAMB16_S1_S1
generic map (
INIT_00 => X"4A302428B824900A128C090A5C1800261500213C005FE812D10420054085A202",
INIT_01 => X"001FFE3440B609703B0427F801A40B8115BC4F655300340288A40D30040E4DD8",
INIT_02 => X"E00424256888D8819801000F9FFFFFFFF149FF1FCA448046C60A0D2437C517F9",
INIT_03 => X"20030640003250640003250F06002CC1740002019824E001CD357832440001FF",
INIT_04 => X"EA2C3FFD400006E04401A8837001FFFC004AEF00080B70E08FB5789421007C5C",
INIT_05 => X"00011A0C40F9FFF80920954FF0F00809DF84A0202879800000F3000029980780",
INIT_06 => X"0805984B7A1FC0A0000101FFF0480080002281F7C3C381F87C03DFFF00009004",
INIT_07 => X"B424068086A205481A60A19000908204A855B000A08A61FF20C3D004D331D340",
INIT_08 => X"1BFA0001600802000023F7FFC08D234B40C2028253000040114200000D0226C0",
INIT_09 => X"EF1F5FF054096C6ADBA169FFC202B1C1FFBEF0440021083DFFCE22DC2880E24D",
INIT_0A => X"45FF0C004041D84862A28C54518DBFF00020004C0A6044901112A0908AA0A300",
INIT_0B => X"018C241102068006C620C03882019480E63180855A492712CC01C49C20201BFE",
INIT_0C => X"08A9464116544302C02D92236488D92236488D92236488D922366446C911B210",
INIT_0D => X"08800444021048034004001890000806002804A0822189000900D80621FFBE00",
INIT_0E => X"060580261013813A2CC396506102C4053FFD5BFF00A04A00200602CA52001100",
INIT_0F => X"080C0B004C202621A85C09411500135844C196D3606941018150098404C1A304",
INIT_10 => X"B02901013416181C96C2C9C600890A2028172192C460D1820302A0130809834A",
INIT_11 => X"9C5E803408250180AC268D185DB3F4350B811068C00049A0A4AA68F05C96A001",
INIT_12 => X"002C006560138F032B1804101244C883052208209040CC849063A747512B7678",
INIT_13 => X"41401E240665750440C9488280254530314080C2C601040420352148A00501B1",
INIT_14 => X"500811204D000700114204A70422016149916011008CAA8858850B00C32591C0",
INIT_15 => X"FFC06E60AC0496022300233104663040808E991765205000070121D41D18D098",
INIT_16 => X"40100401004010040100401004010040102090010008000001C0E010020007DF",
INIT_17 => X"0100401004010040100401004010040100401004010040100401004010040100",
INIT_18 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_19 => X"FFEF9FEEFF7FFDF7FF3E3DFDF7E0000000000000000000000000401004010040",
INIT_1A => X"BEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBFFDFDFFFCF3CF3F",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFEFF7FBFDFEFF7FBFDFEFBEF",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000FFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0001000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E954AA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0004",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA0004154BAFFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"52E974BA0804000AAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0004174BAFF",
INIT_2B => X"FFFFFFFFFFFFFFFFEF552E954AA000400000007FFFFFFFFFFFFFFFFFFFFFFEF5",
INIT_2C => X"A082E95400007FFFFFFFFFFFFFFFFFFFFDFEF5D2E974BA002E97400007FFFFFF",
INIT_2D => X"FFFFFBFDFEF5D2A954AA002E974BA087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFBFDFFF5D2E954BA007FC00BA5D7FFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA000002000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080005000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"A974AA0000104AAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974BA0000174AAFFFF",
INIT_32 => X"FFFFFFFFFFFFDFEF552E954BA080A000AAE3FFFFFFFFFFFFFFFFFFFFFFFEF552",
INIT_33 => X"02A95400087FFFFFFFFFFFFFFFFFFBFDFEF5D2E974AA000A07000007FFFFFFFF",
INIT_34 => X"F7FBFDFFF5D2A954AA082A924281C7FFFFFFFFFFFFFFFFFFBFDFEF5D2A974BA0",
INIT_35 => X"A557FFFFFFFFFFFFFFFF7FBFDFFF552E974BA0020924BA1C7FFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000E3FFFFFFFFFFFFFFEFF7FBFFFFF552E974AA0071C50B",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0000020000000000000000000000000000",
INIT_38 => X"74BA0000174BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954AA080017410FFFFFF",
INIT_39 => X"FFFFFFFFFFDFEF552E954AA0004000AAF7FFFFFFFFFFFFFFFFFFFFFFFEF552A9",
INIT_3A => X"E95410087FFFFFFFFFFFFFFFF7FBFDFEF5D2A954BA082E800AAA2FFFFFFFFFFF",
INIT_3B => X"FBFFFFF552E954BA002E97410087FFFFFFFFFFFFFEFF7FBFDFFF5D2A974AA002",
INIT_3C => X"57FFFFFFFFFFFDFEFF7FBFFFEF552E974AA082A820AA557FFFFFFFFFFFFFEFF7",
INIT_3D => X"5D2E954AA0051554BA5D7FFFFFFFFFBFDFEFF7FFFFFEF5D2A974BA0000020AA5",
INIT_3E => X"0000000000000000000000000000000000000AAFFFFFFFFFFBFDFEFFFFFFDFEF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(2),               -- Port A write enable input
DIA(0)   => data_write_a(21),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(21),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(2),               -- Port B write enable input
DIB(0)   => data_write_b(21),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(21),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_22_10 : RAMB16_S1_S1
generic map (
INIT_00 => X"5290F4CDE914905A14A43D33F488243E17122300F55FEB189B343A1140548380",
INIT_01 => X"A54007B259F6A975386262000C344BA9573C6FF57B18A5FB0ABFCD3C2C5F4F0C",
INIT_02 => X"021DFF8C38B3C009D203551040030071869D0040180AA2DC53DB89BEA8204001",
INIT_03 => X"2603475A969D0475A969D0460EAA401005111011BD506954EDB40F5EF41434C0",
INIT_04 => X"922D9002100ED69E443D988B0D5400103E48003D0800011E803B06B5B9125A15",
INIT_05 => X"281B5A0C06000408F4DF9422010D8802022F2124A8022492580040440002021C",
INIT_06 => X"F780C4C052881ADA0E05440205DA50930FA182010004700083E220800440B588",
INIT_07 => X"049D028B93FB561833D8094A02F5EA92FD7247E10305C40040D136E6A023F7FC",
INIT_08 => X"00028241680A0E002A9400803A884B5B5206B7C2E53CA25144009007A64EBD64",
INIT_09 => X"41008810240240C6694008010392354010000560141801002028A83D2A08E06D",
INIT_0A => X"34000000848BCA6902A29C54539C020E11810098D4067EFF9FF284D483E2AB41",
INIT_0B => X"500001840000C80B410014088040F4A944B1AA313C0022AA0011C0DC00028001",
INIT_0C => X"80B14004D158C8CA24A1C2A870AA1C2A870AA1C2A870AA1C2A872550E1543800",
INIT_0D => X"80A14050A01509E050854498B5281A1C34E506A2C6898B52A154DAC6B6000850",
INIT_0E => X"0B03001A483A4146603050080410089180008800143D83888281A2034A850142",
INIT_0F => X"A4160600349075238473F1210006133835E92273612B3482C090068A0E84AC56",
INIT_10 => X"30060181BA1B13959DC08DA902458870201970B29602562B0581200D141D0959",
INIT_11 => X"E042021C040D0152C8058B3840F044708E7E1C20A0106EA166C13AFC14AA3804",
INIT_12 => X"080E004B0C17C1439A9838301DC1A8438EA32C009DC1A8255300650458A1D588",
INIT_13 => X"018010E186F110A908E3A8CB0026C9A610A908E6A60F0807626610E160589C4C",
INIT_14 => X"2A701667334005800B1605F043858125E0D04110408D2485CA034681E43A1E40",
INIT_15 => X"00646002304244A91102C93A2D608D2A258DF8034188200C050171A41108F084",
INIT_16 => X"110441104411044110441104411044110466C440446CA06951D4EA8010009804",
INIT_17 => X"0040100401004411044110441104411044110441104411044110441104411044",
INIT_18 => X"0401004010040100401004010040100401004010040100401004010040100401",
INIT_19 => X"F7DFBFDEFE8FF1F7DEBDDF7DF7D05122890000000003FFFFFFFF900401004010",
INIT_1A => X"9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7BFFDFD7DDDF7DF7D",
INIT_1B => X"F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE79E7",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000003F9FCFE7F3F9FCFE7F3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA000400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0800",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000002000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2A954BA000015400FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080402010FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2A954BA0004154BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A0004174BAFFFFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0800154AAFFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF552A974AA0000174BAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974A",
INIT_2E => X"000007FFFFFFFFFFFFFFFFFFFFFFEF552E974BA0804000AAA2FFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080400010000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E954AA080005000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000402010FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2A954BA000417410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"804154BAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974BA0000174AAFFFFFFFFFFF",
INIT_34 => X"FFFFFFFEF552A974AA0000104AAE3FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0",
INIT_35 => X"AA2FFFFFFFFFFFFFFFFFFFFFFFEF552E954BA000E124BAE3FFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000007FFFFFFFFFFFFFFFFFFFFDFEF552E954BA080A000A",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804000100000000000000000000000000",
INIT_38 => X"54AA000400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2A954AA080017410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"0174BAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A954BA000415400FFFFFFFFFFFFF",
INIT_3B => X"FFFDFEF552E974AA0804174AAF7FFFFFFFFFFFFFFFFFFFFFFFEF552A974BA000",
INIT_3C => X"2FFFFFFFFFFFFFFFFFFFFFDFEF552E954AA0004000AAA2FFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2A954BA082E800AAAAFFFFFFFFFFFFFFFFFFFBFDFEF5D2E954BA002A820BAA",
INIT_3E => X"0000000000000000000000000000000000000087FFFFFFFFFFFFFFFF7FBFDFEF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(2),               -- Port A write enable input
DIA(0)   => data_write_a(22),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(22),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(2),               -- Port B write enable input
DIB(0)   => data_write_b(22),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(22),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_23_10 : RAMB16_S1_S1
generic map (
INIT_00 => X"EF20906D902424807BC8241BC81801B97D38AD3C0800103362A6741C80A12A02",
INIT_01 => X"001FFF8409F089003B4422000D80C80106804A7951C5B9D1C828043EA28838F9",
INIT_02 => X"E01CEE21649C82C40800000F9FFEFF8E72CA7F5FC2E22809925A0D3611C877F8",
INIT_03 => X"24000400402670400402670D48222DC1764446838624000080007460C40001BF",
INIT_04 => X"68403FFC020560E0443E21037C01FFFC0002EE00628BF0E02FAD781014085014",
INIT_05 => X"0112000202FBFFF00920017FF0F0628BFF8488890979800002F702002BB807A0",
INIT_06 => X"EF85788B681FC000000001FFF0010000000001F7CBC385F87C0BFFFF20040001",
INIT_07 => X"F6E200000000C1440E3AE408009120071070FA07A1CB23FFA403F0C4D23BF7C0",
INIT_08 => X"0BF87CA400804000003FF7FFD8880A034AC09662305AB10555421006891A1089",
INIT_09 => X"BE1F5FEA10092C0896A243FFC0008087FFBEF2000000001DFFC612C0C0400100",
INIT_0A => X"41FF0C2060501000600000000001BFFA800808189A657EF81DD0C00079CC8001",
INIT_0B => X"018C24110A860006C620C0312241C482B20400CC52492710CC80060020A81BFE",
INIT_0C => X"0C08866907048320C20C10030400C10030400C10030400C10030400608018210",
INIT_0D => X"040002000041500300100040000500C000801000C02400000952800001FFBF04",
INIT_0E => X"FC850015385380380CDB86106502C5043FFD5FFF00A04BC010A7724B10000800",
INIT_0F => X"89F90A002A70A710A51C01C05904014861433602A1CAF13F2110055614C72FC0",
INIT_10 => X"E02D02001C1E14981B43253EE50C8220180F1082E06397E07E42200AAC298E57",
INIT_11 => X"8421802400A90022B0070FAE18019214A380344920080B21A58B02AC60BACDF0",
INIT_12 => X"0A2A000C480B0704B54028101AC49C84BB4100009AC49C80857A82D20CE8CB22",
INIT_13 => X"01E00C8103416445C12ED0400027C5292445C12D500B0005A62D344CB241D095",
INIT_14 => X"132C907425604680038706A35132C94BDD011010404428886AC91B11311C8280",
INIT_15 => X"FF000470BE0692020328CA0028042054A92771C50FC070110001C1680809591D",
INIT_16 => X"00802008020080200802008020080200800800200200000000000008004807DF",
INIT_17 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_18 => X"8020080200802008020080200802008020080200802008020080200802008020",
INIT_19 => X"0000000000000000000000000000000000000000000000000000008020080200",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080002010FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974AA000400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000400010FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974AA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080000010FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E954AA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954A",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA000015400FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080002010FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974AA000400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000402010FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E954AA080005000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA080407000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA00041741",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080000010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000402010FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2A954AA080002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954AA080017410FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"552A954BA000415400F7FFFFFFFFFFFFFFFFFFFFFFFFF552A954BA080015410F",
INIT_3E => X"0000000000000000000000000000000000000F7FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(2),               -- Port A write enable input
DIA(0)   => data_write_a(23),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(23),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(2),               -- Port B write enable input
DIB(0)   => data_write_b(23),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(23),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_24_10 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100600007FFF000080108004000800020000840041000080808",
INIT_02 => X"FC5CA803400EB8209000000F9FFEFF8E7240FF1FC22409EA04018E50074017F0",
INIT_03 => X"11100400000000400000000D00002CC07400000090C080019001010A000001BF",
INIT_04 => X"68003FFC00040000000000008001FFFC0002EE00000370E007A100000000E468",
INIT_05 => X"0000000000F8BFF00920004DF0F00001DF8000000079800000F3000029980780",
INIT_06 => X"6E461803081FC000000001FFF0000000000001F7C3C380F87C019FFF00000000",
INIT_07 => X"600C2400013649609C8000980040814210254000A00B21FF2003F2A80D500000",
INIT_08 => X"0BF80000000000000003F7FFD88D2B4A02C0940062EC2804001610020408178B",
INIT_09 => X"8E1F5FE010092C0892A041FFC0000001FFBEF0000000001DFFC002C000000000",
INIT_0A => X"41FF0C0000000000600000000001BFFA0000005501AA00000CE2000009400000",
INIT_0B => X"018C0411020600048620C030020502000200000400490510CC00040020201BF4",
INIT_0C => X"0808064106040300C00C10030400C10030400C10030400C10030400608018210",
INIT_0D => X"0000000000004003000000000000001200580000000000000000000001FFBE00",
INIT_0E => X"0086C022005381380FDB96516140C6043FFD5BFF000041000000004110000000",
INIT_0F => X"80010D804400A7240C840C201D0210840043B4804012500021E0088014C04940",
INIT_10 => X"4109038041021C980200D06410C1924030008142E06024A00043C01100298092",
INIT_11 => X"587CC200002100C14428090A1D02348190814C09C010104025AA40041A0D8005",
INIT_12 => X"022E0030300B0E46177004208000D8C61D7004300000D884817B00011306B2D9",
INIT_13 => X"01E003060344710009875C018100013831000985DC000C20003C310006143B70",
INIT_14 => X"4001850EDC004780144806A64400186CBF8961104000C3807884000846EB9500",
INIT_15 => X"FF0006E08C063C0220002201490418082010A57263E0100008000290161E711C",
INIT_16 => X"00000000000000000000000000000000000000000000000000000000000007DF",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"F2D0AEEAF6E7CC1132CDB4441990000000000000000000000000000000000000",
INIT_1A => X"BEFBE79E79E79E79E79EFBEFBEFBEFBEFBEF9EF9EF9EF9EFA69861219575D75F",
INIT_1B => X"783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1EFBEF",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000783C1E0F0783C1E0F0",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0201000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A000400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA000400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000400000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402010000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"00002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080002010FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000400010FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA00040000",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020100000000000000000000000000",
INIT_38 => X"74BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"000010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA000002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974AA000402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000002010F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(3),               -- Port A write enable input
DIA(0)   => data_write_a(24),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(24),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(3),               -- Port B write enable input
DIB(0)   => data_write_b(24),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(24),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_25_10 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100200002000000080100004000000020000800041000080808",
INIT_02 => X"FC400086000000800000000F9FFEFF8E738FFF1FC204010000000111568DD7F8",
INIT_03 => X"00000400000000400000000D00002CC4740000008000000080000000000001BF",
INIT_04 => X"68003FFF64A564AC000000000001FFFE0082EF00010370E007A1000000004000",
INIT_05 => X"0A00040148F8BFF80920804DF0F00101DFC040000079C92484F30499299837C1",
INIT_06 => X"66041803081FC0E0801101FFFD000E41002299F7E3C380F87C019FFF81200096",
INIT_07 => X"000000080480AE00000080000000000000000000A00B21FF2003E00000000000",
INIT_08 => X"1BF80000400A02000003F7FFFA0008000200A0400008A0000014100200081000",
INIT_09 => X"8E1F5FFA53EFBCACB2E369FFE0010001FFBEF80C40630C7DFFEEBAF000800202",
INIT_0A => X"41FF0C0600000000600000000001BFFE00301000000000000CC020000140000C",
INIT_0B => X"01DCCC31222730A49620C030020100000200000400490D10EC00040220201BF4",
INIT_0C => X"0808064106240300C00C10030400C10030400C10030400C10030400608018210",
INIT_0D => X"0883044582114013412080000000000000000000000000000012800001FFBE00",
INIT_0E => X"00040020000180380FC386106140C6043FFD5BFF00A04B80608003CB120C1106",
INIT_0F => X"0000080040000200040400000100000000009480000240000100080000400900",
INIT_10 => X"0001000000000808000000240000020000000100006004800002001000008012",
INIT_11 => X"0001001808220000002004001900000080800008000000000022400000088000",
INIT_12 => X"0010000000000E00110000000000408009000000000040808063004000008200",
INIT_13 => X"6000000000046100000240000000001021000004400000000010210000001010",
INIT_14 => X"4000000404000800000000060400000088000001800000001084000000088000",
INIT_15 => X"FF800C608C041002000002000006100000002100000000180600000000100018",
INIT_16 => X"4110441104411044110441104411044510629041040D180400000010028047DF",
INIT_17 => X"1104411044110441104411044110441104411044110441104411044110441104",
INIT_18 => X"1044110441104411044110441104411044110441104411044110441104411044",
INIT_19 => X"FBA2894A196A8C5A2932EC15DA080800002FFFFFFFFFFFFFFFFFC11044110441",
INIT_1A => X"2492492492492492492410410410410410410492410492412000531215A69A6B",
INIT_1B => X"158AC562B158AC562B158AC562B158AC562B1588C46231188C46231188C49249",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000B158AC562B158AC562B",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080000010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000010FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08000000",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(3),               -- Port A write enable input
DIA(0)   => data_write_a(25),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(25),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(3),               -- Port B write enable input
DIB(0)   => data_write_b(25),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(25),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_26_10 : RAMB16_S1_S1
generic map (
INIT_00 => X"E9264EAB20190CA3BA4997AA9002AE9C001006B0778015CFA17E0811039879C7",
INIT_01 => X"2FFFF9BB1F773C7F9BB07DFFFDD863FC5FFF3FEFFBBF9FFB22FFFBC7B9F30686",
INIT_02 => X"E06CCC62052E708180F6FFBFFFFCFFFFF9C7FF7FC24332E642090000074037F6",
INIT_03 => X"428003739CD9863739CD9869FE2B7DEAF300029E4E300DFE69A6E644E6FF473F",
INIT_04 => X"7C2FEFFFF5BA124F003DD31EAFFFFFEE9FF7EE6F4C0770FFD7DC7CA53997B2B1",
INIT_05 => X"DFFB5421C1F8BBFAFDBFFACDF0FFCC05DDDBFF3690F9EDB7F5F7AFF639BD7DE3",
INIT_06 => X"EFD044ABC817C3E3A74667FDFFB6FF5727CC3BFEF7C3FAF87FF59F7FFBFEF69F",
INIT_07 => X"00003002132462052E708180EF060C18E5BEFB051225CDFF7002C4EEDE77F6E0",
INIT_08 => X"3FFF7D5000EC75088ED3FF7FC8790E46426CE06CB1F8E041051831FA3068D77E",
INIT_09 => X"C05FD7FF9BEFBDCEFBEE59FEF44F6603EFBEFAFCC2E35E7FDFD147CCF3F583FA",
INIT_0A => X"67FF1C7FBFADEB31E35768E8ED6BFDF3EB3EBF9DDBCE7FDC1DF8A760F3EACC02",
INIT_0B => X"5BDDCC3B336F7C548667D47B7737AF3FD62601EDC25B3533DCEB07F262213FFC",
INIT_0C => X"5F9A06E19F4D93A0EA0F78C35E30D78C35E30D78C35E30D78C35E986BC61AE31",
INIT_0D => X"5FD7AFEFDFFAF59B6FF28FE1D80D73D840607307DCFE1D80EF69A004DFFFF7FF",
INIT_0E => X"0004001F8041897B2FFFC6D86D70CE04FFFFF3FF1F5F5475BD7F72E4D75EBFAF",
INIT_0F => X"F60008003F008237B0040A00010003E020023E0201F45EC0010007E01047D17B",
INIT_10 => X"00010001DC0004C81003DE050A700200001DC0006863E8BD8002000FC0208FA2",
INIT_11 => X"2200E400002801E1A00004C21C0206F60081800800007B00010F02007EC09A0E",
INIT_12 => X"0880007E000807C7C1A612001E0015C7C19C22001E0015C59DFE82011A311AA0",
INIT_13 => X"00001BC00101F60409F0670840070809760409F06984800780097604067D0010",
INIT_14 => X"81019F40042100001F800203D81019EC085614000085C80023D81009CF008A74",
INIT_15 => X"FF802FFDFFAFD082003B032FB987E04021D481D4000819060801E0D00001231D",
INIT_16 => X"EBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEFFBFBFBFBBFCFBB0FFDFEFFEF2DFFFFFB",
INIT_17 => X"BFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAF",
INIT_18 => X"FAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFE",
INIT_19 => X"475B15BCF491E166CC8553F86EDB5C88646FFFFFFFFFFFFFFFFFEBFAFEBFAFEB",
INIT_1A => X"861861861861861861861861861861861861869A69A61861AFBD54D5F871C71D",
INIT_1B => X"984C26130984C26130984C26130984C26130984C26130984C26130984C261861",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000984C26130984C26130",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040201",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(3),               -- Port A write enable input
DIA(0)   => data_write_a(26),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(26),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(3),               -- Port B write enable input
DIB(0)   => data_write_b(26),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(26),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_27_10 : RAMB16_S1_S1
generic map (
INIT_00 => X"00080A40000A41248002029000050A088000008242A0004404480002000A1155",
INIT_01 => X"2FFFF1C11F781C129C107DFFFE0860941E81258CA2B71C2220EC1B86E1A00002",
INIT_02 => X"E1000000810000014400FF6FFFF0FFFFF8007F1FC21110005080200000221FF0",
INIT_03 => X"4080026318C18226318C1821302232EAE00002BE001115FE48620040840A863F",
INIT_04 => X"643D4FFC2530000F003D821C0BFFFF8E9EF79E6D440748FED70060842105B0B0",
INIT_05 => X"D6F39020D1F8A3FAFDBFBACDC8FDC405D1DB7F1490E5EDB7D5CBADB2385D79C3",
INIT_06 => X"6FE000A38007C3032646EFF1F0B6FF46A78C39F8E723F2E47FE59C7F9ADA2612",
INIT_07 => X"00002820000000810000014401060C180190310540118DFF1000C0849673F6C0",
INIT_08 => X"3FF779100062B12A8EC3F47FC80208808210880C00082050000110023068D030",
INIT_09 => X"005F07E09BFFBD07FBAC09F8E42922038F7DF8BEC2E39C5F1FD047CEF1B582D8",
INIT_0A => X"63FF5D5F9FADE911E81C09818109E1F16B16B71092CE7ED81CF403601228C402",
INIT_0B => X"1BFDCC39732F3554866AD57C37BEAF1C152201A4C05B7531D56B05B06A213FF8",
INIT_0C => X"5BCA06F18FC59380F00E34430D10C34430D10C34430D10C34430F0861A2186B5",
INIT_0D => X"5B56ADAB5FAAE58B2F628EA0C80FA3F04040510768EA0C80CC61A0044DFFC6EB",
INIT_0E => X"0004001D800188792CE79715710AE4047FFD23FF315D54358D593474955AB6AD",
INIT_0F => X"520008003B000297B0040200010003E020001F0201E44A400100076000579129",
INIT_10 => X"00010001DC00004A10035E0408300200001DC000086BC8948002000EC000AF22",
INIT_11 => X"02002400002801E1A00000C01E0202F60080800800007B00000782006EC0820A",
INIT_12 => X"0080007E000006A7C10602001E0001A7C10C02001E0001C18DE282010A311AA0",
INIT_13 => X"00001BC00000FE0401F04300400708007E0401F04180800780007E04047D0010",
INIT_14 => X"81011F40040100001F800002F81011EC080604000085C80001F810094F008034",
INIT_15 => X"FF800C6DDDAFD082001B03249887E04001D481D4000009020801E0D00001021F",
INIT_16 => X"AB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6BF1EBDABD8E270BF84A25C6ACB777E3",
INIT_17 => X"B6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6AD",
INIT_18 => X"6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADA",
INIT_19 => X"490E2168100481CA860402104A471688747FFFFFFFFFFFFFFFFFAB6ADAB6ADAB",
INIT_1A => X"000000000000000000000000000000000008200000000000200072F210000001",
INIT_1B => X"05028140A05028140A05028140A05028140A0500804020100804020100800000",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000A05028140A05028140A",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040201",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(3),               -- Port A write enable input
DIA(0)   => data_write_a(27),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(27),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(3),               -- Port B write enable input
DIB(0)   => data_write_b(27),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(27),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_28_10 : RAMB16_S1_S1
generic map (
INIT_00 => X"02200AA400180030808802A900002A08001280A08A801044104A1000001818C3",
INIT_01 => X"0AA00011460214428114180000882214413D0A71592A01D92213D28005210202",
INIT_02 => X"0451110A012100884000AA30200000000C100040104112101100008888200000",
INIT_03 => X"448000318C52A20318C52A20148810200111100C211004AA00034204200A2200",
INIT_04 => X"04004001001A90110000121402AA0000003C00000500000040080421080D0080",
INIT_05 => X"4060000C8001000000002E000000050000001610300000010000802202040012",
INIT_06 => X"1000002080001111001222000425A1040026A008000000000000000009328280",
INIT_07 => X"2491008A00491201210088400122448908A20402000408001000040820000000",
INIT_08 => X"20058310402A160026500000028040101004200C840082115554000112244814",
INIT_09 => X"4140000800000060000720000102028000000490160801020002200011100010",
INIT_0A => X"020000081B34211082B694D4D294000020020381040000000200032040004400",
INIT_0B => X"4800210C19808400500010009110091500020B408810000100200020408B0000",
INIT_0C => X"01028000080118020023604858121604858121604858121604858090B0242C00",
INIT_0D => X"010000800920040804020A6058003108402043058C460580653020005A004039",
INIT_0E => X"00000002800008014004104104420A00C000200005000010040A0020CC000200",
INIT_0F => X"520000000500000010000200000000000000280000040A40000000A000001029",
INIT_10 => X"00000000000000C0000002000830000000000000480008148000000140000020",
INIT_11 => X"020024000000000000000440000000020000800000000000000C00000040020A",
INIT_12 => X"00800000000001804006020000000500400C0200000005400A90000000100000",
INIT_13 => X"0000000000018200001003004000000142000010018080000001420000200000",
INIT_14 => X"8000080000010000000000018800008000060400000000000310000008000034",
INIT_15 => X"000002040080000000110006B081400000400000000009020000000000002200",
INIT_16 => X"802008020080200802008020080200802101210810C39A66A90A85420413A820",
INIT_17 => X"0200802008020080200802008020080200802008020080200802008020080200",
INIT_18 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_19 => X"DE21102C110A00246972BD89A40A0C22E1000000000000000000002008020080",
INIT_1A => X"2082082082082082082082082082082082082082082082080D35050758C30C31",
INIT_1B => X"0582C160B0582C160B0582C160B0582C160B0580C06030180C06030180C08208",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000B0582C160B0582C160B",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(3),               -- Port A write enable input
DIA(0)   => data_write_a(28),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(28),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(3),               -- Port B write enable input
DIB(0)   => data_write_b(28),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(28),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_29_10 : RAMB16_S1_S1
generic map (
INIT_00 => X"79964E4BA01DACAB9E659792D00AAE160002829C7FDFEFCEE97C2815039D70C3",
INIT_01 => X"0ABFF9AB0775343F9AB01DF80D5821FC0FFF3FEFD1AF9FF1207FFBC7B9720586",
INIT_02 => X"002CCC60050E700080F6AAA7BFFC007189C7FF2FC00330E602800000074037F6",
INIT_03 => X"468003210868A63210868A68DA017D207200021C4E200CAA6186A40042FF4300",
INIT_04 => X"7C2FE002F0900001003C5316A6ABFFE21F36E02F0D03701F47D41800109FB281",
INIT_05 => X"4979440580F9B808F49F6A4DF00F8D01DC4B97369078249370F482E62BA41462",
INIT_06 => X"B250442BC81001E1870223FC0BF7F11507C423FE33C078F803F19F00E936721D",
INIT_07 => X"00011080012460050E700080EF020408EC8CFA01122149FF700200665A35D260",
INIT_08 => X"2BFD055040A452000443FF00007906464068406C31F84000000831FA1028575A",
INIT_09 => X"805FD017102690AA694551FE30444681E0820AD40201423FC00122C493500172",
INIT_0A => X"0600002AFFBE2330815568A8AD6ABC02A02A0B0CCB463B4C0748A720B1EA4C00",
INIT_0B => X"0850400A11414C005005000B51158936D20601A98A10200308A002E240010BFC",
INIT_0C => X"05928020194918A22A2268C81A32068C81A32068C81A32068C81A99034640C00",
INIT_0D => X"058102C48970541944B20FA1580561D040406305587A158046282000DBFFF13D",
INIT_0E => X"000000028040890327DCD28928324400DFFFF0001F1F0050342D42A086040B02",
INIT_0F => X"F60000000500802010000A000000000000022A0000141EC0000000A01000507B",
INIT_10 => X"00000000000004C0000082010A700000000000006800283D80000001402000A0",
INIT_11 => X"2200E4000000000000000442040004020001800000000000010D000010401A0E",
INIT_12 => X"08800000000801C040A6120000001540409C2200000015441DAC800010100000",
INIT_13 => X"0000000001019600081027084000000956000810298480000009560002200000",
INIT_14 => X"800088000021000000000201D800088000561400000000002358000088000A74",
INIT_15 => X"00802594A282C0000033010FB181E00020400000000819060000000000002305",
INIT_16 => X"C0B02C0B02C0B02C0B02C0B02C0B02C4B12B312912831A27FCFE7FFB175B6FF8",
INIT_17 => X"0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02",
INIT_18 => X"B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C",
INIT_19 => X"BBCF9F96EE7FFDF7FE783FFDFFEA0C00602FFFFFFFFFFFFFFFFFC0B02C0B02C0",
INIT_1A => X"EFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEEBAEBAEBAEBAEBBFFDF9FBEFFFFFFE",
INIT_1B => X"BFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFBEFB",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000FBFDFEFF7FBFDFEFF7F",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(3),               -- Port A write enable input
DIA(0)   => data_write_a(29),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(29),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(3),               -- Port B write enable input
DIB(0)   => data_write_b(29),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(29),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_30_10 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"F7FFBFFEFF9FE1F7FFBFFFFDFFD0000000000000000000000000000000000000",
INIT_1A => X"9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7AFBD75F5FDF7DF7F",
INIT_1B => X"F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE79E7",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000003F9FCFE7F3F9FCFE7F3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(3),               -- Port A write enable input
DIA(0)   => data_write_a(30),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(30),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(3),               -- Port B write enable input
DIB(0)   => data_write_b(30),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(30),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_31_10 : RAMB16_S1_S1
generic map (
INIT_00 => X"129000008004A00804A40000400800020000000C005FEA005800200400050100",
INIT_01 => X"255FF18019700810180065FFFC0040801E80258CA2951C2200EC0906A0804140",
INIT_02 => X"E0000000000000011000550FDFF0FFFFF0007F1FC200000044000000000817F0",
INIT_03 => X"0000024210A30024210A3001002220C06044469200040154482000408400043F",
INIT_04 => X"602D0FFC2420000E003D80080955FF8E1ECA8E2D400340FE870060842100B030",
INIT_05 => X"0213100040F8A3F8FDBF944DC0FDC001D1CB6904A061EDB6D4C30490281831C1",
INIT_06 => X"6FC000830007C202060445F1F0D25E4207A099F0E303F0E07FE19C7F80402412",
INIT_07 => X"0000200000000000000001100004081001103107000185FF0000C0849673F6C0",
INIT_08 => X"1BF27A00000000000883F47FC800080002008000000820440000100220489020",
INIT_09 => X"011F07E013EFBC06FBA009F8E00120038F3CF82C44630C5D1FC002CCE0808248",
INIT_0A => X"61FF0C06C48BC801600000000001A1F00110101092CE7ED81CF0004012288000",
INIT_0B => X"11DCCC31222730048620C4382204A608142002A440492530C401049020221BF8",
INIT_0C => X"0888066187448380E00C10030400C10030400C10030400C10030600608018210",
INIT_0D => X"080204010200418301208480800D02D00040100240A808008840800405FF8640",
INIT_0E => X"0004001D000180780CE386106100C4043FFD03FF101D40008001304018081004",
INIT_0F => X"000008003A000217A0040000010003E02000160201E040000100074000478100",
INIT_10 => X"00010001DC00000810035C0400000200001DC0000063C0800002000E80008F02",
INIT_11 => X"00000000002801E1A00000801C0202F40080000800007B00000302006E808000",
INIT_12 => X"0000007E00000607810000001E000087810000001E000081846282010A211AA0",
INIT_13 => X"00001BC00000740401E0400000070800340401E04000000780003404045D0010",
INIT_14 => X"01011740040000001F8000025010116C080000000085C80000C8100947008000",
INIT_15 => X"FF800C609C06D082000A03200806A040019481D4000000000801E0D00001001D",
INIT_16 => X"010040100401004010040100401004010060C040040C200950402090128057C3",
INIT_17 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_18 => X"0040100401004010040100401004010040100401004010040100401004010040",
INIT_19 => X"00000000000000000000000000001000802FFFFFFFFFFFFFFFFF810040100401",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(3),               -- Port A write enable input
DIA(0)   => data_write_a(31),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(31),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(3),               -- Port B write enable input
DIB(0)   => data_write_b(31),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(31),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_0_9 : RAMB16_S1_S1
generic map (
INIT_00 => X"ED39BA795990D275FB4A6E96ACC4731DEA4598B0AFB54867F6EE4618C3749803",
INIT_01 => X"8AA0047D8607944AC7DA180001ECA2444042106208408208C20022E9173734B3",
INIT_02 => X"1A7DDD79F9A73E6CCA7DAAF00001000008478020113D98E382FEDF333027C80F",
INIT_03 => X"75D341110C58F31110C58F32A208921F8051500147A0E4AB3493FB3A01EBE240",
INIT_04 => X"86424001531009B100425A97B2AA0001E03501D0A39C8F0078420001106D0C4C",
INIT_05 => X"BCC8CA2EBF03400700402BB20F00239E20341699198600000B08694B16434804",
INIT_06 => X"103FB860B2800161F8432200012DA185F80F24081C3C0707800E600056881308",
INIT_07 => X"B24197ABCDA467F9A73E6CCAFDC3870EEEEC44E2BDFE220094D03022210C011C",
INIT_08 => X"240581B5695EAA80262C080032BF07C7C1FC3F8E94F65B11555EAFFC1C306758",
INIT_09 => X"7E40000BEC004170040DB60017FED1CC0001045002984202003DB931192D60A5",
INIT_0A => X"120071411A74315881A28C141118000C5A85A60444210123820B43B40804674D",
INIT_0B => X"0820008E514045BB514F0106D1D8599581D3A958BC104A89215AC14C48898403",
INIT_0C => X"C261C01C48B1584A0CA3E2687A9A1E2687A9A1E2687A9A1E26870CD061343885",
INIT_0D => X"D274E93A758FA8683AC54B287522E10A74AF4AA59C568752662F5AC218000002",
INIT_0E => X"FF83C002783A0904231C70470C7E0B92800224008AE09FAD4BD48D1FC5D3A4E9",
INIT_0F => X"5BFF078004F075885DFBF7E15C06101C55E921F1F80FAB7FE0F0009E0E903EAD",
INIT_10 => X"F12E0380231F13978FF023FAFDBD9870380230F2D6081F56FFC1E0013C1D207D",
INIT_11 => X"DE7F263C0C8700125C0F8F3C43F1F10BBF7EFC61E01804E1E6C8F8FE807F67FB",
INIT_12 => X"02BE00017C17C1007E5E2E3081C5AC007E6F0E3081C5AC44418D65FE45DEE55B",
INIT_13 => X"61E0042786F103E9F01F9BC3C120C5A703E9F01F978B8C20666703E9F8A0FFED",
INIT_14 => X"FA7E283FFB414F80005F05F10FA7E283F78F6511C048278DCA174FF038FF15B4",
INIT_15 => X"0066A20B61692F293185D8D724E15D3FCC6B7C236FE0691B0700132C1F0EF880",
INIT_16 => X"3A4E93A4E93A4E93A4E93A4E93A4E93A4F942F92E9628540AD2A91442525A000",
INIT_17 => X"A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E9",
INIT_18 => X"4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93",
INIT_19 => X"55F3898E09B56C74DAB15D1CF13501AA495000000000000000003A4E93A4E93A",
INIT_1A => X"082082082082082082082082082082082082082082082082082084E41DC71C71",
INIT_1B => X"E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F82082",
INIT_1C => X"FFFFFFFFFFFFFFF94A5294A5294A5294A5294A52800003E1F0F87C3E1F0F87C3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"3060C183060C187FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"BDEBA0000000000000000000000000000000000000000000003060C183060C18",
INIT_28 => X"168ABA002E82145085155545F7AA975EFFFAABDE00FFAEBDFFF5D2EAAAAAF7AE",
INIT_29 => X"7FFFE10005542145557FD5545FF8000155087FC0155F7D168B55007BFDF45085",
INIT_2A => X"7FFC0010080017555555568AAAFFFFD7545AA8028A00A2802AABAFF8028BEF5D",
INIT_2B => X"FF842AABAA2AE95545FFD168ABAF7AEAAAAAA2FFFDF4500043FE105D2E954BAF",
INIT_2C => X"5007FD7400550415410002E974BA5D5168A00A2D142155005142010FFAE820AA",
INIT_2D => X"FFF780000BA007FE8AAAFF803FFFF5D2A821550000000BA007FD55FF5D7FC014",
INIT_2E => X"000AAFBEAA00007BFDFFF082EBDF455D5142000082E82145FFD17DFEFFFD168B",
INIT_2F => X"DFD75D2AA8A80EA8E2FE3F000000000000000000000000000000000000000000",
INIT_30 => X"68B551475FAF6D1C556F0AA1C24AABEA495FC716F002A975FFE3AA95E00EBAEB",
INIT_31 => X"42A0070071C50BAFEF1FAE0016D56A16D557BC257D415E0216FA3F1E8FC0145B",
INIT_32 => X"8010E004924874825D7FEAA85487FD24AFE3D02DAAAE12BD5545A2803AA00005",
INIT_33 => X"120155EA568E870BAEB8A05A2AEA8B50F55A2F150005A3A438BD04AFAB8F550A",
INIT_34 => X"545E055FFBE81D0BE8EA8A3AA05A2A5504001C74BA42A1571E8028E3DB7816D0",
INIT_35 => X"A5C7E3DFFFE90B45B47ABA497A82FFAFD2A82485FD2415A105C21451ED42A002",
INIT_36 => X"00000000000000000000B55EAAA100AA1D0F6F480B6A555A2A57A002A3D5FDB6",
INIT_37 => X"5EFAAAAB5E1AF3AABFF45592E88A0AFE80A8B0A0000000000000000000000000",
INIT_38 => X"65F520EBE9EF67D7BEA1FD5D556ABEF5D557FEBA55022A3F70C6B405F4D2AE97",
INIT_39 => X"C114728007521170821CE0FDE69411A8DED57CE1055555E5F58EFFC01FE2CACB",
INIT_3A => X"42341D5DEEBEF55080034E0A592A4AD0079C75D6070CC5CBB0280C029ABAA3EB",
INIT_3B => X"7F353AAF6C77F7F20D968BF57812A95E02A2AAB5EB0F280800EFAEE9F5D18F31",
INIT_3C => X"C91565455C141E41887D58AC448B69C30E02116220415A9540AA854140A0A204",
INIT_3D => X"DE6BE93172D7D625B556EEAB157ABEBE1B4D792A4AD1183454180DD3FDCAAAB7",
INIT_3E => X"F0000001FF0000001FF0000001FF0000001FF01EABC4B8014174FF7DA80F52FE",
INIT_3F => X"FF0000001FF0000001FF0000001FF0000001FF0000001FF0000001FF0000001F")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(0),               -- Port A write enable input
DIA(0)   => data_write_a(0),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(0),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(0),               -- Port B write enable input
DIB(0)   => data_write_b(0),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(0),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_1_9 : RAMB16_S1_S1
generic map (
INIT_00 => X"212C001411984004084D000508C53810A03D1450E839B003342114428A000803",
INIT_01 => X"00000019400B100A8196000000CC004400400002000000000000028001340000",
INIT_02 => X"052137AE8031800C0044009000000000061800001CD4019802AD04CCCFC20004",
INIT_03 => X"04514108C60C21008C6042108400000201440020505100000043C30E10E9F000",
INIT_04 => X"02104001011DEFE088805681920000008000004001900800004002108C280008",
INIT_05 => X"040002340105000200000000080001900010000108040000000008411600401C",
INIT_06 => X"1034001042800808201000000001000820020000102000040000000000800180",
INIT_07 => X"64BF81A15EDFDE8031800C00843060C19E030022103600000450020800040004",
INIT_08 => X"00008004691687AA840008000090248CC84E000046000311555521F183060AC5",
INIT_09 => X"0820800D08100171000DB000154440C800400500000852020011200201012021",
INIT_0A => X"02000040001000880A2A04445004000102002041000001008208001440004140",
INIT_0B => X"4820018A1140440078050040511000102000A008183000010002404400000000",
INIT_0C => X"1000C80008000C030030880C2A030A00C28030A80C2A030A00C28018D4061401",
INIT_0D => X"10040802050080200284401C0022880F009E08008205C0020118088018000000",
INIT_0E => X"0F03C00280000000420860C60C0C0B92C0000000004000010042000040102008",
INIT_0F => X"001E078005000108400005E11C0610000000288058000003C0F000A000100000",
INIT_10 => X"F10E0380000000C202300000008D187038000000480800000781E00140002000",
INIT_11 => X"806302380C870010000004400100110800007861E0180000000C400680000001",
INIT_12 => X"023E00000000018000580C308000050000610C30800005000215006800000101",
INIT_13 => X"61E0000000018100B0001843812000014100B00016030C20000141002880026D",
INIT_14 => X"400A20009B404F80000000018400A20044096111C04000000304026000501580",
INIT_15 => X"0046820040082300218450C2800010094000482141E060190700100000002200",
INIT_16 => X"020080200802008020080200802008020080008008600500A82A1100A8000000",
INIT_17 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_18 => X"0080200802008020080200802008020080200802008020080200802008020080",
INIT_19 => X"81328A46BABEFC54A0810C7452B4428A14000000000000000000020080200802",
INIT_1A => X"AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA28A28A28A28A2A8218D2C0C924925",
INIT_1B => X"E974BA5D2E974BA5D2E974BA5D2E974BA5D2E975BADD6EB75BADD6EB75BAAAAA",
INIT_1C => X"FFFFFFFFFFFFFFFD8C6318C6318C6318C6318C63000002E974BA5D2E974BA5D2",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"70E1C3870E1C387FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"5555500000000000000000000000000000000000000000000070E1C3870E1C38",
INIT_28 => X"EBDF455D2EAABEFF7FFE8BFF5D0002155557FFFFFF007FC21EFA2FFD74AAAAD5",
INIT_29 => X"AA95400552AAAABAFFD1574105D7FD75FFAAAA800AAF7AA974BAFFFBE8B45F7A",
INIT_2A => X"0517DF555D2EAAA1055000015500557DF45AAD1400BAA2AE801550051555EFF7",
INIT_2B => X"FFD540155557FD5400F78028BFFFFFBEAB55F780020AAAA80020AA082EAAB550",
INIT_2C => X"AFF842ABEF5D517DF55552A974AAF7AE820AA0851574BAA2D1574AA5D7BFDEBA",
INIT_2D => X"EFAAD1575EF557FFFE10557FFFFFFFFD56AAAAFFFFD7555AAD168B45AAAEAAAB",
INIT_2E => X"0005D7FFDF4500043FE105D2E954BAF7AE80010082A97410557FEABFFAAFBE8B",
INIT_2F => X"51C7A2FBD5490BFD1C056A000000000000000000000000000000000000000000",
INIT_30 => X"974BAF7FFEFB45FFAABDF55492AA8BC2EBDFEAF7F1F840017D4975D2FEF147FC",
INIT_31 => X"080BEF495FC71D54124924385FAAA8AAAE3D145410F7F1D55D71C002DABAEBAA",
INIT_32 => X"002D082082AB8B6DBEDB7DF7F540E2AE85028B40155145F7AF6DBED5450AA1C2",
INIT_33 => X"78E021FF1471FDEAAFFD56F16D5571D2E28E38E0216FA2D1E8E80140F45082B4",
INIT_34 => X"A2DA3FB7DAAD4AAAAF487BC70BFA97F7AF6D417E92482BF84020BA495557E3FF",
INIT_35 => X"55554ADBD7A2FFC7BEFF6FFD7FC7002FD74951D71EDFFABFD16FAAAE92BD5545",
INIT_36 => X"00000000000000000000547AB8F550A8010E00492487482FFFE82A85EBAE2FFC",
INIT_37 => X"1EF005162BEF047FD5545AAFBF7400FBF9424F70000000000000000000000000",
INIT_38 => X"714F8338AAAA1D0AE974AAF7FFFDF55F7AABFF55082CA8B4DF6C1E8F5E540002",
INIT_39 => X"EABEF75550ACBB7582225FF5843404547184164AA5D2EBEEB0A2D555410D3555",
INIT_3A => X"FEAAEB083BC1000FF8409000512AEABFFDF79DCBF755962010BDCBBC21455D7F",
INIT_3B => X"801F8BA0C57740BDAA0688E5405D57D412F7D55F5E50C7F401BAAE8403CF5A3F",
INIT_3C => X"5D16BABAA3EBC3157ABD5FFE55F2AA9FEAFDF7F431A9F7FFE81FF013A8001AFF",
INIT_3D => X"FB863550229BCABEB7DA403FFFDA2FBF7FED2C7F955445079E280A00C56145EF",
INIT_3E => X"0000000000000000000000000000000000000596EBEF55080034E0A592A4AD00",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(0),               -- Port A write enable input
DIA(0)   => data_write_a(1),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(1),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(0),               -- Port B write enable input
DIB(0)   => data_write_b(1),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(1),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_2_9 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10E006600180111284380310006289800480032283E000A34301002001A0817",
INIT_01 => X"0005A00810790848048044A54E404350404000720885800802000906E4910200",
INIT_02 => X"407004208400408044C600C50AA055254010541A110222841200000002402544",
INIT_03 => X"0600011004182401004102408C28414043101000408118000145840440F5C415",
INIT_04 => X"5035855703A2900A000CD3088400F40688C9844409060850925E58A4081A0221",
INIT_05 => X"0200840D1021A15AC50494894850890540D1E12020C6E510818500440A280090",
INIT_06 => X"113044094002801020440090A8011A1224AB9380552102442884882A20004097",
INIT_07 => X"000100880004428400408044860000008C022402102100AA40004404B5075460",
INIT_08 => X"15C23440408C862A2A12382A8A5244145048C06085008010141521F000001240",
INIT_09 => X"400582B9033AA0E7AA4110B0506744810554542450694E710A836188C2C00222",
INIT_0A => X"443518360012C2210B020414109130A28038188096A06B8C120CA440A9C00802",
INIT_0B => X"1345E53300EC68005605002964AF222A5704004D080211121C80024200821780",
INIT_0C => X"181080C1110C882202211488452213C88472213C88472213488441109A442231",
INIT_0D => X"008204440210091341208041000810C00000300220201800A908000038AD0284",
INIT_0E => X"00040002804180300E88D28D206A40000554815500481440300000C44A081100",
INIT_0F => X"000008000500828700000000010000000002380000A00000010000A010050000",
INIT_10 => X"00010000000004CA000214000000020000000000684280000002000140200500",
INIT_11 => X"000000000020000000000442100002840000000800000000010C000026000000",
INIT_12 => X"00000000000805A4800000000000152300000000000015801272000100210020",
INIT_13 => X"000000000101C00000C000000000000940000120000000000009600004050000",
INIT_14 => X"0000130000000000000002018000106000000000000000002380000141000000",
INIT_15 => X"55000190000000000002000280000000011080C0000000000000000000002310",
INIT_16 => X"40902409064190641906419024090244902A9003004800415120D4A190804241",
INIT_17 => X"0900409004090641906419064190240902409024090641906419064190240902",
INIT_18 => X"9044090040900409004190441904419044090040900409004190441904419044",
INIT_19 => X"75960040138D70C030B51C50C7D100A2052F81F81F83F03F03F0419044190441",
INIT_1A => X"0410410410410410410410410410410410410410410410410248602081659659",
INIT_1B => X"5128944A25128944A25128944A25128944A25128944A25128944A25128941041",
INIT_1C => X"FFFFFFFFFFFFFFFE1084210842108421084210843FFF825128944A25128944A2",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"7FD5FF555815607FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"2AA000000000000000000000000000000000000000000000007FD5FF55581560",
INIT_28 => X"FC21EFA2FFD75EFAA8415410AA8415555087BFFF55A2AA800BAFFAE954000800",
INIT_29 => X"84155EFA2AEBDEAAA2FBEAABA5D7FE8B555551421455D0002145552EBFEBA007",
INIT_2A => X"2AEBDF555D2E954BAA2AA974BAFFFFE8B45552EBDF45FFAEAABFFF7FFE8B55F7",
INIT_2B => X"AAAAAAAAAFFD1574105D7FFFF555D2AAAAAA5D2E820BAA2FBEAB5555557DF55A",
INIT_2C => X"50055575EFFF84021555D043DEAA5D04021EF557FC21FFAA8428BFFAAAA954AA",
INIT_2D => X"10085568A00FF80175FFA2D17DFEFF7800215500557DF55AA80001FFAA800015",
INIT_2E => X"0005D00020AAAA80020AA082EAAB5500517DF555D042AA10A284154005D00154",
INIT_2F => X"00AAFFAA9543A080038A2A000000000000000000000000000000000000000000",
INIT_30 => X"0017D5D20B8EAA007FC51C7A2FBD55D2BE800042AFE8E1557D0075D2F45BEAA8",
INIT_31 => X"AA8BC7EBDFEAFEFFD00105FFBC20BDEAAA2FBF8AAA557BE8B6D5D5FFABEF4904",
INIT_32 => X"FFEFB6D555578F7DB6A0BDF7D480E174BFA02A974BAF7F5EFB455D2ABDF55492",
INIT_33 => X"ED1FDE90E3A497492B6AAADAAAE3D155E105571D55D71C002DABA5524820BAB6",
INIT_34 => X"BE8F401D7B6A0001470155C51D0092A071555D5E3AE821D00001FF0871C016DB",
INIT_35 => X"5BE8555400550A38428007FED000E3DA3DFD5E3DFFFBD5A38A021551C5F7AF6D",
INIT_36 => X"00000000000000000000410F45082B4002D082082AB8B6D1C5B7DF7FF78E075C",
INIT_37 => X"5EF005560B55F7AA800AAF7AA954AA00042AAA20000000000000000000000000",
INIT_38 => X"ABEF057D68F5F5A00021EF55042AAAA007FD5555AAFBD7545FBB8020A3F7AE97",
INIT_39 => X"7DF55D7AABFF5428ACA8F45A6C1E8F5EFF84165EFF7802BAB0A2FFEAABA557BE",
INIT_3A => X"CA8AA80800020AAF7FBFFFEF04552ABFFFF841FFE75CA882108202E974AAF7D5",
INIT_3B => X"00151FF0C57401E5F3D1E00A1A884174A8FFAEBFEB0A2D55541051555694F002",
INIT_3C => X"2AA801455D7FE8BFFF680800FFF7AAA155F595542455512A975455D3AA8A0055",
INIT_3D => X"5D79FCAF774AE005BE7895554005D2A8A0B882FFFFE10AAAAAB755A66B6AF56A",
INIT_3E => X"00000000000000000000000000000000000000C3BC1000FF8409000512AEABFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(0),               -- Port A write enable input
DIA(0)   => data_write_a(2),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(2),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(0),               -- Port B write enable input
DIB(0)   => data_write_b(2),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(2),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_3_9 : RAMB16_S1_S1
generic map (
INIT_00 => X"210C00A20020000108430020001600B8156021104940741B3530400E02B92203",
INIT_01 => X"014C9BCA58B1296D24A402C992500B69404040028804A0080A000416A8D90A08",
INIT_02 => X"C12026A484318004404405C9C66E331352180D468B8203980300204442E02B34",
INIT_03 => X"04000748D60D24648D60524C88804D0215011020D15018148040C10A70E1D58C",
INIT_04 => X"18283333240FE41244187308C9104D70944852640901083801750EB0A418C220",
INIT_05 => X"0613142D01912CC2A1B4140528348900C612A104201C689044340ED413A07649",
INIT_06 => X"119000034019881822104C5E68035250A222829710A0A02C18C01A9920842413",
INIT_07 => X"402F00AB0016CA0431800444841020509D038B021230C1990001C644C8273200",
INIT_08 => X"16905000408482088290E8E64010248C4A5AA840C2000110001521F0810A92E7",
INIT_09 => X"0003CE6581BD016342A951AB146C4480530C3B2A8088D3542651670200C1826A",
INIT_0A => X"00735D36209A8A20020894004284B660821030C8990467401218004041020002",
INIT_0B => X"512445B740457154562F957CC08B00093700080D0A4851001D8302D20A0A1530",
INIT_0C => X"00508650008008021021A40861021840869021A408610218C0869810D6043095",
INIT_0D => X"1C8508438450801043A08090380A8834207007022209038080190000999C8F84",
INIT_0E => X"000400200000C0002A48A206204C4205F3304B33004C0041006240140A1C310A",
INIT_0F => X"0000080040000083800400000100000000008400018040000100080000510100",
INIT_10 => X"0001000000000800000244040000020000000100002A0080000200100000A702",
INIT_11 => X"000000000020000000200000080002C000800008000000000022000006808000",
INIT_12 => X"0000000000000A2281000000000040A3810000000000402001400000022002A0",
INIT_13 => X"000000000004200001C0400000000010200001C0400000000010000004490010",
INIT_14 => X"0001070004000000000000060000104C08000000000000001000000903008000",
INIT_15 => X"CC004050CA0C00020220200070040000010401C4000000000000000000100008",
INIT_16 => X"4310E4310A4210A4210A4210A4210A4210A8D0830A68010001B4DA881048061C",
INIT_17 => X"21084290A4210A4210A4210A4210A4210A4210A4210E4310E4310E4310E4310E",
INIT_18 => X"90A421084290A421084390E4310C4390E4310C4390E4310C4290A421084290A4",
INIT_19 => X"015303C0C78C706428A14C586291000A044001FFE000003FFC004290A4210842",
INIT_1A => X"2492492492492492492492492492492492410410410410412821600001249249",
INIT_1B => X"51A8D46A351A8D46A351A8D46A351A8D46A351A9D4EA753A9D4EA753A9D49249",
INIT_1C => X"FFFFFFFFFFFFFFFC00000000000000000000000038F56351A8D46A351A8D46A3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"55AB02055AB0207FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"420000000000000000000000000000000000000000000000007FFFAB57FFFAB5",
INIT_28 => X"A800BAFFAE9554508002AA00AA843DF55FFAA955EFA2D168B55557BEAA000055",
INIT_29 => X"002AB55AAAA955EF005568A00087BE8BFFA2D155410AA8415555087BFFF55A2A",
INIT_2A => X"AAABFF5508003FF555D0002145552ABFEBA007FC21EF007FD75FFAA841541008",
INIT_2B => X"082EBDEAAA2FBEAABA5D7FC0155005168B455D042AB45F7FFD741000042AA10A",
INIT_2C => X"FF7FBEAB55F7AABDEBA5D7FC2010A2D1575FFF7AA975555D2E80145F78415545",
INIT_2D => X"EF5555554AA087BC01FFFFAAAAB55552A954BAFFFFE8B55552EBDE00F7AEAABF",
INIT_2E => X"000082E820BAA2FBEAB5555557DF55A2AEBDF555D2E954BA002EAAABA002A821",
INIT_2F => X"FB7D5D7FEAA3808554203A000000000000000000000000000000000000000000",
INIT_30 => X"1557D1475FAF45BEAA800AAFFAA95578080038A2AA28E3AF55E3A0BA5D7AADB6",
INIT_31 => X"BD55D7BE80004AA1E8E2AB55B6A0925D7085F6AA10087FEABD7AAD57AEBAB68E",
INIT_32 => X"F5D0438140E2FA38B6AEBFF6D1D04AAFFA41040017D5D20B8EAA007FC51C7A2F",
INIT_33 => X"D0A901FFFF801557D1C20B8EAAA2FBE80AA557BE8B6D5D5FFABEF49002FB55FF",
INIT_34 => X"5D20BDE00EBAAA8BC7EBDFEAFEFAB8ABAE925D21C7010EADB525D7FFAE975C75",
INIT_35 => X"F002EADA921420871D74971D24820875C21D5EB8AA8FFF012A954BAFFF5EFB45",
INIT_36 => X"000000000000000000001C24820BAB6FFEFB6D555578F7DB6A0BDF7DEB8E125F",
INIT_37 => X"B55A28408145AAFFFFFFF5D7FEAABA0051400A20000000000000000000000000",
INIT_38 => X"AB55FAD568AA2AFAE975EF555168B55F7AA800BAF7AA955EF00042AAA2A2AEAA",
INIT_39 => X"2AAAA007FD55558A7BD7145FBB8020A35D2ABEF55F7800015F087FEAA00007FE",
INIT_3A => X"968F575D003FF55F7D5420BA5D2ABFEAAF7AE9DFF759A82AEF70800021EF5504",
INIT_3B => X"FFD5145FBAC9755F05040255FFD84175EF55002AAB0A2FFEAABA557BEA3EF057",
INIT_3C => X"82E974AAF7D57DF45552A3FF10AA8429F45A7D5EAF5FFBAEAAA10554155400AA",
INIT_3D => X"FF843FFE77C80825BC052ABFE10550415557085540000005156155FE90A8F5C0",
INIT_3E => X"00000000000000000000000000000000000005500020AAF7FBFFFEF04552ABFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(0),               -- Port A write enable input
DIA(0)   => data_write_a(3),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(3),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(0),               -- Port B write enable input
DIB(0)   => data_write_b(3),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(3),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_4_9 : RAMB16_S1_S1
generic map (
INIT_00 => X"A108400020612C80284210081034849800A00030300004833522C82D04A16002",
INIT_01 => X"2043998A1839284D1CA0650E1E504368403008418984014902030806A0D10200",
INIT_02 => X"C120042200000000044441CE01E80F00A49043118680008002000000026208E4",
INIT_03 => X"040001020019200020011209CC0164C060000000690111040144800042F5C403",
INIT_04 => X"7029AF0F81A00010CCA47700CC513CAC0D0B8E02010740E19754080108988021",
INIT_05 => X"02139405007133C0712244CD20F20105D583000020E9892201D304D42A9835E1",
INIT_06 => X"9190440300078002014405D9EE814C0284A883B6D7038AE079059B7800048092",
INIT_07 => X"000100AA0004408000000004840400008D200102503000782000C00C8025C000",
INIT_08 => X"00728A00408403220811991E02120C044058080004000001101121F220000260",
INIT_09 => X"811001E1185B38AD23C3707AD46440818F3CF80EC423CA7D01D123C80200816A",
INIT_0A => X"45810810A01B40216361056D6150F41200280001900439001FD8A00041400000",
INIT_0B => X"11FC88076266E800D605402962A820211500024808010512C40106D222223B14",
INIT_0C => X"0408804116040B02C02C500B0C02C100B0C02C100B0402C300B0401618058611",
INIT_0D => X"040200050200501301208482200D00D0A0408402C4282200A84800009B878680",
INIT_0E => X"00000020000100024AC88300300060090F0D830F00025400300204D018000804",
INIT_0F => X"8000000040000206A2000800000000000000950002E010000000080000588040",
INIT_10 => X"0000000000000808000554000200000000000100006D0020000000100000BB00",
INIT_11 => X"0000400000000000002000001A0002504001000000000000002280000D800800",
INIT_12 => X"0800000000000E2C802000000000408D801000000000408012440000200110A0",
INIT_13 => X"000000000004680003A0040000000010280003800800000000102800000B0000",
INIT_14 => X"000005C0002000000000000620000158000010000000000010A0000B00000200",
INIT_15 => X"C30146200400104002602600400000000294004000000004000000000010001A",
INIT_16 => X"0080200000008020000000802000000080080000004090014134DA101288C6DB",
INIT_17 => X"0802000000000401806010040180601004018060100000802000000080200000",
INIT_18 => X"8060180601004010040080200802000000000000802008020000000000008020",
INIT_19 => X"C0A28A063807E0500014063450404882846FFE000003FFC00000010040100401",
INIT_1A => X"AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA28A28A28A28A2934C8D0CCD145144",
INIT_1B => X"68341A0D068341A0D068341A0D068341A0D068351A8D46A351A8D46A351AAAAA",
INIT_1C => X"FFFFFFFFFFFFFFFC0000000000000000000000001FE32068341A0D068341A0D0",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"408102040810207FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"800AA00000000000000000000000000000000000000000000040810204081020",
INIT_28 => X"168B55557BEAB4500554200000557FE10FFFBEAA10007FD7410FFAA97555082A",
INIT_29 => X"55574105D2A800AA00043FEBA5D7FEAA00007BE8AAAAA843DF55FFAA955EFA2D",
INIT_2A => X"57BC00AAA2FFEAAAAAA8415555087BFFF55A2AA800BAFFAE9555508002AA0000",
INIT_2B => X"A2AA955EF005568A00087BE8BFFA2D17DE1000517FE10AAAAA8AAA002E975455",
INIT_2C => X"FAA8417410A2D140000F7FBC2010A2D157400AAAE974AAAAAA974BA08002AB55",
INIT_2D => X"EFA2AABDEAA087BEAAAAA2FBD54BA080002145552ABFEAA007FC21EF007FD75F",
INIT_2E => X"00055042AB45F7FFD741000042AA10AAAABFF5508003FF55F7D568A00552EA8B",
INIT_2F => X"5400F7A49057D0824850B8000000000000000000000000000000000000000000",
INIT_30 => X"3AF55F7A0925D7AADB6FB7D5D7FEAB7808554203A145178E00FFFBE8A101475D",
INIT_31 => X"A9557D080038AAA145157428492E8008200043FE925571EFA380871C7028A28E",
INIT_32 => X"AEA8A9200249056D4175C5092AAF5FDA38BE8E1557D1475FAF45BEAA800AAFFA",
INIT_33 => X"AA4954281C0E2FB55B6A0925D7085F6AA10087FEABD7AAD57AEBA08517DE00AA",
INIT_34 => X"007FC51C7007BD55D7BE80004AAFEDB42028EBFBC2028BED152438AAA092492A",
INIT_35 => X"AF7DF6AA00412EAABFFAA803DEBA0875EDA80BEF1C743840040017D5520B8EAA",
INIT_36 => X"0000000000000000000041002FB55FFF5D0438140E2FA38B6AEBFF6DBE84AAEB",
INIT_37 => X"A00FFFFEAA105D5155410FF84021EF0800154B20000000000000000000000000",
INIT_38 => X"DEBA0851574B2AAAEAAB55F78400145AAFFFFFEF5D7FEABFF0051400A25D5568",
INIT_39 => X"68B55F7AA800BAF7AA955EF00042AAA25555410BA082E8201000043FE005D517",
INIT_3A => X"568AA200557DE00AAAAAAA000804001FF005575408AA557FEB2FFAE975EF5551",
INIT_3B => X"D1550AAAA8002010F2AC154B25F2ABFF55F7800015F087FEAA00007FEAB55FAD",
INIT_3C => X"800021EF55042AAAA007FD5555087BD6145FAAC000A2A6FBC00BAAAFBC00BAF7",
INIT_3D => X"F7AEBDFF779A82AA43F7FBE8A00082EA8BFFAA843FEBA08517DE00F3F9574B30",
INIT_3E => X"000000000000000000000000000000000000008003FF55F7D5420BA5D2ABFEAA",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(0),               -- Port A write enable input
DIA(0)   => data_write_a(4),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(4),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(0),               -- Port B write enable input
DIB(0)   => data_write_b(4),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(4),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_5_9 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50DF4A0791B3FCB694379283C81FD996A091832102004A336A20E03C040C002",
INIT_01 => X"805FBDC69830A84D5C6A60000C34C26841280A00084000C8C212892EEAD53235",
INIT_02 => X"3B2026B578918E640A4F01CF8011FF0002080000082CA9998276DF7772C7C80D",
INIT_03 => X"37134108420D700084205702A4008A1D9100002171C0E0051554D93A11F5D140",
INIT_04 => X"8A41A0FC03A56DA000425A819410E3816C086198A388B702A8CA1210844A0C4C",
INIT_05 => X"B1808A062E8BC835F5E84532D708238A282F00A9291224800A2861490343082C",
INIT_06 => X"903FB8483A90581859050424100940825C6184401CDC451B860A6507160C4100",
INIT_07 => X"D26F068BCC96CDF8918E640E96D1A3469D6300E2FFEA27F8E4D23248130E259C",
INIT_08 => X"0BFA82E568442B2A082C0A7E3014250D49DA37A2420619000002AFF48D1222E5",
INIT_09 => X"3F005001E40969289429360416DCD1C46083030604B1CA20C03DF83B0A2C60A5",
INIT_0A => X"14613C71005A10492B888120288F480D58858449026145B3830F449449062B4F",
INIT_0B => X"11AC04934AC648BFD727C031E64170A137D5AA5C3E4B0F8A3C58C34C002290E3",
INIT_0C => X"CA29C6CC50384B6AC6AC86AB31AACA6AB39AAC86AB39AACA6AB3055643559C31",
INIT_0D => X"C673E33CF28F38603855401985228A0614BD30A0A2819852011E5AC2B87F9182",
INIT_0E => X"FF87C002F87A803E460B2516510CA594FF0044FFA4B08BAC4BB2CD0F09CF84E3",
INIT_0F => X"0DFF0F8005F0F5100DFFF5E15D06101C55EB29F1E00BE53FE1F000BE1E802F94",
INIT_10 => X"F12F0380231F17D78FC029FFF58D9A70380230F2FE0017C37FC3E0017C3D005F",
INIT_11 => X"FC7F023C0CA700125C0F8F7E43F1F001BFFE7C69E01804E1E7CCF8FC003FF5F1",
INIT_12 => X"023E00017C1FC1A4BFD82C3081C5BD27BFE30C3081C5BD00C02365D645CEEF5B",
INIT_13 => X"61E0042787F181E9C1EFD8CB8120C5AF41E9C18FD60F0C20666F41E9F009FFFD",
INIT_14 => X"7A7C077FFF404F80005F07F187A7D14BFFC96111C048278DEB074F9930FF9D80",
INIT_15 => X"C064014B8B652E2B3120C81284641D3E8DBF7D636FE860190700132C1F0EFB80",
INIT_16 => X"38CE1384E3384E338CE138CE1384E33C4E3ECE32E128882551349A1CBAA44103",
INIT_17 => X"84E3384E3384E3384E338CE138CE1384E3384E338CE138CE1384E3384E338CE1",
INIT_18 => X"CE138CE138CE138CE1384E3384E3384E3384E338CE138CE138CE138CE1384E33",
INIT_19 => X"F5E5BB4E7F7B9DB7FF3A1B6DB7E8410A8C000000000000000000384E3384E338",
INIT_1A => X"BEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEF9F7CFDFDDCF3CF3D",
INIT_1B => X"BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEFBEF",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000001711C7BBDDEEF77BBDDEEF77",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"FDFFF00000000000000000000000000000000000000000000080000000000000",
INIT_28 => X"FD7410FFAA97410082A800AAAAAE955450055421FFFFFBC0010AAD5574BA557F",
INIT_29 => X"7FD74000055574BA5D7FD7555A2D5575EF55517FF5500557FE10FFFBEAA10007",
INIT_2A => X"0002AABA5D2ABFFFFAA843DF55FFAA955EFA2D168B55557BEAB5500554200000",
INIT_2B => X"5D2A800AA00043FEBA5D7FEAA00007BC00AAAAAEBDF45A28428B45FFD168BFF0",
INIT_2C => X"5080028A00A2FFFDE00F7D57FEBAFF80174BAAAD1555EF555555555005557410",
INIT_2D => X"BA5D2E821FFA2D5554BA557BD75FFAA8415555087BFFF55A2AA800BAFFAE9555",
INIT_2E => X"00000517FE10AAAAA8AAA002E97545557BC00AAA2FFEAAAA082A97545F7D5420",
INIT_2F => X"7010BEDF524AA5571FDFEF000000000000000000000000000000000000000000",
INIT_30 => X"78E00EBFBE8A101475D5400F7A49043D0824850B8A2AE9756D145B401FFFFFFC",
INIT_31 => X"FEAB7D0855420BA1471D74380851524BA5571D757DB6D5525EF555178F6D1451",
INIT_32 => X"8A28B6DEBDF6DBEF1C0A28AAA5524BFFFFA28E3AF55F7A0925D7AADB6FB7D5D7",
INIT_33 => X"5555057D145152428492E8008200043FE925571EFA380871C7028B6AEBDF45B6",
INIT_34 => X"BEAA800AAFFAA9557D080038AAAA2FBF8E10EBD578EAAFF8415482BED1555EF5",
INIT_35 => X"81C209256DFFDF420BA552A821FFB6DF574A85575C55EFBE8E1557D1475FAF45",
INIT_36 => X"0000000000000000000008517DE00AAAEA8A9200249056D4175C50920875FDA3",
INIT_37 => X"5FF5D7BC21EFF7FBD7400F7FBC00BA55557DFF70000000000000000000000000",
INIT_38 => X"01FF5D5568BE7555568A00AAFFEAA105D5155410FF84020AA0800154B2AAAA97",
INIT_39 => X"00145AAFFFFFEF5D7FEABFF0051400A25551554BA0051400BA5551575EFF7D14",
INIT_3A => X"1574B2FFAABFF45FFAAAABFFAAFFFDFFF552EA8AAA55043DFF7AAAEAAB55F784",
INIT_3B => X"8002410FFD5575EF5555421E75555400BA082E8201000043FE005D517DEBA085",
INIT_3C => X"FAE975EF555168B55F7AA800BAF7AA955EF00002AAA2A2FBE8A00A2D16AAAAFF",
INIT_3D => X"0055554088A557FEB25D00021FFFFFFC00BA552A821EFFFFFD74BA5D51575F7F",
INIT_3E => X"000000000000000000000000000000000000000557DE00AAAAAAA000804001FF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(0),               -- Port A write enable input
DIA(0)   => data_write_a(5),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(5),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(0),               -- Port B write enable input
DIB(0)   => data_write_b(5),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(5),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_6_9 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10800B0061A01002840002C03002818000402322520070B313301C4389B2082",
INIT_01 => X"250041CA3839684D18A160000C52426841000000090800090210080008110200",
INIT_02 => X"0020042080010000044654C0000C008010000000001020900200200002620814",
INIT_03 => X"060881021088200021080200E4000A0891000020610111500104C00000F14400",
INIT_04 => X"0880000100000002000052288144004281C050400100280000C8100000080001",
INIT_05 => X"928080840001100A08009000280201000850E022401400002028214043410820",
INIT_06 => X"10100518090012122100C808049310002040000410A0001400000200120840D2",
INIT_07 => X"000100800004400001000000860408108C22000A502010074120044800040001",
INIT_08 => X"50000040D0C4E2088003FD01C01004044058082004000000000121F020408244",
INIT_09 => X"00BF17E9001205A5204911F814444080400100020000D200DFD16400C2A40AA0",
INIT_0A => X"04611C17849000022862A1596C8B5DF04834948900000100220C244840000880",
INIT_0B => X"03AD0413424E4044D665C070C22602291504400D084915020448114080201000",
INIT_0C => X"5E08864011088B22D22C008B0022C408B1022C208B0822C608B1111600458010",
INIT_0D => X"4251A12CD28A300429688001000800000020280204001000A00804309A002182",
INIT_0E => X"0000000280402400420800000000006200FC10002442042429324294014E8CA7",
INIT_0F => X"A40000000500800840000800000000000002280018001480000000A010100052",
INIT_10 => X"00000000000004C2003000010240000000000000680800290000000140202000",
INIT_11 => X"2000C0000000000000000442000001080001000000000000010C000280001804",
INIT_12 => X"08000000000801C300A010000000156000902000000015101200002800000000",
INIT_13 => X"000000000101800038002408000000094000386028040000000940000ED40000",
INIT_14 => X"0003B000002000000000020180002A24005010000000000023000060C7000A40",
INIT_15 => X"3F0280090321000040A410C28108000160008094000810040000000000002300",
INIT_16 => X"284A5284A728CA5284A528CA728CA52C4A5A0A32A300940101349A0408240818",
INIT_17 => X"9CA1294A329CA5284A728CA7284A5284A728CA5284A528CA728CA5284A728CA7",
INIT_18 => X"CA3294A129CA3294A129CA1294A329CA1294A3294A129CA3294A129CA3294A32",
INIT_19 => X"F5F78BCE7F8FF0F4FA955F7CF7F40A80145D55555556AAAAAAAAA94A329CA129",
INIT_1A => X"8E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E39B6CEDECDDF7DF7D",
INIT_1B => X"F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE38E3",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000001A1A33F9FCFE7F3F9FCFE7F3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"555FF00000000000000000000000000000000000000000000080000000000000",
INIT_28 => X"BC0010AAD5574BA557FFDFFF087BFDF45F7AA974AAAAAA97555F784174BAF7D5",
INIT_29 => X"515555508043FE00F7AA97555A2FBD7410AA8428AAAAAAE955450055421FFFFF",
INIT_2A => X"7D1575EFFFAA9555500557FE10FFFBEAA10007FD7410FFAA97400082A800AA08",
INIT_2B => X"0055574BA5D7FD7555A2D5575EF55517FF55A2AA97400552AAAB45082E80155F",
INIT_2C => X"500554200000003DE10FFD5401FFF7AAA8A10082EAAB45A2FFC2000007FD7400",
INIT_2D => X"10AA803FE105D516AABAFF843FFFFAA843DF55FFAA955EFA2D168B55557BEAB5",
INIT_2E => X"000AAAEBDF45A28428B45FFD168BFF00002AABA5D2ABFFFF087BD5545007BFDE",
INIT_2F => X"256DEB84104BAFFD1525FF000000000000000000000000000000000000000000",
INIT_30 => X"9756D145B401FFFFFFC7010BEDF524AA5571FDFEF1C7BFFF55FFA095482B6A49",
INIT_31 => X"4904380824850381C5B5057D1C003DE28F7A49057DAAF5D2428A2842AAAAA2AE",
INIT_32 => X"2AAFB451C2A8017DE3DF525FFFFA49756D145178E00EBFBE8A101475D5400F7A",
INIT_33 => X"2F1C50381471D74380851524BA5571D757DB6D5525EF555178F6DAAA49542841",
INIT_34 => X"AADB6FB7D5D7FEAB7D0855420BA1C0E3FE00E3DB471EFE3AAAAA00082EA8B6DA",
INIT_35 => X"F1C7BD057D1C71FFE10A28038E1049516AAB8FF8428FEFA28E3AF55F7A0925D7",
INIT_36 => X"00000000000000000000B6AEBDF45B68A28B6DEBDF6DBEF1C0A28AAA5524BFFF",
INIT_37 => X"F55F78017400F780001FFAA84000AAFFD1401E70000000000000000000000000",
INIT_38 => X"20BAAA8428AA2AAAA975FF5D7BC21EFF7FBD7400F7FBC00BA55557DFF7557BFD",
INIT_39 => X"EAA105D5155410FF84020AA0800154B2557FC01EF55043FEAAFF80021EFA2D14",
INIT_3A => X"568BE7AA80174AA082ABDF555D2A821EFAAFBC01FFF780155F7555568A00AAFF",
INIT_3B => X"AEA8A10082EA8BEFAAD5554B25551554BA0051400BA5551575EFF7D1401FF5D5",
INIT_3C => X"AAEAAB55F78400145AAFFFFFEF5D7FEABFF0051400A25D2EBFE10AAFFD55EFA2",
INIT_3D => X"552EA8AAA55043DFF7557BC01EF55557DE00AA842AA0000516AABAFF8428BE7A",
INIT_3E => X"0000000000000000000000000000000000000FFAABFF45FFAAAABFFAAFFFDFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(0),               -- Port A write enable input
DIA(0)   => data_write_a(6),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(6),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(0),               -- Port B write enable input
DIB(0)   => data_write_b(6),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(6),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_7_9 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10844B00482258A2842112C02450418800002300500030B313300C418992002",
INIT_01 => X"000009CA3839684D1CA0E0000E51424840000000080000080200080008510204",
INIT_02 => X"0120042086010000044600C00008000004100000000260900200000002402004",
INIT_03 => X"8628A10000082400000002408400080011000000610008000208C00000E14400",
INIT_04 => X"0911800100A000000000524084000040000050001140200100C8100000080102",
INIT_05 => X"0300812401011000000000002000114008008060441000000020024093000000",
INIT_06 => X"9190431C0D4010100000880804010010800000041080081000000200010424B2",
INIT_07 => X"000100AA0004408601000004860000008C02000A103010006928040800062481",
INIT_08 => X"84000048D484C20888000A0002120484C048007004000000000021F000000244",
INIT_09 => X"00A06009881201A520491004106C48A04040002400A15A208001650004001020",
INIT_0A => X"C99E1060201002044809C1040140A001004808810000459033189C0A400118A0",
INIT_0B => X"102000024040484050050041648A0041140C500B08821054C000264120000400",
INIT_0C => X"0404A083260E0832132011880462011880462051881462051881D31018C40620",
INIT_0D => X"0001000080001000813094801A8F80F00A600B52602801A88848011118003700",
INIT_0E => X"000003C007C002808228010410082042C000C000000004001002000400040002",
INIT_0F => X"A4000007800F80C840000800009864038A1200081C0014800000F001F0200052",
INIT_10 => X"00002C0E00E0E4004038000102400002C0E00E0D20100029000001E003E04000",
INIT_11 => X"2000C04031100E0403D0700300080908000100000661801E1900040380001804",
INIT_12 => X"0840878083E8003780A01043203A101780902043203A10082410082880000000",
INIT_13 => X"0601E0187900181035E0240806483248181035E0280410C8198818100DDD0000",
INIT_14 => X"0403774000201021E020FA006040376C00501022131210722060806D47000A40",
INIT_15 => X"00928A0002000110888600C032128201519480D40009902430160403E0E00506",
INIT_16 => X"01000000020080601802000000000405000A0020020081014134928820480010",
INIT_17 => X"0802018040000000006018020080200804010000000000806018020080000004",
INIT_18 => X"0000000001806008020000001006008020080001004008020080201004000020",
INIT_19 => X"0000000000000000000000000000400A004618618618C30C30C3000020180600",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000000B0840000000000000000000",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"1555500000000000000000000000000000000000000000000080000000000000",
INIT_28 => X"A97555F784174BAF7D5555FFF780155EFAAAEA8ABAAAFBFDE0055556AA005D04",
INIT_29 => X"55555EFAAFFFDFEFAAAAAAB455D556AA00FFAE95555087BFDF45F7AA974AAAAA",
INIT_2A => X"02EAAAAA082EA8A00AAAE955450055421FFFFFBC0010AAD5574BA557FFDFFF55",
INIT_2B => X"08043FE00F7AA97555A2FBD7410AA8428AAA557BFDFFF55003DFFFF7FBEAA000",
INIT_2C => X"0082A800AAF7AE975FFA28000010552EBDE00007BEAAAAA2D140000085155555",
INIT_2D => X"45087FEAB455D516AB55557BD55FF00557FE10FFFBEAA10007FD7410FFAA9740",
INIT_2E => X"000A2AA97400552AAAB45082E80155F7D1575EFFFAA955555D51574AAAAFFD55",
INIT_2F => X"AE105D556AA10410E17555000000000000000000000000000000000000000000",
INIT_30 => X"FFF55FFA095482B6A49256DEB84104BAFFD1525FFFF8E175C7A2AAAAA82A2F1F",
INIT_31 => X"F524AA5571FDFEF415B575D7AAF1FFFD7AAAAAFB7D495F6AA10E3AE905551C7B",
INIT_32 => X"003AFEFEBFBEAA001C2EA8A821C2EAAA00A2AE9756D145B401FFFFFFC7010BED",
INIT_33 => X"EDB470101C5B5057D1C003DE28F7A49057DAAF5D2428A2842AAAA497BFAFFF49",
INIT_34 => X"1475D5400F7A490438082485038F7A4905C7A28A070384120BDE100075EAA82B",
INIT_35 => X"D495150492BEF1D2555087BE8B7D555F6AB57417BC05D7145178E00EBFBE8A10",
INIT_36 => X"00000000000000000000AAA495428412AAFB451C2A8017DE3DF525FFFFA49756",
INIT_37 => X"555A2AEA8A10AAD568A00555168A10002E9754D0000000000000000000000000",
INIT_38 => X"8A10AAAE8215D557BFDF55F78017400F780001FFAA84000AAFFD1401E7FFAA97",
INIT_39 => X"C21EFF7FBD7400F7FBC00BA55557DFF7007BD5555AAD57DF55AAAEBDFEF007BE",
INIT_3A => X"428AA2007FE8BFF080028BFFAAFFEAA105D2EAAA005D2AAAA18AAAA975FF5D7B",
INIT_3B => X"043DE0000516AA10F7FBD7408557FC01EF55043FEAAFF80021EFA2D1420BAAA8",
INIT_3C => X"55568A00AAFFEAA105D5155410FF84020AA0800154B2FF8402145A2AA954AA00",
INIT_3D => X"AAFBC01FFF780155F7005140000FFD140145007FE8BEF557BEAB55087FC215D5",
INIT_3E => X"0000000000000000000000000000000000000AA80174AA082ABDF555D2A821EF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(0),               -- Port A write enable input
DIA(0)   => data_write_a(7),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(7),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(0),               -- Port B write enable input
DIB(0)   => data_write_b(7),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(7),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_8_9 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00000648E2840112C00000418000002700500030B3132000400812082",
INIT_01 => X"100008480009004C04A100000252024840000000180800080200010040110204",
INIT_02 => X"0020042000490000004600804008000005100000000024900200000002400004",
INIT_03 => X"0A0C33400008082400000080A4004B0891000020610112000040C00000E5C000",
INIT_04 => X"18800001000000000000512080000040800150400824280110C8100000120200",
INIT_05 => X"908084A10100100200004080280008240810802206940000012C214451610800",
INIT_06 => X"81B000080860109021400008040000202048020414A0021400040200322824C1",
INIT_07 => X"000000080004408049000004860000008402001A50208000630C040800062483",
INIT_08 => X"440000428644212280800A00021004044048002124000000000021F000000244",
INIT_09 => X"00004009001001010008100414644410400102228000D20080114502006409A2",
INIT_0A => X"000051312000042200294429148A4801C80C8C81000045907118040340020832",
INIT_0B => X"4020000240404140004D0544C4AA0001150410090302500011C813428A000400",
INIT_0C => X"46501090008820240240409000240009000240009000240009000120204808A5",
INIT_0D => X"42D1A168D09A301468402480004780F00140080860280004085904309A002196",
INIT_0E => X"00783FC00044340242280000000000020000C0000442106419120004034685A3",
INIT_0F => X"8000F07F800088A80000081EA2F9EC0000064004081010001E0FF00011104040",
INIT_10 => X"0ED0FC7E00000422201080000202658FC7E0000021882020003C1FE000222080",
INIT_11 => X"018059C3F350FE0C00000002A0040500000103961FE780000110010090000800",
INIT_12 => X"FD41FF80000830200021C1CF600012200010D1CF600012121600100810000004",
INIT_13 => X"9E1FE000010A1802100004343ED8000898021000087073D80008980200800002",
INIT_14 => X"0080200000BEB07FE00002086008020000209AEE3F300000246020200000620B",
INIT_15 => X"0088881903210000440610C8000A808040000208901786E4F0FE0C0000000166",
INIT_16 => X"685A1685A769DA368DA368DA769DA36CDA121A11A141800011309284002C0810",
INIT_17 => X"95A5685A1685A5695A368DA368DA769DA368DA368DA7695A1685A1685A5695A1",
INIT_18 => X"5A1695A568DA368DA369DA768DA1685A1695A5685A168DA369DA768DA368DA16",
INIT_19 => X"A4028A0A543EBC57A10A1E75D64108080468618618630C30C30C69DA5685A168",
INIT_1A => X"9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7BF3CCD8DF5B2DB2C",
INIT_1B => X"F87D3E1F4F87D3E1F4F87D3E1F4F87D3E1F4F87C3E1F0F87C3E1F0F87C3E79E7",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000006A6D4F87D3E1F4F87D3E1F4",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"155FF00000000000000000000000000000000000000000000080000000000000",
INIT_28 => X"BFDE0055556AA005D0415555080000000087BEAA10F7803DE00FFAEBFFFF0800",
INIT_29 => X"2AA8AAA557FC0010F780154105D7FC2145005155555F780155EFAAAEA8ABAAAF",
INIT_2A => X"7FFFFF55AA80155FF087BFDF45F7AA974AAAAAA97555F784174BAF7D5555FF55",
INIT_2B => X"AAFFFDFEFAAAAAAB455D556AA00FFAE95555AAFFE8A00552EBFE00F7D17FF45F",
INIT_2C => X"A557FFDFFF5504000AAAAAAA8B55F7D140010552E821EFAAAABDF555555555EF",
INIT_2D => X"55AA8028A00A2D57FF45557BE8A00AAAE955450055421FFFFFBC0010AAD5574B",
INIT_2E => X"000557BFDFFF55003DFFFF7FBEAA00002EAAAAA082EA8A00002AA8A10F784021",
INIT_2F => X"FE10F7AEBAFFF080A175D7000000000000000000000000000000000000000000",
INIT_30 => X"175C7A2AAAAA82A2F1FAE105D556AA10410E17555080E000280071E8A00EB8E3",
INIT_31 => X"4104BAFFD1525FF492EA8AAA5571C2000FF8A17400557FC015514555757DFF8E",
INIT_32 => X"2ABDE10EBDF7AF6DE3FFF8F7DB68A105D71C7BFFF55FFA095482B6A49256DEB8",
INIT_33 => X"AA0BDF6D415B575D7AAF1FFFD7AAAAAFB7D495F6AA10E3AE90555A2FBE8A3849",
INIT_34 => X"FFFFC7010BEDF524AA5571FDFEF550E00082B6A0AFB55F7D1420104124821D7A",
INIT_35 => X"01C2EA8A00F7800017DA2842FA00B6D578F6D557FFDA00A2AE9756D145B401FF",
INIT_36 => X"00000000000000000000497BFAFFF49003AFEFEBFBEAA001C2EA8A821C2EAAA0",
INIT_37 => X"0BA08556AA00AAAABFE00F7AEAABEF082E955450000000000000000000000000",
INIT_38 => X"21555D51575EFFFAA97555A2AEA8A10AAD568A00555168A10002E9754D082E82",
INIT_39 => X"17400F780001FFAA84000AAFFD1401E7082EAAABA5D5140010F7AE974105D7BC",
INIT_3A => X"E8215DA2FFE8ABA082ABFE00AAFBEABFFAAFBEABFFF7AA80145557BFDF55F780",
INIT_3B => X"D540000000402145AA843FFFF007BD5555AAD57DF55AAAEBDFEF007BE8A10AAA",
INIT_3C => X"AAA975FF5D7BC21EFF7FBD7400F7FBC00BA55557DFF75D2E82010F7843DF45FF",
INIT_3D => X"5D2EAAA005D2AAAA185D2AAAA10F780021FFA2803DE10FFD16ABFF5D7BFDE10A",
INIT_3E => X"0000000000000000000000000000000000000007FE8BFF080028BFFAAFFEAA10",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(1),               -- Port A write enable input
DIA(0)   => data_write_a(8),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(8),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(1),               -- Port B write enable input
DIB(0)   => data_write_b(8),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(8),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_9_9 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00018248A2840112C00002C18000002300500030B3132000400812006",
INIT_01 => X"400008000000004C0020000000100248413C0A61590001D90213C10008110204",
INIT_02 => X"01A0042080010000054600C04008000004100000001020900200200002420804",
INIT_03 => X"024003400008012400000010E4004B0891000020610310000144C00000F5C000",
INIT_04 => X"1801800100E000000000510084000040010050020810200000C8900000320200",
INIT_05 => X"918004311104100000000000200008100800002000100000002C234415610820",
INIT_06 => X"81B00008080010100000980804000008800042041080001000100200322C2481",
INIT_07 => X"0000811800044080010000058600000086020002502080006000040800062C80",
INIT_08 => X"0000004001D4618008800A00061004044048002004000000000061F000000244",
INIT_09 => X"000040090802009420409004104444084001022400214A2080014400026401A2",
INIT_0A => X"04000071200000A003CA294140200800C80C8C8100004590111C040040120800",
INIT_0B => X"12210002404848502847040164880021150400080222000200C8034200000000",
INIT_0C => X"4610088010080421021040841021000841021000841021000841010800420820",
INIT_0D => X"42D0A16C529A321068500484000500D10042080040284000084900001A002196",
INIT_0E => X"00000002804000004228010410082002C000C0002400046419120410034285A1",
INIT_0F => X"A00000000500800800000800000000000002290008001080000000A010100042",
INIT_10 => X"00000000000004C2001000000240000000000000680800280000000140202000",
INIT_11 => X"0000C0000000000000000442020001000001000000000000010C800080000804",
INIT_12 => X"08000000000801A7802010000000152780102000000015000600000800000000",
INIT_13 => X"000000000101900011E0240000000009500011E0280000000009500004DD0000",
INIT_14 => X"000137400020000000000201C000136C00101000000000002340002947000240",
INIT_15 => X"0080881901210000000600C280028000419480D4000010040000000000002304",
INIT_16 => X"68DA368DA1685A1685A1685A1685A16C5A121A13A141950051309284A82C0010",
INIT_17 => X"85A1685A1685A1685A368DA368DA368DA368DA368DA368DA368DA368DA368DA3",
INIT_18 => X"5A1685A168DA368DA368DA368DA368DA368DA368DA3685A1685A1685A1685A16",
INIT_19 => X"0157344CCCF48DE68A895C38E2540A8010100000000000000000685A1685A168",
INIT_1A => X"14514514514514514514514514514514514D34D34D34D34D28E1004039248209",
INIT_1B => X"D268341A4D268341A0D069349A0D069349A0D068341A0D068341A0D068345145",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000014D490D069349A0D068341A4",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"EAABA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"03DE00FFAEBFFFF0800155FFAAFBE8B45002A974AAAA803DFFFAA843DF45FFFF",
INIT_29 => X"7BFDE00A2FBD7400F7FBFDFFFA2AEBDE00AAFBEAABA080000000087BEAA10F78",
INIT_2A => X"055401FFF7AEAAA10F780155EFAAAEA8ABAAAFBFDE0055556AA005D041555508",
INIT_2B => X"557FC0010F780154105D7FC2145005155555557BE8BEF007FFDEAAAAD1555EF0",
INIT_2C => X"AF7D5555FFF780154AA5D2AA8A10F7AA974AA082E80010A2AAAAA10552AA8AAA",
INIT_2D => X"BAF7D17FEBAA2AEBDF45002EAAABA087BFDF45F7AA974AAAAAA97555F784174B",
INIT_2E => X"000AAFFE8A00552EBFE00F7D17FF45F7FFFFF55AA80155FF080400145FFFBEAA",
INIT_2F => X"8FC7BE8A3DF7DF7F5E8A92000000000000000000000000000000000000000000",
INIT_30 => X"000280071E8A00EB8E3FE10F7AEBAFFF080A175D7BEF1E8B6D002090482B68E3",
INIT_31 => X"56AA10410E175550871FFE00A2FBD0400FFF5FDFC7B6A0BDE38B6F5E8A92080E",
INIT_32 => X"7BFAE82A2DB555C71C5B451D7FFAAA8A38FF8E175C7A2AAAAA82A2F1FAE105D5",
INIT_33 => X"2AEADA38492EA8AAA5571C2000FF8A17400557FC015514555757D5D71E8BEF14",
INIT_34 => X"B6A49256DEB84104BAFFD1525FFFF84174BA5D20AAA00E3AA904BA142A87010A",
INIT_35 => X"7000400155FFFBEDA82FFD57DEBAAAA0BFF7D0024ADA921C7BFFF55FFA095482",
INIT_36 => X"00000000000000000000A2FBE8A38492ABDE10EBDF7AF6DE3FFF8F7DB68A105D",
INIT_37 => X"BEF080402000F7AAA8B55FFAABDFEFF7D16AA000000000000000000000000000",
INIT_38 => X"FEAAFFD16AA00082E820BA08556AA00AAAABFE00F7AEAABEF082E95545F7D568",
INIT_39 => X"A8A10AAD568A00555168A10002E9754D00517DE00A2FFC2000F7D17FF55FF803",
INIT_3A => X"1575EF555568BEF5D7FE8A10AAFFD55555D7FD5555FFAAA8AAAFFAA97555A2AE",
INIT_3B => X"AE800AA552A97400A2AEBDEAA082EAAABA5D5140010F7AE974105D7BC21555D5",
INIT_3C => X"57BFDF55F78017400F780001FFAA84000AAFFD1401E7FF80174AA5D0028A00AA",
INIT_3D => X"AAFBEABFFF7AA80145080002145F7FBFFE00FFD17FEAAA2803DFEF08043FE005",
INIT_3E => X"0000000000000000000000000000000000000A2FFE8ABA082ABFE00AAFBEABFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(1),               -- Port A write enable input
DIA(0)   => data_write_a(9),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(9),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(1),               -- Port B write enable input
DIB(0)   => data_write_b(9),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(9),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_10_9 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00018248A2840112C00002C18000202300500030B3132000400992006",
INIT_01 => X"254008000000004C002000000010026840000000080000080200010008110204",
INIT_02 => X"0020042000010000004455800008000004100000000000900200000002400004",
INIT_03 => X"020001021089000021081000C400090011000000610001540104C00000F14400",
INIT_04 => X"0811800101A00002000050088554004200C840000000200080C8100000000001",
INIT_05 => X"030080001000100800009400200000000840E020201000000024024001200020",
INIT_06 => X"81B00008080012120004CC080492500280208004148000100000020020042493",
INIT_07 => X"0000000800044080010000048404081085020002502000006000040800062480",
INIT_08 => X"100202400084410808000A00021004044048000004000000000021F020408264",
INIT_09 => X"010040090002008420401004144440004040022484214A2080110108C2C00320",
INIT_0A => X"04004166A48A0001080000000000080080181881000045901118044040020800",
INIT_0B => X"1201000200484910000F0105602622291404020902005002018002400A022000",
INIT_0C => X"0440001011808020120004801120044800120004801120044800110002400884",
INIT_0D => X"008000440210100041308480800F82F00040180260A808008848000018002104",
INIT_0E => X"000000028040000002280104100820020000400020000440100204100A000100",
INIT_0F => X"040000000500800800000000000000000002280008000400000000A010100010",
INIT_10 => X"00000000000004C2001000010000000000000000680800010000000140202000",
INIT_11 => X"200000000000000000000442000001000000000000000000010C000080001000",
INIT_12 => X"00000000000801C0008000000000154000800000000015000410000800000000",
INIT_13 => X"0000000001019800180000080000000958001800000400000009580002800000",
INIT_14 => X"0000A0000000000000000201E0000A0000400000000000002360002080000800",
INIT_15 => X"0080881000000000000600C28102800060000000000800000000000000002306",
INIT_16 => X"401004010040100401004010040100441020D0030008840051309A90BA884010",
INIT_17 => X"0902409024090240900401004010040100401004010040100401004010040100",
INIT_18 => X"1004010040902409024090240902409024090240902409024090240902409024",
INIT_19 => X"F546890A940FE0D3971243555205428290100000000000000000401004010040",
INIT_1A => X"8A28A28A28A28A28A28A28A28A28A28A28A28A28A28A28A29554199854514514",
INIT_1B => X"2B95CAE532994CA6532995CAE572B94CA6532994CA6532994CA6532994CA28A2",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000002718E72B94CA6532994CA657",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"FDE1000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"03DFFFAA843DF45FFFFEAABA007FC2155F7D155545AA80001EFAAFBEAB45557F",
INIT_29 => X"042AB55FFD168B55AA8000010FFFBE8BFFF78402155AAFBE8B45002A974AAAA8",
INIT_2A => X"AD16AABA002ABDE10080000000087BEAA10F7803DE00FFAEBFFFF0800155FF00",
INIT_2B => X"A2FBD7400F7FBFDFFFA2AEBDE00AAFBEAABAA2FFD741055003DFEFF7AA801FFA",
INIT_2C => X"05D0415555007FD74105555555EFF7FBC0145F78028A00A2D142155087BFDE00",
INIT_2D => X"55AAD168ABA002A975FFF7AEBDEBAF780155EFAAAEA8ABAAAFBFDE0055556AA0",
INIT_2E => X"000557BE8BEF007FFDEAAAAD1555EF0055401FFF7AEAAA105D042ABFF5D556AB",
INIT_2F => X"71D7AAFBEFB455D71F8E00000000000000000000000000000000000000000000",
INIT_30 => X"E8B6D002090482B68E38FC7BE8A3DF7DF7F5E8A92007BC217DEBDB55555AA8E0",
INIT_31 => X"EBAFFF080A175D700042AB7DEBDB6DB55BE8E05000EBFFE8BC7E38E07145BEF1",
INIT_32 => X"0A3DFD7F7A4821D7A2D16FA82142EB8E00080E000280071E8A00EB8E3FE10F7A",
INIT_33 => X"ED1421450871FFE00A2FBD0400FFF5FDFC7B6A0BDE38B6F5E8A92B6FBD541049",
INIT_34 => X"A2F1FAE105D556AA10410E175550071D54104951555D7EBF5C5155E3842AA00B",
INIT_35 => X"8410E2ABD749516FB55BED16FA820820955EFE3AEBDEAAFF8E175C7A2AAAAA82",
INIT_36 => X"000000000000000000005D71E8BEF147BFAE82A2DB555C71C5B451D7FFAAA8A3",
INIT_37 => X"1EFA2FFD7545AAAE97555A2FBFDF455D556AA000000000000000000000000000",
INIT_38 => X"8B45AAAA95545F7D568BEF080402000F7AAA8B55FFAABDFEFF7D16AA00087FC0",
INIT_39 => X"6AA00AAAABFE00F7AEAABEF082E9554500042ABFFA2FFFFF45F7AE97400AAFFE",
INIT_3A => X"16AA00FFFBD5400082EBFF45F78400155A2D57FE00552EA8A00082E820BA0855",
INIT_3B => X"D557555A2802AA10FFD54214500517DE00A2FFC2000F7D17FF55FF803FEAAFFD",
INIT_3C => X"FAA97555A2AEA8A10AAD568A00555168A10002E9754D085155410085557555AA",
INIT_3D => X"5D7FD5555FFAAA8AAA002AAAB4508557DF55F7D17FE000804155FFAAAABDEAAF",
INIT_3E => X"0000000000000000000000000000000000000555568BEF5D7FE8A10AAFFD5555",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(1),               -- Port A write enable input
DIA(0)   => data_write_a(10),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(10),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(1),               -- Port B write enable input
DIB(0)   => data_write_b(10),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(10),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_11_9 : RAMB16_S1_S1
generic map (
INIT_00 => X"A101C4B05A0034CA2840712C2D001419000002300500030B31B20084EC992002",
INIT_01 => X"90000986B83028491800E0000C26426040000000080000088200080802512224",
INIT_02 => X"1A2004205E010640024D00800008000004100000040EC090820018003241A00C",
INIT_03 => X"28639100000C5C00000045C08400C8001100000061806A001618C03001E54400",
INIT_04 => X"1A800001000009A0804059A190000040400040008058220008C8100000120D4E",
INIT_05 => X"02000E81080250010000002022000058080400000E1200000020004401000004",
INIT_06 => X"819435143F20101010001008040800B8100102041088011100022200000024B2",
INIT_07 => X"90640D280884453E01064002944180008402001295BA100022E4340800062D82",
INIT_08 => X"400000093204802200280A0012160585C1D808D004000000000323F40C102244",
INIT_09 => X"380040098010001100009204107C5950400000220080C200800900020C006827",
INIT_0A => X"80007100004016EA080801010000080D00200081000045B0511D289940103399",
INIT_0B => X"002000024040410A000D0104408810C115D9C008050042400100D04E88000002",
INIT_0C => X"00655010009264201200C7B421ED0C7B421ED0C7B431ED087B43176843DA1085",
INIT_0D => X"0401020080400A10012494881A4F80F209500BB2602881A488485C1318002000",
INIT_0E => X"6619A540124814800228010410082022C00040002020090020220C9600040802",
INIT_0F => X"ACCC334A802491600C587949B6D0141B4CC600D5761B1599865A500490B86A56",
INIT_10 => X"BAC845542056A61686EC81E3A6CB68AA2C622C9A251C352B330CB4A0092170D8",
INIT_11 => X"BCCAD0B5A81536080CC6B21A21B1FC09CB0F1076D4A200B2AD4068F4101639B5",
INIT_12 => X"4D2CC281E31AA0103AB8D5514066380804B268A2E060901204112566F10AC418",
INIT_13 => X"D551443C47281002540B2C9AAAA8662A1152B202AE3554403028115AA88201A1",
INIT_14 => X"548A20A0492A2724A0621620402A020141F172FB182A32AB6845AB6200251BC9",
INIT_15 => X"00C00A000200074044E6801832728080D00A380B753952C4877E0104DDE4D124",
INIT_16 => X"0080200802008020080200802008020480080022020081010124988800400010",
INIT_17 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_18 => X"0000000000802008020080200802008020080200802008020080200802008020",
INIT_19 => X"55062608804180C0B10A42104201400204000000000000000000000000000000",
INIT_1A => X"00000000000000000000000000000000000820820820820801C4149470000000",
INIT_1B => X"0000000000000000040200000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000007E0F0000000000000100800",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"000AA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0001EFAAFBEAB45557FFDE10082ABDF5508557DF45002ABDFFFF7803DE10AA80",
INIT_29 => X"AEBFF45FFAEBFEAA002A801FFF7FFE8A10A28000000007FC2155F7D155545AA8",
INIT_2A => X"2AABFE10082ABFFEFAAFBE8B45002A974AAAA803DFFFAA843DF45FFFFEAABAA2",
INIT_2B => X"FFD168B55AA8000010FFFBE8BFFF78402155AAD155555A28428BFF002ABDE00A",
INIT_2C => X"F0800155FF00557FF45557FC2010002A80010A2842AAAA007BFFF4500042AB55",
INIT_2D => X"FF5D00154BAF7FBE8BEFFFD540000080000000087BEAA10F7803DE00FFAEBFFF",
INIT_2E => X"000A2FFD741055003DFEFF7AA801FFAAD16AABA002ABDE10A2D168A10A284021",
INIT_2F => X"DFC7F78E3FE28B684070AA000000000000000000000000000000000000000000",
INIT_30 => X"C217DEBDB55555AA8E071D7AAFBEFB455D71F8E00002EBDF6D005B78F7D142AB",
INIT_31 => X"A3DF7DF7F5E8A92BEAEBFF7DEBA0BDEAA1C2A801C7E3FFEFA10B68407038007B",
INIT_32 => X"8A28BFF082ABAE10B6AAB8E280820B8FEFBEF1E8B6D002090482B68E38FC7BE8",
INIT_33 => X"07FF8F7D00042AB7DEBDB6DB55BE8E05000EBFFE8BC7E38E07145B6D15756DA2",
INIT_34 => X"EB8E3FE10F7AEBAFFF080A175D708517DF7D497BC5028142A87000A28A2AA920",
INIT_35 => X"0B6DB6AA28A280001FF5D0A10482FFFFEFBC7E3DF42028080E000280071E8A00",
INIT_36 => X"00000000000000000000B6FBD5410490A3DFD7F7A4821D7A2D16FA82142EB8E0",
INIT_37 => X"FEF007BE8BFF5D2ABDF55F7AABDEAAF784154BA0000000000000000000000000",
INIT_38 => X"DE00FF84154BA087FC01EFA2FFD7545AAAE97555A2FBFDF455D556AA00082EBF",
INIT_39 => X"02000F7AAA8B55FFAABDFEFF7D16AA00FFAEBFFEFAA803DEBA5D2E82155A2FBF",
INIT_3A => X"A95545F7D5555FFAAAAA8BFF002AAAA00FFAAA8AAA080028BFFF7D568BEF0804",
INIT_3B => X"2E95400A2AEA8A00007FEABFF00042ABFFA2FFFFF45F7AE97400AAFFE8B45AAA",
INIT_3C => X"82E820BA08556AA00AAAABFE00F7AEAABEF082E9554508557DFFF007BD54BA5D",
INIT_3D => X"A2D57FE00552EA8A00FFFFE8AAAAA80001FF5D2E82000F7FFFFF45AAFFC20BA0",
INIT_3E => X"0000000000000000000000000000000000000FFFBD5400082EBFF45F78400155",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(1),               -- Port A write enable input
DIA(0)   => data_write_a(11),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(11),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(1),               -- Port B write enable input
DIB(0)   => data_write_b(11),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(11),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_12_9 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50080B01BC002006940202C0DE041196A83183000000023322287E0FC000006",
INIT_01 => X"75400D849830C84C5823E0000C17424840000000080000088200002802153231",
INIT_02 => X"18A026B43ED180040147558040090000061800000C06ED9802768F4472C52005",
INIT_03 => X"2A67E34A528D0524A52850528400C8001100000171C02B550618C91A10E55440",
INIT_04 => X"1BC0000100056C8280825DE98154004300C840800850240080CA921084520A07",
INIT_05 => X"02000F832000500C0000941024000852084060202E100001002000448100000C",
INIT_06 => X"819A1D1C3FE01A1A40045408049A50BA4020C6041090001200006200000000F2",
INIT_07 => X"C26A0719CC96CC6ED18A64019695A854870300FA3968B20068FC06080106249F",
INIT_08 => X"D002024B3E040800008C0A002610240D494A06F3460409000000E3F0AD5282E5",
INIT_09 => X"27A06009200040000400120412445D78400001000410420080218029CC807A27",
INIT_0A => X"18000006848A026F000000000000080000F010C100204593F11A6CDF48003BF8",
INIT_0B => X"000000820040402B28050400400432C9349DF21A31A00ACC0000F04F80020001",
INIT_0C => X"00357804611AE45D05D0833430CD0833420CD0C33420CD0833430668619A1000",
INIT_0D => X"0000000000000A74812DF00E87E80A079F9F90FA0280E87E800C7FF3B8002000",
INIT_0E => X"3B6B0E404D26160682082002000401EA0000C40000800A006002818808000000",
INIT_0F => X"A476D61C809A4DA84272592D6246FC1B17B541F97E1B348EDA93900B2B286C56",
INIT_10 => X"30C669E622DBC325CFD881A962454CFBE5403AB99594362B1DB52720165650D9",
INIT_11 => X"F8D2D39A3745261E4A95A110A3F855000E4B1D32BAB504BB7490FCFF912A3834",
INIT_12 => X"B90E9B018C7530200AB8F8BF41F9A22006B37DC8E1F9A21A70116D4C5080651C",
INIT_13 => X"118780319CCA08AB1001ACDF34B8F1C688AB1002AE3F7B807B6289F368828C4C",
INIT_14 => X"2AF020233376A5ECC016B1A827CDA21160F051DE610A34C50427E6E220323E4A",
INIT_15 => X"0077020000000439FDC05C5806781FAB46095A0B5199B0AC55521524F1864022",
INIT_16 => X"000000000000000000000000000000000026C000002884000130921092804010",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"8020080200000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0051B946088881360A95090CB054420290100000000000000000008020080200",
INIT_1A => X"041041041041041041041041041041041049249249249249200100002D451451",
INIT_1B => X"92C964B2592C964B2592C964B2592C964B2592C86432190C86432190C8641041",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000003800F592C964B2592C964B25",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"7DE1000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"ABDFFFF7803DE10AA80000AAAA843FE0008557DFFF0800020105D557FEAA0055",
INIT_29 => X"D5420000051555FFA2AA8200000557DFFFF7AA80000082ABDF5508557DF45002",
INIT_2A => X"82AA8AAAAAFFC00BA007FC2155F7D155545AA80001EFAAFBEAB45557FFDE10AA",
INIT_2B => X"FFAEBFEAA002A801FFF7FFE8A10A28000000A2D155410F7FFFFEBA08003FE000",
INIT_2C => X"5FFFFEAABA000028A105D2ABFE10A2AABFE1055516ABEF5D517DEAAA2AEBFF45",
INIT_2D => X"55002A820AA08557DFFFF7AA82155AAFBE8B45002A974AAAA803DFFFAA843DF4",
INIT_2E => X"000AAD155555A28428BFF002ABDE00A2AABFE10082ABFFEF0855420000004175",
INIT_2F => X"5010495B7AE921C517DE10000000000000000000000000000000000000000000",
INIT_30 => X"BDF6D005B78F7D142ABDFC7F78E3FE28B684070AABE803AE38145B78FD700000",
INIT_31 => X"BEFB455D71F8E00BED547038145B505FFB6A487000005F7AFD7F7A482038002E",
INIT_32 => X"F1FDE821C003FE001C2EAAAAAB6F5C2082007BC217DEBDB55555AA8E071D7AAF",
INIT_33 => X"D517DEAABEAEBFF7DEBA0BDEAA1C2A801C7E3FFEFA10B68407038B6D550428FF",
INIT_34 => X"B68E38FC7BE8A3DF7DF7F5E8A9200002FA285D20BDE28A2A4B8E10555B68BEF5",
INIT_35 => X"F085F47038140010555142082082005F7DFD7F7A482155BEF1E8B6D002090482",
INIT_36 => X"00000000000000000000B6D15756DA28A28BFF082ABAE10B6AAB8E280820B8FE",
INIT_37 => X"ABA5D7FEAB45080015410007FEAA0055517DE000000000000000000000000000",
INIT_38 => X"AB45F780020BA082EBFFEF007BE8BFF5D2ABDF55F7AABDEAAF784154BAF7802A",
INIT_39 => X"D7545AAAE97555A2FBFDF455D556AA00F7D1554BA5D7BC01FFFF8015410007FE",
INIT_3A => X"4154BAF7D1400BAFFD57FE005D043FE10552EAAAAAFFD140000087FC01EFA2FF",
INIT_3B => X"8428A105D7FEABEF55557DEBAFFAEBFFEFAA803DEBA5D2E82155A2FBFDE00FF8",
INIT_3C => X"7D568BEF080402000F7AAA8B55FFAABDFEFF7D16AA0008003FEBA55003DEBAA2",
INIT_3D => X"FFAAA8AAA080028BFF087BD54AA550402145550000010087FFFF45F78402145F",
INIT_3E => X"0000000000000000000000000000000000000F7D5555FFAAAAA8BFF002AAAA00",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(1),               -- Port A write enable input
DIA(0)   => data_write_a(12),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(12),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(1),               -- Port B write enable input
DIB(0)   => data_write_b(12),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(12),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_13_9 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10154A0441836CA2840512822007C18000E02700500030B31B300040081A042",
INIT_01 => X"00000804A000C04800020000000002404001000008220008A200100802110204",
INIT_02 => X"02200430000104000A4700804008000004100000000420918204D3033240400D",
INIT_03 => X"AA4003400008592400000590C40009141100000C6180C0000000C00001E14000",
INIT_04 => X"0800000102400120088054019000004160004190BAA0270000C8100000600206",
INIT_05 => X"21000012040610050040000227003AA0082400E94C1200000824424005220020",
INIT_06 => X"81963B180C001010580000080400000058000004109C00138000020024142581",
INIT_07 => X"002C8008000441600106400A9600010494020002B8AAA000EF003408000E2580",
INIT_08 => X"000000E48194408000A00A001210040441C80320040210000002ABF004102244",
INIT_09 => X"2A004009640040100400940412D4C4004000022000104200802D983000480120",
INIT_0A => X"8000202020401480000000000000080C90090881000145B0111A14004015080D",
INIT_0B => X"00000002004040AA08050400404040C11444000805200A402090024000008002",
INIT_0C => X"8410000A00280020020040800020040800020000801020000800010020400000",
INIT_0D => X"84A14250A055100050100490000500D00040080040290000084E4000B800610C",
INIT_0E => X"DCD13042BEDA36820228000000000000C000400081A08BC812A2092B02850942",
INIT_0F => X"89B9A260857DB400431969CA985D480949D32804A40AB137341C10B7D6A02EC0",
INIT_10 => X"E6ACA678001CE7D0296C213A460CA4271CA2168AEC1017606E6838216FAD4055",
INIT_11 => X"84AD4961C281B20213073C5FC0058008632D30D522CE80239DCC01AB013A4D20",
INIT_12 => X"2E6B13804A4B01D83461299900F6BD583A519104A0EEBD1A141010B2A4C8E116",
INIT_13 => X"89E5E40913419151EE0E94641828F72B5151EE0D184B321037AF5158BB02D085",
INIT_14 => X"562EC0B42162D68EE0073AE1C562EC13D521921A4170300B2B458B56B01C2280",
INIT_15 => X"00888A120240034000E6DC8285028014B82372011FC1E4F5E0A00929684EAF84",
INIT_16 => X"50942509425094250942509425094254940A1421420082020120908800480030",
INIT_17 => X"0942509425094250942509425094250942509425094250942509425094250942",
INIT_18 => X"9425094250942509425094250942509425094250942509425094250942509425",
INIT_19 => X"F7EFBBEEFF3F7DF7FF3E9F7DF7E2450228000000000000000000509425094250",
INIT_1A => X"BAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBF7DFDFDDD555555",
INIT_1B => X"EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAEBAE",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000000000F7EBF5FAFD7EBF5FAFD7",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"2ABEF00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0020105D557FEAA00557DE10AAD5554BA087FFFF55557BD54AAF7FBC01FFA280",
INIT_29 => X"7BD75EF087FFFFEF557BEAB45552E80155AA802AB45AA843FE0008557DFFF080",
INIT_2A => X"FAE820AA5D5557555082ABDF5508557DF45002ABDFFFF7803DE10AA80000AA08",
INIT_2B => X"0051555FFA2AA8200000557DFFFF7AA80000AAD1420AA087BD7555FFD168AAAF",
INIT_2C => X"5557FFDE10AAAEA8BFFA2FBD7545FFD157555085140010F7AEAABFFAAD542000",
INIT_2D => X"BA557BE8A10A284154BAFFAAAAB45007FC2155F7D155545AA80001EFAAFBEAB4",
INIT_2E => X"000A2D155410F7FFFFEBA08003FE00082AA8AAAAAFFC00BA00002AAAAF7D5574",
INIT_2F => X"0492E3F1C71C7BE8A2ABD7000000000000000000000000000000000000000000",
INIT_30 => X"3AE38145B78FD7000005010495B7AE921C517DE10A2DB50482147FFAF554971D",
INIT_31 => X"E3FE28B684070AA1C71D25D7007FFAFD7497BE8B5555208217DBE8A2AB45BE80",
INIT_32 => X"7FD257DFFD568A82FFA4870BA555F5056D002EBDF6D005B78F7D142ABDFC7F78",
INIT_33 => X"FAAAFBFFBED547038145B505FFB6A487000005F7AFD7F7A482038AADF4709214",
INIT_34 => X"AA8E071D7AAFBEFB455D71F8E00A2A0ADBC7A2FFD257DE3DF52555085142000F",
INIT_35 => X"21C002AA92FFDF574824171EAA10B680124BAFFAAAFB45007BC217DEBDB55555",
INIT_36 => X"00000000000000000000B6D550428FFF1FDE821C003FE001C2EAAAAAB6F5C208",
INIT_37 => X"0105D7BE8B55085142010AAD157545F7AEA8B550000000000000000000000000",
INIT_38 => X"01EFF7AAA8B55F7802AABA5D7FEAB45080015410007FEAA0055517DE00A2FFC0",
INIT_39 => X"E8BFF5D2ABDF55F7AABDEAAF784154BA5D5140145007BE8B55087BEAB555D040",
INIT_3A => X"0020BAA2FFD54105D7FC21EFFFD16AA10FF80174AA557FC21EF082EBFFEF007B",
INIT_3B => X"FBC0155085540000FFAEBFFEFF7D1554BA5D7BC01FFFF8015410007FEAB45F78",
INIT_3C => X"87FC01EFA2FFD7545AAAE97555A2FBFDF455D556AA00A2803FF45AAFFC21EFAA",
INIT_3D => X"552EAAAAAFFD1400005D042AA00F7FBD5410085568A10FF80020AAFFAABFF550",
INIT_3E => X"0000000000000000000000000000000000000F7D1400BAFFD57FE005D043FE10",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(1),               -- Port A write enable input
DIA(0)   => data_write_a(13),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(13),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(1),               -- Port B write enable input
DIB(0)   => data_write_b(13),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(13),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_14_9 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10020A000180000284008280000281800000030000000033022000000580002",
INIT_01 => X"000008020000204D006800000030824840000000084000084200090008510200",
INIT_02 => X"0220043170010A600A4D008040080000041000000028009002000F333240800C",
INIT_03 => X"111813400008002400000000C400090011000000610200001104D83000F14000",
INIT_04 => X"0801800100A000000000540084000040000040000800200000C8100000000748",
INIT_05 => X"0100000000001000000000002000080008000000001000000024024001200020",
INIT_06 => X"819EB84028001010000000080400000000000004108000100000020020040081",
INIT_07 => X"92040608000440100102400A94810206844200021DA2A0002000340800062C80",
INIT_08 => X"000000000084400008800A001214040441481500040000000000A7F408002244",
INIT_09 => X"0A0040090002008420401004104444004000020400214A208001000002400120",
INIT_0A => X"0400002020000000000000000000080C8008088100004590111B480040120000",
INIT_0B => X"1000000200404800000504016000002114000008020000020080024000000000",
INIT_0C => X"0410000010000000000040001000000000000040000000000001000000000000",
INIT_0D => X"04810244825010004010000000000000000000000000000000080000B8002104",
INIT_0E => X"0002C38280001202020800000000001000004000000000401022000002040902",
INIT_0F => X"20000587050001404E8084341CBA3404800828805200008000E0E0A000080002",
INIT_10 => X"4D18178E012010C00224004091C3514072C000444A0400080001C1C140001000",
INIT_11 => X"51709A07424142084458476001003809D0104B01C5710044020C4006010500C5",
INIT_12 => X"C26EE3803180C18006519462A00005001460E4730000050A1011004001060049",
INIT_13 => X"01F9E00660318000000538318740000140000001B4600CE80001400000002B62",
INIT_14 => X"0000000AD89857B0E0684411800000003799EB764D000330C300000000E3554B",
INIT_15 => X"0000021002002C000024008284001A0902000422E3F5960080480A0216A07240",
INIT_16 => X"4090240902409024090240902409024090081021020080015134920800480010",
INIT_17 => X"0902409024090240902409024090240902409024090240902409024090240902",
INIT_18 => X"9024090240902409024090240902409024090240902409024090240902409024",
INIT_19 => X"F5579B4E5C8FF0F7BE9D5F7DF650400200000000000000000000409024090240",
INIT_1A => X"9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7BF7DDDDDFCF3CF3D",
INIT_1B => X"F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE79E7",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000003FFF03F9FCFE7F3F9FCFE7F3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"420BA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"BD54AAF7FBC01FFA2802ABEFA2FBE8B55A2AE80000F7D5555555D2AAAABAAAD1",
INIT_29 => X"AA801FFA28402000AAAE955455500155EF0804155EFAAD5554BA087FFFF55557",
INIT_2A => X"7AEA8B45080417400AA843FE0008557DFFF0800020105D557FEAA00557DE10A2",
INIT_2B => X"087FFFFEF557BEAB45552E80155AA802AB4500516AA00A2AE800BAFFFFC20BAF",
INIT_2C => X"0AA80000AA005568ABAA28402010A2843FEBAFFFBD7410A2D168BFF087BD75EF",
INIT_2D => X"005D7FFDF4555517DFEF00043FEAA082ABDF5508557DF45002ABDFFFF7803DE1",
INIT_2E => X"000AAD1420AA087BD7555FFD168AAAFFAE820AA5D5557555002E80155A280000",
INIT_2F => X"0555412AA8ABAAADB40092000000000000000000000000000000000000000000",
INIT_30 => X"50482147FFAF554971D0492E3F1C71C7BE8A2ABD7A2FFEDB55B6A080038E3DB5",
INIT_31 => X"B7AE921C517DE10A2AE851FFB68402038AAAA955554900105FF0800175D7A2DB",
INIT_32 => X"A0800BAE3F1C0092EBAAADB6D080A12410BE803AE38145B78FD7000005010495",
INIT_33 => X"2D568BC71C71D25D7007FFAFD7497BE8B5555208217DBE8A2AB451C556FA00A2",
INIT_34 => X"142ABDFC7F78E3FE28B684070AA00516DABAA28402038B6803DE82F7F5D5410A",
INIT_35 => X"D002A80155B680000105D7FF8F455D5F78FD7000E3FEAA002EBDF6D005B78F7D",
INIT_36 => X"00000000000000000000AADF47092147FD257DFFD568A82FFA4870BA555F5056",
INIT_37 => X"F55FF84000AAAAFBC0145002AA8AAAAAFFC20000000000000000000000000000",
INIT_38 => X"01EF080417555A2FFC00105D7BE8B55085142010AAD157545F7AEA8B55A2FBFF",
INIT_39 => X"EAB45080015410007FEAA0055517DE00A2AA955FFFF80020BAAAAA9754508000",
INIT_3A => X"AA8B555D557FE00A280020BAAAD140000A2AEBFFEF082A82010F7802AABA5D7F",
INIT_3B => X"803DE00FFD557400AAD56AB455D5140145007BE8B55087BEAB555D04001EFF7A",
INIT_3C => X"82EBFFEF007BE8BFF5D2ABDF55F7AABDEAAF784154BA08557FEAAA284000AAFF",
INIT_3D => X"FF80174AA557FC21EF082A80145F780020105D7BEAB45557BE8B45082EBFEBA0",
INIT_3E => X"0000000000000000000000000000000000000A2FFD54105D7FC21EFFFD16AA10",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(1),               -- Port A write enable input
DIA(0)   => data_write_a(14),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(14),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(1),               -- Port B write enable input
DIB(0)   => data_write_b(14),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(14),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_15_9 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000A000000000284000280000001800020030000000033022000000180002",
INIT_01 => X"8000080000000048000000000000026040000000080000080200000000110200",
INIT_02 => X"0020042004010E60004C0080000800000410000000020090020000300245E005",
INIT_03 => X"0000010000080400000000408400480111000000610008000000C00000E54400",
INIT_04 => X"980000010000000088C2550080000040000040000008A00028C8100000120000",
INIT_05 => X"020004012E025000000001322000000A28008000011000000220004D41000000",
INIT_06 => X"819588000800101000011008040000100001060418800510000A620000000092",
INIT_07 => X"0000000800044004010C20008440810284020002102220002000340800062480",
INIT_08 => X"0000000001140800002C0A001214050540C800400406180000002DF004000244",
INIT_09 => X"1E00400900000000000016041044400440000000000042008001000000000022",
INIT_0A => X"0000000000000220000000000000080C00000081000045901118000040000000",
INIT_0B => X"0000000200404000010500004000000114000009000000000000004200000000",
INIT_0C => X"0000000000000000000040001000040001000000000000000001000020000800",
INIT_0D => X"000000000000001001208000180800000000030200000180800C400030002000",
INIT_0E => X"0000000000002600020800000000001080004000000000000002000000000000",
INIT_0F => X"A400000000000000000008000000000000000000000014800000000000000052",
INIT_10 => X"0000000000000000000000010240000000000000000000290000000000000000",
INIT_11 => X"2001C05838120800000000000000000000010000000000000000000000001804",
INIT_12 => X"081004000000000000A010000000000000902000000000180010002020000000",
INIT_13 => X"6600000000000000000024080000000000000000280400000000000000000000",
INIT_14 => X"0000000000200801000000000000000000501001920000000000000000000A40",
INIT_15 => X"0000020000000000000000003000000000000000000A101C3614000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000080000120980000000010",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000400200000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"28BEF00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"5555555D2AAAABAAAD1420BAFF8000010082A954BA00003DFEF085155400F784",
INIT_29 => X"AE95555A2FBE8BEFA2843DE00AA8015400FF84001EFA2FBE8B55A2AE80000F7D",
INIT_2A => X"2FBEAB45F7D56AABAAAD5554BA087FFFF55557BD54AAF7FBC01FFA2802ABEFF7",
INIT_2B => X"A28402000AAAE955455500155EF0804155EFFFFBE8BFF0800174AA557BFDE10A",
INIT_2C => X"A00557DE10F7D1574AAA2D16AB55FFD568BEF087FE8A1055003FE00A2AA801FF",
INIT_2D => X"00AA802AA00AAAE800BA5D0015545AA843FE0008557DFFF0800020105D557FEA",
INIT_2E => X"00000516AA00A2AE800BAFFFFC20BAF7AEA8B45080417400FFFFC21450800154",
INIT_2F => X"8FD7005150438F78A2DBFF000000000000000000000000000000000000000000",
INIT_30 => X"EDB55B6A080038E3DB50555412AA8ABAAADB40092E38E070280024904AA1C043",
INIT_31 => X"1C71C7BE8A2ABD7E3AA9257DA2FFE8BC7BE8E38E10A28017400E38A051FFA2FF",
INIT_32 => X"00124AA557FFDE10A2FBEDB6DF7D16AABAA2DB50482147FFAF554971D0492E3F",
INIT_33 => X"10038E38A2AE851FFB68402038AAAA955554900105FF0800175D7E3FFEFBD700",
INIT_34 => X"000005010495B7AE921C517DE10FFDF50482A2DB6AB45FFD56DBD7087BEAA384",
INIT_35 => X"0FFF1C017D140410400BE8E28A10AAA085082550A1057DBE803AE38145B78FD7",
INIT_36 => X"000000000000000000001C556FA00A2A0800BAE3F1C0092EBAAADB6D080A1241",
INIT_37 => X"4AA0800020BA550028B550855400AAF7AEBDFEF0000000000000000000000000",
INIT_38 => X"7400AAAE975EFA2FBFFF55FF84000AAAAFBC0145002AA8AAAAAFFC2000AAAA97",
INIT_39 => X"E8B55085142010AAD157545F7AEA8B55AAAE821EFAAFBEAB55F7AAA8A00AA841",
INIT_3A => X"417555AAFFFDF450804020AA557BFFE10A2FFFFFEFF7D568ABAA2FFC00105D7B",
INIT_3B => X"D17DF45007FE8AAA08002AAAAA2AA955FFFF80020BAAAAA975450800001EF080",
INIT_3C => X"7802AABA5D7FEAB45080015410007FEAA0055517DE00FFFBC2000AAFBE8B55F7",
INIT_3D => X"A2AEBFFEF082A82010FFD5421EF5D0000010F7AAA8A10AA8017400552A801EFF",
INIT_3E => X"00000000000000000000000000000000000005D557FE00A280020BAAAD140000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(1),               -- Port A write enable input
DIA(0)   => data_write_a(15),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(15),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(1),               -- Port B write enable input
DIB(0)   => data_write_b(15),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(15),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_16_9 : RAMB16_S1_S1
generic map (
INIT_00 => X"DA22C618B1000482B688B186588884862A400438255FC38381441205BA803003",
INIT_01 => X"7045A80028404C211203A952A90341080B173340412000E1005D628000820484",
INIT_02 => X"428406A4000850848330118D0AAC55001349B108818005460229044001C01784",
INIT_03 => X"092C4020000500020000500986812C405000001A48202050000A214AC0650115",
INIT_04 => X"4804A55440256F504025E003A054F46415A4E62B6FE3307943965A00001A1152",
INIT_05 => X"0000001C40A5B950ADB8EA097057ECE14C86D2B7F85AAD17F4B100000B88148C",
INIT_06 => X"415401DCDCF2C0A8030140BCB0820A200342A1C641C1E8782F508F2B00003584",
INIT_07 => X"002701881A3202080AE00480A2002840BE1480FA004342AA6F12000054004867",
INIT_08 => X"08C54828091002000002B32A8C19064E486A8001510000014140C1E2A14891E0",
INIT_09 => X"015452B103020814004088B64102680B6596594800400413CAC0208944800000",
INIT_0A => X"96AA000484094C000000000000012C9000A0000D0A80000BF8028E87C1B99270",
INIT_0B => X"014808A02004200E540480212000A448C0082024AE50064B44000000000002A2",
INIT_0C => X"0004000D5846256AAEA811150445411150445411150445411150422A088A8200",
INIT_0D => X"00000004010042A204A0C5817D00005034052E40000817D00440004004AD3240",
INIT_0E => X"632B2673FA4587978A2004102800809225545155121740000004900090000000",
INIT_0F => X"00C6564CE7F4EA4B940076D296D003030800462CBD320018CAAAACFE9164C800",
INIT_10 => X"28834ADB1440A114793A4A30A40839AA14910D08DCB2640031955559FD3AC990",
INIT_11 => X"594AB0B1A025371CA0E034E8443C097A800EB090D4AAC91208ED2FA0CE5E09B1",
INIT_12 => X"7B50446083001B94BB38C540EBE61284BB304880E3E4579EDC00992980D58033",
INIT_13 => X"5511121840E7A2CD952ECC12ABC3E6ACB3DFB12ECE315000F61FF1727A85FDBC",
INIT_14 => X"75DEB07F6F2E7084517F126F8395CB2BEFBAB8BA8AF698228CC5E2F08ECA5159",
INIT_15 => X"5580A840A8009F8B108C80A1021B080AFC0DF6422C6077F4A77F20D0C0E21084",
INIT_16 => X"0000000000000000000000000000000000044000102A0001148442A110810359",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"558D11544C690DA64C1C4F68A360400000000000000000000000000000000000",
INIT_1A => X"14D14D14D14D14D14D14D14D14D14D14D14514514514514529E5F87869E79E78",
INIT_1B => X"D1E8F47A3D1E8F47A7D3E9F4FA7D3E9F4FA7D3E9F47A7D1E9F47A7D1E9F4D14D",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000007D3E9F4FA7D3E8F47A3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"C00AA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"03DFEF085155400F78428BEF087FFFFEFF7D168B55AAD17FFFF552EBFE00007F",
INIT_29 => X"2E975EFF7D568BFFFF80175EF0004000BA552A821FFFF8000010082A954BA000",
INIT_2A => X"55540000082EAABFFA2FBE8B55A2AE80000F7D5555555D2AAAABAAAD1420BA5D",
INIT_2B => X"A2FBE8BEFA2843DE00AA8015400FF84001EF0000020AA5D00154005D043FF455",
INIT_2C => X"FA2802ABEF557BEABEF5D0415410087FD74BAAAAEBFFEF557FC00AAF7AE95555",
INIT_2D => X"FFFFAABFEAAFF84001FF002A821FFAAD5554BA087FFFF55557BD54AAF7FBC01F",
INIT_2E => X"000FFFBE8BFF0800174AA557BFDE10A2FBEAB45F7D56AABA082A97545F7D16AB",
INIT_2F => X"FFEF552AB8E38087FC2092000000000000000000000000000000000000000000",
INIT_30 => X"070280024904AA1C0438FD7005150438F78A2DBFF0871F8FC7E3D56AB6DBEDB7",
INIT_31 => X"AA8ABAAADB400924920925EFF7D16ABFFE38E175EF1400000BA412E871FFE38E",
INIT_32 => X"0A1240055003FF6D5551420101C2EAFBD7A2FFEDB55B6A080038E3DB50555412",
INIT_33 => X"57FC00BAE3AA9257DA2FFE8BC7BE8E38E10A28017400E38A051FF0804050BA41",
INIT_34 => X"4971D0492E3F1C71C7BE8A2ABD74975EDBC7550E12410087FD74AAB6AABFFC75",
INIT_35 => X"A08249756DF7D168BC7F7AABAEAAF780051C70824851D7A2DB50482147FFAF55",
INIT_36 => X"00000000000000000000E3FFEFBD70000124AA557FFDE10A2FBEDB6DF7D16AAB",
INIT_37 => X"B55A2D16ABEFFFFBFDFFF552AAAAAA007BC00000000000000000000000000000",
INIT_38 => X"20AA002A955EFAAAA974AA0800020BA550028B550855400AAF7AEBDFEF08516A",
INIT_39 => X"000AAAAFBC0145002AA8AAAAAFFC20000000021EFF7D568BFFA2AA955FF5D040",
INIT_3A => X"E975EF0800174BA002E820105D003DFEF5D51420005D2ABFF45A2FBFFF55FF84",
INIT_3B => X"7BD74AAF7AEBDF455D7BC20BAAAAE821EFAAFBEAB55F7AAA8A00AA8417400AAA",
INIT_3C => X"2FFC00105D7BE8B55085142010AAD157545F7AEA8B5500557DF45552A8200000",
INIT_3D => X"A2FFFFFEFF7D568ABA0804155FFF7D568B55FFAAAAABAFF8415545000015555A",
INIT_3E => X"0000000000000000000000000000000000000AAFFFDF450804020AA557BFFE10",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(2),               -- Port A write enable input
DIA(0)   => data_write_a(16),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(16),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(2),               -- Port B write enable input
DIB(0)   => data_write_b(16),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(16),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_17_9 : RAMB16_S1_S1
generic map (
INIT_00 => X"5284CE4FB7BD2C8994A13392DBD02E14006B82AC7E800D44D3DD2FD5F9B961C0",
INIT_01 => X"2EACD01F7E03FC6793F2199B39FC233C11D93AE6F3BB92B32091DBC339B24542",
INIT_02 => X"E63CCCC00A82C08092A2AFAE667033DB50853379C10BFDC5C6F4044443C817C6",
INIT_03 => X"7FF183635AEF9E3635AEF9E18E237040404446965C0607EE6DB7854AC4DE060C",
INIT_04 => X"D78AC33FB604488B000892EF17BE6D84196482236FE100294152E294350FB697",
INIT_05 => X"081B5F9B409420D0CDB47A05403F6CE0C08A4AB7F840EDB6F48100DFC8081081",
INIT_06 => X"768465354781CBC30316367077B4BDB50646E8D87100A8201ED01C19C020F71A",
INIT_07 => X"4002A110C922480A82D0841147162C48EBB9537A0022DC67987042EE976ABEA7",
INIT_08 => X"DB931BFEF91C00002CC0E019C0C82A4E4820C15A2330E004401891181168C4D1",
INIT_09 => X"09F3A1BC11EFBC66DB65307071477FF1030C397C060B4254064302042F803A69",
INIT_0A => X"3F330802162F3B7EE3F3EC7C7DEF207000F00059D2ED56D7EED2ED3C9A867DC0",
INIT_0B => X"185C44B91BC1740B7605040BE0018CFC7429F326B9E822FFC00074D5A0AB033A",
INIT_0C => X"00367A28FC1B7F7FEFFCFBFF3EFFCFBFF3EFFCFBFF3EFFCFBFF3EFFE7DFF9E00",
INIT_0D => X"0000000008004BA78428C7AD7FC94B533F5B4FFBD2FAD7FCCA786D43FE67C218",
INIT_0E => X"BA494CEBFD4F2667ABB6F68B29760593F33FA0CF170F40006001B1A05C000000",
INIT_0F => X"7F749299D7FAEB237DFE5865B6D2BF23265CBACE542A6FEE92333AFF33E0A9BF",
INIT_10 => X"F6C24B6D18C3C9F8E2881F3F787D776B5DB94A09955054DFDD246675FE7AC153",
INIT_11 => X"BFB349E08FF9A27EDE9FA8AEFD9E7467BFCB195CFEB56A1A70D34D1706FFFA3E",
INIT_12 => X"6FE219CA80725B875EED723FF7FCB2875EDAAFEAF7FD929BFD55BBC71D79F639",
INIT_13 => X"546670D018E7A6E581D7B6AB75FDFCECA6E581D7BB5DDFC6FF0EB7D7E859FDB5",
INIT_14 => X"B978177F6D6AF5ECDB5FB76A5F5FA165B456E0FB308710C49FCFB741598B9C7E",
INIT_15 => X"CFDAAB00AC00A8BBFC8B501CF7A0FED9A540EA1952586CEB54D143ACFF9A3BA9",
INIT_16 => X"000000000000000000000000000000000026E100002F382DBD9ECFE117805F20",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"4372003009EDCC4052E917114F981800C0000000000000000000000000000000",
INIT_1A => X"BA69A69AEBA69AEBA69A69AEBA69AEBA69A69A69A69A69A68698686981D75D74",
INIT_1B => X"6A351A8D46A351A8D068341A0D068341A0D068341A0D46A341A0D46A341A69AE",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000000000046A351A8D46A351A8D4",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"7FEAA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"17FFFF552EBFE00007FC00AA087FFFFFFFFFFFFFEFF7FBEAB450804001EFAAD5",
INIT_29 => X"D168A000004020AA5D7BE8B450051401EF087FD74AA087FFFFEFF7D168B55AAD",
INIT_2A => X"D7FEAB55FF80175EFFF8000010082A954BA00003DFEF085155400F78428BEFAA",
INIT_2B => X"F7D568BFFFF80175EF0004000BA552A821FF5D00020BA552A82000552A821555",
INIT_2C => X"AAAD1420BAFFFFFDF45AAD17FFFFAAFBC01EF5D0015555557BFDEBA5D2E975EF",
INIT_2D => X"BA007FEABEF005555555A2D1554BAA2FBE8B55A2AE80000F7D5555555D2AAAAB",
INIT_2E => X"0000000020AA5D00154005D043FF45555540000082EAABFF00516AA10552E820",
INIT_2F => X"8B550000071EFB6DF7AE92000000000000000000000000000000000000000000",
INIT_30 => X"F8FC7E3D56AB6DBEDB7FFEF552AB8E38087FC2092147FFFFFFFFFBFDFC7EBF5E",
INIT_31 => X"150438F78A2DBFFBED16AA381C0A07082497FEFB6D1451471EF007BD04920871",
INIT_32 => X"2A850105D2A80155417BEFB6DEB8E175FFE38E070280024904AA1C0438FD7005",
INIT_33 => X"D7BFAEBA4920925EFF7D16ABFFE38E175EF1400000BA412E871FF550A0009249",
INIT_34 => X"E3DB50555412AA8ABAAADB40092FFF5FFF6DAADF7FFD7B6F1C71EF55001756D5",
INIT_35 => X"7145B6AA28492487082007FEDBD700515556DA2DF50492A2FFEDB55B6A080038",
INIT_36 => X"000000000000000000000804050BA410A1240055003FF6D5551420101C2EAFBD",
INIT_37 => X"FEFF7FBFFF55A2D16AB550000175EFFFFBEAA000000000000000000000000000",
INIT_38 => X"55EF087FC200008516AB55A2D16ABEFFFFBFDFFF552AAAAAA007BC0000557FFD",
INIT_39 => X"020BA550028B550855400AAF7AEBDFEFF7D568AAA5D2A97410007BFFFFF55515",
INIT_3A => X"A955EF5D2E80010002A954005D2A82155087FFFFEFAAAA975EFAAAA974AA0800",
INIT_3B => X"D1575FF5504175EF5D7FEAAAA0000021EFF7D568BFFA2AA955FF5D04020AA002",
INIT_3C => X"2FBFFF55FF84000AAAAFBC0145002AA8AAAAAFFC2000FFD57DFFFAAFFFDF55FF",
INIT_3D => X"5D51420005D2ABFF45557FE8AAA000415410007BFFF450051555EFA2FBC0000A",
INIT_3E => X"00000000000000000000000000000000000000800174BA002E820105D003DFEF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(2),               -- Port A write enable input
DIA(0)   => data_write_a(17),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(17),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(2),               -- Port B write enable input
DIB(0)   => data_write_b(17),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(17),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_18_9 : RAMB16_S1_S1
generic map (
INIT_00 => X"69844019080000A21A611406840014122A641074155FC28A2024001001801003",
INIT_01 => X"7443D920034004180005E9E3C90360C0041C0181002001602025800008440084",
INIT_02 => X"E2DCCCE61D5C008103F2000781FC0FEDEAC2161B0B8FB0008620044443006010",
INIT_03 => X"884E300802006900802006995C896D605200000856E24A040000640052141103",
INIT_04 => X"480520FC026125AC0025C9122644E3E40EC8E2001001302281841A009038A86A",
INIT_05 => X"432000040089983070019400F01010004C8DB841405A80A100B586200FAC24AE",
INIT_06 => X"09044359DC7040000000002C109B0E0A00A1104641C0803804000707284600E1",
INIT_07 => X"400D10100400481D5EB08501620000007500CE801241021FE78E404860140060",
INIT_08 => X"00880C0106A0528020019307CC082A0A4A6A01ED725021400040D028000A9729",
INIT_09 => X"00117063038000282081402E4106400B6186128040600C10C1C0200950508110",
INIT_0A => X"C0C30C2E21580C874004008080003C32A10A19090C02010E1022944061688000",
INIT_0B => X"0180A8062026000DC425C0301311324AA2373088479105D044A1022000001835",
INIT_0C => X"0D89844703649000000200000000000000000000000000000000000000000010",
INIT_0D => X"0D8306C182701404C1973010802020404084001E00010802046092B5001FB365",
INIT_0E => X"528EB314068AB8B803DB00002900800400FC503F08180050942E4200020C1B06",
INIT_0F => X"40A51D66280D6032C5F96D3C51555D5D7D5AA87285820814A3CCC501C2A60820",
INIT_10 => X"8B35A3FEBF1FEDFD9C2B30E0468AAAD5D48F37E8FC1304102947998A03984C10",
INIT_11 => X"440FE1DD772D37A0A321BC6968F32658BF2D4F2A80BF8FE3F9FE3AC362080529",
INIT_12 => X"5487910D7E5A6D961A28456A1832E5161A100DD5182BC54020EA67A189C6ED36",
INIT_13 => X"AA444CAF91EDD1B725868403BE06323551B725868A100ABD119753B70964122B",
INIT_14 => X"EDC259048ACD868EE3803D65CEDC258A8F80D55E007C3F8EBB56F4C5362C978F",
INIT_15 => X"3F240014BE84370001B6922070440556B15F7FABBC0031BCF2257C41634B14D4",
INIT_16 => X"C1B06C1B06C1B06C1B06C1B06C1B06C1B0491069068000004060300A005A0118",
INIT_17 => X"1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06",
INIT_18 => X"B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C",
INIT_19 => X"B28BBECEB80EE173C2300F7DF16000000000000000000000000041B06C1B06C1",
INIT_1A => X"8A28A28AAAAAAA28A28A28AAAAAAA28A28A28A28A28A28A2910591505C104104",
INIT_1B => X"28944A25128944A25128944A25128944A25128944A2552A954AA5128944AAAA2",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000128944A25128944A251",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"9540000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"BEAB450804001EFAAD57FEAA087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974BA082E",
INIT_29 => X"7FFFFFFFFFBFDF45AAD568B55080028B55002E82000087FFFFFFFFFFFFFEFF7F",
INIT_2A => X"0043DE10AA843DE00087FFFFEFF7D168B55AAD17FFFF552EBFE00007FC00AA08",
INIT_2B => X"0004020AA5D7BE8B450051401EF087FD74AAAAFFFDF45A2D16AB55F7FFFFFFF0",
INIT_2C => X"0F78428BEFAA80000000804154BA55042ABEF5D7FD75FFAAD540145AAD168A00",
INIT_2D => X"00082E95555085168A10557FD7545FF8000010082A954BA00003DFEF08515540",
INIT_2E => X"0005D00020BA552A82000552A821555D7FEAB55FF80175EF5D00020105D2A974",
INIT_2F => X"DFFF5D2A954AA082A92428000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFBFDFC7EBF5E8B550000071EFB6DF7AE921C7FFFFFFFFFFFFFFFF7FBF",
INIT_31 => X"AB8E38087FC2092087FFDFC7E3F1FAF55A2DF6DB7D1C002AB7D002A82028147F",
INIT_32 => X"DF6DB7DE3F5FAFC708003DE28B68E38E280871F8FC7E3D56AB6DBEDB7FFEF552",
INIT_33 => X"ADF4516DBED16AA381C0A07082497FEFB6D1451471EF007BD0492B6F1F8F55AA",
INIT_34 => X"1C0438FD7005150438F78A2DBFFA28407038140410492550A2ABC7497BD25FFA",
INIT_35 => X"F5D0E05000492097428002E9557D1C516FA28417BD5545E38E070280024904AA",
INIT_36 => X"00000000000000000000550A00092492A850105D2A80155417BEFB6DEB8E175F",
INIT_37 => X"FFFFFFFFDFEFF7FBFFFEF552E974AA082A820AA0000000000000000000000000",
INIT_38 => X"ABEF002A800AA557FFDFEFF7FBFFF55A2D16AB550000175EFFFFBEAA00557FFF",
INIT_39 => X"6ABEFFFFBFDFFF552AAAAAA007BC0000087BFDF45AAD568B55AAFBFDFEF55042",
INIT_3A => X"FC2000FFD56AB45A2FFFDFFFAAD16AB4500043DEAAFFAEAAAAA08516AB55A2D1",
INIT_3B => X"2AA8B45087FC01EFA2FFD55EFF7D568AAA5D2A97410007BFFFFF5551555EF087",
INIT_3C => X"AAA974AA0800020BA550028B550855400AAF7AEBDFEFA280154BA55040000055",
INIT_3D => X"087FFFFEFAAAA975EF5D2E974000804154BA082A975EF5D517DEAA007BD5545A",
INIT_3E => X"00000000000000000000000000000000000005D2E80010002A954005D2A82155",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(2),               -- Port A write enable input
DIA(0)   => data_write_a(18),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(18),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(2),               -- Port B write enable input
DIB(0)   => data_write_b(18),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(18),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_19_9 : RAMB16_S1_S1
generic map (
INIT_00 => X"042200000000000041088001001AA00000000000000000000000500802000003",
INIT_01 => X"040048000024000000000404000000000A22000800000800004A200000000001",
INIT_02 => X"200C8840085EB00480060000001C008002489E0F000405EA0004040404000000",
INIT_03 => X"24004000000000000000000900002C4050000000000069500208400002E14100",
INIT_04 => X"4800200C0000000044002000C80020E40000E200000130200188000000800100",
INIT_05 => X"000000000080181000000000701000004C8000000058800000B1000009880480",
INIT_06 => X"80500081081040000000002C100040400000004641C080380400070100000000",
INIT_07 => X"4020109801A4CE005C00048380142810010564C4100114012002402028044808",
INIT_08 => X"0070700000000000000083004C3902420062000020E0000100004082A140102B",
INIT_09 => X"001150200000000000000026400000016186100000000010C04002C000000000",
INIT_0A => X"007C00008082C0002000000000002C3000000004050001030102040000000000",
INIT_0B => X"0000000000000000000000000000010000800011000000000000000000000BC0",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"000000000000000000000000000000042000760000000000000000010004B200",
INIT_0E => X"0D74002280300F0002FB069040000060000C5003000800000000000000000000",
INIT_0F => X"C01AE8004500744C780687DBA828008080A5FC0D385598035D0008A00C015660",
INIT_10 => X"39D8140040201BF861F0E7D693E6170022408116DFE0AB3006BA0011401D02AC",
INIT_11 => X"5412E4997F5249FD005043B8680CC98F00D0F2DD0140100406FE053A98F6ECC7",
INIT_12 => X"7418663001858040E153888000010840E165D0000000285C246A181C03FE4662",
INIT_13 => X"8199830066F0020858385974000001260208583854E2200000660208D6B1423F",
INIT_14 => X"8235AC508FCE8811042040F008235AE04420C040CF00C031C80009B8F224978B",
INIT_15 => X"030004E00000C220010808C10D9A92A74CD7CF4A09051110AD5A3C9200B7F280",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000118",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"07208BBA3F0C7010C660C7441920000000000000000000000000000000000000",
INIT_1A => X"861869A61861861861869A61861861861861861861861861A8208C4C1534D34C",
INIT_1B => X"984C26130984C26130984C26130984C26130984D26930984C26130984C261861",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000984C26130984C26130",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"174BA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFDFEF5D2A974BA082E95400F7FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0004",
INIT_29 => X"FFFFFFFFFFFFFFFFF7FBFDFFF552E974BAA2FFFFE10087FFFFFFFFFFFFFFFFFF",
INIT_2A => X"004001EFAAAEA8ABA087FFFFFFFFFFFFFEFF7FBEAB450804001EFAAD57FEAAF7",
INIT_2B => X"FFFBFDF45AAD568B55080028B55002E82000F7FFFFFFFFFFFFDFEFA2D568B550",
INIT_2C => X"0007FC00AAF7FFFFFFFF7FBE8B55AAD16ABEF5D2ABFF55080402010087FFFFFF",
INIT_2D => X"55A2FFFDFEF5D2EBFE00AAFFFFEBA087FFFFEFF7D168B55AAD17FFFF552EBFE0",
INIT_2E => X"000AAFFFDF45A2D16AB55F7FFFFFFF00043DE10AA843DE00557FFDFEFA2D16AB",
INIT_2F => X"FFEF552A974AA0000104AA000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFF7FBFDFFF5D2A954AA082A92428E3FFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"0071EFB6DF7AE92EBFFFFFFFFFFFFDFEFF7F5FAFC7492A974AAB6F5F8E101C7F",
INIT_32 => X"F1F8FD7AAD16AB450000001FFBEA4A8AAA147FFFFFFFFFBFDFC7EBF5E8B55000",
INIT_33 => X"00000010087FFDFC7E3F1FAF55A2DF6DB7D1C002AB7D002A82028FFFFFFFEFF7",
INIT_34 => X"BEDB7FFEF552AB8E38087FC2092F7FBF8FC7E3F5EAB45B6DF6FBEF5D2AB8F7D0",
INIT_35 => X"84971F8FC7AAD56DB6DBEF5F8FD7412ABFE28B6F5F8E820871F8FC7E3D56AB6D",
INIT_36 => X"00000000000000000000B6F1F8F55AADF6DB7DE3F5FAFC708003DE28B68E38E2",
INIT_37 => X"FFFFFFFFFFFFFFFFFDFEF552E954AA0004000AA0000000000000000000000000",
INIT_38 => X"54AAF7D568A00557FFFFFFFFFFFDFEFF7FBFFFEF552E974AA082A820AAA2FFFF",
INIT_39 => X"FFF55A2D16AB550000175EFFFFBEAA00A2FFFFFFFF7FBFDFFFFFD568B55002A9",
INIT_3A => X"A800AAF7FBFDFEFF7D56AB45AAD56AB450004001EFFF842AAAA557FFDFEFF7FB",
INIT_3B => X"FFFFFFF552AA8BEF080402000087BFDF45AAD568B55AAFBFDFEF55042ABEF002",
INIT_3C => X"8516AB55A2D16ABEFFFFBFDFFF552AAAAAA007BC0000FFFBE8B55AAD168B55F7",
INIT_3D => X"00043DEAAFFAEAAAAA08556AB55A2D57FFFFF7D568B45002ABDEAAFFD16AA000",
INIT_3E => X"0000000000000000000000000000000000000FFD56AB45A2FFFDFFFAAD16AB45",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(2),               -- Port A write enable input
DIA(0)   => data_write_a(19),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(19),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(2),               -- Port B write enable input
DIB(0)   => data_write_b(19),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(19),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_20_9 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000003",
INIT_01 => X"F55FF80000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"E05022020800008400F655001FFCFF80018FA804400000000000004400000001",
INIT_03 => X"00000000000000000000000900002CC07000000000000000000000000000013F",
INIT_04 => X"68002FFE40900010000180000001FFEC0012EE0C001370F40780000000000000",
INIT_05 => X"0840000880FCBBF0100E204DF0F88311DD8005080679800000F3000029980580",
INIT_06 => X"001000030817C8E8840155FDF9001001050023F6C3C3D0F87FA19F7F011000E4",
INIT_07 => X"000000090492260800008000EE00000000000000002101FF2002C00000004018",
INIT_08 => X"2A040001071004000013FF7FCA302C0C0008214800002101554031F800000000",
INIT_09 => X"801F57F200000090000489FEC0000001EFBEF0040008023FDFC0000000004006",
INIT_0A => X"0000000008000000000000000000ADF000000200000008000008028300110230",
INIT_0B => X"0000000000000800080000000000000000000000000000000800800A40000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"000000040900005C848538000020000000800000080000020000800101FFB600",
INIT_0E => X"00800000003A010003000000000000600FFC53FF001800000002004080000000",
INIT_0F => X"0001000000007408040000004000000004E9000008020000200000000E800800",
INIT_10 => X"00200000000313100010002000008000000000129600040000400000001D0010",
INIT_11 => X"81C012060000000000218F7840000100800004000000000066C0000080080000",
INIT_12 => X"800000000017C000100000000001A800080000000001A8040000002840008185",
INIT_13 => X"0000000006F00000100200000000012600001004000000000066000000801040",
INIT_14 => X"0000200410100000000005F00000020080090A0000000085C800002000586000",
INIT_15 => X"FF00400000000000020020020001000040283024E4F2860400008000030ED080",
INIT_16 => X"00000000000000000000000000000004010201001003020200000000000127DB",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"A0700030038200010089120104D2040020000000000000000000000000000000",
INIT_1A => X"2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2C30C30C30C30C306982121A1E79E79",
INIT_1B => X"32190C86432190C86432190C86432190C86432190C86432190C86432190CB2CB",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000432190C86432190C864",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0201000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF552A974AA0004174BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA0804",
INIT_29 => X"7FFFFFFFFFFFFFFFFFFFFFFEF552E954AA000400000F7FFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E954BA007FC00BA087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974BA082E9540000",
INIT_2B => X"FFFFFFFFFF7FBFDFFF552E974BAA2FFFFE10FFFFFFFFFFFFFFFFFFFFFBFDFFF5",
INIT_2C => X"FAAD57FEAA007FFFFFFFFFFFFFEFF7FBFFF550800020BAAAD56AAAAF7FFFFFFF",
INIT_2D => X"EFF7D56AB450000021EFA2D57DE10087FFFFFFFFFFFFFEFF7FBEAB450804001E",
INIT_2E => X"000F7FFFFFFFFFFFFDFEFA2D568B550004001EFAAAEA8ABA5D7FFFFFFFFFFFDF",
INIT_2F => X"FFFF5D2E954AA080005000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFEF552A974AA0000104AAFFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"A954AA082A92428087FFFFFFFFFFFFFFFFFFBFDFEF5D2E974AA000A07000E3FF",
INIT_32 => X"FFFFFEFF7FBFFFFF552E974AA0071C50BA1C7FFFFFFFFFFFFFFFF7FBFDFFF5D2",
INIT_33 => X"EDF6FABAEBFFFFFFFFFFFFDFEFF7F5FAFC7492A974AAB6F5F8E10E3FFFFFFFFF",
INIT_34 => X"EBF5E8B550000071EFB6DF7AE921C7FFFFFFFFFBFDFEFE3F5F8F450004050AAB",
INIT_35 => X"A497FFFFFFF7FBF8FC7EBD168B450804021FFB6D57DE28147FFFFFFFFFBFDFC7",
INIT_36 => X"00000000000000000000FFFFFFFEFF7F1F8FD7AAD16AB450000001FFBEA4A8AA",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2A954AA0800174100000000000000000000000000",
INIT_38 => X"74AA002E95410A2FFFFFFFFFFFFFFFFFFFFFDFEF552E954AA0004000AAFFFFFF",
INIT_39 => X"FDFEFF7FBFFFEF552E974AA082A820AA087FFFFFFFFFFFFFEFF7FBFDFFF5D2A9",
INIT_3A => X"568A00AAFFFFFFFFFFBFDFEFFFFFFDFEF5D2E954AA0051554BA557FFFFFFFFFF",
INIT_3B => X"D16AB450804174AAFFFFFFEBAA2FFFFFFFF7FBFDFFFFFD568B55002A954AAF7D",
INIT_3C => X"57FFDFEFF7FBFFF55A2D16AB550000175EFFFFBEAA005D7FFFFEFF7FBFDFFFAA",
INIT_3D => X"0004001EFFF842AAAA087BFDFEFF7FFEAB45A2D568B550804001EFF7D57DEBA5",
INIT_3E => X"0000000000000000000000000000000000000F7FBFDFEFF7D56AB45AAD56AB45",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(2),               -- Port A write enable input
DIA(0)   => data_write_a(20),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(20),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(2),               -- Port B write enable input
DIB(0)   => data_write_b(20),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(20),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_21_9 : RAMB16_S1_S1
generic map (
INIT_00 => X"4A302428B824900A128C090A5C1800261500213C005FE812D10420054085A202",
INIT_01 => X"001FFE3440B609703B0427F801A40B8115BC4F655300340288A40D30040E4DD8",
INIT_02 => X"E00424256888D8819801000F9FFFFFFFF149FF1FCA448046C60A0D2437C517F9",
INIT_03 => X"20030640003250640003250F06002CC1740002019824E001CD357832440001FF",
INIT_04 => X"EA2C3FFD400006E04401A8837001FFFC004AEF00080B70E08FB5789421007C5C",
INIT_05 => X"00011A0C40F9FFF80920954FF0F00809DF84A0202879800000F3000029980780",
INIT_06 => X"0805984B7A1FC0A0000101FFF0480080002281F7C3C381F87C03DFFF00009004",
INIT_07 => X"B424068086A205481A60A19000908204A855B000A08A61FF20C3D004D331D340",
INIT_08 => X"1BFA0001600802000023F7FFC08D234B40C2028253000040114200000D0226C0",
INIT_09 => X"EF1F5FF054096C6ADBA169FFC202B1C1FFBEF0440021083DFFCE22DC2880E24D",
INIT_0A => X"45FF0C004041D84862A28C54518DBFF00020004C0A6044901112A0908AA0A300",
INIT_0B => X"018C241102068006C620C03882019480E63180855A492712CC01C49C20201BFE",
INIT_0C => X"08A9464116544302C02D92236488D92236488D92236488D922366446C911B210",
INIT_0D => X"08800444021048034004001890000806002804A0822189000900D80621FFBE00",
INIT_0E => X"060580261013813A2CC396506102C4053FFD5BFF00A04A00200602CA52001100",
INIT_0F => X"080C0B004C202621A85C09411500135844C196D3606941018150098404C1A304",
INIT_10 => X"B02901013416181C96C2C9C600890A2028172192C460D1820302A0130809834A",
INIT_11 => X"9C5E803408250180AC268D185DB3F4350B811068C00049A0A4AA68F05C96A001",
INIT_12 => X"002C006560138F032B1804101244C883052208209040CC849063A747512B7678",
INIT_13 => X"41401E240665750440C9488280254530314080C2C601040420352148A00501B1",
INIT_14 => X"500811204D000700114204A70422016149916011008CAA8858850B00C32591C0",
INIT_15 => X"FFC06E60AC0496022300233104663040808E991765205000070121D41D18D098",
INIT_16 => X"40100401004010040100401004010040102090010008000001C0E010020007DF",
INIT_17 => X"0100401004010040100401004010040100401004010040100401004010040100",
INIT_18 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_19 => X"FFEF9FEEFF7FFDF7FF3E3DFDF7E0000000000000000000000000401004010040",
INIT_1A => X"BEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBFFDFDFFFCF3CF3F",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFEFF7FBFDFEFF7FBFDFEFBEF",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000FFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0001000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E954AA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0004",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA0004154BAFFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"52E974BA0804000AAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0004174BAFF",
INIT_2B => X"FFFFFFFFFFFFFFFFEF552E954AA000400000007FFFFFFFFFFFFFFFFFFFFFFEF5",
INIT_2C => X"A082E95400007FFFFFFFFFFFFFFFFFFFFDFEF5D2E974BA002E97400007FFFFFF",
INIT_2D => X"FFFFFBFDFEF5D2A954AA002E974BA087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFBFDFFF5D2E954BA007FC00BA5D7FFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA000002000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080005000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"A974AA0000104AAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974BA0000174AAFFFF",
INIT_32 => X"FFFFFFFFFFFFDFEF552E954BA080A000AAE3FFFFFFFFFFFFFFFFFFFFFFFEF552",
INIT_33 => X"02A95400087FFFFFFFFFFFFFFFFFFBFDFEF5D2E974AA000A07000007FFFFFFFF",
INIT_34 => X"F7FBFDFFF5D2A954AA082A924281C7FFFFFFFFFFFFFFFFFFBFDFEF5D2A974BA0",
INIT_35 => X"A557FFFFFFFFFFFFFFFF7FBFDFFF552E974BA0020924BA1C7FFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000E3FFFFFFFFFFFFFFEFF7FBFFFFF552E974AA0071C50B",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0000020000000000000000000000000000",
INIT_38 => X"74BA0000174BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954AA080017410FFFFFF",
INIT_39 => X"FFFFFFFFFFDFEF552E954AA0004000AAF7FFFFFFFFFFFFFFFFFFFFFFFEF552A9",
INIT_3A => X"E95410087FFFFFFFFFFFFFFFF7FBFDFEF5D2A954BA082E800AAA2FFFFFFFFFFF",
INIT_3B => X"FBFFFFF552E954BA002E97410087FFFFFFFFFFFFFEFF7FBFDFFF5D2A974AA002",
INIT_3C => X"57FFFFFFFFFFFDFEFF7FBFFFEF552E974AA082A820AA557FFFFFFFFFFFFFEFF7",
INIT_3D => X"5D2E954AA0051554BA5D7FFFFFFFFFBFDFEFF7FFFFFEF5D2A974BA0000020AA5",
INIT_3E => X"0000000000000000000000000000000000000AAFFFFFFFFFFBFDFEFFFFFFDFEF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(2),               -- Port A write enable input
DIA(0)   => data_write_a(21),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(21),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(2),               -- Port B write enable input
DIB(0)   => data_write_b(21),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(21),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_22_9 : RAMB16_S1_S1
generic map (
INIT_00 => X"5290F4CDE914905A14A43D33F488243E17122300F55FEB189B343A1140548380",
INIT_01 => X"A54007B259F6A975386262000C344BA9573C6FF57B18A5FB0ABFCD3C2C5F4F0C",
INIT_02 => X"021DFF8C38B3C009D203551040030071869D0040180AA2DC53DB89BEA8204001",
INIT_03 => X"2603475A969D0475A969D0460EAA401005111011BD506954EDB40F5EF41434C0",
INIT_04 => X"922D9002100ED69E443D988B0D5400103E48003D0800011E803B06B5B9125A15",
INIT_05 => X"281B5A0C06000408F4DF9422010D8802022F2124A8022492580040440002021C",
INIT_06 => X"F780C4C052881ADA0E05440205DA50930FA182010004700083E220800440B588",
INIT_07 => X"049D028B93FB561833D8094A02F5EA92FD7247E10305C40040D136E6A023F7FC",
INIT_08 => X"00028241680A0E002A9400803A884B5B5206B7C2E53CA25144009007A64EBD64",
INIT_09 => X"41008810240240C6694008010392354010000560141801002028A83D2A08E06D",
INIT_0A => X"34000000848BCA6902A29C54539C020E11810098D4067EFF9FF284D483E2AB41",
INIT_0B => X"500001840000C80B410014088040F4A944B1AA313C0022AA0011C0DC00028001",
INIT_0C => X"80B14004D158C8CA24A1C2A870AA1C2A870AA1C2A870AA1C2A872550E1543800",
INIT_0D => X"80A14050A01509E050854498B5281A1C34E506A2C6898B52A154DAC6B6000850",
INIT_0E => X"0B03001A483A4146603050080410089180008800143D83888281A2034A850142",
INIT_0F => X"A4160600349075238473F1210006133835E92273612B3482C090068A0E84AC56",
INIT_10 => X"30060181BA1B13959DC08DA902458870201970B29602562B0581200D141D0959",
INIT_11 => X"E042021C040D0152C8058B3840F044708E7E1C20A0106EA166C13AFC14AA3804",
INIT_12 => X"080E004B0C17C1439A9838301DC1A8438EA32C009DC1A8255300650458A1D588",
INIT_13 => X"018010E186F110A908E3A8CB0026C9A610A908E6A60F0807626610E160589C4C",
INIT_14 => X"2A701667334005800B1605F043858125E0D04110408D2485CA034681E43A1E40",
INIT_15 => X"00646002304244A91102C93A2D608D2A258DF8034188200C050171A41108F084",
INIT_16 => X"110441104411044110441104411044110466C440446CA06951D4EA8010009804",
INIT_17 => X"0040100401004411044110441104411044110441104411044110441104411044",
INIT_18 => X"0401004010040100401004010040100401004010040100401004010040100401",
INIT_19 => X"F7DFBFDEFE8FF1F7DEBDDF7DF7D05122890000000003FFFFFFFF900401004010",
INIT_1A => X"9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7BFFDFD7DDDF7DF7D",
INIT_1B => X"F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE79E7",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000003F9FCFE7F3F9FCFE7F3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA000400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0800",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000002000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2A954BA000015400FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080402010FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2A954BA0004154BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A0004174BAFFFFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0800154AAFFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF552A974AA0000174BAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974A",
INIT_2E => X"000007FFFFFFFFFFFFFFFFFFFFFFEF552E974BA0804000AAA2FFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080400010000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E954AA080005000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000402010FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2A954BA000417410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"804154BAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974BA0000174AAFFFFFFFFFFF",
INIT_34 => X"FFFFFFFEF552A974AA0000104AAE3FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0",
INIT_35 => X"AA2FFFFFFFFFFFFFFFFFFFFFFFEF552E954BA000E124BAE3FFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000007FFFFFFFFFFFFFFFFFFFFDFEF552E954BA080A000A",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804000100000000000000000000000000",
INIT_38 => X"54AA000400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2A954AA080017410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"0174BAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A954BA000415400FFFFFFFFFFFFF",
INIT_3B => X"FFFDFEF552E974AA0804174AAF7FFFFFFFFFFFFFFFFFFFFFFFEF552A974BA000",
INIT_3C => X"2FFFFFFFFFFFFFFFFFFFFFDFEF552E954AA0004000AAA2FFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2A954BA082E800AAAAFFFFFFFFFFFFFFFFFFFBFDFEF5D2E954BA002A820BAA",
INIT_3E => X"0000000000000000000000000000000000000087FFFFFFFFFFFFFFFF7FBFDFEF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(2),               -- Port A write enable input
DIA(0)   => data_write_a(22),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(22),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(2),               -- Port B write enable input
DIB(0)   => data_write_b(22),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(22),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_23_9 : RAMB16_S1_S1
generic map (
INIT_00 => X"EF20906D902424807BC8241BC81801B97D38AD3C0800103362A6741C80A12A02",
INIT_01 => X"001FFF8409F089003B4422000D80C80106804A7951C5B9D1C828043EA28838F9",
INIT_02 => X"E01CEE21649C82C40800000F9FFEFF8E72CA7F5FC2E22809925A0D3611C877F8",
INIT_03 => X"24000400402670400402670D48222DC1764446838624000080007460C40001BF",
INIT_04 => X"68403FFC020560E0443E21037C01FFFC0002EE00628BF0E02FAD781014085014",
INIT_05 => X"0112000202FBFFF00920017FF0F0628BFF8488890979800002F702002BB807A0",
INIT_06 => X"EF85788B681FC000000001FFF0010000000001F7CBC385F87C0BFFFF20040001",
INIT_07 => X"F6E200000000C1440E3AE408009120071070FA07A1CB23FFA403F0C4D23BF7C0",
INIT_08 => X"0BF87CA400804000003FF7FFD8880A034AC09662305AB10555421006891A1089",
INIT_09 => X"BE1F5FEA10092C0896A243FFC0008087FFBEF2000000001DFFC612C0C0400100",
INIT_0A => X"41FF0C2060501000600000000001BFFA800808189A657EF81DD0C00079CC8001",
INIT_0B => X"018C24110A860006C620C0312241C482B20400CC52492710CC80060020A81BFE",
INIT_0C => X"0C08866907048320C20C10030400C10030400C10030400C10030400608018210",
INIT_0D => X"040002000041500300100040000500C000801000C02400000952800001FFBF04",
INIT_0E => X"FC850015385380380CDB86106502C5043FFD5FFF00A04BC010A7724B10000800",
INIT_0F => X"89F90A002A70A710A51C01C05904014861433602A1CAF13F2110055614C72FC0",
INIT_10 => X"E02D02001C1E14981B43253EE50C8220180F1082E06397E07E42200AAC298E57",
INIT_11 => X"8421802400A90022B0070FAE18019214A380344920080B21A58B02AC60BACDF0",
INIT_12 => X"0A2A000C480B0704B54028101AC49C84BB4100009AC49C80857A82D20CE8CB22",
INIT_13 => X"01E00C8103416445C12ED0400027C5292445C12D500B0005A62D344CB241D095",
INIT_14 => X"132C907425604680038706A35132C94BDD011010404428886AC91B11311C8280",
INIT_15 => X"FF000470BE0692020328CA0028042054A92771C50FC070110001C1680809591D",
INIT_16 => X"00802008020080200802008020080200800800200200000000000008004807DF",
INIT_17 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_18 => X"8020080200802008020080200802008020080200802008020080200802008020",
INIT_19 => X"0000000000000000000000000000000000000000000000000000008020080200",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080002010FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974AA000400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000400010FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974AA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080000010FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E954AA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954A",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA000015400FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080002010FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974AA000400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000402010FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E954AA080005000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA080407000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA00041741",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080000010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000402010FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2A954AA080002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954AA080017410FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"552A954BA000415400F7FFFFFFFFFFFFFFFFFFFFFFFFF552A954BA080015410F",
INIT_3E => X"0000000000000000000000000000000000000F7FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(2),               -- Port A write enable input
DIA(0)   => data_write_a(23),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(23),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(2),               -- Port B write enable input
DIB(0)   => data_write_b(23),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(23),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_24_9 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100600007FFF000080108004000800020000840041000080808",
INIT_02 => X"FC5CA803400EB8209000000F9FFEFF8E7240FF1FC22409EA04018E50074017F0",
INIT_03 => X"11100400000000400000000D00002CC07400000090C080019001010A000001BF",
INIT_04 => X"68003FFC00040000000000008001FFFC0002EE00000370E007A100000000E468",
INIT_05 => X"0000000000F8BFF00920004DF0F00001DF8000000079800000F3000029980780",
INIT_06 => X"6E461803081FC000000001FFF0000000000001F7C3C380F87C019FFF00000000",
INIT_07 => X"600C2400013649609C8000980040814210254000A00B21FF2003F2A80D500000",
INIT_08 => X"0BF80000000000000003F7FFD88D2B4A02C0940062EC2804001610020408178B",
INIT_09 => X"8E1F5FE010092C0892A041FFC0000001FFBEF0000000001DFFC002C000000000",
INIT_0A => X"41FF0C0000000000600000000001BFFA0000005501AA00000CE2000009400000",
INIT_0B => X"018C0411020600048620C030020502000200000400490510CC00040020201BF4",
INIT_0C => X"0808064106040300C00C10030400C10030400C10030400C10030400608018210",
INIT_0D => X"0000000000004003000000000000001200580000000000000000000001FFBE00",
INIT_0E => X"0086C022005381380FDB96516140C6043FFD5BFF000041000000004110000000",
INIT_0F => X"80010D804400A7240C840C201D0210840043B4804012500021E0088014C04940",
INIT_10 => X"4109038041021C980200D06410C1924030008142E06024A00043C01100298092",
INIT_11 => X"587CC200002100C14428090A1D02348190814C09C010104025AA40041A0D8005",
INIT_12 => X"022E0030300B0E46177004208000D8C61D7004300000D884817B00011306B2D9",
INIT_13 => X"01E003060344710009875C018100013831000985DC000C20003C310006143B70",
INIT_14 => X"4001850EDC004780144806A64400186CBF8961104000C3807884000846EB9500",
INIT_15 => X"FF0006E08C063C0220002201490418082010A57263E0100008000290161E711C",
INIT_16 => X"00000000000000000000000000000000000000000000000000000000000007DF",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"F2D0AEEAF6E7CC1132CDB4441990000000000000000000000000000000000000",
INIT_1A => X"BEFBE79E79E79E79E79EFBEFBEFBEFBEFBEF9EF9EF9EF9EFA69861219575D75F",
INIT_1B => X"783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1EFBEF",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000783C1E0F0783C1E0F0",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0201000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A000400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA000400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000400000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402010000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"00002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080002010FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000400010FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA00040000",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020100000000000000000000000000",
INIT_38 => X"74BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"000010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA000002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974AA000402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000002010F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(3),               -- Port A write enable input
DIA(0)   => data_write_a(24),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(24),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(3),               -- Port B write enable input
DIB(0)   => data_write_b(24),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(24),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_25_9 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100200002000000080100004000000020000800041000080808",
INIT_02 => X"FC400086000000800000000F9FFEFF8E738FFF1FC204010000000111568DD7F8",
INIT_03 => X"00000400000000400000000D00002CC4740000008000000080000000000001BF",
INIT_04 => X"68003FFF64A564AC000000000001FFFE0082EF00010370E007A1000000004000",
INIT_05 => X"0A00040148F8BFF80920804DF0F00101DFC040000079C92484F30499299837C1",
INIT_06 => X"66041803081FC0E0801101FFFD000E41002299F7E3C380F87C019FFF81200096",
INIT_07 => X"000000080480AE00000080000000000000000000A00B21FF2003E00000000000",
INIT_08 => X"1BF80000400A02000003F7FFFA0008000200A0400008A0000014100200081000",
INIT_09 => X"8E1F5FFA53EFBCACB2E369FFE0010001FFBEF80C40630C7DFFEEBAF000800202",
INIT_0A => X"41FF0C0600000000600000000001BFFE00301000000000000CC020000140000C",
INIT_0B => X"01DCCC31222730A49620C030020100000200000400490D10EC00040220201BF4",
INIT_0C => X"0808064106240300C00C10030400C10030400C10030400C10030400608018210",
INIT_0D => X"0883044582114013412080000000000000000000000000000012800001FFBE00",
INIT_0E => X"00040020000180380FC386106140C6043FFD5BFF00A04B80608003CB120C1106",
INIT_0F => X"0000080040000200040400000100000000009480000240000100080000400900",
INIT_10 => X"0001000000000808000000240000020000000100006004800002001000008012",
INIT_11 => X"0001001808220000002004001900000080800008000000000022400000088000",
INIT_12 => X"0010000000000E00110000000000408009000000000040808063004000008200",
INIT_13 => X"6000000000046100000240000000001021000004400000000010210000001010",
INIT_14 => X"4000000404000800000000060400000088000001800000001084000000088000",
INIT_15 => X"FF800C608C041002000002000006100000002100000000180600000000100018",
INIT_16 => X"4110441104411044110441104411044510629041040D180400000010028047DF",
INIT_17 => X"1104411044110441104411044110441104411044110441104411044110441104",
INIT_18 => X"1044110441104411044110441104411044110441104411044110441104411044",
INIT_19 => X"FBA2894A196A8C5A2932EC15DA080800002FFFFFFFFFFFFFFFFFC11044110441",
INIT_1A => X"2492492492492492492410410410410410410492410492412000531215A69A6B",
INIT_1B => X"158AC562B158AC562B158AC562B158AC562B1588C46231188C46231188C49249",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000B158AC562B158AC562B",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080000010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000010FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08000000",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(3),               -- Port A write enable input
DIA(0)   => data_write_a(25),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(25),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(3),               -- Port B write enable input
DIB(0)   => data_write_b(25),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(25),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_26_9 : RAMB16_S1_S1
generic map (
INIT_00 => X"E9264EAB20190CA3BA4997AA9002AE9C001006B0778015CFA17E0811039879C7",
INIT_01 => X"2FFFF9BB1F773C7F9BB07DFFFDD863FC5FFF3FEFFBBF9FFB22FFFBC7B9F30686",
INIT_02 => X"E06CCC62052E708180F6FFBFFFFCFFFFF9C7FF7FC24332E642090000074037F6",
INIT_03 => X"428003739CD9863739CD9869FE2B7DEAF300029E4E300DFE69A6E644E6FF473F",
INIT_04 => X"7C2FEFFFF5BA124F003DD31EAFFFFFEE9FF7EE6F4C0770FFD7DC7CA53997B2B1",
INIT_05 => X"DFFB5421C1F8BBFAFDBFFACDF0FFCC05DDDBFF3690F9EDB7F5F7AFF639BD7DE3",
INIT_06 => X"EFD044ABC817C3E3A74667FDFFB6FF5727CC3BFEF7C3FAF87FF59F7FFBFEF69F",
INIT_07 => X"00003002132462052E708180EF060C18E5BEFB051225CDFF7002C4EEDE77F6E0",
INIT_08 => X"3FFF7D5000EC75088ED3FF7FC8790E46426CE06CB1F8E041051831FA3068D77E",
INIT_09 => X"C05FD7FF9BEFBDCEFBEE59FEF44F6603EFBEFAFCC2E35E7FDFD147CCF3F583FA",
INIT_0A => X"67FF1C7FBFADEB31E35768E8ED6BFDF3EB3EBF9DDBCE7FDC1DF8A760F3EACC02",
INIT_0B => X"5BDDCC3B336F7C548667D47B7737AF3FD62601EDC25B3533DCEB07F262213FFC",
INIT_0C => X"5F9A06E19F4D93A0EA0F78C35E30D78C35E30D78C35E30D78C35E986BC61AE31",
INIT_0D => X"5FD7AFEFDFFAF59B6FF28FE1D80D73D840607307DCFE1D80EF69A004DFFFF7FF",
INIT_0E => X"0004001F8041897B2FFFC6D86D70CE04FFFFF3FF1F5F5475BD7F72E4D75EBFAF",
INIT_0F => X"F60008003F008237B0040A00010003E020023E0201F45EC0010007E01047D17B",
INIT_10 => X"00010001DC0004C81003DE050A700200001DC0006863E8BD8002000FC0208FA2",
INIT_11 => X"2200E400002801E1A00004C21C0206F60081800800007B00010F02007EC09A0E",
INIT_12 => X"0880007E000807C7C1A612001E0015C7C19C22001E0015C59DFE82011A311AA0",
INIT_13 => X"00001BC00101F60409F0670840070809760409F06984800780097604067D0010",
INIT_14 => X"81019F40042100001F800203D81019EC085614000085C80023D81009CF008A74",
INIT_15 => X"FF802FFDFFAFD082003B032FB987E04021D481D4000819060801E0D00001231D",
INIT_16 => X"EBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEFFBFBFBFBBFCFBB0FFDFEFFEF2DFFFFFB",
INIT_17 => X"BFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAF",
INIT_18 => X"FAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFE",
INIT_19 => X"475B15BCF491E166CC8553F86EDB5C88646FFFFFFFFFFFFFFFFFEBFAFEBFAFEB",
INIT_1A => X"861861861861861861861861861861861861869A69A61861AFBD54D5F871C71D",
INIT_1B => X"984C26130984C26130984C26130984C26130984C26130984C26130984C261861",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000984C26130984C26130",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040201",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(3),               -- Port A write enable input
DIA(0)   => data_write_a(26),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(26),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(3),               -- Port B write enable input
DIB(0)   => data_write_b(26),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(26),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_27_9 : RAMB16_S1_S1
generic map (
INIT_00 => X"00080A40000A41248002029000050A088000008242A0004404480002000A1155",
INIT_01 => X"2FFFF1C11F781C129C107DFFFE0860941E81258CA2B71C2220EC1B86E1A00002",
INIT_02 => X"E1000000810000014400FF6FFFF0FFFFF8007F1FC21110005080200000221FF0",
INIT_03 => X"4080026318C18226318C1821302232EAE00002BE001115FE48620040840A863F",
INIT_04 => X"643D4FFC2530000F003D821C0BFFFF8E9EF79E6D440748FED70060842105B0B0",
INIT_05 => X"D6F39020D1F8A3FAFDBFBACDC8FDC405D1DB7F1490E5EDB7D5CBADB2385D79C3",
INIT_06 => X"6FE000A38007C3032646EFF1F0B6FF46A78C39F8E723F2E47FE59C7F9ADA2612",
INIT_07 => X"00002820000000810000014401060C180190310540118DFF1000C0849673F6C0",
INIT_08 => X"3FF779100062B12A8EC3F47FC80208808210880C00082050000110023068D030",
INIT_09 => X"005F07E09BFFBD07FBAC09F8E42922038F7DF8BEC2E39C5F1FD047CEF1B582D8",
INIT_0A => X"63FF5D5F9FADE911E81C09818109E1F16B16B71092CE7ED81CF403601228C402",
INIT_0B => X"1BFDCC39732F3554866AD57C37BEAF1C152201A4C05B7531D56B05B06A213FF8",
INIT_0C => X"5BCA06F18FC59380F00E34430D10C34430D10C34430D10C34430F0861A2186B5",
INIT_0D => X"5B56ADAB5FAAE58B2F628EA0C80FA3F04040510768EA0C80CC61A0044DFFC6EB",
INIT_0E => X"0004001D800188792CE79715710AE4047FFD23FF315D54358D593474955AB6AD",
INIT_0F => X"520008003B000297B0040200010003E020001F0201E44A400100076000579129",
INIT_10 => X"00010001DC00004A10035E0408300200001DC000086BC8948002000EC000AF22",
INIT_11 => X"02002400002801E1A00000C01E0202F60080800800007B00000782006EC0820A",
INIT_12 => X"0080007E000006A7C10602001E0001A7C10C02001E0001C18DE282010A311AA0",
INIT_13 => X"00001BC00000FE0401F04300400708007E0401F04180800780007E04047D0010",
INIT_14 => X"81011F40040100001F800002F81011EC080604000085C80001F810094F008034",
INIT_15 => X"FF800C6DDDAFD082001B03249887E04001D481D4000009020801E0D00001021F",
INIT_16 => X"AB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6BF1EBDABD8E270BF84A25C6ACB777E3",
INIT_17 => X"B6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6AD",
INIT_18 => X"6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADA",
INIT_19 => X"490E2168100481CA860402104A471688747FFFFFFFFFFFFFFFFFAB6ADAB6ADAB",
INIT_1A => X"000000000000000000000000000000000008200000000000200072F210000001",
INIT_1B => X"05028140A05028140A05028140A05028140A0500804020100804020100800000",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000A05028140A05028140A",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040201",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(3),               -- Port A write enable input
DIA(0)   => data_write_a(27),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(27),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(3),               -- Port B write enable input
DIB(0)   => data_write_b(27),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(27),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_28_9 : RAMB16_S1_S1
generic map (
INIT_00 => X"02200AA400180030808802A900002A08001280A08A801044104A1000001818C3",
INIT_01 => X"0AA00011460214428114180000882214413D0A71592A01D92213D28005210202",
INIT_02 => X"0451110A012100884000AA30200000000C100040104112101100008888200000",
INIT_03 => X"448000318C52A20318C52A20148810200111100C211004AA00034204200A2200",
INIT_04 => X"04004001001A90110000121402AA0000003C00000500000040080421080D0080",
INIT_05 => X"4060000C8001000000002E000000050000001610300000010000802202040012",
INIT_06 => X"1000002080001111001222000425A1040026A008000000000000000009328280",
INIT_07 => X"2491008A00491201210088400122448908A20402000408001000040820000000",
INIT_08 => X"20058310402A160026500000028040101004200C840082115554000112244814",
INIT_09 => X"4140000800000060000720000102028000000490160801020002200011100010",
INIT_0A => X"020000081B34211082B694D4D294000020020381040000000200032040004400",
INIT_0B => X"4800210C19808400500010009110091500020B408810000100200020408B0000",
INIT_0C => X"01028000080118020023604858121604858121604858121604858090B0242C00",
INIT_0D => X"010000800920040804020A6058003108402043058C460580653020005A004039",
INIT_0E => X"00000002800008014004104104420A00C000200005000010040A0020CC000200",
INIT_0F => X"520000000500000010000200000000000000280000040A40000000A000001029",
INIT_10 => X"00000000000000C0000002000830000000000000480008148000000140000020",
INIT_11 => X"020024000000000000000440000000020000800000000000000C00000040020A",
INIT_12 => X"00800000000001804006020000000500400C0200000005400A90000000100000",
INIT_13 => X"0000000000018200001003004000000142000010018080000001420000200000",
INIT_14 => X"8000080000010000000000018800008000060400000000000310000008000034",
INIT_15 => X"000002040080000000110006B081400000400000000009020000000000002200",
INIT_16 => X"802008020080200802008020080200802101210810C39A66A90A85420413A820",
INIT_17 => X"0200802008020080200802008020080200802008020080200802008020080200",
INIT_18 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_19 => X"DE21102C110A00246972BD89A40A0C22E1000000000000000000002008020080",
INIT_1A => X"2082082082082082082082082082082082082082082082080D35050758C30C31",
INIT_1B => X"0582C160B0582C160B0582C160B0582C160B0580C06030180C06030180C08208",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000B0582C160B0582C160B",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(3),               -- Port A write enable input
DIA(0)   => data_write_a(28),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(28),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(3),               -- Port B write enable input
DIB(0)   => data_write_b(28),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(28),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_29_9 : RAMB16_S1_S1
generic map (
INIT_00 => X"79964E4BA01DACAB9E659792D00AAE160002829C7FDFEFCEE97C2815039D70C3",
INIT_01 => X"0ABFF9AB0775343F9AB01DF80D5821FC0FFF3FEFD1AF9FF1207FFBC7B9720586",
INIT_02 => X"002CCC60050E700080F6AAA7BFFC007189C7FF2FC00330E602800000074037F6",
INIT_03 => X"468003210868A63210868A68DA017D207200021C4E200CAA6186A40042FF4300",
INIT_04 => X"7C2FE002F0900001003C5316A6ABFFE21F36E02F0D03701F47D41800109FB281",
INIT_05 => X"4979440580F9B808F49F6A4DF00F8D01DC4B97369078249370F482E62BA41462",
INIT_06 => X"B250442BC81001E1870223FC0BF7F11507C423FE33C078F803F19F00E936721D",
INIT_07 => X"00011080012460050E700080EF020408EC8CFA01122149FF700200665A35D260",
INIT_08 => X"2BFD055040A452000443FF00007906464068406C31F84000000831FA1028575A",
INIT_09 => X"805FD017102690AA694551FE30444681E0820AD40201423FC00122C493500172",
INIT_0A => X"0600002AFFBE2330815568A8AD6ABC02A02A0B0CCB463B4C0748A720B1EA4C00",
INIT_0B => X"0850400A11414C005005000B51158936D20601A98A10200308A002E240010BFC",
INIT_0C => X"05928020194918A22A2268C81A32068C81A32068C81A32068C81A99034640C00",
INIT_0D => X"058102C48970541944B20FA1580561D040406305587A158046282000DBFFF13D",
INIT_0E => X"000000028040890327DCD28928324400DFFFF0001F1F0050342D42A086040B02",
INIT_0F => X"F60000000500802010000A000000000000022A0000141EC0000000A01000507B",
INIT_10 => X"00000000000004C0000082010A700000000000006800283D80000001402000A0",
INIT_11 => X"2200E4000000000000000442040004020001800000000000010D000010401A0E",
INIT_12 => X"08800000000801C040A6120000001540409C2200000015441DAC800010100000",
INIT_13 => X"0000000001019600081027084000000956000810298480000009560002200000",
INIT_14 => X"800088000021000000000201D800088000561400000000002358000088000A74",
INIT_15 => X"00802594A282C0000033010FB181E00020400000000819060000000000002305",
INIT_16 => X"C0B02C0B02C0B02C0B02C0B02C0B02C4B12B312912831A27FCFE7FFB175B6FF8",
INIT_17 => X"0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02",
INIT_18 => X"B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C",
INIT_19 => X"BBCF9F96EE7FFDF7FE783FFDFFEA0C00602FFFFFFFFFFFFFFFFFC0B02C0B02C0",
INIT_1A => X"EFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEEBAEBAEBAEBAEBBFFDF9FBEFFFFFFE",
INIT_1B => X"BFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFBEFB",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000FBFDFEFF7FBFDFEFF7F",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(3),               -- Port A write enable input
DIA(0)   => data_write_a(29),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(29),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(3),               -- Port B write enable input
DIB(0)   => data_write_b(29),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(29),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_30_9 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"F7FFBFFEFF9FE1F7FFBFFFFDFFD0000000000000000000000000000000000000",
INIT_1A => X"9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7AFBD75F5FDF7DF7F",
INIT_1B => X"F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE79E7",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000003F9FCFE7F3F9FCFE7F3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(3),               -- Port A write enable input
DIA(0)   => data_write_a(30),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(30),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(3),               -- Port B write enable input
DIB(0)   => data_write_b(30),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(30),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_31_9 : RAMB16_S1_S1
generic map (
INIT_00 => X"129000008004A00804A40000400800020000000C005FEA005800200400050100",
INIT_01 => X"255FF18019700810180065FFFC0040801E80258CA2951C2200EC0906A0804140",
INIT_02 => X"E0000000000000011000550FDFF0FFFFF0007F1FC200000044000000000817F0",
INIT_03 => X"0000024210A30024210A3001002220C06044469200040154482000408400043F",
INIT_04 => X"602D0FFC2420000E003D80080955FF8E1ECA8E2D400340FE870060842100B030",
INIT_05 => X"0213100040F8A3F8FDBF944DC0FDC001D1CB6904A061EDB6D4C30490281831C1",
INIT_06 => X"6FC000830007C202060445F1F0D25E4207A099F0E303F0E07FE19C7F80402412",
INIT_07 => X"0000200000000000000001100004081001103107000185FF0000C0849673F6C0",
INIT_08 => X"1BF27A00000000000883F47FC800080002008000000820440000100220489020",
INIT_09 => X"011F07E013EFBC06FBA009F8E00120038F3CF82C44630C5D1FC002CCE0808248",
INIT_0A => X"61FF0C06C48BC801600000000001A1F00110101092CE7ED81CF0004012288000",
INIT_0B => X"11DCCC31222730048620C4382204A608142002A440492530C401049020221BF8",
INIT_0C => X"0888066187448380E00C10030400C10030400C10030400C10030600608018210",
INIT_0D => X"080204010200418301208480800D02D00040100240A808008840800405FF8640",
INIT_0E => X"0004001D000180780CE386106100C4043FFD03FF101D40008001304018081004",
INIT_0F => X"000008003A000217A0040000010003E02000160201E040000100074000478100",
INIT_10 => X"00010001DC00000810035C0400000200001DC0000063C0800002000E80008F02",
INIT_11 => X"00000000002801E1A00000801C0202F40080000800007B00000302006E808000",
INIT_12 => X"0000007E00000607810000001E000087810000001E000081846282010A211AA0",
INIT_13 => X"00001BC00000740401E0400000070800340401E04000000780003404045D0010",
INIT_14 => X"01011740040000001F8000025010116C080000000085C80000C8100947008000",
INIT_15 => X"FF800C609C06D082000A03200806A040019481D4000000000801E0D00001001D",
INIT_16 => X"010040100401004010040100401004010060C040040C200950402090128057C3",
INIT_17 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_18 => X"0040100401004010040100401004010040100401004010040100401004010040",
INIT_19 => X"00000000000000000000000000001000802FFFFFFFFFFFFFFFFF810040100401",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(3),               -- Port A write enable input
DIA(0)   => data_write_a(31),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(31),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(3),               -- Port B write enable input
DIB(0)   => data_write_b(31),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(31),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_0_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"ED39BA795990D275FB4A6E96ACC4731DEA4598B0AFB54867F6EE4618C3749803",
INIT_01 => X"8AA0047D8607944AC7DA180001ECA2444042106208408208C20022E9173734B3",
INIT_02 => X"1A7DDD79F9A73E6CCA7DAAF00001000008478020113D98E382FEDF333027C80F",
INIT_03 => X"75D341110C58F31110C58F32A208921F8051500147A0E4AB3493FB3A01EBE240",
INIT_04 => X"86424001531009B100425A97B2AA0001E03501D0A39C8F0078420001106D0C4C",
INIT_05 => X"BCC8CA2EBF03400700402BB20F00239E20341699198600000B08694B16434804",
INIT_06 => X"103FB860B2800161F8432200012DA185F80F24081C3C0707800E600056881308",
INIT_07 => X"B24197ABCDA467F9A73E6CCAFDC3870EEEEC44E2BDFE220094D03022210C011C",
INIT_08 => X"240581B5695EAA80262C080032BF07C7C1FC3F8E94F65B11555EAFFC1C306758",
INIT_09 => X"7E40000BEC004170040DB60017FED1CC0001045002984202003DB931192D60A5",
INIT_0A => X"120071411A74315881A28C141118000C5A85A60444210123820B43B40804674D",
INIT_0B => X"0820008E514045BB514F0106D1D8599581D3A958BC104A89215AC14C48898403",
INIT_0C => X"C261C01C48B1584A0CA3E2687A9A1E2687A9A1E2687A9A1E26870CD061343885",
INIT_0D => X"D274E93A758FA8683AC54B287522E10A74AF4AA59C568752662F5AC218000002",
INIT_0E => X"FF83C002783A0904231C70470C7E0B92800224008AE09FAD4BD48D1FC5D3A4E9",
INIT_0F => X"5BFF078004F075885DFBF7E15C06101C55E921F1F80FAB7FE0F0009E0E903EAD",
INIT_10 => X"F12E0380231F13978FF023FAFDBD9870380230F2D6081F56FFC1E0013C1D207D",
INIT_11 => X"DE7F263C0C8700125C0F8F3C43F1F10BBF7EFC61E01804E1E6C8F8FE807F67FB",
INIT_12 => X"02BE00017C17C1007E5E2E3081C5AC007E6F0E3081C5AC44418D65FE45DEE55B",
INIT_13 => X"61E0042786F103E9F01F9BC3C120C5A703E9F01F978B8C20666703E9F8A0FFED",
INIT_14 => X"FA7E283FFB414F80005F05F10FA7E283F78F6511C048278DCA174FF038FF15B4",
INIT_15 => X"0066A20B61692F293185D8D724E15D3FCC6B7C236FE0691B0700132C1F0EF880",
INIT_16 => X"3A4E93A4E93A4E93A4E93A4E93A4E93A4F942F92E9628540AD2A91442525A000",
INIT_17 => X"A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E9",
INIT_18 => X"4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93",
INIT_19 => X"55F3898E09B56C74DAB15D1CF13501AA495000000000000000003A4E93A4E93A",
INIT_1A => X"082082082082082082082082082082082082082082082082082084E41DC71C71",
INIT_1B => X"E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F82082",
INIT_1C => X"FFFFFFFFFFFFFFF94A5294A5294A5294A5294A52800003E1F0F87C3E1F0F87C3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"3060C183060C187FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"BDEBA0000000000000000000000000000000000000000000003060C183060C18",
INIT_28 => X"168ABA002E82145085155545F7AA975EFFFAABDE00FFAEBDFFF5D2EAAAAAF7AE",
INIT_29 => X"7FFFE10005542145557FD5545FF8000155087FC0155F7D168B55007BFDF45085",
INIT_2A => X"7FFC0010080017555555568AAAFFFFD7545AA8028A00A2802AABAFF8028BEF5D",
INIT_2B => X"FF842AABAA2AE95545FFD168ABAF7AEAAAAAA2FFFDF4500043FE105D2E954BAF",
INIT_2C => X"5007FD7400550415410002E974BA5D5168A00A2D142155005142010FFAE820AA",
INIT_2D => X"FFF780000BA007FE8AAAFF803FFFF5D2A821550000000BA007FD55FF5D7FC014",
INIT_2E => X"000AAFBEAA00007BFDFFF082EBDF455D5142000082E82145FFD17DFEFFFD168B",
INIT_2F => X"DFD75D2AA8A80EA8E2FE3F000000000000000000000000000000000000000000",
INIT_30 => X"68B551475FAF6D1C556F0AA1C24AABEA495FC716F002A975FFE3AA95E00EBAEB",
INIT_31 => X"42A0070071C50BAFEF1FAE0016D56A16D557BC257D415E0216FA3F1E8FC0145B",
INIT_32 => X"8010E004924874825D7FEAA85487FD24AFE3D02DAAAE12BD5545A2803AA00005",
INIT_33 => X"120155EA568E870BAEB8A05A2AEA8B50F55A2F150005A3A438BD04AFAB8F550A",
INIT_34 => X"545E055FFBE81D0BE8EA8A3AA05A2A5504001C74BA42A1571E8028E3DB7816D0",
INIT_35 => X"A5C7E3DFFFE90B45B47ABA497A82FFAFD2A82485FD2415A105C21451ED42A002",
INIT_36 => X"00000000000000000000B55EAAA100AA1D0F6F480B6A555A2A57A002A3D5FDB6",
INIT_37 => X"5EFAAAAB5E1AF3AABFF45592E88A0AFE80A8B0A0000000000000000000000000",
INIT_38 => X"65F520EBE9EF67D7BEA1FD5D556ABEF5D557FEBA55022A3F70C6B405F4D2AE97",
INIT_39 => X"C114728007521170821CE0FDE69411A8DED57CE1055555E5F58EFFC01FE2CACB",
INIT_3A => X"42341D5DEEBEF55080034E0A592A4AD0079C75D6070CC5CBB0280C029ABAA3EB",
INIT_3B => X"7F353AAF6C77F7F20D968BF57812A95E02A2AAB5EB0F280800EFAEE9F5D18F31",
INIT_3C => X"C91565455C141E41887D58AC448B69C30E02116220415A9540AA854140A0A204",
INIT_3D => X"DE6BE93172D7D625B556EEAB157ABEBE1B4D792A4AD1183454180DD3FDCAAAB7",
INIT_3E => X"F0000001FF0000001FF0000001FF0000001FF01EABC4B8014174FF7DA80F52FE",
INIT_3F => X"FF0000001FF0000001FF0000001FF0000001FF0000001FF0000001FF0000001F")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024,               -- Port A enable input
WEA      => wbe_a_lo_1024(0),               -- Port A write enable input
DIA(0)   => data_write_a(0),        -- Port A data input
DOA(0)   => data_read_a_lo_1024(0),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024,               -- Port B enable input
WEB      => wbe_b_lo_1024(0),               -- Port B write enable input
DIB(0)   => data_write_b(0),        -- Port B data input
DOB(0)   => data_read_b_lo_1024(0),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_1_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"212C001411984004084D000508C53810A03D1450E839B003342114428A000803",
INIT_01 => X"00000019400B100A8196000000CC004400400002000000000000028001340000",
INIT_02 => X"052137AE8031800C0044009000000000061800001CD4019802AD04CCCFC20004",
INIT_03 => X"04514108C60C21008C6042108400000201440020505100000043C30E10E9F000",
INIT_04 => X"02104001011DEFE088805681920000008000004001900800004002108C280008",
INIT_05 => X"040002340105000200000000080001900010000108040000000008411600401C",
INIT_06 => X"1034001042800808201000000001000820020000102000040000000000800180",
INIT_07 => X"64BF81A15EDFDE8031800C00843060C19E030022103600000450020800040004",
INIT_08 => X"00008004691687AA840008000090248CC84E000046000311555521F183060AC5",
INIT_09 => X"0820800D08100171000DB000154440C800400500000852020011200201012021",
INIT_0A => X"02000040001000880A2A04445004000102002041000001008208001440004140",
INIT_0B => X"4820018A1140440078050040511000102000A008183000010002404400000000",
INIT_0C => X"1000C80008000C030030880C2A030A00C28030A80C2A030A00C28018D4061401",
INIT_0D => X"10040802050080200284401C0022880F009E08008205C0020118088018000000",
INIT_0E => X"0F03C00280000000420860C60C0C0B92C0000000004000010042000040102008",
INIT_0F => X"001E078005000108400005E11C0610000000288058000003C0F000A000100000",
INIT_10 => X"F10E0380000000C202300000008D187038000000480800000781E00140002000",
INIT_11 => X"806302380C870010000004400100110800007861E0180000000C400680000001",
INIT_12 => X"023E00000000018000580C308000050000610C30800005000215006800000101",
INIT_13 => X"61E0000000018100B0001843812000014100B00016030C20000141002880026D",
INIT_14 => X"400A20009B404F80000000018400A20044096111C04000000304026000501580",
INIT_15 => X"0046820040082300218450C2800010094000482141E060190700100000002200",
INIT_16 => X"020080200802008020080200802008020080008008600500A82A1100A8000000",
INIT_17 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_18 => X"0080200802008020080200802008020080200802008020080200802008020080",
INIT_19 => X"81328A46BABEFC54A0810C7452B4428A14000000000000000000020080200802",
INIT_1A => X"AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA28A28A28A28A2A8218D2C0C924925",
INIT_1B => X"E974BA5D2E974BA5D2E974BA5D2E974BA5D2E975BADD6EB75BADD6EB75BAAAAA",
INIT_1C => X"FFFFFFFFFFFFFFFD8C6318C6318C6318C6318C63000002E974BA5D2E974BA5D2",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"70E1C3870E1C387FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"5555500000000000000000000000000000000000000000000070E1C3870E1C38",
INIT_28 => X"EBDF455D2EAABEFF7FFE8BFF5D0002155557FFFFFF007FC21EFA2FFD74AAAAD5",
INIT_29 => X"AA95400552AAAABAFFD1574105D7FD75FFAAAA800AAF7AA974BAFFFBE8B45F7A",
INIT_2A => X"0517DF555D2EAAA1055000015500557DF45AAD1400BAA2AE801550051555EFF7",
INIT_2B => X"FFD540155557FD5400F78028BFFFFFBEAB55F780020AAAA80020AA082EAAB550",
INIT_2C => X"AFF842ABEF5D517DF55552A974AAF7AE820AA0851574BAA2D1574AA5D7BFDEBA",
INIT_2D => X"EFAAD1575EF557FFFE10557FFFFFFFFD56AAAAFFFFD7555AAD168B45AAAEAAAB",
INIT_2E => X"0005D7FFDF4500043FE105D2E954BAF7AE80010082A97410557FEABFFAAFBE8B",
INIT_2F => X"51C7A2FBD5490BFD1C056A000000000000000000000000000000000000000000",
INIT_30 => X"974BAF7FFEFB45FFAABDF55492AA8BC2EBDFEAF7F1F840017D4975D2FEF147FC",
INIT_31 => X"080BEF495FC71D54124924385FAAA8AAAE3D145410F7F1D55D71C002DABAEBAA",
INIT_32 => X"002D082082AB8B6DBEDB7DF7F540E2AE85028B40155145F7AF6DBED5450AA1C2",
INIT_33 => X"78E021FF1471FDEAAFFD56F16D5571D2E28E38E0216FA2D1E8E80140F45082B4",
INIT_34 => X"A2DA3FB7DAAD4AAAAF487BC70BFA97F7AF6D417E92482BF84020BA495557E3FF",
INIT_35 => X"55554ADBD7A2FFC7BEFF6FFD7FC7002FD74951D71EDFFABFD16FAAAE92BD5545",
INIT_36 => X"00000000000000000000547AB8F550A8010E00492487482FFFE82A85EBAE2FFC",
INIT_37 => X"1EF005162BEF047FD5545AAFBF7400FBF9424F70000000000000000000000000",
INIT_38 => X"714F8338AAAA1D0AE974AAF7FFFDF55F7AABFF55082CA8B4DF6C1E8F5E540002",
INIT_39 => X"EABEF75550ACBB7582225FF5843404547184164AA5D2EBEEB0A2D555410D3555",
INIT_3A => X"FEAAEB083BC1000FF8409000512AEABFFDF79DCBF755962010BDCBBC21455D7F",
INIT_3B => X"801F8BA0C57740BDAA0688E5405D57D412F7D55F5E50C7F401BAAE8403CF5A3F",
INIT_3C => X"5D16BABAA3EBC3157ABD5FFE55F2AA9FEAFDF7F431A9F7FFE81FF013A8001AFF",
INIT_3D => X"FB863550229BCABEB7DA403FFFDA2FBF7FED2C7F955445079E280A00C56145EF",
INIT_3E => X"0000000000000000000000000000000000000596EBEF55080034E0A592A4AD00",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024,               -- Port A enable input
WEA      => wbe_a_lo_1024(0),               -- Port A write enable input
DIA(0)   => data_write_a(1),        -- Port A data input
DOA(0)   => data_read_a_lo_1024(1),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024,               -- Port B enable input
WEB      => wbe_b_lo_1024(0),               -- Port B write enable input
DIB(0)   => data_write_b(1),        -- Port B data input
DOB(0)   => data_read_b_lo_1024(1),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_2_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10E006600180111284380310006289800480032283E000A34301002001A0817",
INIT_01 => X"0005A00810790848048044A54E404350404000720885800802000906E4910200",
INIT_02 => X"407004208400408044C600C50AA055254010541A110222841200000002402544",
INIT_03 => X"0600011004182401004102408C28414043101000408118000145840440F5C415",
INIT_04 => X"5035855703A2900A000CD3088400F40688C9844409060850925E58A4081A0221",
INIT_05 => X"0200840D1021A15AC50494894850890540D1E12020C6E510818500440A280090",
INIT_06 => X"113044094002801020440090A8011A1224AB9380552102442884882A20004097",
INIT_07 => X"000100880004428400408044860000008C022402102100AA40004404B5075460",
INIT_08 => X"15C23440408C862A2A12382A8A5244145048C06085008010141521F000001240",
INIT_09 => X"400582B9033AA0E7AA4110B0506744810554542450694E710A836188C2C00222",
INIT_0A => X"443518360012C2210B020414109130A28038188096A06B8C120CA440A9C00802",
INIT_0B => X"1345E53300EC68005605002964AF222A5704004D080211121C80024200821780",
INIT_0C => X"181080C1110C882202211488452213C88472213C88472213488441109A442231",
INIT_0D => X"008204440210091341208041000810C00000300220201800A908000038AD0284",
INIT_0E => X"00040002804180300E88D28D206A40000554815500481440300000C44A081100",
INIT_0F => X"000008000500828700000000010000000002380000A00000010000A010050000",
INIT_10 => X"00010000000004CA000214000000020000000000684280000002000140200500",
INIT_11 => X"000000000020000000000442100002840000000800000000010C000026000000",
INIT_12 => X"00000000000805A4800000000000152300000000000015801272000100210020",
INIT_13 => X"000000000101C00000C000000000000940000120000000000009600004050000",
INIT_14 => X"0000130000000000000002018000106000000000000000002380000141000000",
INIT_15 => X"55000190000000000002000280000000011080C0000000000000000000002310",
INIT_16 => X"40902409064190641906419024090244902A9003004800415120D4A190804241",
INIT_17 => X"0900409004090641906419064190240902409024090641906419064190240902",
INIT_18 => X"9044090040900409004190441904419044090040900409004190441904419044",
INIT_19 => X"75960040138D70C030B51C50C7D100A2052F81F81F83F03F03F0419044190441",
INIT_1A => X"0410410410410410410410410410410410410410410410410248602081659659",
INIT_1B => X"5128944A25128944A25128944A25128944A25128944A25128944A25128941041",
INIT_1C => X"FFFFFFFFFFFFFFFE1084210842108421084210843FFF825128944A25128944A2",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"7FD5FF555815607FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"2AA000000000000000000000000000000000000000000000007FD5FF55581560",
INIT_28 => X"FC21EFA2FFD75EFAA8415410AA8415555087BFFF55A2AA800BAFFAE954000800",
INIT_29 => X"84155EFA2AEBDEAAA2FBEAABA5D7FE8B555551421455D0002145552EBFEBA007",
INIT_2A => X"2AEBDF555D2E954BAA2AA974BAFFFFE8B45552EBDF45FFAEAABFFF7FFE8B55F7",
INIT_2B => X"AAAAAAAAAFFD1574105D7FFFF555D2AAAAAA5D2E820BAA2FBEAB5555557DF55A",
INIT_2C => X"50055575EFFF84021555D043DEAA5D04021EF557FC21FFAA8428BFFAAAA954AA",
INIT_2D => X"10085568A00FF80175FFA2D17DFEFF7800215500557DF55AA80001FFAA800015",
INIT_2E => X"0005D00020AAAA80020AA082EAAB5500517DF555D042AA10A284154005D00154",
INIT_2F => X"00AAFFAA9543A080038A2A000000000000000000000000000000000000000000",
INIT_30 => X"0017D5D20B8EAA007FC51C7A2FBD55D2BE800042AFE8E1557D0075D2F45BEAA8",
INIT_31 => X"AA8BC7EBDFEAFEFFD00105FFBC20BDEAAA2FBF8AAA557BE8B6D5D5FFABEF4904",
INIT_32 => X"FFEFB6D555578F7DB6A0BDF7D480E174BFA02A974BAF7F5EFB455D2ABDF55492",
INIT_33 => X"ED1FDE90E3A497492B6AAADAAAE3D155E105571D55D71C002DABA5524820BAB6",
INIT_34 => X"BE8F401D7B6A0001470155C51D0092A071555D5E3AE821D00001FF0871C016DB",
INIT_35 => X"5BE8555400550A38428007FED000E3DA3DFD5E3DFFFBD5A38A021551C5F7AF6D",
INIT_36 => X"00000000000000000000410F45082B4002D082082AB8B6D1C5B7DF7FF78E075C",
INIT_37 => X"5EF005560B55F7AA800AAF7AA954AA00042AAA20000000000000000000000000",
INIT_38 => X"ABEF057D68F5F5A00021EF55042AAAA007FD5555AAFBD7545FBB8020A3F7AE97",
INIT_39 => X"7DF55D7AABFF5428ACA8F45A6C1E8F5EFF84165EFF7802BAB0A2FFEAABA557BE",
INIT_3A => X"CA8AA80800020AAF7FBFFFEF04552ABFFFF841FFE75CA882108202E974AAF7D5",
INIT_3B => X"00151FF0C57401E5F3D1E00A1A884174A8FFAEBFEB0A2D55541051555694F002",
INIT_3C => X"2AA801455D7FE8BFFF680800FFF7AAA155F595542455512A975455D3AA8A0055",
INIT_3D => X"5D79FCAF774AE005BE7895554005D2A8A0B882FFFFE10AAAAAB755A66B6AF56A",
INIT_3E => X"00000000000000000000000000000000000000C3BC1000FF8409000512AEABFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024,               -- Port A enable input
WEA      => wbe_a_lo_1024(0),               -- Port A write enable input
DIA(0)   => data_write_a(2),        -- Port A data input
DOA(0)   => data_read_a_lo_1024(2),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024,               -- Port B enable input
WEB      => wbe_b_lo_1024(0),               -- Port B write enable input
DIB(0)   => data_write_b(2),        -- Port B data input
DOB(0)   => data_read_b_lo_1024(2),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_3_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"210C00A20020000108430020001600B8156021104940741B3530400E02B92203",
INIT_01 => X"014C9BCA58B1296D24A402C992500B69404040028804A0080A000416A8D90A08",
INIT_02 => X"C12026A484318004404405C9C66E331352180D468B8203980300204442E02B34",
INIT_03 => X"04000748D60D24648D60524C88804D0215011020D15018148040C10A70E1D58C",
INIT_04 => X"18283333240FE41244187308C9104D70944852640901083801750EB0A418C220",
INIT_05 => X"0613142D01912CC2A1B4140528348900C612A104201C689044340ED413A07649",
INIT_06 => X"119000034019881822104C5E68035250A222829710A0A02C18C01A9920842413",
INIT_07 => X"402F00AB0016CA0431800444841020509D038B021230C1990001C644C8273200",
INIT_08 => X"16905000408482088290E8E64010248C4A5AA840C2000110001521F0810A92E7",
INIT_09 => X"0003CE6581BD016342A951AB146C4480530C3B2A8088D3542651670200C1826A",
INIT_0A => X"00735D36209A8A20020894004284B660821030C8990467401218004041020002",
INIT_0B => X"512445B740457154562F957CC08B00093700080D0A4851001D8302D20A0A1530",
INIT_0C => X"00508650008008021021A40861021840869021A408610218C0869810D6043095",
INIT_0D => X"1C8508438450801043A08090380A8834207007022209038080190000999C8F84",
INIT_0E => X"000400200000C0002A48A206204C4205F3304B33004C0041006240140A1C310A",
INIT_0F => X"0000080040000083800400000100000000008400018040000100080000510100",
INIT_10 => X"0001000000000800000244040000020000000100002A0080000200100000A702",
INIT_11 => X"000000000020000000200000080002C000800008000000000022000006808000",
INIT_12 => X"0000000000000A2281000000000040A3810000000000402001400000022002A0",
INIT_13 => X"000000000004200001C0400000000010200001C0400000000010000004490010",
INIT_14 => X"0001070004000000000000060000104C08000000000000001000000903008000",
INIT_15 => X"CC004050CA0C00020220200070040000010401C4000000000000000000100008",
INIT_16 => X"4310E4310A4210A4210A4210A4210A4210A8D0830A68010001B4DA881048061C",
INIT_17 => X"21084290A4210A4210A4210A4210A4210A4210A4210E4310E4310E4310E4310E",
INIT_18 => X"90A421084290A421084390E4310C4390E4310C4390E4310C4290A421084290A4",
INIT_19 => X"015303C0C78C706428A14C586291000A044001FFE000003FFC004290A4210842",
INIT_1A => X"2492492492492492492492492492492492410410410410412821600001249249",
INIT_1B => X"51A8D46A351A8D46A351A8D46A351A8D46A351A9D4EA753A9D4EA753A9D49249",
INIT_1C => X"FFFFFFFFFFFFFFFC00000000000000000000000038F56351A8D46A351A8D46A3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"55AB02055AB0207FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"420000000000000000000000000000000000000000000000007FFFAB57FFFAB5",
INIT_28 => X"A800BAFFAE9554508002AA00AA843DF55FFAA955EFA2D168B55557BEAA000055",
INIT_29 => X"002AB55AAAA955EF005568A00087BE8BFFA2D155410AA8415555087BFFF55A2A",
INIT_2A => X"AAABFF5508003FF555D0002145552ABFEBA007FC21EF007FD75FFAA841541008",
INIT_2B => X"082EBDEAAA2FBEAABA5D7FC0155005168B455D042AB45F7FFD741000042AA10A",
INIT_2C => X"FF7FBEAB55F7AABDEBA5D7FC2010A2D1575FFF7AA975555D2E80145F78415545",
INIT_2D => X"EF5555554AA087BC01FFFFAAAAB55552A954BAFFFFE8B55552EBDE00F7AEAABF",
INIT_2E => X"000082E820BAA2FBEAB5555557DF55A2AEBDF555D2E954BA002EAAABA002A821",
INIT_2F => X"FB7D5D7FEAA3808554203A000000000000000000000000000000000000000000",
INIT_30 => X"1557D1475FAF45BEAA800AAFFAA95578080038A2AA28E3AF55E3A0BA5D7AADB6",
INIT_31 => X"BD55D7BE80004AA1E8E2AB55B6A0925D7085F6AA10087FEABD7AAD57AEBAB68E",
INIT_32 => X"F5D0438140E2FA38B6AEBFF6D1D04AAFFA41040017D5D20B8EAA007FC51C7A2F",
INIT_33 => X"D0A901FFFF801557D1C20B8EAAA2FBE80AA557BE8B6D5D5FFABEF49002FB55FF",
INIT_34 => X"5D20BDE00EBAAA8BC7EBDFEAFEFAB8ABAE925D21C7010EADB525D7FFAE975C75",
INIT_35 => X"F002EADA921420871D74971D24820875C21D5EB8AA8FFF012A954BAFFF5EFB45",
INIT_36 => X"000000000000000000001C24820BAB6FFEFB6D555578F7DB6A0BDF7DEB8E125F",
INIT_37 => X"B55A28408145AAFFFFFFF5D7FEAABA0051400A20000000000000000000000000",
INIT_38 => X"AB55FAD568AA2AFAE975EF555168B55F7AA800BAF7AA955EF00042AAA2A2AEAA",
INIT_39 => X"2AAAA007FD55558A7BD7145FBB8020A35D2ABEF55F7800015F087FEAA00007FE",
INIT_3A => X"968F575D003FF55F7D5420BA5D2ABFEAAF7AE9DFF759A82AEF70800021EF5504",
INIT_3B => X"FFD5145FBAC9755F05040255FFD84175EF55002AAB0A2FFEAABA557BEA3EF057",
INIT_3C => X"82E974AAF7D57DF45552A3FF10AA8429F45A7D5EAF5FFBAEAAA10554155400AA",
INIT_3D => X"FF843FFE77C80825BC052ABFE10550415557085540000005156155FE90A8F5C0",
INIT_3E => X"00000000000000000000000000000000000005500020AAF7FBFFFEF04552ABFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024,               -- Port A enable input
WEA      => wbe_a_lo_1024(0),               -- Port A write enable input
DIA(0)   => data_write_a(3),        -- Port A data input
DOA(0)   => data_read_a_lo_1024(3),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024,               -- Port B enable input
WEB      => wbe_b_lo_1024(0),               -- Port B write enable input
DIB(0)   => data_write_b(3),        -- Port B data input
DOB(0)   => data_read_b_lo_1024(3),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_4_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"A108400020612C80284210081034849800A00030300004833522C82D04A16002",
INIT_01 => X"2043998A1839284D1CA0650E1E504368403008418984014902030806A0D10200",
INIT_02 => X"C120042200000000044441CE01E80F00A49043118680008002000000026208E4",
INIT_03 => X"040001020019200020011209CC0164C060000000690111040144800042F5C403",
INIT_04 => X"7029AF0F81A00010CCA47700CC513CAC0D0B8E02010740E19754080108988021",
INIT_05 => X"02139405007133C0712244CD20F20105D583000020E9892201D304D42A9835E1",
INIT_06 => X"9190440300078002014405D9EE814C0284A883B6D7038AE079059B7800048092",
INIT_07 => X"000100AA0004408000000004840400008D200102503000782000C00C8025C000",
INIT_08 => X"00728A00408403220811991E02120C044058080004000001101121F220000260",
INIT_09 => X"811001E1185B38AD23C3707AD46440818F3CF80EC423CA7D01D123C80200816A",
INIT_0A => X"45810810A01B40216361056D6150F41200280001900439001FD8A00041400000",
INIT_0B => X"11FC88076266E800D605402962A820211500024808010512C40106D222223B14",
INIT_0C => X"0408804116040B02C02C500B0C02C100B0C02C100B0402C300B0401618058611",
INIT_0D => X"040200050200501301208482200D00D0A0408402C4282200A84800009B878680",
INIT_0E => X"00000020000100024AC88300300060090F0D830F00025400300204D018000804",
INIT_0F => X"8000000040000206A2000800000000000000950002E010000000080000588040",
INIT_10 => X"0000000000000808000554000200000000000100006D0020000000100000BB00",
INIT_11 => X"0000400000000000002000001A0002504001000000000000002280000D800800",
INIT_12 => X"0800000000000E2C802000000000408D801000000000408012440000200110A0",
INIT_13 => X"000000000004680003A0040000000010280003800800000000102800000B0000",
INIT_14 => X"000005C0002000000000000620000158000010000000000010A0000B00000200",
INIT_15 => X"C30146200400104002602600400000000294004000000004000000000010001A",
INIT_16 => X"0080200000008020000000802000000080080000004090014134DA101288C6DB",
INIT_17 => X"0802000000000401806010040180601004018060100000802000000080200000",
INIT_18 => X"8060180601004010040080200802000000000000802008020000000000008020",
INIT_19 => X"C0A28A063807E0500014063450404882846FFE000003FFC00000010040100401",
INIT_1A => X"AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA28A28A28A28A2934C8D0CCD145144",
INIT_1B => X"68341A0D068341A0D068341A0D068341A0D068351A8D46A351A8D46A351AAAAA",
INIT_1C => X"FFFFFFFFFFFFFFFC0000000000000000000000001FE32068341A0D068341A0D0",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"408102040810207FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"800AA00000000000000000000000000000000000000000000040810204081020",
INIT_28 => X"168B55557BEAB4500554200000557FE10FFFBEAA10007FD7410FFAA97555082A",
INIT_29 => X"55574105D2A800AA00043FEBA5D7FEAA00007BE8AAAAA843DF55FFAA955EFA2D",
INIT_2A => X"57BC00AAA2FFEAAAAAA8415555087BFFF55A2AA800BAFFAE9555508002AA0000",
INIT_2B => X"A2AA955EF005568A00087BE8BFFA2D17DE1000517FE10AAAAA8AAA002E975455",
INIT_2C => X"FAA8417410A2D140000F7FBC2010A2D157400AAAE974AAAAAA974BA08002AB55",
INIT_2D => X"EFA2AABDEAA087BEAAAAA2FBD54BA080002145552ABFEAA007FC21EF007FD75F",
INIT_2E => X"00055042AB45F7FFD741000042AA10AAAABFF5508003FF55F7D568A00552EA8B",
INIT_2F => X"5400F7A49057D0824850B8000000000000000000000000000000000000000000",
INIT_30 => X"3AF55F7A0925D7AADB6FB7D5D7FEAB7808554203A145178E00FFFBE8A101475D",
INIT_31 => X"A9557D080038AAA145157428492E8008200043FE925571EFA380871C7028A28E",
INIT_32 => X"AEA8A9200249056D4175C5092AAF5FDA38BE8E1557D1475FAF45BEAA800AAFFA",
INIT_33 => X"AA4954281C0E2FB55B6A0925D7085F6AA10087FEABD7AAD57AEBA08517DE00AA",
INIT_34 => X"007FC51C7007BD55D7BE80004AAFEDB42028EBFBC2028BED152438AAA092492A",
INIT_35 => X"AF7DF6AA00412EAABFFAA803DEBA0875EDA80BEF1C743840040017D5520B8EAA",
INIT_36 => X"0000000000000000000041002FB55FFF5D0438140E2FA38B6AEBFF6DBE84AAEB",
INIT_37 => X"A00FFFFEAA105D5155410FF84021EF0800154B20000000000000000000000000",
INIT_38 => X"DEBA0851574B2AAAEAAB55F78400145AAFFFFFEF5D7FEABFF0051400A25D5568",
INIT_39 => X"68B55F7AA800BAF7AA955EF00042AAA25555410BA082E8201000043FE005D517",
INIT_3A => X"568AA200557DE00AAAAAAA000804001FF005575408AA557FEB2FFAE975EF5551",
INIT_3B => X"D1550AAAA8002010F2AC154B25F2ABFF55F7800015F087FEAA00007FEAB55FAD",
INIT_3C => X"800021EF55042AAAA007FD5555087BD6145FAAC000A2A6FBC00BAAAFBC00BAF7",
INIT_3D => X"F7AEBDFF779A82AA43F7FBE8A00082EA8BFFAA843FEBA08517DE00F3F9574B30",
INIT_3E => X"000000000000000000000000000000000000008003FF55F7D5420BA5D2ABFEAA",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024,               -- Port A enable input
WEA      => wbe_a_lo_1024(0),               -- Port A write enable input
DIA(0)   => data_write_a(4),        -- Port A data input
DOA(0)   => data_read_a_lo_1024(4),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024,               -- Port B enable input
WEB      => wbe_b_lo_1024(0),               -- Port B write enable input
DIB(0)   => data_write_b(4),        -- Port B data input
DOB(0)   => data_read_b_lo_1024(4),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_5_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50DF4A0791B3FCB694379283C81FD996A091832102004A336A20E03C040C002",
INIT_01 => X"805FBDC69830A84D5C6A60000C34C26841280A00084000C8C212892EEAD53235",
INIT_02 => X"3B2026B578918E640A4F01CF8011FF0002080000082CA9998276DF7772C7C80D",
INIT_03 => X"37134108420D700084205702A4008A1D9100002171C0E0051554D93A11F5D140",
INIT_04 => X"8A41A0FC03A56DA000425A819410E3816C086198A388B702A8CA1210844A0C4C",
INIT_05 => X"B1808A062E8BC835F5E84532D708238A282F00A9291224800A2861490343082C",
INIT_06 => X"903FB8483A90581859050424100940825C6184401CDC451B860A6507160C4100",
INIT_07 => X"D26F068BCC96CDF8918E640E96D1A3469D6300E2FFEA27F8E4D23248130E259C",
INIT_08 => X"0BFA82E568442B2A082C0A7E3014250D49DA37A2420619000002AFF48D1222E5",
INIT_09 => X"3F005001E40969289429360416DCD1C46083030604B1CA20C03DF83B0A2C60A5",
INIT_0A => X"14613C71005A10492B888120288F480D58858449026145B3830F449449062B4F",
INIT_0B => X"11AC04934AC648BFD727C031E64170A137D5AA5C3E4B0F8A3C58C34C002290E3",
INIT_0C => X"CA29C6CC50384B6AC6AC86AB31AACA6AB39AAC86AB39AACA6AB3055643559C31",
INIT_0D => X"C673E33CF28F38603855401985228A0614BD30A0A2819852011E5AC2B87F9182",
INIT_0E => X"FF87C002F87A803E460B2516510CA594FF0044FFA4B08BAC4BB2CD0F09CF84E3",
INIT_0F => X"0DFF0F8005F0F5100DFFF5E15D06101C55EB29F1E00BE53FE1F000BE1E802F94",
INIT_10 => X"F12F0380231F17D78FC029FFF58D9A70380230F2FE0017C37FC3E0017C3D005F",
INIT_11 => X"FC7F023C0CA700125C0F8F7E43F1F001BFFE7C69E01804E1E7CCF8FC003FF5F1",
INIT_12 => X"023E00017C1FC1A4BFD82C3081C5BD27BFE30C3081C5BD00C02365D645CEEF5B",
INIT_13 => X"61E0042787F181E9C1EFD8CB8120C5AF41E9C18FD60F0C20666F41E9F009FFFD",
INIT_14 => X"7A7C077FFF404F80005F07F187A7D14BFFC96111C048278DEB074F9930FF9D80",
INIT_15 => X"C064014B8B652E2B3120C81284641D3E8DBF7D636FE860190700132C1F0EFB80",
INIT_16 => X"38CE1384E3384E338CE138CE1384E33C4E3ECE32E128882551349A1CBAA44103",
INIT_17 => X"84E3384E3384E3384E338CE138CE1384E3384E338CE138CE1384E3384E338CE1",
INIT_18 => X"CE138CE138CE138CE1384E3384E3384E3384E338CE138CE138CE138CE1384E33",
INIT_19 => X"F5E5BB4E7F7B9DB7FF3A1B6DB7E8410A8C000000000000000000384E3384E338",
INIT_1A => X"BEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEF9F7CFDFDDCF3CF3D",
INIT_1B => X"BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEFBEF",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000001711C7BBDDEEF77BBDDEEF77",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"FDFFF00000000000000000000000000000000000000000000080000000000000",
INIT_28 => X"FD7410FFAA97410082A800AAAAAE955450055421FFFFFBC0010AAD5574BA557F",
INIT_29 => X"7FD74000055574BA5D7FD7555A2D5575EF55517FF5500557FE10FFFBEAA10007",
INIT_2A => X"0002AABA5D2ABFFFFAA843DF55FFAA955EFA2D168B55557BEAB5500554200000",
INIT_2B => X"5D2A800AA00043FEBA5D7FEAA00007BC00AAAAAEBDF45A28428B45FFD168BFF0",
INIT_2C => X"5080028A00A2FFFDE00F7D57FEBAFF80174BAAAD1555EF555555555005557410",
INIT_2D => X"BA5D2E821FFA2D5554BA557BD75FFAA8415555087BFFF55A2AA800BAFFAE9555",
INIT_2E => X"00000517FE10AAAAA8AAA002E97545557BC00AAA2FFEAAAA082A97545F7D5420",
INIT_2F => X"7010BEDF524AA5571FDFEF000000000000000000000000000000000000000000",
INIT_30 => X"78E00EBFBE8A101475D5400F7A49043D0824850B8A2AE9756D145B401FFFFFFC",
INIT_31 => X"FEAB7D0855420BA1471D74380851524BA5571D757DB6D5525EF555178F6D1451",
INIT_32 => X"8A28B6DEBDF6DBEF1C0A28AAA5524BFFFFA28E3AF55F7A0925D7AADB6FB7D5D7",
INIT_33 => X"5555057D145152428492E8008200043FE925571EFA380871C7028B6AEBDF45B6",
INIT_34 => X"BEAA800AAFFAA9557D080038AAAA2FBF8E10EBD578EAAFF8415482BED1555EF5",
INIT_35 => X"81C209256DFFDF420BA552A821FFB6DF574A85575C55EFBE8E1557D1475FAF45",
INIT_36 => X"0000000000000000000008517DE00AAAEA8A9200249056D4175C50920875FDA3",
INIT_37 => X"5FF5D7BC21EFF7FBD7400F7FBC00BA55557DFF70000000000000000000000000",
INIT_38 => X"01FF5D5568BE7555568A00AAFFEAA105D5155410FF84020AA0800154B2AAAA97",
INIT_39 => X"00145AAFFFFFEF5D7FEABFF0051400A25551554BA0051400BA5551575EFF7D14",
INIT_3A => X"1574B2FFAABFF45FFAAAABFFAAFFFDFFF552EA8AAA55043DFF7AAAEAAB55F784",
INIT_3B => X"8002410FFD5575EF5555421E75555400BA082E8201000043FE005D517DEBA085",
INIT_3C => X"FAE975EF555168B55F7AA800BAF7AA955EF00002AAA2A2FBE8A00A2D16AAAAFF",
INIT_3D => X"0055554088A557FEB25D00021FFFFFFC00BA552A821EFFFFFD74BA5D51575F7F",
INIT_3E => X"000000000000000000000000000000000000000557DE00AAAAAAA000804001FF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024,               -- Port A enable input
WEA      => wbe_a_lo_1024(0),               -- Port A write enable input
DIA(0)   => data_write_a(5),        -- Port A data input
DOA(0)   => data_read_a_lo_1024(5),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024,               -- Port B enable input
WEB      => wbe_b_lo_1024(0),               -- Port B write enable input
DIB(0)   => data_write_b(5),        -- Port B data input
DOB(0)   => data_read_b_lo_1024(5),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_6_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10800B0061A01002840002C03002818000402322520070B313301C4389B2082",
INIT_01 => X"250041CA3839684D18A160000C52426841000000090800090210080008110200",
INIT_02 => X"0020042080010000044654C0000C008010000000001020900200200002620814",
INIT_03 => X"060881021088200021080200E4000A0891000020610111500104C00000F14400",
INIT_04 => X"0880000100000002000052288144004281C050400100280000C8100000080001",
INIT_05 => X"928080840001100A08009000280201000850E022401400002028214043410820",
INIT_06 => X"10100518090012122100C808049310002040000410A0001400000200120840D2",
INIT_07 => X"000100800004400001000000860408108C22000A502010074120044800040001",
INIT_08 => X"50000040D0C4E2088003FD01C01004044058082004000000000121F020408244",
INIT_09 => X"00BF17E9001205A5204911F814444080400100020000D200DFD16400C2A40AA0",
INIT_0A => X"04611C17849000022862A1596C8B5DF04834948900000100220C244840000880",
INIT_0B => X"03AD0413424E4044D665C070C22602291504400D084915020448114080201000",
INIT_0C => X"5E08864011088B22D22C008B0022C408B1022C208B0822C608B1111600458010",
INIT_0D => X"4251A12CD28A300429688001000800000020280204001000A00804309A002182",
INIT_0E => X"0000000280402400420800000000006200FC10002442042429324294014E8CA7",
INIT_0F => X"A40000000500800840000800000000000002280018001480000000A010100052",
INIT_10 => X"00000000000004C2003000010240000000000000680800290000000140202000",
INIT_11 => X"2000C0000000000000000442000001080001000000000000010C000280001804",
INIT_12 => X"08000000000801C300A010000000156000902000000015101200002800000000",
INIT_13 => X"000000000101800038002408000000094000386028040000000940000ED40000",
INIT_14 => X"0003B000002000000000020180002A24005010000000000023000060C7000A40",
INIT_15 => X"3F0280090321000040A410C28108000160008094000810040000000000002300",
INIT_16 => X"284A5284A728CA5284A528CA728CA52C4A5A0A32A300940101349A0408240818",
INIT_17 => X"9CA1294A329CA5284A728CA7284A5284A728CA5284A528CA728CA5284A728CA7",
INIT_18 => X"CA3294A129CA3294A129CA1294A329CA1294A3294A129CA3294A129CA3294A32",
INIT_19 => X"F5F78BCE7F8FF0F4FA955F7CF7F40A80145D55555556AAAAAAAAA94A329CA129",
INIT_1A => X"8E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E39B6CEDECDDF7DF7D",
INIT_1B => X"F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE38E3",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000001A1A33F9FCFE7F3F9FCFE7F3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"555FF00000000000000000000000000000000000000000000080000000000000",
INIT_28 => X"BC0010AAD5574BA557FFDFFF087BFDF45F7AA974AAAAAA97555F784174BAF7D5",
INIT_29 => X"515555508043FE00F7AA97555A2FBD7410AA8428AAAAAAE955450055421FFFFF",
INIT_2A => X"7D1575EFFFAA9555500557FE10FFFBEAA10007FD7410FFAA97400082A800AA08",
INIT_2B => X"0055574BA5D7FD7555A2D5575EF55517FF55A2AA97400552AAAB45082E80155F",
INIT_2C => X"500554200000003DE10FFD5401FFF7AAA8A10082EAAB45A2FFC2000007FD7400",
INIT_2D => X"10AA803FE105D516AABAFF843FFFFAA843DF55FFAA955EFA2D168B55557BEAB5",
INIT_2E => X"000AAAEBDF45A28428B45FFD168BFF00002AABA5D2ABFFFF087BD5545007BFDE",
INIT_2F => X"256DEB84104BAFFD1525FF000000000000000000000000000000000000000000",
INIT_30 => X"9756D145B401FFFFFFC7010BEDF524AA5571FDFEF1C7BFFF55FFA095482B6A49",
INIT_31 => X"4904380824850381C5B5057D1C003DE28F7A49057DAAF5D2428A2842AAAAA2AE",
INIT_32 => X"2AAFB451C2A8017DE3DF525FFFFA49756D145178E00EBFBE8A101475D5400F7A",
INIT_33 => X"2F1C50381471D74380851524BA5571D757DB6D5525EF555178F6DAAA49542841",
INIT_34 => X"AADB6FB7D5D7FEAB7D0855420BA1C0E3FE00E3DB471EFE3AAAAA00082EA8B6DA",
INIT_35 => X"F1C7BD057D1C71FFE10A28038E1049516AAB8FF8428FEFA28E3AF55F7A0925D7",
INIT_36 => X"00000000000000000000B6AEBDF45B68A28B6DEBDF6DBEF1C0A28AAA5524BFFF",
INIT_37 => X"F55F78017400F780001FFAA84000AAFFD1401E70000000000000000000000000",
INIT_38 => X"20BAAA8428AA2AAAA975FF5D7BC21EFF7FBD7400F7FBC00BA55557DFF7557BFD",
INIT_39 => X"EAA105D5155410FF84020AA0800154B2557FC01EF55043FEAAFF80021EFA2D14",
INIT_3A => X"568BE7AA80174AA082ABDF555D2A821EFAAFBC01FFF780155F7555568A00AAFF",
INIT_3B => X"AEA8A10082EA8BEFAAD5554B25551554BA0051400BA5551575EFF7D1401FF5D5",
INIT_3C => X"AAEAAB55F78400145AAFFFFFEF5D7FEABFF0051400A25D2EBFE10AAFFD55EFA2",
INIT_3D => X"552EA8AAA55043DFF7557BC01EF55557DE00AA842AA0000516AABAFF8428BE7A",
INIT_3E => X"0000000000000000000000000000000000000FFAABFF45FFAAAABFFAAFFFDFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024,               -- Port A enable input
WEA      => wbe_a_lo_1024(0),               -- Port A write enable input
DIA(0)   => data_write_a(6),        -- Port A data input
DOA(0)   => data_read_a_lo_1024(6),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024,               -- Port B enable input
WEB      => wbe_b_lo_1024(0),               -- Port B write enable input
DIB(0)   => data_write_b(6),        -- Port B data input
DOB(0)   => data_read_b_lo_1024(6),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_7_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10844B00482258A2842112C02450418800002300500030B313300C418992002",
INIT_01 => X"000009CA3839684D1CA0E0000E51424840000000080000080200080008510204",
INIT_02 => X"0120042086010000044600C00008000004100000000260900200000002402004",
INIT_03 => X"8628A10000082400000002408400080011000000610008000208C00000E14400",
INIT_04 => X"0911800100A000000000524084000040000050001140200100C8100000080102",
INIT_05 => X"0300812401011000000000002000114008008060441000000020024093000000",
INIT_06 => X"9190431C0D4010100000880804010010800000041080081000000200010424B2",
INIT_07 => X"000100AA0004408601000004860000008C02000A103010006928040800062481",
INIT_08 => X"84000048D484C20888000A0002120484C048007004000000000021F000000244",
INIT_09 => X"00A06009881201A520491004106C48A04040002400A15A208001650004001020",
INIT_0A => X"C99E1060201002044809C1040140A001004808810000459033189C0A400118A0",
INIT_0B => X"102000024040484050050041648A0041140C500B08821054C000264120000400",
INIT_0C => X"0404A083260E0832132011880462011880462051881462051881D31018C40620",
INIT_0D => X"0001000080001000813094801A8F80F00A600B52602801A88848011118003700",
INIT_0E => X"000003C007C002808228010410082042C000C000000004001002000400040002",
INIT_0F => X"A4000007800F80C840000800009864038A1200081C0014800000F001F0200052",
INIT_10 => X"00002C0E00E0E4004038000102400002C0E00E0D20100029000001E003E04000",
INIT_11 => X"2000C04031100E0403D0700300080908000100000661801E1900040380001804",
INIT_12 => X"0840878083E8003780A01043203A101780902043203A10082410082880000000",
INIT_13 => X"0601E0187900181035E0240806483248181035E0280410C8198818100DDD0000",
INIT_14 => X"0403774000201021E020FA006040376C00501022131210722060806D47000A40",
INIT_15 => X"00928A0002000110888600C032128201519480D40009902430160403E0E00506",
INIT_16 => X"01000000020080601802000000000405000A0020020081014134928820480010",
INIT_17 => X"0802018040000000006018020080200804010000000000806018020080000004",
INIT_18 => X"0000000001806008020000001006008020080001004008020080201004000020",
INIT_19 => X"0000000000000000000000000000400A004618618618C30C30C3000020180600",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000000B0840000000000000000000",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"1555500000000000000000000000000000000000000000000080000000000000",
INIT_28 => X"A97555F784174BAF7D5555FFF780155EFAAAEA8ABAAAFBFDE0055556AA005D04",
INIT_29 => X"55555EFAAFFFDFEFAAAAAAB455D556AA00FFAE95555087BFDF45F7AA974AAAAA",
INIT_2A => X"02EAAAAA082EA8A00AAAE955450055421FFFFFBC0010AAD5574BA557FFDFFF55",
INIT_2B => X"08043FE00F7AA97555A2FBD7410AA8428AAA557BFDFFF55003DFFFF7FBEAA000",
INIT_2C => X"0082A800AAF7AE975FFA28000010552EBDE00007BEAAAAA2D140000085155555",
INIT_2D => X"45087FEAB455D516AB55557BD55FF00557FE10FFFBEAA10007FD7410FFAA9740",
INIT_2E => X"000A2AA97400552AAAB45082E80155F7D1575EFFFAA955555D51574AAAAFFD55",
INIT_2F => X"AE105D556AA10410E17555000000000000000000000000000000000000000000",
INIT_30 => X"FFF55FFA095482B6A49256DEB84104BAFFD1525FFFF8E175C7A2AAAAA82A2F1F",
INIT_31 => X"F524AA5571FDFEF415B575D7AAF1FFFD7AAAAAFB7D495F6AA10E3AE905551C7B",
INIT_32 => X"003AFEFEBFBEAA001C2EA8A821C2EAAA00A2AE9756D145B401FFFFFFC7010BED",
INIT_33 => X"EDB470101C5B5057D1C003DE28F7A49057DAAF5D2428A2842AAAA497BFAFFF49",
INIT_34 => X"1475D5400F7A490438082485038F7A4905C7A28A070384120BDE100075EAA82B",
INIT_35 => X"D495150492BEF1D2555087BE8B7D555F6AB57417BC05D7145178E00EBFBE8A10",
INIT_36 => X"00000000000000000000AAA495428412AAFB451C2A8017DE3DF525FFFFA49756",
INIT_37 => X"555A2AEA8A10AAD568A00555168A10002E9754D0000000000000000000000000",
INIT_38 => X"8A10AAAE8215D557BFDF55F78017400F780001FFAA84000AAFFD1401E7FFAA97",
INIT_39 => X"C21EFF7FBD7400F7FBC00BA55557DFF7007BD5555AAD57DF55AAAEBDFEF007BE",
INIT_3A => X"428AA2007FE8BFF080028BFFAAFFEAA105D2EAAA005D2AAAA18AAAA975FF5D7B",
INIT_3B => X"043DE0000516AA10F7FBD7408557FC01EF55043FEAAFF80021EFA2D1420BAAA8",
INIT_3C => X"55568A00AAFFEAA105D5155410FF84020AA0800154B2FF8402145A2AA954AA00",
INIT_3D => X"AAFBC01FFF780155F7005140000FFD140145007FE8BEF557BEAB55087FC215D5",
INIT_3E => X"0000000000000000000000000000000000000AA80174AA082ABDF555D2A821EF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024,               -- Port A enable input
WEA      => wbe_a_lo_1024(0),               -- Port A write enable input
DIA(0)   => data_write_a(7),        -- Port A data input
DOA(0)   => data_read_a_lo_1024(7),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024,               -- Port B enable input
WEB      => wbe_b_lo_1024(0),               -- Port B write enable input
DIB(0)   => data_write_b(7),        -- Port B data input
DOB(0)   => data_read_b_lo_1024(7),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_8_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00000648E2840112C00000418000002700500030B3132000400812082",
INIT_01 => X"100008480009004C04A100000252024840000000180800080200010040110204",
INIT_02 => X"0020042000490000004600804008000005100000000024900200000002400004",
INIT_03 => X"0A0C33400008082400000080A4004B0891000020610112000040C00000E5C000",
INIT_04 => X"18800001000000000000512080000040800150400824280110C8100000120200",
INIT_05 => X"908084A10100100200004080280008240810802206940000012C214451610800",
INIT_06 => X"81B000080860109021400008040000202048020414A0021400040200322824C1",
INIT_07 => X"000000080004408049000004860000008402001A50208000630C040800062483",
INIT_08 => X"440000428644212280800A00021004044048002124000000000021F000000244",
INIT_09 => X"00004009001001010008100414644410400102228000D20080114502006409A2",
INIT_0A => X"000051312000042200294429148A4801C80C8C81000045907118040340020832",
INIT_0B => X"4020000240404140004D0544C4AA0001150410090302500011C813428A000400",
INIT_0C => X"46501090008820240240409000240009000240009000240009000120204808A5",
INIT_0D => X"42D1A168D09A301468402480004780F00140080860280004085904309A002196",
INIT_0E => X"00783FC00044340242280000000000020000C0000442106419120004034685A3",
INIT_0F => X"8000F07F800088A80000081EA2F9EC0000064004081010001E0FF00011104040",
INIT_10 => X"0ED0FC7E00000422201080000202658FC7E0000021882020003C1FE000222080",
INIT_11 => X"018059C3F350FE0C00000002A0040500000103961FE780000110010090000800",
INIT_12 => X"FD41FF80000830200021C1CF600012200010D1CF600012121600100810000004",
INIT_13 => X"9E1FE000010A1802100004343ED8000898021000087073D80008980200800002",
INIT_14 => X"0080200000BEB07FE00002086008020000209AEE3F300000246020200000620B",
INIT_15 => X"0088881903210000440610C8000A808040000208901786E4F0FE0C0000000166",
INIT_16 => X"685A1685A769DA368DA368DA769DA36CDA121A11A141800011309284002C0810",
INIT_17 => X"95A5685A1685A5695A368DA368DA769DA368DA368DA7695A1685A1685A5695A1",
INIT_18 => X"5A1695A568DA368DA369DA768DA1685A1695A5685A168DA369DA768DA368DA16",
INIT_19 => X"A4028A0A543EBC57A10A1E75D64108080468618618630C30C30C69DA5685A168",
INIT_1A => X"9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7BF3CCD8DF5B2DB2C",
INIT_1B => X"F87D3E1F4F87D3E1F4F87D3E1F4F87D3E1F4F87C3E1F0F87C3E1F0F87C3E79E7",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000006A6D4F87D3E1F4F87D3E1F4",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"155FF00000000000000000000000000000000000000000000080000000000000",
INIT_28 => X"BFDE0055556AA005D0415555080000000087BEAA10F7803DE00FFAEBFFFF0800",
INIT_29 => X"2AA8AAA557FC0010F780154105D7FC2145005155555F780155EFAAAEA8ABAAAF",
INIT_2A => X"7FFFFF55AA80155FF087BFDF45F7AA974AAAAAA97555F784174BAF7D5555FF55",
INIT_2B => X"AAFFFDFEFAAAAAAB455D556AA00FFAE95555AAFFE8A00552EBFE00F7D17FF45F",
INIT_2C => X"A557FFDFFF5504000AAAAAAA8B55F7D140010552E821EFAAAABDF555555555EF",
INIT_2D => X"55AA8028A00A2D57FF45557BE8A00AAAE955450055421FFFFFBC0010AAD5574B",
INIT_2E => X"000557BFDFFF55003DFFFF7FBEAA00002EAAAAA082EA8A00002AA8A10F784021",
INIT_2F => X"FE10F7AEBAFFF080A175D7000000000000000000000000000000000000000000",
INIT_30 => X"175C7A2AAAAA82A2F1FAE105D556AA10410E17555080E000280071E8A00EB8E3",
INIT_31 => X"4104BAFFD1525FF492EA8AAA5571C2000FF8A17400557FC015514555757DFF8E",
INIT_32 => X"2ABDE10EBDF7AF6DE3FFF8F7DB68A105D71C7BFFF55FFA095482B6A49256DEB8",
INIT_33 => X"AA0BDF6D415B575D7AAF1FFFD7AAAAAFB7D495F6AA10E3AE90555A2FBE8A3849",
INIT_34 => X"FFFFC7010BEDF524AA5571FDFEF550E00082B6A0AFB55F7D1420104124821D7A",
INIT_35 => X"01C2EA8A00F7800017DA2842FA00B6D578F6D557FFDA00A2AE9756D145B401FF",
INIT_36 => X"00000000000000000000497BFAFFF49003AFEFEBFBEAA001C2EA8A821C2EAAA0",
INIT_37 => X"0BA08556AA00AAAABFE00F7AEAABEF082E955450000000000000000000000000",
INIT_38 => X"21555D51575EFFFAA97555A2AEA8A10AAD568A00555168A10002E9754D082E82",
INIT_39 => X"17400F780001FFAA84000AAFFD1401E7082EAAABA5D5140010F7AE974105D7BC",
INIT_3A => X"E8215DA2FFE8ABA082ABFE00AAFBEABFFAAFBEABFFF7AA80145557BFDF55F780",
INIT_3B => X"D540000000402145AA843FFFF007BD5555AAD57DF55AAAEBDFEF007BE8A10AAA",
INIT_3C => X"AAA975FF5D7BC21EFF7FBD7400F7FBC00BA55557DFF75D2E82010F7843DF45FF",
INIT_3D => X"5D2EAAA005D2AAAA185D2AAAA10F780021FFA2803DE10FFD16ABFF5D7BFDE10A",
INIT_3E => X"0000000000000000000000000000000000000007FE8BFF080028BFFAAFFEAA10",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024,               -- Port A enable input
WEA      => wbe_a_lo_1024(1),               -- Port A write enable input
DIA(0)   => data_write_a(8),        -- Port A data input
DOA(0)   => data_read_a_lo_1024(8),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024,               -- Port B enable input
WEB      => wbe_b_lo_1024(1),               -- Port B write enable input
DIB(0)   => data_write_b(8),        -- Port B data input
DOB(0)   => data_read_b_lo_1024(8),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_9_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00018248A2840112C00002C18000002300500030B3132000400812006",
INIT_01 => X"400008000000004C0020000000100248413C0A61590001D90213C10008110204",
INIT_02 => X"01A0042080010000054600C04008000004100000001020900200200002420804",
INIT_03 => X"024003400008012400000010E4004B0891000020610310000144C00000F5C000",
INIT_04 => X"1801800100E000000000510084000040010050020810200000C8900000320200",
INIT_05 => X"918004311104100000000000200008100800002000100000002C234415610820",
INIT_06 => X"81B00008080010100000980804000008800042041080001000100200322C2481",
INIT_07 => X"0000811800044080010000058600000086020002502080006000040800062C80",
INIT_08 => X"0000004001D4618008800A00061004044048002004000000000061F000000244",
INIT_09 => X"000040090802009420409004104444084001022400214A2080014400026401A2",
INIT_0A => X"04000071200000A003CA294140200800C80C8C8100004590111C040040120800",
INIT_0B => X"12210002404848502847040164880021150400080222000200C8034200000000",
INIT_0C => X"4610088010080421021040841021000841021000841021000841010800420820",
INIT_0D => X"42D0A16C529A321068500484000500D10042080040284000084900001A002196",
INIT_0E => X"00000002804000004228010410082002C000C0002400046419120410034285A1",
INIT_0F => X"A00000000500800800000800000000000002290008001080000000A010100042",
INIT_10 => X"00000000000004C2001000000240000000000000680800280000000140202000",
INIT_11 => X"0000C0000000000000000442020001000001000000000000010C800080000804",
INIT_12 => X"08000000000801A7802010000000152780102000000015000600000800000000",
INIT_13 => X"000000000101900011E0240000000009500011E0280000000009500004DD0000",
INIT_14 => X"000137400020000000000201C000136C00101000000000002340002947000240",
INIT_15 => X"0080881901210000000600C280028000419480D4000010040000000000002304",
INIT_16 => X"68DA368DA1685A1685A1685A1685A16C5A121A13A141950051309284A82C0010",
INIT_17 => X"85A1685A1685A1685A368DA368DA368DA368DA368DA368DA368DA368DA368DA3",
INIT_18 => X"5A1685A168DA368DA368DA368DA368DA368DA368DA3685A1685A1685A1685A16",
INIT_19 => X"0157344CCCF48DE68A895C38E2540A8010100000000000000000685A1685A168",
INIT_1A => X"14514514514514514514514514514514514D34D34D34D34D28E1004039248209",
INIT_1B => X"D268341A4D268341A0D069349A0D069349A0D068341A0D068341A0D068345145",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000014D490D069349A0D068341A4",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"EAABA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"03DE00FFAEBFFFF0800155FFAAFBE8B45002A974AAAA803DFFFAA843DF45FFFF",
INIT_29 => X"7BFDE00A2FBD7400F7FBFDFFFA2AEBDE00AAFBEAABA080000000087BEAA10F78",
INIT_2A => X"055401FFF7AEAAA10F780155EFAAAEA8ABAAAFBFDE0055556AA005D041555508",
INIT_2B => X"557FC0010F780154105D7FC2145005155555557BE8BEF007FFDEAAAAD1555EF0",
INIT_2C => X"AF7D5555FFF780154AA5D2AA8A10F7AA974AA082E80010A2AAAAA10552AA8AAA",
INIT_2D => X"BAF7D17FEBAA2AEBDF45002EAAABA087BFDF45F7AA974AAAAAA97555F784174B",
INIT_2E => X"000AAFFE8A00552EBFE00F7D17FF45F7FFFFF55AA80155FF080400145FFFBEAA",
INIT_2F => X"8FC7BE8A3DF7DF7F5E8A92000000000000000000000000000000000000000000",
INIT_30 => X"000280071E8A00EB8E3FE10F7AEBAFFF080A175D7BEF1E8B6D002090482B68E3",
INIT_31 => X"56AA10410E175550871FFE00A2FBD0400FFF5FDFC7B6A0BDE38B6F5E8A92080E",
INIT_32 => X"7BFAE82A2DB555C71C5B451D7FFAAA8A38FF8E175C7A2AAAAA82A2F1FAE105D5",
INIT_33 => X"2AEADA38492EA8AAA5571C2000FF8A17400557FC015514555757D5D71E8BEF14",
INIT_34 => X"B6A49256DEB84104BAFFD1525FFFF84174BA5D20AAA00E3AA904BA142A87010A",
INIT_35 => X"7000400155FFFBEDA82FFD57DEBAAAA0BFF7D0024ADA921C7BFFF55FFA095482",
INIT_36 => X"00000000000000000000A2FBE8A38492ABDE10EBDF7AF6DE3FFF8F7DB68A105D",
INIT_37 => X"BEF080402000F7AAA8B55FFAABDFEFF7D16AA000000000000000000000000000",
INIT_38 => X"FEAAFFD16AA00082E820BA08556AA00AAAABFE00F7AEAABEF082E95545F7D568",
INIT_39 => X"A8A10AAD568A00555168A10002E9754D00517DE00A2FFC2000F7D17FF55FF803",
INIT_3A => X"1575EF555568BEF5D7FE8A10AAFFD55555D7FD5555FFAAA8AAAFFAA97555A2AE",
INIT_3B => X"AE800AA552A97400A2AEBDEAA082EAAABA5D5140010F7AE974105D7BC21555D5",
INIT_3C => X"57BFDF55F78017400F780001FFAA84000AAFFD1401E7FF80174AA5D0028A00AA",
INIT_3D => X"AAFBEABFFF7AA80145080002145F7FBFFE00FFD17FEAAA2803DFEF08043FE005",
INIT_3E => X"0000000000000000000000000000000000000A2FFE8ABA082ABFE00AAFBEABFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024,               -- Port A enable input
WEA      => wbe_a_lo_1024(1),               -- Port A write enable input
DIA(0)   => data_write_a(9),        -- Port A data input
DOA(0)   => data_read_a_lo_1024(9),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024,               -- Port B enable input
WEB      => wbe_b_lo_1024(1),               -- Port B write enable input
DIB(0)   => data_write_b(9),        -- Port B data input
DOB(0)   => data_read_b_lo_1024(9),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_10_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00018248A2840112C00002C18000202300500030B3132000400992006",
INIT_01 => X"254008000000004C002000000010026840000000080000080200010008110204",
INIT_02 => X"0020042000010000004455800008000004100000000000900200000002400004",
INIT_03 => X"020001021089000021081000C400090011000000610001540104C00000F14400",
INIT_04 => X"0811800101A00002000050088554004200C840000000200080C8100000000001",
INIT_05 => X"030080001000100800009400200000000840E020201000000024024001200020",
INIT_06 => X"81B00008080012120004CC080492500280208004148000100000020020042493",
INIT_07 => X"0000000800044080010000048404081085020002502000006000040800062480",
INIT_08 => X"100202400084410808000A00021004044048000004000000000021F020408264",
INIT_09 => X"010040090002008420401004144440004040022484214A2080110108C2C00320",
INIT_0A => X"04004166A48A0001080000000000080080181881000045901118044040020800",
INIT_0B => X"1201000200484910000F0105602622291404020902005002018002400A022000",
INIT_0C => X"0440001011808020120004801120044800120004801120044800110002400884",
INIT_0D => X"008000440210100041308480800F82F00040180260A808008848000018002104",
INIT_0E => X"000000028040000002280104100820020000400020000440100204100A000100",
INIT_0F => X"040000000500800800000000000000000002280008000400000000A010100010",
INIT_10 => X"00000000000004C2001000010000000000000000680800010000000140202000",
INIT_11 => X"200000000000000000000442000001000000000000000000010C000080001000",
INIT_12 => X"00000000000801C0008000000000154000800000000015000410000800000000",
INIT_13 => X"0000000001019800180000080000000958001800000400000009580002800000",
INIT_14 => X"0000A0000000000000000201E0000A0000400000000000002360002080000800",
INIT_15 => X"0080881000000000000600C28102800060000000000800000000000000002306",
INIT_16 => X"401004010040100401004010040100441020D0030008840051309A90BA884010",
INIT_17 => X"0902409024090240900401004010040100401004010040100401004010040100",
INIT_18 => X"1004010040902409024090240902409024090240902409024090240902409024",
INIT_19 => X"F546890A940FE0D3971243555205428290100000000000000000401004010040",
INIT_1A => X"8A28A28A28A28A28A28A28A28A28A28A28A28A28A28A28A29554199854514514",
INIT_1B => X"2B95CAE532994CA6532995CAE572B94CA6532994CA6532994CA6532994CA28A2",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000002718E72B94CA6532994CA657",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"FDE1000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"03DFFFAA843DF45FFFFEAABA007FC2155F7D155545AA80001EFAAFBEAB45557F",
INIT_29 => X"042AB55FFD168B55AA8000010FFFBE8BFFF78402155AAFBE8B45002A974AAAA8",
INIT_2A => X"AD16AABA002ABDE10080000000087BEAA10F7803DE00FFAEBFFFF0800155FF00",
INIT_2B => X"A2FBD7400F7FBFDFFFA2AEBDE00AAFBEAABAA2FFD741055003DFEFF7AA801FFA",
INIT_2C => X"05D0415555007FD74105555555EFF7FBC0145F78028A00A2D142155087BFDE00",
INIT_2D => X"55AAD168ABA002A975FFF7AEBDEBAF780155EFAAAEA8ABAAAFBFDE0055556AA0",
INIT_2E => X"000557BE8BEF007FFDEAAAAD1555EF0055401FFF7AEAAA105D042ABFF5D556AB",
INIT_2F => X"71D7AAFBEFB455D71F8E00000000000000000000000000000000000000000000",
INIT_30 => X"E8B6D002090482B68E38FC7BE8A3DF7DF7F5E8A92007BC217DEBDB55555AA8E0",
INIT_31 => X"EBAFFF080A175D700042AB7DEBDB6DB55BE8E05000EBFFE8BC7E38E07145BEF1",
INIT_32 => X"0A3DFD7F7A4821D7A2D16FA82142EB8E00080E000280071E8A00EB8E3FE10F7A",
INIT_33 => X"ED1421450871FFE00A2FBD0400FFF5FDFC7B6A0BDE38B6F5E8A92B6FBD541049",
INIT_34 => X"A2F1FAE105D556AA10410E175550071D54104951555D7EBF5C5155E3842AA00B",
INIT_35 => X"8410E2ABD749516FB55BED16FA820820955EFE3AEBDEAAFF8E175C7A2AAAAA82",
INIT_36 => X"000000000000000000005D71E8BEF147BFAE82A2DB555C71C5B451D7FFAAA8A3",
INIT_37 => X"1EFA2FFD7545AAAE97555A2FBFDF455D556AA000000000000000000000000000",
INIT_38 => X"8B45AAAA95545F7D568BEF080402000F7AAA8B55FFAABDFEFF7D16AA00087FC0",
INIT_39 => X"6AA00AAAABFE00F7AEAABEF082E9554500042ABFFA2FFFFF45F7AE97400AAFFE",
INIT_3A => X"16AA00FFFBD5400082EBFF45F78400155A2D57FE00552EA8A00082E820BA0855",
INIT_3B => X"D557555A2802AA10FFD54214500517DE00A2FFC2000F7D17FF55FF803FEAAFFD",
INIT_3C => X"FAA97555A2AEA8A10AAD568A00555168A10002E9754D085155410085557555AA",
INIT_3D => X"5D7FD5555FFAAA8AAA002AAAB4508557DF55F7D17FE000804155FFAAAABDEAAF",
INIT_3E => X"0000000000000000000000000000000000000555568BEF5D7FE8A10AAFFD5555",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024,               -- Port A enable input
WEA      => wbe_a_lo_1024(1),               -- Port A write enable input
DIA(0)   => data_write_a(10),        -- Port A data input
DOA(0)   => data_read_a_lo_1024(10),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024,               -- Port B enable input
WEB      => wbe_b_lo_1024(1),               -- Port B write enable input
DIB(0)   => data_write_b(10),        -- Port B data input
DOB(0)   => data_read_b_lo_1024(10),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_11_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"A101C4B05A0034CA2840712C2D001419000002300500030B31B20084EC992002",
INIT_01 => X"90000986B83028491800E0000C26426040000000080000088200080802512224",
INIT_02 => X"1A2004205E010640024D00800008000004100000040EC090820018003241A00C",
INIT_03 => X"28639100000C5C00000045C08400C8001100000061806A001618C03001E54400",
INIT_04 => X"1A800001000009A0804059A190000040400040008058220008C8100000120D4E",
INIT_05 => X"02000E81080250010000002022000058080400000E1200000020004401000004",
INIT_06 => X"819435143F20101010001008040800B8100102041088011100022200000024B2",
INIT_07 => X"90640D280884453E01064002944180008402001295BA100022E4340800062D82",
INIT_08 => X"400000093204802200280A0012160585C1D808D004000000000323F40C102244",
INIT_09 => X"380040098010001100009204107C5950400000220080C200800900020C006827",
INIT_0A => X"80007100004016EA080801010000080D00200081000045B0511D289940103399",
INIT_0B => X"002000024040410A000D0104408810C115D9C008050042400100D04E88000002",
INIT_0C => X"00655010009264201200C7B421ED0C7B421ED0C7B431ED087B43176843DA1085",
INIT_0D => X"0401020080400A10012494881A4F80F209500BB2602881A488485C1318002000",
INIT_0E => X"6619A540124814800228010410082022C00040002020090020220C9600040802",
INIT_0F => X"ACCC334A802491600C587949B6D0141B4CC600D5761B1599865A500490B86A56",
INIT_10 => X"BAC845542056A61686EC81E3A6CB68AA2C622C9A251C352B330CB4A0092170D8",
INIT_11 => X"BCCAD0B5A81536080CC6B21A21B1FC09CB0F1076D4A200B2AD4068F4101639B5",
INIT_12 => X"4D2CC281E31AA0103AB8D5514066380804B268A2E060901204112566F10AC418",
INIT_13 => X"D551443C47281002540B2C9AAAA8662A1152B202AE3554403028115AA88201A1",
INIT_14 => X"548A20A0492A2724A0621620402A020141F172FB182A32AB6845AB6200251BC9",
INIT_15 => X"00C00A000200074044E6801832728080D00A380B753952C4877E0104DDE4D124",
INIT_16 => X"0080200802008020080200802008020480080022020081010124988800400010",
INIT_17 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_18 => X"0000000000802008020080200802008020080200802008020080200802008020",
INIT_19 => X"55062608804180C0B10A42104201400204000000000000000000000000000000",
INIT_1A => X"00000000000000000000000000000000000820820820820801C4149470000000",
INIT_1B => X"0000000000000000040200000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000007E0F0000000000000100800",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"000AA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0001EFAAFBEAB45557FFDE10082ABDF5508557DF45002ABDFFFF7803DE10AA80",
INIT_29 => X"AEBFF45FFAEBFEAA002A801FFF7FFE8A10A28000000007FC2155F7D155545AA8",
INIT_2A => X"2AABFE10082ABFFEFAAFBE8B45002A974AAAA803DFFFAA843DF45FFFFEAABAA2",
INIT_2B => X"FFD168B55AA8000010FFFBE8BFFF78402155AAD155555A28428BFF002ABDE00A",
INIT_2C => X"F0800155FF00557FF45557FC2010002A80010A2842AAAA007BFFF4500042AB55",
INIT_2D => X"FF5D00154BAF7FBE8BEFFFD540000080000000087BEAA10F7803DE00FFAEBFFF",
INIT_2E => X"000A2FFD741055003DFEFF7AA801FFAAD16AABA002ABDE10A2D168A10A284021",
INIT_2F => X"DFC7F78E3FE28B684070AA000000000000000000000000000000000000000000",
INIT_30 => X"C217DEBDB55555AA8E071D7AAFBEFB455D71F8E00002EBDF6D005B78F7D142AB",
INIT_31 => X"A3DF7DF7F5E8A92BEAEBFF7DEBA0BDEAA1C2A801C7E3FFEFA10B68407038007B",
INIT_32 => X"8A28BFF082ABAE10B6AAB8E280820B8FEFBEF1E8B6D002090482B68E38FC7BE8",
INIT_33 => X"07FF8F7D00042AB7DEBDB6DB55BE8E05000EBFFE8BC7E38E07145B6D15756DA2",
INIT_34 => X"EB8E3FE10F7AEBAFFF080A175D708517DF7D497BC5028142A87000A28A2AA920",
INIT_35 => X"0B6DB6AA28A280001FF5D0A10482FFFFEFBC7E3DF42028080E000280071E8A00",
INIT_36 => X"00000000000000000000B6FBD5410490A3DFD7F7A4821D7A2D16FA82142EB8E0",
INIT_37 => X"FEF007BE8BFF5D2ABDF55F7AABDEAAF784154BA0000000000000000000000000",
INIT_38 => X"DE00FF84154BA087FC01EFA2FFD7545AAAE97555A2FBFDF455D556AA00082EBF",
INIT_39 => X"02000F7AAA8B55FFAABDFEFF7D16AA00FFAEBFFEFAA803DEBA5D2E82155A2FBF",
INIT_3A => X"A95545F7D5555FFAAAAA8BFF002AAAA00FFAAA8AAA080028BFFF7D568BEF0804",
INIT_3B => X"2E95400A2AEA8A00007FEABFF00042ABFFA2FFFFF45F7AE97400AAFFE8B45AAA",
INIT_3C => X"82E820BA08556AA00AAAABFE00F7AEAABEF082E9554508557DFFF007BD54BA5D",
INIT_3D => X"A2D57FE00552EA8A00FFFFE8AAAAA80001FF5D2E82000F7FFFFF45AAFFC20BA0",
INIT_3E => X"0000000000000000000000000000000000000FFFBD5400082EBFF45F78400155",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024,               -- Port A enable input
WEA      => wbe_a_lo_1024(1),               -- Port A write enable input
DIA(0)   => data_write_a(11),        -- Port A data input
DOA(0)   => data_read_a_lo_1024(11),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024,               -- Port B enable input
WEB      => wbe_b_lo_1024(1),               -- Port B write enable input
DIB(0)   => data_write_b(11),        -- Port B data input
DOB(0)   => data_read_b_lo_1024(11),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_12_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50080B01BC002006940202C0DE041196A83183000000023322287E0FC000006",
INIT_01 => X"75400D849830C84C5823E0000C17424840000000080000088200002802153231",
INIT_02 => X"18A026B43ED180040147558040090000061800000C06ED9802768F4472C52005",
INIT_03 => X"2A67E34A528D0524A52850528400C8001100000171C02B550618C91A10E55440",
INIT_04 => X"1BC0000100056C8280825DE98154004300C840800850240080CA921084520A07",
INIT_05 => X"02000F832000500C0000941024000852084060202E100001002000448100000C",
INIT_06 => X"819A1D1C3FE01A1A40045408049A50BA4020C6041090001200006200000000F2",
INIT_07 => X"C26A0719CC96CC6ED18A64019695A854870300FA3968B20068FC06080106249F",
INIT_08 => X"D002024B3E040800008C0A002610240D494A06F3460409000000E3F0AD5282E5",
INIT_09 => X"27A06009200040000400120412445D78400001000410420080218029CC807A27",
INIT_0A => X"18000006848A026F000000000000080000F010C100204593F11A6CDF48003BF8",
INIT_0B => X"000000820040402B28050400400432C9349DF21A31A00ACC0000F04F80020001",
INIT_0C => X"00357804611AE45D05D0833430CD0833420CD0C33420CD0833430668619A1000",
INIT_0D => X"0000000000000A74812DF00E87E80A079F9F90FA0280E87E800C7FF3B8002000",
INIT_0E => X"3B6B0E404D26160682082002000401EA0000C40000800A006002818808000000",
INIT_0F => X"A476D61C809A4DA84272592D6246FC1B17B541F97E1B348EDA93900B2B286C56",
INIT_10 => X"30C669E622DBC325CFD881A962454CFBE5403AB99594362B1DB52720165650D9",
INIT_11 => X"F8D2D39A3745261E4A95A110A3F855000E4B1D32BAB504BB7490FCFF912A3834",
INIT_12 => X"B90E9B018C7530200AB8F8BF41F9A22006B37DC8E1F9A21A70116D4C5080651C",
INIT_13 => X"118780319CCA08AB1001ACDF34B8F1C688AB1002AE3F7B807B6289F368828C4C",
INIT_14 => X"2AF020233376A5ECC016B1A827CDA21160F051DE610A34C50427E6E220323E4A",
INIT_15 => X"0077020000000439FDC05C5806781FAB46095A0B5199B0AC55521524F1864022",
INIT_16 => X"000000000000000000000000000000000026C000002884000130921092804010",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"8020080200000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0051B946088881360A95090CB054420290100000000000000000008020080200",
INIT_1A => X"041041041041041041041041041041041049249249249249200100002D451451",
INIT_1B => X"92C964B2592C964B2592C964B2592C964B2592C86432190C86432190C8641041",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000003800F592C964B2592C964B25",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"7DE1000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"ABDFFFF7803DE10AA80000AAAA843FE0008557DFFF0800020105D557FEAA0055",
INIT_29 => X"D5420000051555FFA2AA8200000557DFFFF7AA80000082ABDF5508557DF45002",
INIT_2A => X"82AA8AAAAAFFC00BA007FC2155F7D155545AA80001EFAAFBEAB45557FFDE10AA",
INIT_2B => X"FFAEBFEAA002A801FFF7FFE8A10A28000000A2D155410F7FFFFEBA08003FE000",
INIT_2C => X"5FFFFEAABA000028A105D2ABFE10A2AABFE1055516ABEF5D517DEAAA2AEBFF45",
INIT_2D => X"55002A820AA08557DFFFF7AA82155AAFBE8B45002A974AAAA803DFFFAA843DF4",
INIT_2E => X"000AAD155555A28428BFF002ABDE00A2AABFE10082ABFFEF0855420000004175",
INIT_2F => X"5010495B7AE921C517DE10000000000000000000000000000000000000000000",
INIT_30 => X"BDF6D005B78F7D142ABDFC7F78E3FE28B684070AABE803AE38145B78FD700000",
INIT_31 => X"BEFB455D71F8E00BED547038145B505FFB6A487000005F7AFD7F7A482038002E",
INIT_32 => X"F1FDE821C003FE001C2EAAAAAB6F5C2082007BC217DEBDB55555AA8E071D7AAF",
INIT_33 => X"D517DEAABEAEBFF7DEBA0BDEAA1C2A801C7E3FFEFA10B68407038B6D550428FF",
INIT_34 => X"B68E38FC7BE8A3DF7DF7F5E8A9200002FA285D20BDE28A2A4B8E10555B68BEF5",
INIT_35 => X"F085F47038140010555142082082005F7DFD7F7A482155BEF1E8B6D002090482",
INIT_36 => X"00000000000000000000B6D15756DA28A28BFF082ABAE10B6AAB8E280820B8FE",
INIT_37 => X"ABA5D7FEAB45080015410007FEAA0055517DE000000000000000000000000000",
INIT_38 => X"AB45F780020BA082EBFFEF007BE8BFF5D2ABDF55F7AABDEAAF784154BAF7802A",
INIT_39 => X"D7545AAAE97555A2FBFDF455D556AA00F7D1554BA5D7BC01FFFF8015410007FE",
INIT_3A => X"4154BAF7D1400BAFFD57FE005D043FE10552EAAAAAFFD140000087FC01EFA2FF",
INIT_3B => X"8428A105D7FEABEF55557DEBAFFAEBFFEFAA803DEBA5D2E82155A2FBFDE00FF8",
INIT_3C => X"7D568BEF080402000F7AAA8B55FFAABDFEFF7D16AA0008003FEBA55003DEBAA2",
INIT_3D => X"FFAAA8AAA080028BFF087BD54AA550402145550000010087FFFF45F78402145F",
INIT_3E => X"0000000000000000000000000000000000000F7D5555FFAAAAA8BFF002AAAA00",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024,               -- Port A enable input
WEA      => wbe_a_lo_1024(1),               -- Port A write enable input
DIA(0)   => data_write_a(12),        -- Port A data input
DOA(0)   => data_read_a_lo_1024(12),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024,               -- Port B enable input
WEB      => wbe_b_lo_1024(1),               -- Port B write enable input
DIB(0)   => data_write_b(12),        -- Port B data input
DOB(0)   => data_read_b_lo_1024(12),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_13_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10154A0441836CA2840512822007C18000E02700500030B31B300040081A042",
INIT_01 => X"00000804A000C04800020000000002404001000008220008A200100802110204",
INIT_02 => X"02200430000104000A4700804008000004100000000420918204D3033240400D",
INIT_03 => X"AA4003400008592400000590C40009141100000C6180C0000000C00001E14000",
INIT_04 => X"0800000102400120088054019000004160004190BAA0270000C8100000600206",
INIT_05 => X"21000012040610050040000227003AA0082400E94C1200000824424005220020",
INIT_06 => X"81963B180C001010580000080400000058000004109C00138000020024142581",
INIT_07 => X"002C8008000441600106400A9600010494020002B8AAA000EF003408000E2580",
INIT_08 => X"000000E48194408000A00A001210040441C80320040210000002ABF004102244",
INIT_09 => X"2A004009640040100400940412D4C4004000022000104200802D983000480120",
INIT_0A => X"8000202020401480000000000000080C90090881000145B0111A14004015080D",
INIT_0B => X"00000002004040AA08050400404040C11444000805200A402090024000008002",
INIT_0C => X"8410000A00280020020040800020040800020000801020000800010020400000",
INIT_0D => X"84A14250A055100050100490000500D00040080040290000084E4000B800610C",
INIT_0E => X"DCD13042BEDA36820228000000000000C000400081A08BC812A2092B02850942",
INIT_0F => X"89B9A260857DB400431969CA985D480949D32804A40AB137341C10B7D6A02EC0",
INIT_10 => X"E6ACA678001CE7D0296C213A460CA4271CA2168AEC1017606E6838216FAD4055",
INIT_11 => X"84AD4961C281B20213073C5FC0058008632D30D522CE80239DCC01AB013A4D20",
INIT_12 => X"2E6B13804A4B01D83461299900F6BD583A519104A0EEBD1A141010B2A4C8E116",
INIT_13 => X"89E5E40913419151EE0E94641828F72B5151EE0D184B321037AF5158BB02D085",
INIT_14 => X"562EC0B42162D68EE0073AE1C562EC13D521921A4170300B2B458B56B01C2280",
INIT_15 => X"00888A120240034000E6DC8285028014B82372011FC1E4F5E0A00929684EAF84",
INIT_16 => X"50942509425094250942509425094254940A1421420082020120908800480030",
INIT_17 => X"0942509425094250942509425094250942509425094250942509425094250942",
INIT_18 => X"9425094250942509425094250942509425094250942509425094250942509425",
INIT_19 => X"F7EFBBEEFF3F7DF7FF3E9F7DF7E2450228000000000000000000509425094250",
INIT_1A => X"BAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBF7DFDFDDD555555",
INIT_1B => X"EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAEBAE",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000000000F7EBF5FAFD7EBF5FAFD7",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"2ABEF00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0020105D557FEAA00557DE10AAD5554BA087FFFF55557BD54AAF7FBC01FFA280",
INIT_29 => X"7BD75EF087FFFFEF557BEAB45552E80155AA802AB45AA843FE0008557DFFF080",
INIT_2A => X"FAE820AA5D5557555082ABDF5508557DF45002ABDFFFF7803DE10AA80000AA08",
INIT_2B => X"0051555FFA2AA8200000557DFFFF7AA80000AAD1420AA087BD7555FFD168AAAF",
INIT_2C => X"5557FFDE10AAAEA8BFFA2FBD7545FFD157555085140010F7AEAABFFAAD542000",
INIT_2D => X"BA557BE8A10A284154BAFFAAAAB45007FC2155F7D155545AA80001EFAAFBEAB4",
INIT_2E => X"000A2D155410F7FFFFEBA08003FE00082AA8AAAAAFFC00BA00002AAAAF7D5574",
INIT_2F => X"0492E3F1C71C7BE8A2ABD7000000000000000000000000000000000000000000",
INIT_30 => X"3AE38145B78FD7000005010495B7AE921C517DE10A2DB50482147FFAF554971D",
INIT_31 => X"E3FE28B684070AA1C71D25D7007FFAFD7497BE8B5555208217DBE8A2AB45BE80",
INIT_32 => X"7FD257DFFD568A82FFA4870BA555F5056D002EBDF6D005B78F7D142ABDFC7F78",
INIT_33 => X"FAAAFBFFBED547038145B505FFB6A487000005F7AFD7F7A482038AADF4709214",
INIT_34 => X"AA8E071D7AAFBEFB455D71F8E00A2A0ADBC7A2FFD257DE3DF52555085142000F",
INIT_35 => X"21C002AA92FFDF574824171EAA10B680124BAFFAAAFB45007BC217DEBDB55555",
INIT_36 => X"00000000000000000000B6D550428FFF1FDE821C003FE001C2EAAAAAB6F5C208",
INIT_37 => X"0105D7BE8B55085142010AAD157545F7AEA8B550000000000000000000000000",
INIT_38 => X"01EFF7AAA8B55F7802AABA5D7FEAB45080015410007FEAA0055517DE00A2FFC0",
INIT_39 => X"E8BFF5D2ABDF55F7AABDEAAF784154BA5D5140145007BE8B55087BEAB555D040",
INIT_3A => X"0020BAA2FFD54105D7FC21EFFFD16AA10FF80174AA557FC21EF082EBFFEF007B",
INIT_3B => X"FBC0155085540000FFAEBFFEFF7D1554BA5D7BC01FFFF8015410007FEAB45F78",
INIT_3C => X"87FC01EFA2FFD7545AAAE97555A2FBFDF455D556AA00A2803FF45AAFFC21EFAA",
INIT_3D => X"552EAAAAAFFD1400005D042AA00F7FBD5410085568A10FF80020AAFFAABFF550",
INIT_3E => X"0000000000000000000000000000000000000F7D1400BAFFD57FE005D043FE10",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024,               -- Port A enable input
WEA      => wbe_a_lo_1024(1),               -- Port A write enable input
DIA(0)   => data_write_a(13),        -- Port A data input
DOA(0)   => data_read_a_lo_1024(13),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024,               -- Port B enable input
WEB      => wbe_b_lo_1024(1),               -- Port B write enable input
DIB(0)   => data_write_b(13),        -- Port B data input
DOB(0)   => data_read_b_lo_1024(13),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_14_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10020A000180000284008280000281800000030000000033022000000580002",
INIT_01 => X"000008020000204D006800000030824840000000084000084200090008510200",
INIT_02 => X"0220043170010A600A4D008040080000041000000028009002000F333240800C",
INIT_03 => X"111813400008002400000000C400090011000000610200001104D83000F14000",
INIT_04 => X"0801800100A000000000540084000040000040000800200000C8100000000748",
INIT_05 => X"0100000000001000000000002000080008000000001000000024024001200020",
INIT_06 => X"819EB84028001010000000080400000000000004108000100000020020040081",
INIT_07 => X"92040608000440100102400A94810206844200021DA2A0002000340800062C80",
INIT_08 => X"000000000084400008800A001214040441481500040000000000A7F408002244",
INIT_09 => X"0A0040090002008420401004104444004000020400214A208001000002400120",
INIT_0A => X"0400002020000000000000000000080C8008088100004590111B480040120000",
INIT_0B => X"1000000200404800000504016000002114000008020000020080024000000000",
INIT_0C => X"0410000010000000000040001000000000000040000000000001000000000000",
INIT_0D => X"04810244825010004010000000000000000000000000000000080000B8002104",
INIT_0E => X"0002C38280001202020800000000001000004000000000401022000002040902",
INIT_0F => X"20000587050001404E8084341CBA3404800828805200008000E0E0A000080002",
INIT_10 => X"4D18178E012010C00224004091C3514072C000444A0400080001C1C140001000",
INIT_11 => X"51709A07424142084458476001003809D0104B01C5710044020C4006010500C5",
INIT_12 => X"C26EE3803180C18006519462A00005001460E4730000050A1011004001060049",
INIT_13 => X"01F9E00660318000000538318740000140000001B4600CE80001400000002B62",
INIT_14 => X"0000000AD89857B0E0684411800000003799EB764D000330C300000000E3554B",
INIT_15 => X"0000021002002C000024008284001A0902000422E3F5960080480A0216A07240",
INIT_16 => X"4090240902409024090240902409024090081021020080015134920800480010",
INIT_17 => X"0902409024090240902409024090240902409024090240902409024090240902",
INIT_18 => X"9024090240902409024090240902409024090240902409024090240902409024",
INIT_19 => X"F5579B4E5C8FF0F7BE9D5F7DF650400200000000000000000000409024090240",
INIT_1A => X"9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7BF7DDDDDFCF3CF3D",
INIT_1B => X"F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE79E7",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000003FFF03F9FCFE7F3F9FCFE7F3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"420BA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"BD54AAF7FBC01FFA2802ABEFA2FBE8B55A2AE80000F7D5555555D2AAAABAAAD1",
INIT_29 => X"AA801FFA28402000AAAE955455500155EF0804155EFAAD5554BA087FFFF55557",
INIT_2A => X"7AEA8B45080417400AA843FE0008557DFFF0800020105D557FEAA00557DE10A2",
INIT_2B => X"087FFFFEF557BEAB45552E80155AA802AB4500516AA00A2AE800BAFFFFC20BAF",
INIT_2C => X"0AA80000AA005568ABAA28402010A2843FEBAFFFBD7410A2D168BFF087BD75EF",
INIT_2D => X"005D7FFDF4555517DFEF00043FEAA082ABDF5508557DF45002ABDFFFF7803DE1",
INIT_2E => X"000AAD1420AA087BD7555FFD168AAAFFAE820AA5D5557555002E80155A280000",
INIT_2F => X"0555412AA8ABAAADB40092000000000000000000000000000000000000000000",
INIT_30 => X"50482147FFAF554971D0492E3F1C71C7BE8A2ABD7A2FFEDB55B6A080038E3DB5",
INIT_31 => X"B7AE921C517DE10A2AE851FFB68402038AAAA955554900105FF0800175D7A2DB",
INIT_32 => X"A0800BAE3F1C0092EBAAADB6D080A12410BE803AE38145B78FD7000005010495",
INIT_33 => X"2D568BC71C71D25D7007FFAFD7497BE8B5555208217DBE8A2AB451C556FA00A2",
INIT_34 => X"142ABDFC7F78E3FE28B684070AA00516DABAA28402038B6803DE82F7F5D5410A",
INIT_35 => X"D002A80155B680000105D7FF8F455D5F78FD7000E3FEAA002EBDF6D005B78F7D",
INIT_36 => X"00000000000000000000AADF47092147FD257DFFD568A82FFA4870BA555F5056",
INIT_37 => X"F55FF84000AAAAFBC0145002AA8AAAAAFFC20000000000000000000000000000",
INIT_38 => X"01EF080417555A2FFC00105D7BE8B55085142010AAD157545F7AEA8B55A2FBFF",
INIT_39 => X"EAB45080015410007FEAA0055517DE00A2AA955FFFF80020BAAAAA9754508000",
INIT_3A => X"AA8B555D557FE00A280020BAAAD140000A2AEBFFEF082A82010F7802AABA5D7F",
INIT_3B => X"803DE00FFD557400AAD56AB455D5140145007BE8B55087BEAB555D04001EFF7A",
INIT_3C => X"82EBFFEF007BE8BFF5D2ABDF55F7AABDEAAF784154BA08557FEAAA284000AAFF",
INIT_3D => X"FF80174AA557FC21EF082A80145F780020105D7BEAB45557BE8B45082EBFEBA0",
INIT_3E => X"0000000000000000000000000000000000000A2FFD54105D7FC21EFFFD16AA10",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024,               -- Port A enable input
WEA      => wbe_a_lo_1024(1),               -- Port A write enable input
DIA(0)   => data_write_a(14),        -- Port A data input
DOA(0)   => data_read_a_lo_1024(14),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024,               -- Port B enable input
WEB      => wbe_b_lo_1024(1),               -- Port B write enable input
DIB(0)   => data_write_b(14),        -- Port B data input
DOB(0)   => data_read_b_lo_1024(14),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_15_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000A000000000284000280000001800020030000000033022000000180002",
INIT_01 => X"8000080000000048000000000000026040000000080000080200000000110200",
INIT_02 => X"0020042004010E60004C0080000800000410000000020090020000300245E005",
INIT_03 => X"0000010000080400000000408400480111000000610008000000C00000E54400",
INIT_04 => X"980000010000000088C2550080000040000040000008A00028C8100000120000",
INIT_05 => X"020004012E025000000001322000000A28008000011000000220004D41000000",
INIT_06 => X"819588000800101000011008040000100001060418800510000A620000000092",
INIT_07 => X"0000000800044004010C20008440810284020002102220002000340800062480",
INIT_08 => X"0000000001140800002C0A001214050540C800400406180000002DF004000244",
INIT_09 => X"1E00400900000000000016041044400440000000000042008001000000000022",
INIT_0A => X"0000000000000220000000000000080C00000081000045901118000040000000",
INIT_0B => X"0000000200404000010500004000000114000009000000000000004200000000",
INIT_0C => X"0000000000000000000040001000040001000000000000000001000020000800",
INIT_0D => X"000000000000001001208000180800000000030200000180800C400030002000",
INIT_0E => X"0000000000002600020800000000001080004000000000000002000000000000",
INIT_0F => X"A400000000000000000008000000000000000000000014800000000000000052",
INIT_10 => X"0000000000000000000000010240000000000000000000290000000000000000",
INIT_11 => X"2001C05838120800000000000000000000010000000000000000000000001804",
INIT_12 => X"081004000000000000A010000000000000902000000000180010002020000000",
INIT_13 => X"6600000000000000000024080000000000000000280400000000000000000000",
INIT_14 => X"0000000000200801000000000000000000501001920000000000000000000A40",
INIT_15 => X"0000020000000000000000003000000000000000000A101C3614000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000080000120980000000010",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000400200000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"28BEF00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"5555555D2AAAABAAAD1420BAFF8000010082A954BA00003DFEF085155400F784",
INIT_29 => X"AE95555A2FBE8BEFA2843DE00AA8015400FF84001EFA2FBE8B55A2AE80000F7D",
INIT_2A => X"2FBEAB45F7D56AABAAAD5554BA087FFFF55557BD54AAF7FBC01FFA2802ABEFF7",
INIT_2B => X"A28402000AAAE955455500155EF0804155EFFFFBE8BFF0800174AA557BFDE10A",
INIT_2C => X"A00557DE10F7D1574AAA2D16AB55FFD568BEF087FE8A1055003FE00A2AA801FF",
INIT_2D => X"00AA802AA00AAAE800BA5D0015545AA843FE0008557DFFF0800020105D557FEA",
INIT_2E => X"00000516AA00A2AE800BAFFFFC20BAF7AEA8B45080417400FFFFC21450800154",
INIT_2F => X"8FD7005150438F78A2DBFF000000000000000000000000000000000000000000",
INIT_30 => X"EDB55B6A080038E3DB50555412AA8ABAAADB40092E38E070280024904AA1C043",
INIT_31 => X"1C71C7BE8A2ABD7E3AA9257DA2FFE8BC7BE8E38E10A28017400E38A051FFA2FF",
INIT_32 => X"00124AA557FFDE10A2FBEDB6DF7D16AABAA2DB50482147FFAF554971D0492E3F",
INIT_33 => X"10038E38A2AE851FFB68402038AAAA955554900105FF0800175D7E3FFEFBD700",
INIT_34 => X"000005010495B7AE921C517DE10FFDF50482A2DB6AB45FFD56DBD7087BEAA384",
INIT_35 => X"0FFF1C017D140410400BE8E28A10AAA085082550A1057DBE803AE38145B78FD7",
INIT_36 => X"000000000000000000001C556FA00A2A0800BAE3F1C0092EBAAADB6D080A1241",
INIT_37 => X"4AA0800020BA550028B550855400AAF7AEBDFEF0000000000000000000000000",
INIT_38 => X"7400AAAE975EFA2FBFFF55FF84000AAAAFBC0145002AA8AAAAAFFC2000AAAA97",
INIT_39 => X"E8B55085142010AAD157545F7AEA8B55AAAE821EFAAFBEAB55F7AAA8A00AA841",
INIT_3A => X"417555AAFFFDF450804020AA557BFFE10A2FFFFFEFF7D568ABAA2FFC00105D7B",
INIT_3B => X"D17DF45007FE8AAA08002AAAAA2AA955FFFF80020BAAAAA975450800001EF080",
INIT_3C => X"7802AABA5D7FEAB45080015410007FEAA0055517DE00FFFBC2000AAFBE8B55F7",
INIT_3D => X"A2AEBFFEF082A82010FFD5421EF5D0000010F7AAA8A10AA8017400552A801EFF",
INIT_3E => X"00000000000000000000000000000000000005D557FE00A280020BAAAD140000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024,               -- Port A enable input
WEA      => wbe_a_lo_1024(1),               -- Port A write enable input
DIA(0)   => data_write_a(15),        -- Port A data input
DOA(0)   => data_read_a_lo_1024(15),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024,               -- Port B enable input
WEB      => wbe_b_lo_1024(1),               -- Port B write enable input
DIB(0)   => data_write_b(15),        -- Port B data input
DOB(0)   => data_read_b_lo_1024(15),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_16_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"DA22C618B1000482B688B186588884862A400438255FC38381441205BA803003",
INIT_01 => X"7045A80028404C211203A952A90341080B173340412000E1005D628000820484",
INIT_02 => X"428406A4000850848330118D0AAC55001349B108818005460229044001C01784",
INIT_03 => X"092C4020000500020000500986812C405000001A48202050000A214AC0650115",
INIT_04 => X"4804A55440256F504025E003A054F46415A4E62B6FE3307943965A00001A1152",
INIT_05 => X"0000001C40A5B950ADB8EA097057ECE14C86D2B7F85AAD17F4B100000B88148C",
INIT_06 => X"415401DCDCF2C0A8030140BCB0820A200342A1C641C1E8782F508F2B00003584",
INIT_07 => X"002701881A3202080AE00480A2002840BE1480FA004342AA6F12000054004867",
INIT_08 => X"08C54828091002000002B32A8C19064E486A8001510000014140C1E2A14891E0",
INIT_09 => X"015452B103020814004088B64102680B6596594800400413CAC0208944800000",
INIT_0A => X"96AA000484094C000000000000012C9000A0000D0A80000BF8028E87C1B99270",
INIT_0B => X"014808A02004200E540480212000A448C0082024AE50064B44000000000002A2",
INIT_0C => X"0004000D5846256AAEA811150445411150445411150445411150422A088A8200",
INIT_0D => X"00000004010042A204A0C5817D00005034052E40000817D00440004004AD3240",
INIT_0E => X"632B2673FA4587978A2004102800809225545155121740000004900090000000",
INIT_0F => X"00C6564CE7F4EA4B940076D296D003030800462CBD320018CAAAACFE9164C800",
INIT_10 => X"28834ADB1440A114793A4A30A40839AA14910D08DCB2640031955559FD3AC990",
INIT_11 => X"594AB0B1A025371CA0E034E8443C097A800EB090D4AAC91208ED2FA0CE5E09B1",
INIT_12 => X"7B50446083001B94BB38C540EBE61284BB304880E3E4579EDC00992980D58033",
INIT_13 => X"5511121840E7A2CD952ECC12ABC3E6ACB3DFB12ECE315000F61FF1727A85FDBC",
INIT_14 => X"75DEB07F6F2E7084517F126F8395CB2BEFBAB8BA8AF698228CC5E2F08ECA5159",
INIT_15 => X"5580A840A8009F8B108C80A1021B080AFC0DF6422C6077F4A77F20D0C0E21084",
INIT_16 => X"0000000000000000000000000000000000044000102A0001148442A110810359",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"558D11544C690DA64C1C4F68A360400000000000000000000000000000000000",
INIT_1A => X"14D14D14D14D14D14D14D14D14D14D14D14514514514514529E5F87869E79E78",
INIT_1B => X"D1E8F47A3D1E8F47A7D3E9F4FA7D3E9F4FA7D3E9F47A7D1E9F47A7D1E9F4D14D",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000007D3E9F4FA7D3E8F47A3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"C00AA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"03DFEF085155400F78428BEF087FFFFEFF7D168B55AAD17FFFF552EBFE00007F",
INIT_29 => X"2E975EFF7D568BFFFF80175EF0004000BA552A821FFFF8000010082A954BA000",
INIT_2A => X"55540000082EAABFFA2FBE8B55A2AE80000F7D5555555D2AAAABAAAD1420BA5D",
INIT_2B => X"A2FBE8BEFA2843DE00AA8015400FF84001EF0000020AA5D00154005D043FF455",
INIT_2C => X"FA2802ABEF557BEABEF5D0415410087FD74BAAAAEBFFEF557FC00AAF7AE95555",
INIT_2D => X"FFFFAABFEAAFF84001FF002A821FFAAD5554BA087FFFF55557BD54AAF7FBC01F",
INIT_2E => X"000FFFBE8BFF0800174AA557BFDE10A2FBEAB45F7D56AABA082A97545F7D16AB",
INIT_2F => X"FFEF552AB8E38087FC2092000000000000000000000000000000000000000000",
INIT_30 => X"070280024904AA1C0438FD7005150438F78A2DBFF0871F8FC7E3D56AB6DBEDB7",
INIT_31 => X"AA8ABAAADB400924920925EFF7D16ABFFE38E175EF1400000BA412E871FFE38E",
INIT_32 => X"0A1240055003FF6D5551420101C2EAFBD7A2FFEDB55B6A080038E3DB50555412",
INIT_33 => X"57FC00BAE3AA9257DA2FFE8BC7BE8E38E10A28017400E38A051FF0804050BA41",
INIT_34 => X"4971D0492E3F1C71C7BE8A2ABD74975EDBC7550E12410087FD74AAB6AABFFC75",
INIT_35 => X"A08249756DF7D168BC7F7AABAEAAF780051C70824851D7A2DB50482147FFAF55",
INIT_36 => X"00000000000000000000E3FFEFBD70000124AA557FFDE10A2FBEDB6DF7D16AAB",
INIT_37 => X"B55A2D16ABEFFFFBFDFFF552AAAAAA007BC00000000000000000000000000000",
INIT_38 => X"20AA002A955EFAAAA974AA0800020BA550028B550855400AAF7AEBDFEF08516A",
INIT_39 => X"000AAAAFBC0145002AA8AAAAAFFC20000000021EFF7D568BFFA2AA955FF5D040",
INIT_3A => X"E975EF0800174BA002E820105D003DFEF5D51420005D2ABFF45A2FBFFF55FF84",
INIT_3B => X"7BD74AAF7AEBDF455D7BC20BAAAAE821EFAAFBEAB55F7AAA8A00AA8417400AAA",
INIT_3C => X"2FFC00105D7BE8B55085142010AAD157545F7AEA8B5500557DF45552A8200000",
INIT_3D => X"A2FFFFFEFF7D568ABA0804155FFF7D568B55FFAAAAABAFF8415545000015555A",
INIT_3E => X"0000000000000000000000000000000000000AAFFFDF450804020AA557BFFE10",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024,               -- Port A enable input
WEA      => wbe_a_lo_1024(2),               -- Port A write enable input
DIA(0)   => data_write_a(16),        -- Port A data input
DOA(0)   => data_read_a_lo_1024(16),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024,               -- Port B enable input
WEB      => wbe_b_lo_1024(2),               -- Port B write enable input
DIB(0)   => data_write_b(16),        -- Port B data input
DOB(0)   => data_read_b_lo_1024(16),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_17_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"5284CE4FB7BD2C8994A13392DBD02E14006B82AC7E800D44D3DD2FD5F9B961C0",
INIT_01 => X"2EACD01F7E03FC6793F2199B39FC233C11D93AE6F3BB92B32091DBC339B24542",
INIT_02 => X"E63CCCC00A82C08092A2AFAE667033DB50853379C10BFDC5C6F4044443C817C6",
INIT_03 => X"7FF183635AEF9E3635AEF9E18E237040404446965C0607EE6DB7854AC4DE060C",
INIT_04 => X"D78AC33FB604488B000892EF17BE6D84196482236FE100294152E294350FB697",
INIT_05 => X"081B5F9B409420D0CDB47A05403F6CE0C08A4AB7F840EDB6F48100DFC8081081",
INIT_06 => X"768465354781CBC30316367077B4BDB50646E8D87100A8201ED01C19C020F71A",
INIT_07 => X"4002A110C922480A82D0841147162C48EBB9537A0022DC67987042EE976ABEA7",
INIT_08 => X"DB931BFEF91C00002CC0E019C0C82A4E4820C15A2330E004401891181168C4D1",
INIT_09 => X"09F3A1BC11EFBC66DB65307071477FF1030C397C060B4254064302042F803A69",
INIT_0A => X"3F330802162F3B7EE3F3EC7C7DEF207000F00059D2ED56D7EED2ED3C9A867DC0",
INIT_0B => X"185C44B91BC1740B7605040BE0018CFC7429F326B9E822FFC00074D5A0AB033A",
INIT_0C => X"00367A28FC1B7F7FEFFCFBFF3EFFCFBFF3EFFCFBFF3EFFCFBFF3EFFE7DFF9E00",
INIT_0D => X"0000000008004BA78428C7AD7FC94B533F5B4FFBD2FAD7FCCA786D43FE67C218",
INIT_0E => X"BA494CEBFD4F2667ABB6F68B29760593F33FA0CF170F40006001B1A05C000000",
INIT_0F => X"7F749299D7FAEB237DFE5865B6D2BF23265CBACE542A6FEE92333AFF33E0A9BF",
INIT_10 => X"F6C24B6D18C3C9F8E2881F3F787D776B5DB94A09955054DFDD246675FE7AC153",
INIT_11 => X"BFB349E08FF9A27EDE9FA8AEFD9E7467BFCB195CFEB56A1A70D34D1706FFFA3E",
INIT_12 => X"6FE219CA80725B875EED723FF7FCB2875EDAAFEAF7FD929BFD55BBC71D79F639",
INIT_13 => X"546670D018E7A6E581D7B6AB75FDFCECA6E581D7BB5DDFC6FF0EB7D7E859FDB5",
INIT_14 => X"B978177F6D6AF5ECDB5FB76A5F5FA165B456E0FB308710C49FCFB741598B9C7E",
INIT_15 => X"CFDAAB00AC00A8BBFC8B501CF7A0FED9A540EA1952586CEB54D143ACFF9A3BA9",
INIT_16 => X"000000000000000000000000000000000026E100002F382DBD9ECFE117805F20",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"4372003009EDCC4052E917114F981800C0000000000000000000000000000000",
INIT_1A => X"BA69A69AEBA69AEBA69A69AEBA69AEBA69A69A69A69A69A68698686981D75D74",
INIT_1B => X"6A351A8D46A351A8D068341A0D068341A0D068341A0D46A341A0D46A341A69AE",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000000000046A351A8D46A351A8D4",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"7FEAA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"17FFFF552EBFE00007FC00AA087FFFFFFFFFFFFFEFF7FBEAB450804001EFAAD5",
INIT_29 => X"D168A000004020AA5D7BE8B450051401EF087FD74AA087FFFFEFF7D168B55AAD",
INIT_2A => X"D7FEAB55FF80175EFFF8000010082A954BA00003DFEF085155400F78428BEFAA",
INIT_2B => X"F7D568BFFFF80175EF0004000BA552A821FF5D00020BA552A82000552A821555",
INIT_2C => X"AAAD1420BAFFFFFDF45AAD17FFFFAAFBC01EF5D0015555557BFDEBA5D2E975EF",
INIT_2D => X"BA007FEABEF005555555A2D1554BAA2FBE8B55A2AE80000F7D5555555D2AAAAB",
INIT_2E => X"0000000020AA5D00154005D043FF45555540000082EAABFF00516AA10552E820",
INIT_2F => X"8B550000071EFB6DF7AE92000000000000000000000000000000000000000000",
INIT_30 => X"F8FC7E3D56AB6DBEDB7FFEF552AB8E38087FC2092147FFFFFFFFFBFDFC7EBF5E",
INIT_31 => X"150438F78A2DBFFBED16AA381C0A07082497FEFB6D1451471EF007BD04920871",
INIT_32 => X"2A850105D2A80155417BEFB6DEB8E175FFE38E070280024904AA1C0438FD7005",
INIT_33 => X"D7BFAEBA4920925EFF7D16ABFFE38E175EF1400000BA412E871FF550A0009249",
INIT_34 => X"E3DB50555412AA8ABAAADB40092FFF5FFF6DAADF7FFD7B6F1C71EF55001756D5",
INIT_35 => X"7145B6AA28492487082007FEDBD700515556DA2DF50492A2FFEDB55B6A080038",
INIT_36 => X"000000000000000000000804050BA410A1240055003FF6D5551420101C2EAFBD",
INIT_37 => X"FEFF7FBFFF55A2D16AB550000175EFFFFBEAA000000000000000000000000000",
INIT_38 => X"55EF087FC200008516AB55A2D16ABEFFFFBFDFFF552AAAAAA007BC0000557FFD",
INIT_39 => X"020BA550028B550855400AAF7AEBDFEFF7D568AAA5D2A97410007BFFFFF55515",
INIT_3A => X"A955EF5D2E80010002A954005D2A82155087FFFFEFAAAA975EFAAAA974AA0800",
INIT_3B => X"D1575FF5504175EF5D7FEAAAA0000021EFF7D568BFFA2AA955FF5D04020AA002",
INIT_3C => X"2FBFFF55FF84000AAAAFBC0145002AA8AAAAAFFC2000FFD57DFFFAAFFFDF55FF",
INIT_3D => X"5D51420005D2ABFF45557FE8AAA000415410007BFFF450051555EFA2FBC0000A",
INIT_3E => X"00000000000000000000000000000000000000800174BA002E820105D003DFEF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024,               -- Port A enable input
WEA      => wbe_a_lo_1024(2),               -- Port A write enable input
DIA(0)   => data_write_a(17),        -- Port A data input
DOA(0)   => data_read_a_lo_1024(17),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024,               -- Port B enable input
WEB      => wbe_b_lo_1024(2),               -- Port B write enable input
DIB(0)   => data_write_b(17),        -- Port B data input
DOB(0)   => data_read_b_lo_1024(17),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_18_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"69844019080000A21A611406840014122A641074155FC28A2024001001801003",
INIT_01 => X"7443D920034004180005E9E3C90360C0041C0181002001602025800008440084",
INIT_02 => X"E2DCCCE61D5C008103F2000781FC0FEDEAC2161B0B8FB0008620044443006010",
INIT_03 => X"884E300802006900802006995C896D605200000856E24A040000640052141103",
INIT_04 => X"480520FC026125AC0025C9122644E3E40EC8E2001001302281841A009038A86A",
INIT_05 => X"432000040089983070019400F01010004C8DB841405A80A100B586200FAC24AE",
INIT_06 => X"09044359DC7040000000002C109B0E0A00A1104641C0803804000707284600E1",
INIT_07 => X"400D10100400481D5EB08501620000007500CE801241021FE78E404860140060",
INIT_08 => X"00880C0106A0528020019307CC082A0A4A6A01ED725021400040D028000A9729",
INIT_09 => X"00117063038000282081402E4106400B6186128040600C10C1C0200950508110",
INIT_0A => X"C0C30C2E21580C874004008080003C32A10A19090C02010E1022944061688000",
INIT_0B => X"0180A8062026000DC425C0301311324AA2373088479105D044A1022000001835",
INIT_0C => X"0D89844703649000000200000000000000000000000000000000000000000010",
INIT_0D => X"0D8306C182701404C1973010802020404084001E00010802046092B5001FB365",
INIT_0E => X"528EB314068AB8B803DB00002900800400FC503F08180050942E4200020C1B06",
INIT_0F => X"40A51D66280D6032C5F96D3C51555D5D7D5AA87285820814A3CCC501C2A60820",
INIT_10 => X"8B35A3FEBF1FEDFD9C2B30E0468AAAD5D48F37E8FC1304102947998A03984C10",
INIT_11 => X"440FE1DD772D37A0A321BC6968F32658BF2D4F2A80BF8FE3F9FE3AC362080529",
INIT_12 => X"5487910D7E5A6D961A28456A1832E5161A100DD5182BC54020EA67A189C6ED36",
INIT_13 => X"AA444CAF91EDD1B725868403BE06323551B725868A100ABD119753B70964122B",
INIT_14 => X"EDC259048ACD868EE3803D65CEDC258A8F80D55E007C3F8EBB56F4C5362C978F",
INIT_15 => X"3F240014BE84370001B6922070440556B15F7FABBC0031BCF2257C41634B14D4",
INIT_16 => X"C1B06C1B06C1B06C1B06C1B06C1B06C1B0491069068000004060300A005A0118",
INIT_17 => X"1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06",
INIT_18 => X"B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C",
INIT_19 => X"B28BBECEB80EE173C2300F7DF16000000000000000000000000041B06C1B06C1",
INIT_1A => X"8A28A28AAAAAAA28A28A28AAAAAAA28A28A28A28A28A28A2910591505C104104",
INIT_1B => X"28944A25128944A25128944A25128944A25128944A2552A954AA5128944AAAA2",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000128944A25128944A251",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"9540000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"BEAB450804001EFAAD57FEAA087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974BA082E",
INIT_29 => X"7FFFFFFFFFBFDF45AAD568B55080028B55002E82000087FFFFFFFFFFFFFEFF7F",
INIT_2A => X"0043DE10AA843DE00087FFFFEFF7D168B55AAD17FFFF552EBFE00007FC00AA08",
INIT_2B => X"0004020AA5D7BE8B450051401EF087FD74AAAAFFFDF45A2D16AB55F7FFFFFFF0",
INIT_2C => X"0F78428BEFAA80000000804154BA55042ABEF5D7FD75FFAAD540145AAD168A00",
INIT_2D => X"00082E95555085168A10557FD7545FF8000010082A954BA00003DFEF08515540",
INIT_2E => X"0005D00020BA552A82000552A821555D7FEAB55FF80175EF5D00020105D2A974",
INIT_2F => X"DFFF5D2A954AA082A92428000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFBFDFC7EBF5E8B550000071EFB6DF7AE921C7FFFFFFFFFFFFFFFF7FBF",
INIT_31 => X"AB8E38087FC2092087FFDFC7E3F1FAF55A2DF6DB7D1C002AB7D002A82028147F",
INIT_32 => X"DF6DB7DE3F5FAFC708003DE28B68E38E280871F8FC7E3D56AB6DBEDB7FFEF552",
INIT_33 => X"ADF4516DBED16AA381C0A07082497FEFB6D1451471EF007BD0492B6F1F8F55AA",
INIT_34 => X"1C0438FD7005150438F78A2DBFFA28407038140410492550A2ABC7497BD25FFA",
INIT_35 => X"F5D0E05000492097428002E9557D1C516FA28417BD5545E38E070280024904AA",
INIT_36 => X"00000000000000000000550A00092492A850105D2A80155417BEFB6DEB8E175F",
INIT_37 => X"FFFFFFFFDFEFF7FBFFFEF552E974AA082A820AA0000000000000000000000000",
INIT_38 => X"ABEF002A800AA557FFDFEFF7FBFFF55A2D16AB550000175EFFFFBEAA00557FFF",
INIT_39 => X"6ABEFFFFBFDFFF552AAAAAA007BC0000087BFDF45AAD568B55AAFBFDFEF55042",
INIT_3A => X"FC2000FFD56AB45A2FFFDFFFAAD16AB4500043DEAAFFAEAAAAA08516AB55A2D1",
INIT_3B => X"2AA8B45087FC01EFA2FFD55EFF7D568AAA5D2A97410007BFFFFF5551555EF087",
INIT_3C => X"AAA974AA0800020BA550028B550855400AAF7AEBDFEFA280154BA55040000055",
INIT_3D => X"087FFFFEFAAAA975EF5D2E974000804154BA082A975EF5D517DEAA007BD5545A",
INIT_3E => X"00000000000000000000000000000000000005D2E80010002A954005D2A82155",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024,               -- Port A enable input
WEA      => wbe_a_lo_1024(2),               -- Port A write enable input
DIA(0)   => data_write_a(18),        -- Port A data input
DOA(0)   => data_read_a_lo_1024(18),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024,               -- Port B enable input
WEB      => wbe_b_lo_1024(2),               -- Port B write enable input
DIB(0)   => data_write_b(18),        -- Port B data input
DOB(0)   => data_read_b_lo_1024(18),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_19_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"042200000000000041088001001AA00000000000000000000000500802000003",
INIT_01 => X"040048000024000000000404000000000A22000800000800004A200000000001",
INIT_02 => X"200C8840085EB00480060000001C008002489E0F000405EA0004040404000000",
INIT_03 => X"24004000000000000000000900002C4050000000000069500208400002E14100",
INIT_04 => X"4800200C0000000044002000C80020E40000E200000130200188000000800100",
INIT_05 => X"000000000080181000000000701000004C8000000058800000B1000009880480",
INIT_06 => X"80500081081040000000002C100040400000004641C080380400070100000000",
INIT_07 => X"4020109801A4CE005C00048380142810010564C4100114012002402028044808",
INIT_08 => X"0070700000000000000083004C3902420062000020E0000100004082A140102B",
INIT_09 => X"001150200000000000000026400000016186100000000010C04002C000000000",
INIT_0A => X"007C00008082C0002000000000002C3000000004050001030102040000000000",
INIT_0B => X"0000000000000000000000000000010000800011000000000000000000000BC0",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"000000000000000000000000000000042000760000000000000000010004B200",
INIT_0E => X"0D74002280300F0002FB069040000060000C5003000800000000000000000000",
INIT_0F => X"C01AE8004500744C780687DBA828008080A5FC0D385598035D0008A00C015660",
INIT_10 => X"39D8140040201BF861F0E7D693E6170022408116DFE0AB3006BA0011401D02AC",
INIT_11 => X"5412E4997F5249FD005043B8680CC98F00D0F2DD0140100406FE053A98F6ECC7",
INIT_12 => X"7418663001858040E153888000010840E165D0000000285C246A181C03FE4662",
INIT_13 => X"8199830066F0020858385974000001260208583854E2200000660208D6B1423F",
INIT_14 => X"8235AC508FCE8811042040F008235AE04420C040CF00C031C80009B8F224978B",
INIT_15 => X"030004E00000C220010808C10D9A92A74CD7CF4A09051110AD5A3C9200B7F280",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000118",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"07208BBA3F0C7010C660C7441920000000000000000000000000000000000000",
INIT_1A => X"861869A61861861861869A61861861861861861861861861A8208C4C1534D34C",
INIT_1B => X"984C26130984C26130984C26130984C26130984D26930984C26130984C261861",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000984C26130984C26130",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"174BA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFDFEF5D2A974BA082E95400F7FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0004",
INIT_29 => X"FFFFFFFFFFFFFFFFF7FBFDFFF552E974BAA2FFFFE10087FFFFFFFFFFFFFFFFFF",
INIT_2A => X"004001EFAAAEA8ABA087FFFFFFFFFFFFFEFF7FBEAB450804001EFAAD57FEAAF7",
INIT_2B => X"FFFBFDF45AAD568B55080028B55002E82000F7FFFFFFFFFFFFDFEFA2D568B550",
INIT_2C => X"0007FC00AAF7FFFFFFFF7FBE8B55AAD16ABEF5D2ABFF55080402010087FFFFFF",
INIT_2D => X"55A2FFFDFEF5D2EBFE00AAFFFFEBA087FFFFEFF7D168B55AAD17FFFF552EBFE0",
INIT_2E => X"000AAFFFDF45A2D16AB55F7FFFFFFF00043DE10AA843DE00557FFDFEFA2D16AB",
INIT_2F => X"FFEF552A974AA0000104AA000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFF7FBFDFFF5D2A954AA082A92428E3FFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"0071EFB6DF7AE92EBFFFFFFFFFFFFDFEFF7F5FAFC7492A974AAB6F5F8E101C7F",
INIT_32 => X"F1F8FD7AAD16AB450000001FFBEA4A8AAA147FFFFFFFFFBFDFC7EBF5E8B55000",
INIT_33 => X"00000010087FFDFC7E3F1FAF55A2DF6DB7D1C002AB7D002A82028FFFFFFFEFF7",
INIT_34 => X"BEDB7FFEF552AB8E38087FC2092F7FBF8FC7E3F5EAB45B6DF6FBEF5D2AB8F7D0",
INIT_35 => X"84971F8FC7AAD56DB6DBEF5F8FD7412ABFE28B6F5F8E820871F8FC7E3D56AB6D",
INIT_36 => X"00000000000000000000B6F1F8F55AADF6DB7DE3F5FAFC708003DE28B68E38E2",
INIT_37 => X"FFFFFFFFFFFFFFFFFDFEF552E954AA0004000AA0000000000000000000000000",
INIT_38 => X"54AAF7D568A00557FFFFFFFFFFFDFEFF7FBFFFEF552E974AA082A820AAA2FFFF",
INIT_39 => X"FFF55A2D16AB550000175EFFFFBEAA00A2FFFFFFFF7FBFDFFFFFD568B55002A9",
INIT_3A => X"A800AAF7FBFDFEFF7D56AB45AAD56AB450004001EFFF842AAAA557FFDFEFF7FB",
INIT_3B => X"FFFFFFF552AA8BEF080402000087BFDF45AAD568B55AAFBFDFEF55042ABEF002",
INIT_3C => X"8516AB55A2D16ABEFFFFBFDFFF552AAAAAA007BC0000FFFBE8B55AAD168B55F7",
INIT_3D => X"00043DEAAFFAEAAAAA08556AB55A2D57FFFFF7D568B45002ABDEAAFFD16AA000",
INIT_3E => X"0000000000000000000000000000000000000FFD56AB45A2FFFDFFFAAD16AB45",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024,               -- Port A enable input
WEA      => wbe_a_lo_1024(2),               -- Port A write enable input
DIA(0)   => data_write_a(19),        -- Port A data input
DOA(0)   => data_read_a_lo_1024(19),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024,               -- Port B enable input
WEB      => wbe_b_lo_1024(2),               -- Port B write enable input
DIB(0)   => data_write_b(19),        -- Port B data input
DOB(0)   => data_read_b_lo_1024(19),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_20_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000003",
INIT_01 => X"F55FF80000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"E05022020800008400F655001FFCFF80018FA804400000000000004400000001",
INIT_03 => X"00000000000000000000000900002CC07000000000000000000000000000013F",
INIT_04 => X"68002FFE40900010000180000001FFEC0012EE0C001370F40780000000000000",
INIT_05 => X"0840000880FCBBF0100E204DF0F88311DD8005080679800000F3000029980580",
INIT_06 => X"001000030817C8E8840155FDF9001001050023F6C3C3D0F87FA19F7F011000E4",
INIT_07 => X"000000090492260800008000EE00000000000000002101FF2002C00000004018",
INIT_08 => X"2A040001071004000013FF7FCA302C0C0008214800002101554031F800000000",
INIT_09 => X"801F57F200000090000489FEC0000001EFBEF0040008023FDFC0000000004006",
INIT_0A => X"0000000008000000000000000000ADF000000200000008000008028300110230",
INIT_0B => X"0000000000000800080000000000000000000000000000000800800A40000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"000000040900005C848538000020000000800000080000020000800101FFB600",
INIT_0E => X"00800000003A010003000000000000600FFC53FF001800000002004080000000",
INIT_0F => X"0001000000007408040000004000000004E9000008020000200000000E800800",
INIT_10 => X"00200000000313100010002000008000000000129600040000400000001D0010",
INIT_11 => X"81C012060000000000218F7840000100800004000000000066C0000080080000",
INIT_12 => X"800000000017C000100000000001A800080000000001A8040000002840008185",
INIT_13 => X"0000000006F00000100200000000012600001004000000000066000000801040",
INIT_14 => X"0000200410100000000005F00000020080090A0000000085C800002000586000",
INIT_15 => X"FF00400000000000020020020001000040283024E4F2860400008000030ED080",
INIT_16 => X"00000000000000000000000000000004010201001003020200000000000127DB",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"A0700030038200010089120104D2040020000000000000000000000000000000",
INIT_1A => X"2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2C30C30C30C30C306982121A1E79E79",
INIT_1B => X"32190C86432190C86432190C86432190C86432190C86432190C86432190CB2CB",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000432190C86432190C864",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0201000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF552A974AA0004174BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA0804",
INIT_29 => X"7FFFFFFFFFFFFFFFFFFFFFFEF552E954AA000400000F7FFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E954BA007FC00BA087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974BA082E9540000",
INIT_2B => X"FFFFFFFFFF7FBFDFFF552E974BAA2FFFFE10FFFFFFFFFFFFFFFFFFFFFBFDFFF5",
INIT_2C => X"FAAD57FEAA007FFFFFFFFFFFFFEFF7FBFFF550800020BAAAD56AAAAF7FFFFFFF",
INIT_2D => X"EFF7D56AB450000021EFA2D57DE10087FFFFFFFFFFFFFEFF7FBEAB450804001E",
INIT_2E => X"000F7FFFFFFFFFFFFDFEFA2D568B550004001EFAAAEA8ABA5D7FFFFFFFFFFFDF",
INIT_2F => X"FFFF5D2E954AA080005000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFEF552A974AA0000104AAFFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"A954AA082A92428087FFFFFFFFFFFFFFFFFFBFDFEF5D2E974AA000A07000E3FF",
INIT_32 => X"FFFFFEFF7FBFFFFF552E974AA0071C50BA1C7FFFFFFFFFFFFFFFF7FBFDFFF5D2",
INIT_33 => X"EDF6FABAEBFFFFFFFFFFFFDFEFF7F5FAFC7492A974AAB6F5F8E10E3FFFFFFFFF",
INIT_34 => X"EBF5E8B550000071EFB6DF7AE921C7FFFFFFFFFBFDFEFE3F5F8F450004050AAB",
INIT_35 => X"A497FFFFFFF7FBF8FC7EBD168B450804021FFB6D57DE28147FFFFFFFFFBFDFC7",
INIT_36 => X"00000000000000000000FFFFFFFEFF7F1F8FD7AAD16AB450000001FFBEA4A8AA",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2A954AA0800174100000000000000000000000000",
INIT_38 => X"74AA002E95410A2FFFFFFFFFFFFFFFFFFFFFDFEF552E954AA0004000AAFFFFFF",
INIT_39 => X"FDFEFF7FBFFFEF552E974AA082A820AA087FFFFFFFFFFFFFEFF7FBFDFFF5D2A9",
INIT_3A => X"568A00AAFFFFFFFFFFBFDFEFFFFFFDFEF5D2E954AA0051554BA557FFFFFFFFFF",
INIT_3B => X"D16AB450804174AAFFFFFFEBAA2FFFFFFFF7FBFDFFFFFD568B55002A954AAF7D",
INIT_3C => X"57FFDFEFF7FBFFF55A2D16AB550000175EFFFFBEAA005D7FFFFEFF7FBFDFFFAA",
INIT_3D => X"0004001EFFF842AAAA087BFDFEFF7FFEAB45A2D568B550804001EFF7D57DEBA5",
INIT_3E => X"0000000000000000000000000000000000000F7FBFDFEFF7D56AB45AAD56AB45",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024,               -- Port A enable input
WEA      => wbe_a_lo_1024(2),               -- Port A write enable input
DIA(0)   => data_write_a(20),        -- Port A data input
DOA(0)   => data_read_a_lo_1024(20),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024,               -- Port B enable input
WEB      => wbe_b_lo_1024(2),               -- Port B write enable input
DIB(0)   => data_write_b(20),        -- Port B data input
DOB(0)   => data_read_b_lo_1024(20),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_21_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"4A302428B824900A128C090A5C1800261500213C005FE812D10420054085A202",
INIT_01 => X"001FFE3440B609703B0427F801A40B8115BC4F655300340288A40D30040E4DD8",
INIT_02 => X"E00424256888D8819801000F9FFFFFFFF149FF1FCA448046C60A0D2437C517F9",
INIT_03 => X"20030640003250640003250F06002CC1740002019824E001CD357832440001FF",
INIT_04 => X"EA2C3FFD400006E04401A8837001FFFC004AEF00080B70E08FB5789421007C5C",
INIT_05 => X"00011A0C40F9FFF80920954FF0F00809DF84A0202879800000F3000029980780",
INIT_06 => X"0805984B7A1FC0A0000101FFF0480080002281F7C3C381F87C03DFFF00009004",
INIT_07 => X"B424068086A205481A60A19000908204A855B000A08A61FF20C3D004D331D340",
INIT_08 => X"1BFA0001600802000023F7FFC08D234B40C2028253000040114200000D0226C0",
INIT_09 => X"EF1F5FF054096C6ADBA169FFC202B1C1FFBEF0440021083DFFCE22DC2880E24D",
INIT_0A => X"45FF0C004041D84862A28C54518DBFF00020004C0A6044901112A0908AA0A300",
INIT_0B => X"018C241102068006C620C03882019480E63180855A492712CC01C49C20201BFE",
INIT_0C => X"08A9464116544302C02D92236488D92236488D92236488D922366446C911B210",
INIT_0D => X"08800444021048034004001890000806002804A0822189000900D80621FFBE00",
INIT_0E => X"060580261013813A2CC396506102C4053FFD5BFF00A04A00200602CA52001100",
INIT_0F => X"080C0B004C202621A85C09411500135844C196D3606941018150098404C1A304",
INIT_10 => X"B02901013416181C96C2C9C600890A2028172192C460D1820302A0130809834A",
INIT_11 => X"9C5E803408250180AC268D185DB3F4350B811068C00049A0A4AA68F05C96A001",
INIT_12 => X"002C006560138F032B1804101244C883052208209040CC849063A747512B7678",
INIT_13 => X"41401E240665750440C9488280254530314080C2C601040420352148A00501B1",
INIT_14 => X"500811204D000700114204A70422016149916011008CAA8858850B00C32591C0",
INIT_15 => X"FFC06E60AC0496022300233104663040808E991765205000070121D41D18D098",
INIT_16 => X"40100401004010040100401004010040102090010008000001C0E010020007DF",
INIT_17 => X"0100401004010040100401004010040100401004010040100401004010040100",
INIT_18 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_19 => X"FFEF9FEEFF7FFDF7FF3E3DFDF7E0000000000000000000000000401004010040",
INIT_1A => X"BEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBFFDFDFFFCF3CF3F",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFEFF7FBFDFEFF7FBFDFEFBEF",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000FFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0001000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E954AA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0004",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA0004154BAFFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"52E974BA0804000AAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0004174BAFF",
INIT_2B => X"FFFFFFFFFFFFFFFFEF552E954AA000400000007FFFFFFFFFFFFFFFFFFFFFFEF5",
INIT_2C => X"A082E95400007FFFFFFFFFFFFFFFFFFFFDFEF5D2E974BA002E97400007FFFFFF",
INIT_2D => X"FFFFFBFDFEF5D2A954AA002E974BA087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFBFDFFF5D2E954BA007FC00BA5D7FFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA000002000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080005000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"A974AA0000104AAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974BA0000174AAFFFF",
INIT_32 => X"FFFFFFFFFFFFDFEF552E954BA080A000AAE3FFFFFFFFFFFFFFFFFFFFFFFEF552",
INIT_33 => X"02A95400087FFFFFFFFFFFFFFFFFFBFDFEF5D2E974AA000A07000007FFFFFFFF",
INIT_34 => X"F7FBFDFFF5D2A954AA082A924281C7FFFFFFFFFFFFFFFFFFBFDFEF5D2A974BA0",
INIT_35 => X"A557FFFFFFFFFFFFFFFF7FBFDFFF552E974BA0020924BA1C7FFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000E3FFFFFFFFFFFFFFEFF7FBFFFFF552E974AA0071C50B",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0000020000000000000000000000000000",
INIT_38 => X"74BA0000174BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954AA080017410FFFFFF",
INIT_39 => X"FFFFFFFFFFDFEF552E954AA0004000AAF7FFFFFFFFFFFFFFFFFFFFFFFEF552A9",
INIT_3A => X"E95410087FFFFFFFFFFFFFFFF7FBFDFEF5D2A954BA082E800AAA2FFFFFFFFFFF",
INIT_3B => X"FBFFFFF552E954BA002E97410087FFFFFFFFFFFFFEFF7FBFDFFF5D2A974AA002",
INIT_3C => X"57FFFFFFFFFFFDFEFF7FBFFFEF552E974AA082A820AA557FFFFFFFFFFFFFEFF7",
INIT_3D => X"5D2E954AA0051554BA5D7FFFFFFFFFBFDFEFF7FFFFFEF5D2A974BA0000020AA5",
INIT_3E => X"0000000000000000000000000000000000000AAFFFFFFFFFFBFDFEFFFFFFDFEF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024,               -- Port A enable input
WEA      => wbe_a_lo_1024(2),               -- Port A write enable input
DIA(0)   => data_write_a(21),        -- Port A data input
DOA(0)   => data_read_a_lo_1024(21),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024,               -- Port B enable input
WEB      => wbe_b_lo_1024(2),               -- Port B write enable input
DIB(0)   => data_write_b(21),        -- Port B data input
DOB(0)   => data_read_b_lo_1024(21),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_22_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"5290F4CDE914905A14A43D33F488243E17122300F55FEB189B343A1140548380",
INIT_01 => X"A54007B259F6A975386262000C344BA9573C6FF57B18A5FB0ABFCD3C2C5F4F0C",
INIT_02 => X"021DFF8C38B3C009D203551040030071869D0040180AA2DC53DB89BEA8204001",
INIT_03 => X"2603475A969D0475A969D0460EAA401005111011BD506954EDB40F5EF41434C0",
INIT_04 => X"922D9002100ED69E443D988B0D5400103E48003D0800011E803B06B5B9125A15",
INIT_05 => X"281B5A0C06000408F4DF9422010D8802022F2124A8022492580040440002021C",
INIT_06 => X"F780C4C052881ADA0E05440205DA50930FA182010004700083E220800440B588",
INIT_07 => X"049D028B93FB561833D8094A02F5EA92FD7247E10305C40040D136E6A023F7FC",
INIT_08 => X"00028241680A0E002A9400803A884B5B5206B7C2E53CA25144009007A64EBD64",
INIT_09 => X"41008810240240C6694008010392354010000560141801002028A83D2A08E06D",
INIT_0A => X"34000000848BCA6902A29C54539C020E11810098D4067EFF9FF284D483E2AB41",
INIT_0B => X"500001840000C80B410014088040F4A944B1AA313C0022AA0011C0DC00028001",
INIT_0C => X"80B14004D158C8CA24A1C2A870AA1C2A870AA1C2A870AA1C2A872550E1543800",
INIT_0D => X"80A14050A01509E050854498B5281A1C34E506A2C6898B52A154DAC6B6000850",
INIT_0E => X"0B03001A483A4146603050080410089180008800143D83888281A2034A850142",
INIT_0F => X"A4160600349075238473F1210006133835E92273612B3482C090068A0E84AC56",
INIT_10 => X"30060181BA1B13959DC08DA902458870201970B29602562B0581200D141D0959",
INIT_11 => X"E042021C040D0152C8058B3840F044708E7E1C20A0106EA166C13AFC14AA3804",
INIT_12 => X"080E004B0C17C1439A9838301DC1A8438EA32C009DC1A8255300650458A1D588",
INIT_13 => X"018010E186F110A908E3A8CB0026C9A610A908E6A60F0807626610E160589C4C",
INIT_14 => X"2A701667334005800B1605F043858125E0D04110408D2485CA034681E43A1E40",
INIT_15 => X"00646002304244A91102C93A2D608D2A258DF8034188200C050171A41108F084",
INIT_16 => X"110441104411044110441104411044110466C440446CA06951D4EA8010009804",
INIT_17 => X"0040100401004411044110441104411044110441104411044110441104411044",
INIT_18 => X"0401004010040100401004010040100401004010040100401004010040100401",
INIT_19 => X"F7DFBFDEFE8FF1F7DEBDDF7DF7D05122890000000003FFFFFFFF900401004010",
INIT_1A => X"9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7BFFDFD7DDDF7DF7D",
INIT_1B => X"F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE79E7",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000003F9FCFE7F3F9FCFE7F3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA000400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0800",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000002000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2A954BA000015400FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080402010FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2A954BA0004154BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A0004174BAFFFFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0800154AAFFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF552A974AA0000174BAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974A",
INIT_2E => X"000007FFFFFFFFFFFFFFFFFFFFFFEF552E974BA0804000AAA2FFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080400010000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E954AA080005000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000402010FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2A954BA000417410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"804154BAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974BA0000174AAFFFFFFFFFFF",
INIT_34 => X"FFFFFFFEF552A974AA0000104AAE3FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0",
INIT_35 => X"AA2FFFFFFFFFFFFFFFFFFFFFFFEF552E954BA000E124BAE3FFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000007FFFFFFFFFFFFFFFFFFFFDFEF552E954BA080A000A",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804000100000000000000000000000000",
INIT_38 => X"54AA000400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2A954AA080017410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"0174BAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A954BA000415400FFFFFFFFFFFFF",
INIT_3B => X"FFFDFEF552E974AA0804174AAF7FFFFFFFFFFFFFFFFFFFFFFFEF552A974BA000",
INIT_3C => X"2FFFFFFFFFFFFFFFFFFFFFDFEF552E954AA0004000AAA2FFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2A954BA082E800AAAAFFFFFFFFFFFFFFFFFFFBFDFEF5D2E954BA002A820BAA",
INIT_3E => X"0000000000000000000000000000000000000087FFFFFFFFFFFFFFFF7FBFDFEF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024,               -- Port A enable input
WEA      => wbe_a_lo_1024(2),               -- Port A write enable input
DIA(0)   => data_write_a(22),        -- Port A data input
DOA(0)   => data_read_a_lo_1024(22),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024,               -- Port B enable input
WEB      => wbe_b_lo_1024(2),               -- Port B write enable input
DIB(0)   => data_write_b(22),        -- Port B data input
DOB(0)   => data_read_b_lo_1024(22),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_23_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"EF20906D902424807BC8241BC81801B97D38AD3C0800103362A6741C80A12A02",
INIT_01 => X"001FFF8409F089003B4422000D80C80106804A7951C5B9D1C828043EA28838F9",
INIT_02 => X"E01CEE21649C82C40800000F9FFEFF8E72CA7F5FC2E22809925A0D3611C877F8",
INIT_03 => X"24000400402670400402670D48222DC1764446838624000080007460C40001BF",
INIT_04 => X"68403FFC020560E0443E21037C01FFFC0002EE00628BF0E02FAD781014085014",
INIT_05 => X"0112000202FBFFF00920017FF0F0628BFF8488890979800002F702002BB807A0",
INIT_06 => X"EF85788B681FC000000001FFF0010000000001F7CBC385F87C0BFFFF20040001",
INIT_07 => X"F6E200000000C1440E3AE408009120071070FA07A1CB23FFA403F0C4D23BF7C0",
INIT_08 => X"0BF87CA400804000003FF7FFD8880A034AC09662305AB10555421006891A1089",
INIT_09 => X"BE1F5FEA10092C0896A243FFC0008087FFBEF2000000001DFFC612C0C0400100",
INIT_0A => X"41FF0C2060501000600000000001BFFA800808189A657EF81DD0C00079CC8001",
INIT_0B => X"018C24110A860006C620C0312241C482B20400CC52492710CC80060020A81BFE",
INIT_0C => X"0C08866907048320C20C10030400C10030400C10030400C10030400608018210",
INIT_0D => X"040002000041500300100040000500C000801000C02400000952800001FFBF04",
INIT_0E => X"FC850015385380380CDB86106502C5043FFD5FFF00A04BC010A7724B10000800",
INIT_0F => X"89F90A002A70A710A51C01C05904014861433602A1CAF13F2110055614C72FC0",
INIT_10 => X"E02D02001C1E14981B43253EE50C8220180F1082E06397E07E42200AAC298E57",
INIT_11 => X"8421802400A90022B0070FAE18019214A380344920080B21A58B02AC60BACDF0",
INIT_12 => X"0A2A000C480B0704B54028101AC49C84BB4100009AC49C80857A82D20CE8CB22",
INIT_13 => X"01E00C8103416445C12ED0400027C5292445C12D500B0005A62D344CB241D095",
INIT_14 => X"132C907425604680038706A35132C94BDD011010404428886AC91B11311C8280",
INIT_15 => X"FF000470BE0692020328CA0028042054A92771C50FC070110001C1680809591D",
INIT_16 => X"00802008020080200802008020080200800800200200000000000008004807DF",
INIT_17 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_18 => X"8020080200802008020080200802008020080200802008020080200802008020",
INIT_19 => X"0000000000000000000000000000000000000000000000000000008020080200",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080002010FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974AA000400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000400010FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974AA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080000010FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E954AA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954A",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA000015400FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080002010FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974AA000400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000402010FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E954AA080005000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA080407000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA00041741",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080000010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000402010FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2A954AA080002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954AA080017410FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"552A954BA000415400F7FFFFFFFFFFFFFFFFFFFFFFFFF552A954BA080015410F",
INIT_3E => X"0000000000000000000000000000000000000F7FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024,               -- Port A enable input
WEA      => wbe_a_lo_1024(2),               -- Port A write enable input
DIA(0)   => data_write_a(23),        -- Port A data input
DOA(0)   => data_read_a_lo_1024(23),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024,               -- Port B enable input
WEB      => wbe_b_lo_1024(2),               -- Port B write enable input
DIB(0)   => data_write_b(23),        -- Port B data input
DOB(0)   => data_read_b_lo_1024(23),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_24_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100600007FFF000080108004000800020000840041000080808",
INIT_02 => X"FC5CA803400EB8209000000F9FFEFF8E7240FF1FC22409EA04018E50074017F0",
INIT_03 => X"11100400000000400000000D00002CC07400000090C080019001010A000001BF",
INIT_04 => X"68003FFC00040000000000008001FFFC0002EE00000370E007A100000000E468",
INIT_05 => X"0000000000F8BFF00920004DF0F00001DF8000000079800000F3000029980780",
INIT_06 => X"6E461803081FC000000001FFF0000000000001F7C3C380F87C019FFF00000000",
INIT_07 => X"600C2400013649609C8000980040814210254000A00B21FF2003F2A80D500000",
INIT_08 => X"0BF80000000000000003F7FFD88D2B4A02C0940062EC2804001610020408178B",
INIT_09 => X"8E1F5FE010092C0892A041FFC0000001FFBEF0000000001DFFC002C000000000",
INIT_0A => X"41FF0C0000000000600000000001BFFA0000005501AA00000CE2000009400000",
INIT_0B => X"018C0411020600048620C030020502000200000400490510CC00040020201BF4",
INIT_0C => X"0808064106040300C00C10030400C10030400C10030400C10030400608018210",
INIT_0D => X"0000000000004003000000000000001200580000000000000000000001FFBE00",
INIT_0E => X"0086C022005381380FDB96516140C6043FFD5BFF000041000000004110000000",
INIT_0F => X"80010D804400A7240C840C201D0210840043B4804012500021E0088014C04940",
INIT_10 => X"4109038041021C980200D06410C1924030008142E06024A00043C01100298092",
INIT_11 => X"587CC200002100C14428090A1D02348190814C09C010104025AA40041A0D8005",
INIT_12 => X"022E0030300B0E46177004208000D8C61D7004300000D884817B00011306B2D9",
INIT_13 => X"01E003060344710009875C018100013831000985DC000C20003C310006143B70",
INIT_14 => X"4001850EDC004780144806A64400186CBF8961104000C3807884000846EB9500",
INIT_15 => X"FF0006E08C063C0220002201490418082010A57263E0100008000290161E711C",
INIT_16 => X"00000000000000000000000000000000000000000000000000000000000007DF",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"F2D0AEEAF6E7CC1132CDB4441990000000000000000000000000000000000000",
INIT_1A => X"BEFBE79E79E79E79E79EFBEFBEFBEFBEFBEF9EF9EF9EF9EFA69861219575D75F",
INIT_1B => X"783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1EFBEF",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000783C1E0F0783C1E0F0",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0201000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A000400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA000400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000400000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402010000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"00002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080002010FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000400010FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA00040000",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020100000000000000000000000000",
INIT_38 => X"74BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"000010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA000002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974AA000402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000002010F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024,               -- Port A enable input
WEA      => wbe_a_lo_1024(3),               -- Port A write enable input
DIA(0)   => data_write_a(24),        -- Port A data input
DOA(0)   => data_read_a_lo_1024(24),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024,               -- Port B enable input
WEB      => wbe_b_lo_1024(3),               -- Port B write enable input
DIB(0)   => data_write_b(24),        -- Port B data input
DOB(0)   => data_read_b_lo_1024(24),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_25_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100200002000000080100004000000020000800041000080808",
INIT_02 => X"FC400086000000800000000F9FFEFF8E738FFF1FC204010000000111568DD7F8",
INIT_03 => X"00000400000000400000000D00002CC4740000008000000080000000000001BF",
INIT_04 => X"68003FFF64A564AC000000000001FFFE0082EF00010370E007A1000000004000",
INIT_05 => X"0A00040148F8BFF80920804DF0F00101DFC040000079C92484F30499299837C1",
INIT_06 => X"66041803081FC0E0801101FFFD000E41002299F7E3C380F87C019FFF81200096",
INIT_07 => X"000000080480AE00000080000000000000000000A00B21FF2003E00000000000",
INIT_08 => X"1BF80000400A02000003F7FFFA0008000200A0400008A0000014100200081000",
INIT_09 => X"8E1F5FFA53EFBCACB2E369FFE0010001FFBEF80C40630C7DFFEEBAF000800202",
INIT_0A => X"41FF0C0600000000600000000001BFFE00301000000000000CC020000140000C",
INIT_0B => X"01DCCC31222730A49620C030020100000200000400490D10EC00040220201BF4",
INIT_0C => X"0808064106240300C00C10030400C10030400C10030400C10030400608018210",
INIT_0D => X"0883044582114013412080000000000000000000000000000012800001FFBE00",
INIT_0E => X"00040020000180380FC386106140C6043FFD5BFF00A04B80608003CB120C1106",
INIT_0F => X"0000080040000200040400000100000000009480000240000100080000400900",
INIT_10 => X"0001000000000808000000240000020000000100006004800002001000008012",
INIT_11 => X"0001001808220000002004001900000080800008000000000022400000088000",
INIT_12 => X"0010000000000E00110000000000408009000000000040808063004000008200",
INIT_13 => X"6000000000046100000240000000001021000004400000000010210000001010",
INIT_14 => X"4000000404000800000000060400000088000001800000001084000000088000",
INIT_15 => X"FF800C608C041002000002000006100000002100000000180600000000100018",
INIT_16 => X"4110441104411044110441104411044510629041040D180400000010028047DF",
INIT_17 => X"1104411044110441104411044110441104411044110441104411044110441104",
INIT_18 => X"1044110441104411044110441104411044110441104411044110441104411044",
INIT_19 => X"FBA2894A196A8C5A2932EC15DA080800002FFFFFFFFFFFFFFFFFC11044110441",
INIT_1A => X"2492492492492492492410410410410410410492410492412000531215A69A6B",
INIT_1B => X"158AC562B158AC562B158AC562B158AC562B1588C46231188C46231188C49249",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000B158AC562B158AC562B",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080000010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000010FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08000000",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024,               -- Port A enable input
WEA      => wbe_a_lo_1024(3),               -- Port A write enable input
DIA(0)   => data_write_a(25),        -- Port A data input
DOA(0)   => data_read_a_lo_1024(25),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024,               -- Port B enable input
WEB      => wbe_b_lo_1024(3),               -- Port B write enable input
DIB(0)   => data_write_b(25),        -- Port B data input
DOB(0)   => data_read_b_lo_1024(25),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_26_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"E9264EAB20190CA3BA4997AA9002AE9C001006B0778015CFA17E0811039879C7",
INIT_01 => X"2FFFF9BB1F773C7F9BB07DFFFDD863FC5FFF3FEFFBBF9FFB22FFFBC7B9F30686",
INIT_02 => X"E06CCC62052E708180F6FFBFFFFCFFFFF9C7FF7FC24332E642090000074037F6",
INIT_03 => X"428003739CD9863739CD9869FE2B7DEAF300029E4E300DFE69A6E644E6FF473F",
INIT_04 => X"7C2FEFFFF5BA124F003DD31EAFFFFFEE9FF7EE6F4C0770FFD7DC7CA53997B2B1",
INIT_05 => X"DFFB5421C1F8BBFAFDBFFACDF0FFCC05DDDBFF3690F9EDB7F5F7AFF639BD7DE3",
INIT_06 => X"EFD044ABC817C3E3A74667FDFFB6FF5727CC3BFEF7C3FAF87FF59F7FFBFEF69F",
INIT_07 => X"00003002132462052E708180EF060C18E5BEFB051225CDFF7002C4EEDE77F6E0",
INIT_08 => X"3FFF7D5000EC75088ED3FF7FC8790E46426CE06CB1F8E041051831FA3068D77E",
INIT_09 => X"C05FD7FF9BEFBDCEFBEE59FEF44F6603EFBEFAFCC2E35E7FDFD147CCF3F583FA",
INIT_0A => X"67FF1C7FBFADEB31E35768E8ED6BFDF3EB3EBF9DDBCE7FDC1DF8A760F3EACC02",
INIT_0B => X"5BDDCC3B336F7C548667D47B7737AF3FD62601EDC25B3533DCEB07F262213FFC",
INIT_0C => X"5F9A06E19F4D93A0EA0F78C35E30D78C35E30D78C35E30D78C35E986BC61AE31",
INIT_0D => X"5FD7AFEFDFFAF59B6FF28FE1D80D73D840607307DCFE1D80EF69A004DFFFF7FF",
INIT_0E => X"0004001F8041897B2FFFC6D86D70CE04FFFFF3FF1F5F5475BD7F72E4D75EBFAF",
INIT_0F => X"F60008003F008237B0040A00010003E020023E0201F45EC0010007E01047D17B",
INIT_10 => X"00010001DC0004C81003DE050A700200001DC0006863E8BD8002000FC0208FA2",
INIT_11 => X"2200E400002801E1A00004C21C0206F60081800800007B00010F02007EC09A0E",
INIT_12 => X"0880007E000807C7C1A612001E0015C7C19C22001E0015C59DFE82011A311AA0",
INIT_13 => X"00001BC00101F60409F0670840070809760409F06984800780097604067D0010",
INIT_14 => X"81019F40042100001F800203D81019EC085614000085C80023D81009CF008A74",
INIT_15 => X"FF802FFDFFAFD082003B032FB987E04021D481D4000819060801E0D00001231D",
INIT_16 => X"EBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEFFBFBFBFBBFCFBB0FFDFEFFEF2DFFFFFB",
INIT_17 => X"BFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAF",
INIT_18 => X"FAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFE",
INIT_19 => X"475B15BCF491E166CC8553F86EDB5C88646FFFFFFFFFFFFFFFFFEBFAFEBFAFEB",
INIT_1A => X"861861861861861861861861861861861861869A69A61861AFBD54D5F871C71D",
INIT_1B => X"984C26130984C26130984C26130984C26130984C26130984C26130984C261861",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000984C26130984C26130",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040201",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024,               -- Port A enable input
WEA      => wbe_a_lo_1024(3),               -- Port A write enable input
DIA(0)   => data_write_a(26),        -- Port A data input
DOA(0)   => data_read_a_lo_1024(26),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024,               -- Port B enable input
WEB      => wbe_b_lo_1024(3),               -- Port B write enable input
DIB(0)   => data_write_b(26),        -- Port B data input
DOB(0)   => data_read_b_lo_1024(26),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_27_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"00080A40000A41248002029000050A088000008242A0004404480002000A1155",
INIT_01 => X"2FFFF1C11F781C129C107DFFFE0860941E81258CA2B71C2220EC1B86E1A00002",
INIT_02 => X"E1000000810000014400FF6FFFF0FFFFF8007F1FC21110005080200000221FF0",
INIT_03 => X"4080026318C18226318C1821302232EAE00002BE001115FE48620040840A863F",
INIT_04 => X"643D4FFC2530000F003D821C0BFFFF8E9EF79E6D440748FED70060842105B0B0",
INIT_05 => X"D6F39020D1F8A3FAFDBFBACDC8FDC405D1DB7F1490E5EDB7D5CBADB2385D79C3",
INIT_06 => X"6FE000A38007C3032646EFF1F0B6FF46A78C39F8E723F2E47FE59C7F9ADA2612",
INIT_07 => X"00002820000000810000014401060C180190310540118DFF1000C0849673F6C0",
INIT_08 => X"3FF779100062B12A8EC3F47FC80208808210880C00082050000110023068D030",
INIT_09 => X"005F07E09BFFBD07FBAC09F8E42922038F7DF8BEC2E39C5F1FD047CEF1B582D8",
INIT_0A => X"63FF5D5F9FADE911E81C09818109E1F16B16B71092CE7ED81CF403601228C402",
INIT_0B => X"1BFDCC39732F3554866AD57C37BEAF1C152201A4C05B7531D56B05B06A213FF8",
INIT_0C => X"5BCA06F18FC59380F00E34430D10C34430D10C34430D10C34430F0861A2186B5",
INIT_0D => X"5B56ADAB5FAAE58B2F628EA0C80FA3F04040510768EA0C80CC61A0044DFFC6EB",
INIT_0E => X"0004001D800188792CE79715710AE4047FFD23FF315D54358D593474955AB6AD",
INIT_0F => X"520008003B000297B0040200010003E020001F0201E44A400100076000579129",
INIT_10 => X"00010001DC00004A10035E0408300200001DC000086BC8948002000EC000AF22",
INIT_11 => X"02002400002801E1A00000C01E0202F60080800800007B00000782006EC0820A",
INIT_12 => X"0080007E000006A7C10602001E0001A7C10C02001E0001C18DE282010A311AA0",
INIT_13 => X"00001BC00000FE0401F04300400708007E0401F04180800780007E04047D0010",
INIT_14 => X"81011F40040100001F800002F81011EC080604000085C80001F810094F008034",
INIT_15 => X"FF800C6DDDAFD082001B03249887E04001D481D4000009020801E0D00001021F",
INIT_16 => X"AB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6BF1EBDABD8E270BF84A25C6ACB777E3",
INIT_17 => X"B6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6AD",
INIT_18 => X"6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADA",
INIT_19 => X"490E2168100481CA860402104A471688747FFFFFFFFFFFFFFFFFAB6ADAB6ADAB",
INIT_1A => X"000000000000000000000000000000000008200000000000200072F210000001",
INIT_1B => X"05028140A05028140A05028140A05028140A0500804020100804020100800000",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000A05028140A05028140A",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040201",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024,               -- Port A enable input
WEA      => wbe_a_lo_1024(3),               -- Port A write enable input
DIA(0)   => data_write_a(27),        -- Port A data input
DOA(0)   => data_read_a_lo_1024(27),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024,               -- Port B enable input
WEB      => wbe_b_lo_1024(3),               -- Port B write enable input
DIB(0)   => data_write_b(27),        -- Port B data input
DOB(0)   => data_read_b_lo_1024(27),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_28_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"02200AA400180030808802A900002A08001280A08A801044104A1000001818C3",
INIT_01 => X"0AA00011460214428114180000882214413D0A71592A01D92213D28005210202",
INIT_02 => X"0451110A012100884000AA30200000000C100040104112101100008888200000",
INIT_03 => X"448000318C52A20318C52A20148810200111100C211004AA00034204200A2200",
INIT_04 => X"04004001001A90110000121402AA0000003C00000500000040080421080D0080",
INIT_05 => X"4060000C8001000000002E000000050000001610300000010000802202040012",
INIT_06 => X"1000002080001111001222000425A1040026A008000000000000000009328280",
INIT_07 => X"2491008A00491201210088400122448908A20402000408001000040820000000",
INIT_08 => X"20058310402A160026500000028040101004200C840082115554000112244814",
INIT_09 => X"4140000800000060000720000102028000000490160801020002200011100010",
INIT_0A => X"020000081B34211082B694D4D294000020020381040000000200032040004400",
INIT_0B => X"4800210C19808400500010009110091500020B408810000100200020408B0000",
INIT_0C => X"01028000080118020023604858121604858121604858121604858090B0242C00",
INIT_0D => X"010000800920040804020A6058003108402043058C460580653020005A004039",
INIT_0E => X"00000002800008014004104104420A00C000200005000010040A0020CC000200",
INIT_0F => X"520000000500000010000200000000000000280000040A40000000A000001029",
INIT_10 => X"00000000000000C0000002000830000000000000480008148000000140000020",
INIT_11 => X"020024000000000000000440000000020000800000000000000C00000040020A",
INIT_12 => X"00800000000001804006020000000500400C0200000005400A90000000100000",
INIT_13 => X"0000000000018200001003004000000142000010018080000001420000200000",
INIT_14 => X"8000080000010000000000018800008000060400000000000310000008000034",
INIT_15 => X"000002040080000000110006B081400000400000000009020000000000002200",
INIT_16 => X"802008020080200802008020080200802101210810C39A66A90A85420413A820",
INIT_17 => X"0200802008020080200802008020080200802008020080200802008020080200",
INIT_18 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_19 => X"DE21102C110A00246972BD89A40A0C22E1000000000000000000002008020080",
INIT_1A => X"2082082082082082082082082082082082082082082082080D35050758C30C31",
INIT_1B => X"0582C160B0582C160B0582C160B0582C160B0580C06030180C06030180C08208",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000B0582C160B0582C160B",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024,               -- Port A enable input
WEA      => wbe_a_lo_1024(3),               -- Port A write enable input
DIA(0)   => data_write_a(28),        -- Port A data input
DOA(0)   => data_read_a_lo_1024(28),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024,               -- Port B enable input
WEB      => wbe_b_lo_1024(3),               -- Port B write enable input
DIB(0)   => data_write_b(28),        -- Port B data input
DOB(0)   => data_read_b_lo_1024(28),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_29_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"79964E4BA01DACAB9E659792D00AAE160002829C7FDFEFCEE97C2815039D70C3",
INIT_01 => X"0ABFF9AB0775343F9AB01DF80D5821FC0FFF3FEFD1AF9FF1207FFBC7B9720586",
INIT_02 => X"002CCC60050E700080F6AAA7BFFC007189C7FF2FC00330E602800000074037F6",
INIT_03 => X"468003210868A63210868A68DA017D207200021C4E200CAA6186A40042FF4300",
INIT_04 => X"7C2FE002F0900001003C5316A6ABFFE21F36E02F0D03701F47D41800109FB281",
INIT_05 => X"4979440580F9B808F49F6A4DF00F8D01DC4B97369078249370F482E62BA41462",
INIT_06 => X"B250442BC81001E1870223FC0BF7F11507C423FE33C078F803F19F00E936721D",
INIT_07 => X"00011080012460050E700080EF020408EC8CFA01122149FF700200665A35D260",
INIT_08 => X"2BFD055040A452000443FF00007906464068406C31F84000000831FA1028575A",
INIT_09 => X"805FD017102690AA694551FE30444681E0820AD40201423FC00122C493500172",
INIT_0A => X"0600002AFFBE2330815568A8AD6ABC02A02A0B0CCB463B4C0748A720B1EA4C00",
INIT_0B => X"0850400A11414C005005000B51158936D20601A98A10200308A002E240010BFC",
INIT_0C => X"05928020194918A22A2268C81A32068C81A32068C81A32068C81A99034640C00",
INIT_0D => X"058102C48970541944B20FA1580561D040406305587A158046282000DBFFF13D",
INIT_0E => X"000000028040890327DCD28928324400DFFFF0001F1F0050342D42A086040B02",
INIT_0F => X"F60000000500802010000A000000000000022A0000141EC0000000A01000507B",
INIT_10 => X"00000000000004C0000082010A700000000000006800283D80000001402000A0",
INIT_11 => X"2200E4000000000000000442040004020001800000000000010D000010401A0E",
INIT_12 => X"08800000000801C040A6120000001540409C2200000015441DAC800010100000",
INIT_13 => X"0000000001019600081027084000000956000810298480000009560002200000",
INIT_14 => X"800088000021000000000201D800088000561400000000002358000088000A74",
INIT_15 => X"00802594A282C0000033010FB181E00020400000000819060000000000002305",
INIT_16 => X"C0B02C0B02C0B02C0B02C0B02C0B02C4B12B312912831A27FCFE7FFB175B6FF8",
INIT_17 => X"0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02",
INIT_18 => X"B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C",
INIT_19 => X"BBCF9F96EE7FFDF7FE783FFDFFEA0C00602FFFFFFFFFFFFFFFFFC0B02C0B02C0",
INIT_1A => X"EFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEEBAEBAEBAEBAEBBFFDF9FBEFFFFFFE",
INIT_1B => X"BFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFBEFB",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000FBFDFEFF7FBFDFEFF7F",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024,               -- Port A enable input
WEA      => wbe_a_lo_1024(3),               -- Port A write enable input
DIA(0)   => data_write_a(29),        -- Port A data input
DOA(0)   => data_read_a_lo_1024(29),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024,               -- Port B enable input
WEB      => wbe_b_lo_1024(3),               -- Port B write enable input
DIB(0)   => data_write_b(29),        -- Port B data input
DOB(0)   => data_read_b_lo_1024(29),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_30_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"F7FFBFFEFF9FE1F7FFBFFFFDFFD0000000000000000000000000000000000000",
INIT_1A => X"9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7AFBD75F5FDF7DF7F",
INIT_1B => X"F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE79E7",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000003F9FCFE7F3F9FCFE7F3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024,               -- Port A enable input
WEA      => wbe_a_lo_1024(3),               -- Port A write enable input
DIA(0)   => data_write_a(30),        -- Port A data input
DOA(0)   => data_read_a_lo_1024(30),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024,               -- Port B enable input
WEB      => wbe_b_lo_1024(3),               -- Port B write enable input
DIB(0)   => data_write_b(30),        -- Port B data input
DOB(0)   => data_read_b_lo_1024(30),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_31_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"129000008004A00804A40000400800020000000C005FEA005800200400050100",
INIT_01 => X"255FF18019700810180065FFFC0040801E80258CA2951C2200EC0906A0804140",
INIT_02 => X"E0000000000000011000550FDFF0FFFFF0007F1FC200000044000000000817F0",
INIT_03 => X"0000024210A30024210A3001002220C06044469200040154482000408400043F",
INIT_04 => X"602D0FFC2420000E003D80080955FF8E1ECA8E2D400340FE870060842100B030",
INIT_05 => X"0213100040F8A3F8FDBF944DC0FDC001D1CB6904A061EDB6D4C30490281831C1",
INIT_06 => X"6FC000830007C202060445F1F0D25E4207A099F0E303F0E07FE19C7F80402412",
INIT_07 => X"0000200000000000000001100004081001103107000185FF0000C0849673F6C0",
INIT_08 => X"1BF27A00000000000883F47FC800080002008000000820440000100220489020",
INIT_09 => X"011F07E013EFBC06FBA009F8E00120038F3CF82C44630C5D1FC002CCE0808248",
INIT_0A => X"61FF0C06C48BC801600000000001A1F00110101092CE7ED81CF0004012288000",
INIT_0B => X"11DCCC31222730048620C4382204A608142002A440492530C401049020221BF8",
INIT_0C => X"0888066187448380E00C10030400C10030400C10030400C10030600608018210",
INIT_0D => X"080204010200418301208480800D02D00040100240A808008840800405FF8640",
INIT_0E => X"0004001D000180780CE386106100C4043FFD03FF101D40008001304018081004",
INIT_0F => X"000008003A000217A0040000010003E02000160201E040000100074000478100",
INIT_10 => X"00010001DC00000810035C0400000200001DC0000063C0800002000E80008F02",
INIT_11 => X"00000000002801E1A00000801C0202F40080000800007B00000302006E808000",
INIT_12 => X"0000007E00000607810000001E000087810000001E000081846282010A211AA0",
INIT_13 => X"00001BC00000740401E0400000070800340401E04000000780003404045D0010",
INIT_14 => X"01011740040000001F8000025010116C080000000085C80000C8100947008000",
INIT_15 => X"FF800C609C06D082000A03200806A040019481D4000000000801E0D00001001D",
INIT_16 => X"010040100401004010040100401004010060C040040C200950402090128057C3",
INIT_17 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_18 => X"0040100401004010040100401004010040100401004010040100401004010040",
INIT_19 => X"00000000000000000000000000001000802FFFFFFFFFFFFFFFFF810040100401",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024,               -- Port A enable input
WEA      => wbe_a_lo_1024(3),               -- Port A write enable input
DIA(0)   => data_write_a(31),        -- Port A data input
DOA(0)   => data_read_a_lo_1024(31),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024,               -- Port B enable input
WEB      => wbe_b_lo_1024(3),               -- Port B write enable input
DIB(0)   => data_write_b(31),        -- Port B data input
DOB(0)   => data_read_b_lo_1024(31),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_0_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"ED39BA795990D275FB4A6E96ACC4731DEA4598B0AFB54867F6EE4618C3749803",
INIT_01 => X"8AA0047D8607944AC7DA180001ECA2444042106208408208C20022E9173734B3",
INIT_02 => X"1A7DDD79F9A73E6CCA7DAAF00001000008478020113D98E382FEDF333027C80F",
INIT_03 => X"75D341110C58F31110C58F32A208921F8051500147A0E4AB3493FB3A01EBE240",
INIT_04 => X"86424001531009B100425A97B2AA0001E03501D0A39C8F0078420001106D0C4C",
INIT_05 => X"BCC8CA2EBF03400700402BB20F00239E20341699198600000B08694B16434804",
INIT_06 => X"103FB860B2800161F8432200012DA185F80F24081C3C0707800E600056881308",
INIT_07 => X"B24197ABCDA467F9A73E6CCAFDC3870EEEEC44E2BDFE220094D03022210C011C",
INIT_08 => X"240581B5695EAA80262C080032BF07C7C1FC3F8E94F65B11555EAFFC1C306758",
INIT_09 => X"7E40000BEC004170040DB60017FED1CC0001045002984202003DB931192D60A5",
INIT_0A => X"120071411A74315881A28C141118000C5A85A60444210123820B43B40804674D",
INIT_0B => X"0820008E514045BB514F0106D1D8599581D3A958BC104A89215AC14C48898403",
INIT_0C => X"C261C01C48B1584A0CA3E2687A9A1E2687A9A1E2687A9A1E26870CD061343885",
INIT_0D => X"D274E93A758FA8683AC54B287522E10A74AF4AA59C568752662F5AC218000002",
INIT_0E => X"FF83C002783A0904231C70470C7E0B92800224008AE09FAD4BD48D1FC5D3A4E9",
INIT_0F => X"5BFF078004F075885DFBF7E15C06101C55E921F1F80FAB7FE0F0009E0E903EAD",
INIT_10 => X"F12E0380231F13978FF023FAFDBD9870380230F2D6081F56FFC1E0013C1D207D",
INIT_11 => X"DE7F263C0C8700125C0F8F3C43F1F10BBF7EFC61E01804E1E6C8F8FE807F67FB",
INIT_12 => X"02BE00017C17C1007E5E2E3081C5AC007E6F0E3081C5AC44418D65FE45DEE55B",
INIT_13 => X"61E0042786F103E9F01F9BC3C120C5A703E9F01F978B8C20666703E9F8A0FFED",
INIT_14 => X"FA7E283FFB414F80005F05F10FA7E283F78F6511C048278DCA174FF038FF15B4",
INIT_15 => X"0066A20B61692F293185D8D724E15D3FCC6B7C236FE0691B0700132C1F0EF880",
INIT_16 => X"3A4E93A4E93A4E93A4E93A4E93A4E93A4F942F92E9628540AD2A91442525A000",
INIT_17 => X"A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E9",
INIT_18 => X"4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93",
INIT_19 => X"55F3898E09B56C74DAB15D1CF13501AA495000000000000000003A4E93A4E93A",
INIT_1A => X"082082082082082082082082082082082082082082082082082084E41DC71C71",
INIT_1B => X"E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F82082",
INIT_1C => X"FFFFFFFFFFFFFFF94A5294A5294A5294A5294A52800003E1F0F87C3E1F0F87C3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"3060C183060C187FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"BDEBA0000000000000000000000000000000000000000000003060C183060C18",
INIT_28 => X"168ABA002E82145085155545F7AA975EFFFAABDE00FFAEBDFFF5D2EAAAAAF7AE",
INIT_29 => X"7FFFE10005542145557FD5545FF8000155087FC0155F7D168B55007BFDF45085",
INIT_2A => X"7FFC0010080017555555568AAAFFFFD7545AA8028A00A2802AABAFF8028BEF5D",
INIT_2B => X"FF842AABAA2AE95545FFD168ABAF7AEAAAAAA2FFFDF4500043FE105D2E954BAF",
INIT_2C => X"5007FD7400550415410002E974BA5D5168A00A2D142155005142010FFAE820AA",
INIT_2D => X"FFF780000BA007FE8AAAFF803FFFF5D2A821550000000BA007FD55FF5D7FC014",
INIT_2E => X"000AAFBEAA00007BFDFFF082EBDF455D5142000082E82145FFD17DFEFFFD168B",
INIT_2F => X"DFD75D2AA8A80EA8E2FE3F000000000000000000000000000000000000000000",
INIT_30 => X"68B551475FAF6D1C556F0AA1C24AABEA495FC716F002A975FFE3AA95E00EBAEB",
INIT_31 => X"42A0070071C50BAFEF1FAE0016D56A16D557BC257D415E0216FA3F1E8FC0145B",
INIT_32 => X"8010E004924874825D7FEAA85487FD24AFE3D02DAAAE12BD5545A2803AA00005",
INIT_33 => X"120155EA568E870BAEB8A05A2AEA8B50F55A2F150005A3A438BD04AFAB8F550A",
INIT_34 => X"545E055FFBE81D0BE8EA8A3AA05A2A5504001C74BA42A1571E8028E3DB7816D0",
INIT_35 => X"A5C7E3DFFFE90B45B47ABA497A82FFAFD2A82485FD2415A105C21451ED42A002",
INIT_36 => X"00000000000000000000B55EAAA100AA1D0F6F480B6A555A2A57A002A3D5FDB6",
INIT_37 => X"5EFAAAAB5E1AF3AABFF45592E88A0AFE80A8B0A0000000000000000000000000",
INIT_38 => X"65F520EBE9EF67D7BEA1FD5D556ABEF5D557FEBA55022A3F70C6B405F4D2AE97",
INIT_39 => X"C114728007521170821CE0FDE69411A8DED57CE1055555E5F58EFFC01FE2CACB",
INIT_3A => X"42341D5DEEBEF55080034E0A592A4AD0079C75D6070CC5CBB0280C029ABAA3EB",
INIT_3B => X"7F353AAF6C77F7F20D968BF57812A95E02A2AAB5EB0F280800EFAEE9F5D18F31",
INIT_3C => X"C91565455C141E41887D58AC448B69C30E02116220415A9540AA854140A0A204",
INIT_3D => X"DE6BE93172D7D625B556EEAB157ABEBE1B4D792A4AD1183454180DD3FDCAAAB7",
INIT_3E => X"F0000001FF0000001FF0000001FF0000001FF01EABC4B8014174FF7DA80F52FE",
INIT_3F => X"FF0000001FF0000001FF0000001FF0000001FF0000001FF0000001FF0000001F")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024,               -- Port A enable input
WEA      => wbe_a_hi_1024(0),               -- Port A write enable input
DIA(0)   => data_write_a(0),        -- Port A data input
DOA(0)   => data_read_a_hi_1024(0),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024,               -- Port B enable input
WEB      => wbe_b_hi_1024(0),               -- Port B write enable input
DIB(0)   => data_write_b(0),        -- Port B data input
DOB(0)   => data_read_b_hi_1024(0),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_1_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"212C001411984004084D000508C53810A03D1450E839B003342114428A000803",
INIT_01 => X"00000019400B100A8196000000CC004400400002000000000000028001340000",
INIT_02 => X"052137AE8031800C0044009000000000061800001CD4019802AD04CCCFC20004",
INIT_03 => X"04514108C60C21008C6042108400000201440020505100000043C30E10E9F000",
INIT_04 => X"02104001011DEFE088805681920000008000004001900800004002108C280008",
INIT_05 => X"040002340105000200000000080001900010000108040000000008411600401C",
INIT_06 => X"1034001042800808201000000001000820020000102000040000000000800180",
INIT_07 => X"64BF81A15EDFDE8031800C00843060C19E030022103600000450020800040004",
INIT_08 => X"00008004691687AA840008000090248CC84E000046000311555521F183060AC5",
INIT_09 => X"0820800D08100171000DB000154440C800400500000852020011200201012021",
INIT_0A => X"02000040001000880A2A04445004000102002041000001008208001440004140",
INIT_0B => X"4820018A1140440078050040511000102000A008183000010002404400000000",
INIT_0C => X"1000C80008000C030030880C2A030A00C28030A80C2A030A00C28018D4061401",
INIT_0D => X"10040802050080200284401C0022880F009E08008205C0020118088018000000",
INIT_0E => X"0F03C00280000000420860C60C0C0B92C0000000004000010042000040102008",
INIT_0F => X"001E078005000108400005E11C0610000000288058000003C0F000A000100000",
INIT_10 => X"F10E0380000000C202300000008D187038000000480800000781E00140002000",
INIT_11 => X"806302380C870010000004400100110800007861E0180000000C400680000001",
INIT_12 => X"023E00000000018000580C308000050000610C30800005000215006800000101",
INIT_13 => X"61E0000000018100B0001843812000014100B00016030C20000141002880026D",
INIT_14 => X"400A20009B404F80000000018400A20044096111C04000000304026000501580",
INIT_15 => X"0046820040082300218450C2800010094000482141E060190700100000002200",
INIT_16 => X"020080200802008020080200802008020080008008600500A82A1100A8000000",
INIT_17 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_18 => X"0080200802008020080200802008020080200802008020080200802008020080",
INIT_19 => X"81328A46BABEFC54A0810C7452B4428A14000000000000000000020080200802",
INIT_1A => X"AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA28A28A28A28A2A8218D2C0C924925",
INIT_1B => X"E974BA5D2E974BA5D2E974BA5D2E974BA5D2E975BADD6EB75BADD6EB75BAAAAA",
INIT_1C => X"FFFFFFFFFFFFFFFD8C6318C6318C6318C6318C63000002E974BA5D2E974BA5D2",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"70E1C3870E1C387FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"5555500000000000000000000000000000000000000000000070E1C3870E1C38",
INIT_28 => X"EBDF455D2EAABEFF7FFE8BFF5D0002155557FFFFFF007FC21EFA2FFD74AAAAD5",
INIT_29 => X"AA95400552AAAABAFFD1574105D7FD75FFAAAA800AAF7AA974BAFFFBE8B45F7A",
INIT_2A => X"0517DF555D2EAAA1055000015500557DF45AAD1400BAA2AE801550051555EFF7",
INIT_2B => X"FFD540155557FD5400F78028BFFFFFBEAB55F780020AAAA80020AA082EAAB550",
INIT_2C => X"AFF842ABEF5D517DF55552A974AAF7AE820AA0851574BAA2D1574AA5D7BFDEBA",
INIT_2D => X"EFAAD1575EF557FFFE10557FFFFFFFFD56AAAAFFFFD7555AAD168B45AAAEAAAB",
INIT_2E => X"0005D7FFDF4500043FE105D2E954BAF7AE80010082A97410557FEABFFAAFBE8B",
INIT_2F => X"51C7A2FBD5490BFD1C056A000000000000000000000000000000000000000000",
INIT_30 => X"974BAF7FFEFB45FFAABDF55492AA8BC2EBDFEAF7F1F840017D4975D2FEF147FC",
INIT_31 => X"080BEF495FC71D54124924385FAAA8AAAE3D145410F7F1D55D71C002DABAEBAA",
INIT_32 => X"002D082082AB8B6DBEDB7DF7F540E2AE85028B40155145F7AF6DBED5450AA1C2",
INIT_33 => X"78E021FF1471FDEAAFFD56F16D5571D2E28E38E0216FA2D1E8E80140F45082B4",
INIT_34 => X"A2DA3FB7DAAD4AAAAF487BC70BFA97F7AF6D417E92482BF84020BA495557E3FF",
INIT_35 => X"55554ADBD7A2FFC7BEFF6FFD7FC7002FD74951D71EDFFABFD16FAAAE92BD5545",
INIT_36 => X"00000000000000000000547AB8F550A8010E00492487482FFFE82A85EBAE2FFC",
INIT_37 => X"1EF005162BEF047FD5545AAFBF7400FBF9424F70000000000000000000000000",
INIT_38 => X"714F8338AAAA1D0AE974AAF7FFFDF55F7AABFF55082CA8B4DF6C1E8F5E540002",
INIT_39 => X"EABEF75550ACBB7582225FF5843404547184164AA5D2EBEEB0A2D555410D3555",
INIT_3A => X"FEAAEB083BC1000FF8409000512AEABFFDF79DCBF755962010BDCBBC21455D7F",
INIT_3B => X"801F8BA0C57740BDAA0688E5405D57D412F7D55F5E50C7F401BAAE8403CF5A3F",
INIT_3C => X"5D16BABAA3EBC3157ABD5FFE55F2AA9FEAFDF7F431A9F7FFE81FF013A8001AFF",
INIT_3D => X"FB863550229BCABEB7DA403FFFDA2FBF7FED2C7F955445079E280A00C56145EF",
INIT_3E => X"0000000000000000000000000000000000000596EBEF55080034E0A592A4AD00",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024,               -- Port A enable input
WEA      => wbe_a_hi_1024(0),               -- Port A write enable input
DIA(0)   => data_write_a(1),        -- Port A data input
DOA(0)   => data_read_a_hi_1024(1),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024,               -- Port B enable input
WEB      => wbe_b_hi_1024(0),               -- Port B write enable input
DIB(0)   => data_write_b(1),        -- Port B data input
DOB(0)   => data_read_b_hi_1024(1),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_2_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10E006600180111284380310006289800480032283E000A34301002001A0817",
INIT_01 => X"0005A00810790848048044A54E404350404000720885800802000906E4910200",
INIT_02 => X"407004208400408044C600C50AA055254010541A110222841200000002402544",
INIT_03 => X"0600011004182401004102408C28414043101000408118000145840440F5C415",
INIT_04 => X"5035855703A2900A000CD3088400F40688C9844409060850925E58A4081A0221",
INIT_05 => X"0200840D1021A15AC50494894850890540D1E12020C6E510818500440A280090",
INIT_06 => X"113044094002801020440090A8011A1224AB9380552102442884882A20004097",
INIT_07 => X"000100880004428400408044860000008C022402102100AA40004404B5075460",
INIT_08 => X"15C23440408C862A2A12382A8A5244145048C06085008010141521F000001240",
INIT_09 => X"400582B9033AA0E7AA4110B0506744810554542450694E710A836188C2C00222",
INIT_0A => X"443518360012C2210B020414109130A28038188096A06B8C120CA440A9C00802",
INIT_0B => X"1345E53300EC68005605002964AF222A5704004D080211121C80024200821780",
INIT_0C => X"181080C1110C882202211488452213C88472213C88472213488441109A442231",
INIT_0D => X"008204440210091341208041000810C00000300220201800A908000038AD0284",
INIT_0E => X"00040002804180300E88D28D206A40000554815500481440300000C44A081100",
INIT_0F => X"000008000500828700000000010000000002380000A00000010000A010050000",
INIT_10 => X"00010000000004CA000214000000020000000000684280000002000140200500",
INIT_11 => X"000000000020000000000442100002840000000800000000010C000026000000",
INIT_12 => X"00000000000805A4800000000000152300000000000015801272000100210020",
INIT_13 => X"000000000101C00000C000000000000940000120000000000009600004050000",
INIT_14 => X"0000130000000000000002018000106000000000000000002380000141000000",
INIT_15 => X"55000190000000000002000280000000011080C0000000000000000000002310",
INIT_16 => X"40902409064190641906419024090244902A9003004800415120D4A190804241",
INIT_17 => X"0900409004090641906419064190240902409024090641906419064190240902",
INIT_18 => X"9044090040900409004190441904419044090040900409004190441904419044",
INIT_19 => X"75960040138D70C030B51C50C7D100A2052F81F81F83F03F03F0419044190441",
INIT_1A => X"0410410410410410410410410410410410410410410410410248602081659659",
INIT_1B => X"5128944A25128944A25128944A25128944A25128944A25128944A25128941041",
INIT_1C => X"FFFFFFFFFFFFFFFE1084210842108421084210843FFF825128944A25128944A2",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"7FD5FF555815607FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"2AA000000000000000000000000000000000000000000000007FD5FF55581560",
INIT_28 => X"FC21EFA2FFD75EFAA8415410AA8415555087BFFF55A2AA800BAFFAE954000800",
INIT_29 => X"84155EFA2AEBDEAAA2FBEAABA5D7FE8B555551421455D0002145552EBFEBA007",
INIT_2A => X"2AEBDF555D2E954BAA2AA974BAFFFFE8B45552EBDF45FFAEAABFFF7FFE8B55F7",
INIT_2B => X"AAAAAAAAAFFD1574105D7FFFF555D2AAAAAA5D2E820BAA2FBEAB5555557DF55A",
INIT_2C => X"50055575EFFF84021555D043DEAA5D04021EF557FC21FFAA8428BFFAAAA954AA",
INIT_2D => X"10085568A00FF80175FFA2D17DFEFF7800215500557DF55AA80001FFAA800015",
INIT_2E => X"0005D00020AAAA80020AA082EAAB5500517DF555D042AA10A284154005D00154",
INIT_2F => X"00AAFFAA9543A080038A2A000000000000000000000000000000000000000000",
INIT_30 => X"0017D5D20B8EAA007FC51C7A2FBD55D2BE800042AFE8E1557D0075D2F45BEAA8",
INIT_31 => X"AA8BC7EBDFEAFEFFD00105FFBC20BDEAAA2FBF8AAA557BE8B6D5D5FFABEF4904",
INIT_32 => X"FFEFB6D555578F7DB6A0BDF7D480E174BFA02A974BAF7F5EFB455D2ABDF55492",
INIT_33 => X"ED1FDE90E3A497492B6AAADAAAE3D155E105571D55D71C002DABA5524820BAB6",
INIT_34 => X"BE8F401D7B6A0001470155C51D0092A071555D5E3AE821D00001FF0871C016DB",
INIT_35 => X"5BE8555400550A38428007FED000E3DA3DFD5E3DFFFBD5A38A021551C5F7AF6D",
INIT_36 => X"00000000000000000000410F45082B4002D082082AB8B6D1C5B7DF7FF78E075C",
INIT_37 => X"5EF005560B55F7AA800AAF7AA954AA00042AAA20000000000000000000000000",
INIT_38 => X"ABEF057D68F5F5A00021EF55042AAAA007FD5555AAFBD7545FBB8020A3F7AE97",
INIT_39 => X"7DF55D7AABFF5428ACA8F45A6C1E8F5EFF84165EFF7802BAB0A2FFEAABA557BE",
INIT_3A => X"CA8AA80800020AAF7FBFFFEF04552ABFFFF841FFE75CA882108202E974AAF7D5",
INIT_3B => X"00151FF0C57401E5F3D1E00A1A884174A8FFAEBFEB0A2D55541051555694F002",
INIT_3C => X"2AA801455D7FE8BFFF680800FFF7AAA155F595542455512A975455D3AA8A0055",
INIT_3D => X"5D79FCAF774AE005BE7895554005D2A8A0B882FFFFE10AAAAAB755A66B6AF56A",
INIT_3E => X"00000000000000000000000000000000000000C3BC1000FF8409000512AEABFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024,               -- Port A enable input
WEA      => wbe_a_hi_1024(0),               -- Port A write enable input
DIA(0)   => data_write_a(2),        -- Port A data input
DOA(0)   => data_read_a_hi_1024(2),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024,               -- Port B enable input
WEB      => wbe_b_hi_1024(0),               -- Port B write enable input
DIB(0)   => data_write_b(2),        -- Port B data input
DOB(0)   => data_read_b_hi_1024(2),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_3_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"210C00A20020000108430020001600B8156021104940741B3530400E02B92203",
INIT_01 => X"014C9BCA58B1296D24A402C992500B69404040028804A0080A000416A8D90A08",
INIT_02 => X"C12026A484318004404405C9C66E331352180D468B8203980300204442E02B34",
INIT_03 => X"04000748D60D24648D60524C88804D0215011020D15018148040C10A70E1D58C",
INIT_04 => X"18283333240FE41244187308C9104D70944852640901083801750EB0A418C220",
INIT_05 => X"0613142D01912CC2A1B4140528348900C612A104201C689044340ED413A07649",
INIT_06 => X"119000034019881822104C5E68035250A222829710A0A02C18C01A9920842413",
INIT_07 => X"402F00AB0016CA0431800444841020509D038B021230C1990001C644C8273200",
INIT_08 => X"16905000408482088290E8E64010248C4A5AA840C2000110001521F0810A92E7",
INIT_09 => X"0003CE6581BD016342A951AB146C4480530C3B2A8088D3542651670200C1826A",
INIT_0A => X"00735D36209A8A20020894004284B660821030C8990467401218004041020002",
INIT_0B => X"512445B740457154562F957CC08B00093700080D0A4851001D8302D20A0A1530",
INIT_0C => X"00508650008008021021A40861021840869021A408610218C0869810D6043095",
INIT_0D => X"1C8508438450801043A08090380A8834207007022209038080190000999C8F84",
INIT_0E => X"000400200000C0002A48A206204C4205F3304B33004C0041006240140A1C310A",
INIT_0F => X"0000080040000083800400000100000000008400018040000100080000510100",
INIT_10 => X"0001000000000800000244040000020000000100002A0080000200100000A702",
INIT_11 => X"000000000020000000200000080002C000800008000000000022000006808000",
INIT_12 => X"0000000000000A2281000000000040A3810000000000402001400000022002A0",
INIT_13 => X"000000000004200001C0400000000010200001C0400000000010000004490010",
INIT_14 => X"0001070004000000000000060000104C08000000000000001000000903008000",
INIT_15 => X"CC004050CA0C00020220200070040000010401C4000000000000000000100008",
INIT_16 => X"4310E4310A4210A4210A4210A4210A4210A8D0830A68010001B4DA881048061C",
INIT_17 => X"21084290A4210A4210A4210A4210A4210A4210A4210E4310E4310E4310E4310E",
INIT_18 => X"90A421084290A421084390E4310C4390E4310C4390E4310C4290A421084290A4",
INIT_19 => X"015303C0C78C706428A14C586291000A044001FFE000003FFC004290A4210842",
INIT_1A => X"2492492492492492492492492492492492410410410410412821600001249249",
INIT_1B => X"51A8D46A351A8D46A351A8D46A351A8D46A351A9D4EA753A9D4EA753A9D49249",
INIT_1C => X"FFFFFFFFFFFFFFFC00000000000000000000000038F56351A8D46A351A8D46A3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"55AB02055AB0207FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"420000000000000000000000000000000000000000000000007FFFAB57FFFAB5",
INIT_28 => X"A800BAFFAE9554508002AA00AA843DF55FFAA955EFA2D168B55557BEAA000055",
INIT_29 => X"002AB55AAAA955EF005568A00087BE8BFFA2D155410AA8415555087BFFF55A2A",
INIT_2A => X"AAABFF5508003FF555D0002145552ABFEBA007FC21EF007FD75FFAA841541008",
INIT_2B => X"082EBDEAAA2FBEAABA5D7FC0155005168B455D042AB45F7FFD741000042AA10A",
INIT_2C => X"FF7FBEAB55F7AABDEBA5D7FC2010A2D1575FFF7AA975555D2E80145F78415545",
INIT_2D => X"EF5555554AA087BC01FFFFAAAAB55552A954BAFFFFE8B55552EBDE00F7AEAABF",
INIT_2E => X"000082E820BAA2FBEAB5555557DF55A2AEBDF555D2E954BA002EAAABA002A821",
INIT_2F => X"FB7D5D7FEAA3808554203A000000000000000000000000000000000000000000",
INIT_30 => X"1557D1475FAF45BEAA800AAFFAA95578080038A2AA28E3AF55E3A0BA5D7AADB6",
INIT_31 => X"BD55D7BE80004AA1E8E2AB55B6A0925D7085F6AA10087FEABD7AAD57AEBAB68E",
INIT_32 => X"F5D0438140E2FA38B6AEBFF6D1D04AAFFA41040017D5D20B8EAA007FC51C7A2F",
INIT_33 => X"D0A901FFFF801557D1C20B8EAAA2FBE80AA557BE8B6D5D5FFABEF49002FB55FF",
INIT_34 => X"5D20BDE00EBAAA8BC7EBDFEAFEFAB8ABAE925D21C7010EADB525D7FFAE975C75",
INIT_35 => X"F002EADA921420871D74971D24820875C21D5EB8AA8FFF012A954BAFFF5EFB45",
INIT_36 => X"000000000000000000001C24820BAB6FFEFB6D555578F7DB6A0BDF7DEB8E125F",
INIT_37 => X"B55A28408145AAFFFFFFF5D7FEAABA0051400A20000000000000000000000000",
INIT_38 => X"AB55FAD568AA2AFAE975EF555168B55F7AA800BAF7AA955EF00042AAA2A2AEAA",
INIT_39 => X"2AAAA007FD55558A7BD7145FBB8020A35D2ABEF55F7800015F087FEAA00007FE",
INIT_3A => X"968F575D003FF55F7D5420BA5D2ABFEAAF7AE9DFF759A82AEF70800021EF5504",
INIT_3B => X"FFD5145FBAC9755F05040255FFD84175EF55002AAB0A2FFEAABA557BEA3EF057",
INIT_3C => X"82E974AAF7D57DF45552A3FF10AA8429F45A7D5EAF5FFBAEAAA10554155400AA",
INIT_3D => X"FF843FFE77C80825BC052ABFE10550415557085540000005156155FE90A8F5C0",
INIT_3E => X"00000000000000000000000000000000000005500020AAF7FBFFFEF04552ABFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024,               -- Port A enable input
WEA      => wbe_a_hi_1024(0),               -- Port A write enable input
DIA(0)   => data_write_a(3),        -- Port A data input
DOA(0)   => data_read_a_hi_1024(3),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024,               -- Port B enable input
WEB      => wbe_b_hi_1024(0),               -- Port B write enable input
DIB(0)   => data_write_b(3),        -- Port B data input
DOB(0)   => data_read_b_hi_1024(3),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_4_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"A108400020612C80284210081034849800A00030300004833522C82D04A16002",
INIT_01 => X"2043998A1839284D1CA0650E1E504368403008418984014902030806A0D10200",
INIT_02 => X"C120042200000000044441CE01E80F00A49043118680008002000000026208E4",
INIT_03 => X"040001020019200020011209CC0164C060000000690111040144800042F5C403",
INIT_04 => X"7029AF0F81A00010CCA47700CC513CAC0D0B8E02010740E19754080108988021",
INIT_05 => X"02139405007133C0712244CD20F20105D583000020E9892201D304D42A9835E1",
INIT_06 => X"9190440300078002014405D9EE814C0284A883B6D7038AE079059B7800048092",
INIT_07 => X"000100AA0004408000000004840400008D200102503000782000C00C8025C000",
INIT_08 => X"00728A00408403220811991E02120C044058080004000001101121F220000260",
INIT_09 => X"811001E1185B38AD23C3707AD46440818F3CF80EC423CA7D01D123C80200816A",
INIT_0A => X"45810810A01B40216361056D6150F41200280001900439001FD8A00041400000",
INIT_0B => X"11FC88076266E800D605402962A820211500024808010512C40106D222223B14",
INIT_0C => X"0408804116040B02C02C500B0C02C100B0C02C100B0402C300B0401618058611",
INIT_0D => X"040200050200501301208482200D00D0A0408402C4282200A84800009B878680",
INIT_0E => X"00000020000100024AC88300300060090F0D830F00025400300204D018000804",
INIT_0F => X"8000000040000206A2000800000000000000950002E010000000080000588040",
INIT_10 => X"0000000000000808000554000200000000000100006D0020000000100000BB00",
INIT_11 => X"0000400000000000002000001A0002504001000000000000002280000D800800",
INIT_12 => X"0800000000000E2C802000000000408D801000000000408012440000200110A0",
INIT_13 => X"000000000004680003A0040000000010280003800800000000102800000B0000",
INIT_14 => X"000005C0002000000000000620000158000010000000000010A0000B00000200",
INIT_15 => X"C30146200400104002602600400000000294004000000004000000000010001A",
INIT_16 => X"0080200000008020000000802000000080080000004090014134DA101288C6DB",
INIT_17 => X"0802000000000401806010040180601004018060100000802000000080200000",
INIT_18 => X"8060180601004010040080200802000000000000802008020000000000008020",
INIT_19 => X"C0A28A063807E0500014063450404882846FFE000003FFC00000010040100401",
INIT_1A => X"AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA28A28A28A28A2934C8D0CCD145144",
INIT_1B => X"68341A0D068341A0D068341A0D068341A0D068351A8D46A351A8D46A351AAAAA",
INIT_1C => X"FFFFFFFFFFFFFFFC0000000000000000000000001FE32068341A0D068341A0D0",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"408102040810207FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"800AA00000000000000000000000000000000000000000000040810204081020",
INIT_28 => X"168B55557BEAB4500554200000557FE10FFFBEAA10007FD7410FFAA97555082A",
INIT_29 => X"55574105D2A800AA00043FEBA5D7FEAA00007BE8AAAAA843DF55FFAA955EFA2D",
INIT_2A => X"57BC00AAA2FFEAAAAAA8415555087BFFF55A2AA800BAFFAE9555508002AA0000",
INIT_2B => X"A2AA955EF005568A00087BE8BFFA2D17DE1000517FE10AAAAA8AAA002E975455",
INIT_2C => X"FAA8417410A2D140000F7FBC2010A2D157400AAAE974AAAAAA974BA08002AB55",
INIT_2D => X"EFA2AABDEAA087BEAAAAA2FBD54BA080002145552ABFEAA007FC21EF007FD75F",
INIT_2E => X"00055042AB45F7FFD741000042AA10AAAABFF5508003FF55F7D568A00552EA8B",
INIT_2F => X"5400F7A49057D0824850B8000000000000000000000000000000000000000000",
INIT_30 => X"3AF55F7A0925D7AADB6FB7D5D7FEAB7808554203A145178E00FFFBE8A101475D",
INIT_31 => X"A9557D080038AAA145157428492E8008200043FE925571EFA380871C7028A28E",
INIT_32 => X"AEA8A9200249056D4175C5092AAF5FDA38BE8E1557D1475FAF45BEAA800AAFFA",
INIT_33 => X"AA4954281C0E2FB55B6A0925D7085F6AA10087FEABD7AAD57AEBA08517DE00AA",
INIT_34 => X"007FC51C7007BD55D7BE80004AAFEDB42028EBFBC2028BED152438AAA092492A",
INIT_35 => X"AF7DF6AA00412EAABFFAA803DEBA0875EDA80BEF1C743840040017D5520B8EAA",
INIT_36 => X"0000000000000000000041002FB55FFF5D0438140E2FA38B6AEBFF6DBE84AAEB",
INIT_37 => X"A00FFFFEAA105D5155410FF84021EF0800154B20000000000000000000000000",
INIT_38 => X"DEBA0851574B2AAAEAAB55F78400145AAFFFFFEF5D7FEABFF0051400A25D5568",
INIT_39 => X"68B55F7AA800BAF7AA955EF00042AAA25555410BA082E8201000043FE005D517",
INIT_3A => X"568AA200557DE00AAAAAAA000804001FF005575408AA557FEB2FFAE975EF5551",
INIT_3B => X"D1550AAAA8002010F2AC154B25F2ABFF55F7800015F087FEAA00007FEAB55FAD",
INIT_3C => X"800021EF55042AAAA007FD5555087BD6145FAAC000A2A6FBC00BAAAFBC00BAF7",
INIT_3D => X"F7AEBDFF779A82AA43F7FBE8A00082EA8BFFAA843FEBA08517DE00F3F9574B30",
INIT_3E => X"000000000000000000000000000000000000008003FF55F7D5420BA5D2ABFEAA",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024,               -- Port A enable input
WEA      => wbe_a_hi_1024(0),               -- Port A write enable input
DIA(0)   => data_write_a(4),        -- Port A data input
DOA(0)   => data_read_a_hi_1024(4),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024,               -- Port B enable input
WEB      => wbe_b_hi_1024(0),               -- Port B write enable input
DIB(0)   => data_write_b(4),        -- Port B data input
DOB(0)   => data_read_b_hi_1024(4),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_5_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50DF4A0791B3FCB694379283C81FD996A091832102004A336A20E03C040C002",
INIT_01 => X"805FBDC69830A84D5C6A60000C34C26841280A00084000C8C212892EEAD53235",
INIT_02 => X"3B2026B578918E640A4F01CF8011FF0002080000082CA9998276DF7772C7C80D",
INIT_03 => X"37134108420D700084205702A4008A1D9100002171C0E0051554D93A11F5D140",
INIT_04 => X"8A41A0FC03A56DA000425A819410E3816C086198A388B702A8CA1210844A0C4C",
INIT_05 => X"B1808A062E8BC835F5E84532D708238A282F00A9291224800A2861490343082C",
INIT_06 => X"903FB8483A90581859050424100940825C6184401CDC451B860A6507160C4100",
INIT_07 => X"D26F068BCC96CDF8918E640E96D1A3469D6300E2FFEA27F8E4D23248130E259C",
INIT_08 => X"0BFA82E568442B2A082C0A7E3014250D49DA37A2420619000002AFF48D1222E5",
INIT_09 => X"3F005001E40969289429360416DCD1C46083030604B1CA20C03DF83B0A2C60A5",
INIT_0A => X"14613C71005A10492B888120288F480D58858449026145B3830F449449062B4F",
INIT_0B => X"11AC04934AC648BFD727C031E64170A137D5AA5C3E4B0F8A3C58C34C002290E3",
INIT_0C => X"CA29C6CC50384B6AC6AC86AB31AACA6AB39AAC86AB39AACA6AB3055643559C31",
INIT_0D => X"C673E33CF28F38603855401985228A0614BD30A0A2819852011E5AC2B87F9182",
INIT_0E => X"FF87C002F87A803E460B2516510CA594FF0044FFA4B08BAC4BB2CD0F09CF84E3",
INIT_0F => X"0DFF0F8005F0F5100DFFF5E15D06101C55EB29F1E00BE53FE1F000BE1E802F94",
INIT_10 => X"F12F0380231F17D78FC029FFF58D9A70380230F2FE0017C37FC3E0017C3D005F",
INIT_11 => X"FC7F023C0CA700125C0F8F7E43F1F001BFFE7C69E01804E1E7CCF8FC003FF5F1",
INIT_12 => X"023E00017C1FC1A4BFD82C3081C5BD27BFE30C3081C5BD00C02365D645CEEF5B",
INIT_13 => X"61E0042787F181E9C1EFD8CB8120C5AF41E9C18FD60F0C20666F41E9F009FFFD",
INIT_14 => X"7A7C077FFF404F80005F07F187A7D14BFFC96111C048278DEB074F9930FF9D80",
INIT_15 => X"C064014B8B652E2B3120C81284641D3E8DBF7D636FE860190700132C1F0EFB80",
INIT_16 => X"38CE1384E3384E338CE138CE1384E33C4E3ECE32E128882551349A1CBAA44103",
INIT_17 => X"84E3384E3384E3384E338CE138CE1384E3384E338CE138CE1384E3384E338CE1",
INIT_18 => X"CE138CE138CE138CE1384E3384E3384E3384E338CE138CE138CE138CE1384E33",
INIT_19 => X"F5E5BB4E7F7B9DB7FF3A1B6DB7E8410A8C000000000000000000384E3384E338",
INIT_1A => X"BEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEF9F7CFDFDDCF3CF3D",
INIT_1B => X"BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEFBEF",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000001711C7BBDDEEF77BBDDEEF77",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"FDFFF00000000000000000000000000000000000000000000080000000000000",
INIT_28 => X"FD7410FFAA97410082A800AAAAAE955450055421FFFFFBC0010AAD5574BA557F",
INIT_29 => X"7FD74000055574BA5D7FD7555A2D5575EF55517FF5500557FE10FFFBEAA10007",
INIT_2A => X"0002AABA5D2ABFFFFAA843DF55FFAA955EFA2D168B55557BEAB5500554200000",
INIT_2B => X"5D2A800AA00043FEBA5D7FEAA00007BC00AAAAAEBDF45A28428B45FFD168BFF0",
INIT_2C => X"5080028A00A2FFFDE00F7D57FEBAFF80174BAAAD1555EF555555555005557410",
INIT_2D => X"BA5D2E821FFA2D5554BA557BD75FFAA8415555087BFFF55A2AA800BAFFAE9555",
INIT_2E => X"00000517FE10AAAAA8AAA002E97545557BC00AAA2FFEAAAA082A97545F7D5420",
INIT_2F => X"7010BEDF524AA5571FDFEF000000000000000000000000000000000000000000",
INIT_30 => X"78E00EBFBE8A101475D5400F7A49043D0824850B8A2AE9756D145B401FFFFFFC",
INIT_31 => X"FEAB7D0855420BA1471D74380851524BA5571D757DB6D5525EF555178F6D1451",
INIT_32 => X"8A28B6DEBDF6DBEF1C0A28AAA5524BFFFFA28E3AF55F7A0925D7AADB6FB7D5D7",
INIT_33 => X"5555057D145152428492E8008200043FE925571EFA380871C7028B6AEBDF45B6",
INIT_34 => X"BEAA800AAFFAA9557D080038AAAA2FBF8E10EBD578EAAFF8415482BED1555EF5",
INIT_35 => X"81C209256DFFDF420BA552A821FFB6DF574A85575C55EFBE8E1557D1475FAF45",
INIT_36 => X"0000000000000000000008517DE00AAAEA8A9200249056D4175C50920875FDA3",
INIT_37 => X"5FF5D7BC21EFF7FBD7400F7FBC00BA55557DFF70000000000000000000000000",
INIT_38 => X"01FF5D5568BE7555568A00AAFFEAA105D5155410FF84020AA0800154B2AAAA97",
INIT_39 => X"00145AAFFFFFEF5D7FEABFF0051400A25551554BA0051400BA5551575EFF7D14",
INIT_3A => X"1574B2FFAABFF45FFAAAABFFAAFFFDFFF552EA8AAA55043DFF7AAAEAAB55F784",
INIT_3B => X"8002410FFD5575EF5555421E75555400BA082E8201000043FE005D517DEBA085",
INIT_3C => X"FAE975EF555168B55F7AA800BAF7AA955EF00002AAA2A2FBE8A00A2D16AAAAFF",
INIT_3D => X"0055554088A557FEB25D00021FFFFFFC00BA552A821EFFFFFD74BA5D51575F7F",
INIT_3E => X"000000000000000000000000000000000000000557DE00AAAAAAA000804001FF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024,               -- Port A enable input
WEA      => wbe_a_hi_1024(0),               -- Port A write enable input
DIA(0)   => data_write_a(5),        -- Port A data input
DOA(0)   => data_read_a_hi_1024(5),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024,               -- Port B enable input
WEB      => wbe_b_hi_1024(0),               -- Port B write enable input
DIB(0)   => data_write_b(5),        -- Port B data input
DOB(0)   => data_read_b_hi_1024(5),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_6_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10800B0061A01002840002C03002818000402322520070B313301C4389B2082",
INIT_01 => X"250041CA3839684D18A160000C52426841000000090800090210080008110200",
INIT_02 => X"0020042080010000044654C0000C008010000000001020900200200002620814",
INIT_03 => X"060881021088200021080200E4000A0891000020610111500104C00000F14400",
INIT_04 => X"0880000100000002000052288144004281C050400100280000C8100000080001",
INIT_05 => X"928080840001100A08009000280201000850E022401400002028214043410820",
INIT_06 => X"10100518090012122100C808049310002040000410A0001400000200120840D2",
INIT_07 => X"000100800004400001000000860408108C22000A502010074120044800040001",
INIT_08 => X"50000040D0C4E2088003FD01C01004044058082004000000000121F020408244",
INIT_09 => X"00BF17E9001205A5204911F814444080400100020000D200DFD16400C2A40AA0",
INIT_0A => X"04611C17849000022862A1596C8B5DF04834948900000100220C244840000880",
INIT_0B => X"03AD0413424E4044D665C070C22602291504400D084915020448114080201000",
INIT_0C => X"5E08864011088B22D22C008B0022C408B1022C208B0822C608B1111600458010",
INIT_0D => X"4251A12CD28A300429688001000800000020280204001000A00804309A002182",
INIT_0E => X"0000000280402400420800000000006200FC10002442042429324294014E8CA7",
INIT_0F => X"A40000000500800840000800000000000002280018001480000000A010100052",
INIT_10 => X"00000000000004C2003000010240000000000000680800290000000140202000",
INIT_11 => X"2000C0000000000000000442000001080001000000000000010C000280001804",
INIT_12 => X"08000000000801C300A010000000156000902000000015101200002800000000",
INIT_13 => X"000000000101800038002408000000094000386028040000000940000ED40000",
INIT_14 => X"0003B000002000000000020180002A24005010000000000023000060C7000A40",
INIT_15 => X"3F0280090321000040A410C28108000160008094000810040000000000002300",
INIT_16 => X"284A5284A728CA5284A528CA728CA52C4A5A0A32A300940101349A0408240818",
INIT_17 => X"9CA1294A329CA5284A728CA7284A5284A728CA5284A528CA728CA5284A728CA7",
INIT_18 => X"CA3294A129CA3294A129CA1294A329CA1294A3294A129CA3294A129CA3294A32",
INIT_19 => X"F5F78BCE7F8FF0F4FA955F7CF7F40A80145D55555556AAAAAAAAA94A329CA129",
INIT_1A => X"8E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E39B6CEDECDDF7DF7D",
INIT_1B => X"F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE38E3",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000001A1A33F9FCFE7F3F9FCFE7F3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"555FF00000000000000000000000000000000000000000000080000000000000",
INIT_28 => X"BC0010AAD5574BA557FFDFFF087BFDF45F7AA974AAAAAA97555F784174BAF7D5",
INIT_29 => X"515555508043FE00F7AA97555A2FBD7410AA8428AAAAAAE955450055421FFFFF",
INIT_2A => X"7D1575EFFFAA9555500557FE10FFFBEAA10007FD7410FFAA97400082A800AA08",
INIT_2B => X"0055574BA5D7FD7555A2D5575EF55517FF55A2AA97400552AAAB45082E80155F",
INIT_2C => X"500554200000003DE10FFD5401FFF7AAA8A10082EAAB45A2FFC2000007FD7400",
INIT_2D => X"10AA803FE105D516AABAFF843FFFFAA843DF55FFAA955EFA2D168B55557BEAB5",
INIT_2E => X"000AAAEBDF45A28428B45FFD168BFF00002AABA5D2ABFFFF087BD5545007BFDE",
INIT_2F => X"256DEB84104BAFFD1525FF000000000000000000000000000000000000000000",
INIT_30 => X"9756D145B401FFFFFFC7010BEDF524AA5571FDFEF1C7BFFF55FFA095482B6A49",
INIT_31 => X"4904380824850381C5B5057D1C003DE28F7A49057DAAF5D2428A2842AAAAA2AE",
INIT_32 => X"2AAFB451C2A8017DE3DF525FFFFA49756D145178E00EBFBE8A101475D5400F7A",
INIT_33 => X"2F1C50381471D74380851524BA5571D757DB6D5525EF555178F6DAAA49542841",
INIT_34 => X"AADB6FB7D5D7FEAB7D0855420BA1C0E3FE00E3DB471EFE3AAAAA00082EA8B6DA",
INIT_35 => X"F1C7BD057D1C71FFE10A28038E1049516AAB8FF8428FEFA28E3AF55F7A0925D7",
INIT_36 => X"00000000000000000000B6AEBDF45B68A28B6DEBDF6DBEF1C0A28AAA5524BFFF",
INIT_37 => X"F55F78017400F780001FFAA84000AAFFD1401E70000000000000000000000000",
INIT_38 => X"20BAAA8428AA2AAAA975FF5D7BC21EFF7FBD7400F7FBC00BA55557DFF7557BFD",
INIT_39 => X"EAA105D5155410FF84020AA0800154B2557FC01EF55043FEAAFF80021EFA2D14",
INIT_3A => X"568BE7AA80174AA082ABDF555D2A821EFAAFBC01FFF780155F7555568A00AAFF",
INIT_3B => X"AEA8A10082EA8BEFAAD5554B25551554BA0051400BA5551575EFF7D1401FF5D5",
INIT_3C => X"AAEAAB55F78400145AAFFFFFEF5D7FEABFF0051400A25D2EBFE10AAFFD55EFA2",
INIT_3D => X"552EA8AAA55043DFF7557BC01EF55557DE00AA842AA0000516AABAFF8428BE7A",
INIT_3E => X"0000000000000000000000000000000000000FFAABFF45FFAAAABFFAAFFFDFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024,               -- Port A enable input
WEA      => wbe_a_hi_1024(0),               -- Port A write enable input
DIA(0)   => data_write_a(6),        -- Port A data input
DOA(0)   => data_read_a_hi_1024(6),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024,               -- Port B enable input
WEB      => wbe_b_hi_1024(0),               -- Port B write enable input
DIB(0)   => data_write_b(6),        -- Port B data input
DOB(0)   => data_read_b_hi_1024(6),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_7_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10844B00482258A2842112C02450418800002300500030B313300C418992002",
INIT_01 => X"000009CA3839684D1CA0E0000E51424840000000080000080200080008510204",
INIT_02 => X"0120042086010000044600C00008000004100000000260900200000002402004",
INIT_03 => X"8628A10000082400000002408400080011000000610008000208C00000E14400",
INIT_04 => X"0911800100A000000000524084000040000050001140200100C8100000080102",
INIT_05 => X"0300812401011000000000002000114008008060441000000020024093000000",
INIT_06 => X"9190431C0D4010100000880804010010800000041080081000000200010424B2",
INIT_07 => X"000100AA0004408601000004860000008C02000A103010006928040800062481",
INIT_08 => X"84000048D484C20888000A0002120484C048007004000000000021F000000244",
INIT_09 => X"00A06009881201A520491004106C48A04040002400A15A208001650004001020",
INIT_0A => X"C99E1060201002044809C1040140A001004808810000459033189C0A400118A0",
INIT_0B => X"102000024040484050050041648A0041140C500B08821054C000264120000400",
INIT_0C => X"0404A083260E0832132011880462011880462051881462051881D31018C40620",
INIT_0D => X"0001000080001000813094801A8F80F00A600B52602801A88848011118003700",
INIT_0E => X"000003C007C002808228010410082042C000C000000004001002000400040002",
INIT_0F => X"A4000007800F80C840000800009864038A1200081C0014800000F001F0200052",
INIT_10 => X"00002C0E00E0E4004038000102400002C0E00E0D20100029000001E003E04000",
INIT_11 => X"2000C04031100E0403D0700300080908000100000661801E1900040380001804",
INIT_12 => X"0840878083E8003780A01043203A101780902043203A10082410082880000000",
INIT_13 => X"0601E0187900181035E0240806483248181035E0280410C8198818100DDD0000",
INIT_14 => X"0403774000201021E020FA006040376C00501022131210722060806D47000A40",
INIT_15 => X"00928A0002000110888600C032128201519480D40009902430160403E0E00506",
INIT_16 => X"01000000020080601802000000000405000A0020020081014134928820480010",
INIT_17 => X"0802018040000000006018020080200804010000000000806018020080000004",
INIT_18 => X"0000000001806008020000001006008020080001004008020080201004000020",
INIT_19 => X"0000000000000000000000000000400A004618618618C30C30C3000020180600",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000000B0840000000000000000000",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"1555500000000000000000000000000000000000000000000080000000000000",
INIT_28 => X"A97555F784174BAF7D5555FFF780155EFAAAEA8ABAAAFBFDE0055556AA005D04",
INIT_29 => X"55555EFAAFFFDFEFAAAAAAB455D556AA00FFAE95555087BFDF45F7AA974AAAAA",
INIT_2A => X"02EAAAAA082EA8A00AAAE955450055421FFFFFBC0010AAD5574BA557FFDFFF55",
INIT_2B => X"08043FE00F7AA97555A2FBD7410AA8428AAA557BFDFFF55003DFFFF7FBEAA000",
INIT_2C => X"0082A800AAF7AE975FFA28000010552EBDE00007BEAAAAA2D140000085155555",
INIT_2D => X"45087FEAB455D516AB55557BD55FF00557FE10FFFBEAA10007FD7410FFAA9740",
INIT_2E => X"000A2AA97400552AAAB45082E80155F7D1575EFFFAA955555D51574AAAAFFD55",
INIT_2F => X"AE105D556AA10410E17555000000000000000000000000000000000000000000",
INIT_30 => X"FFF55FFA095482B6A49256DEB84104BAFFD1525FFFF8E175C7A2AAAAA82A2F1F",
INIT_31 => X"F524AA5571FDFEF415B575D7AAF1FFFD7AAAAAFB7D495F6AA10E3AE905551C7B",
INIT_32 => X"003AFEFEBFBEAA001C2EA8A821C2EAAA00A2AE9756D145B401FFFFFFC7010BED",
INIT_33 => X"EDB470101C5B5057D1C003DE28F7A49057DAAF5D2428A2842AAAA497BFAFFF49",
INIT_34 => X"1475D5400F7A490438082485038F7A4905C7A28A070384120BDE100075EAA82B",
INIT_35 => X"D495150492BEF1D2555087BE8B7D555F6AB57417BC05D7145178E00EBFBE8A10",
INIT_36 => X"00000000000000000000AAA495428412AAFB451C2A8017DE3DF525FFFFA49756",
INIT_37 => X"555A2AEA8A10AAD568A00555168A10002E9754D0000000000000000000000000",
INIT_38 => X"8A10AAAE8215D557BFDF55F78017400F780001FFAA84000AAFFD1401E7FFAA97",
INIT_39 => X"C21EFF7FBD7400F7FBC00BA55557DFF7007BD5555AAD57DF55AAAEBDFEF007BE",
INIT_3A => X"428AA2007FE8BFF080028BFFAAFFEAA105D2EAAA005D2AAAA18AAAA975FF5D7B",
INIT_3B => X"043DE0000516AA10F7FBD7408557FC01EF55043FEAAFF80021EFA2D1420BAAA8",
INIT_3C => X"55568A00AAFFEAA105D5155410FF84020AA0800154B2FF8402145A2AA954AA00",
INIT_3D => X"AAFBC01FFF780155F7005140000FFD140145007FE8BEF557BEAB55087FC215D5",
INIT_3E => X"0000000000000000000000000000000000000AA80174AA082ABDF555D2A821EF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024,               -- Port A enable input
WEA      => wbe_a_hi_1024(0),               -- Port A write enable input
DIA(0)   => data_write_a(7),        -- Port A data input
DOA(0)   => data_read_a_hi_1024(7),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024,               -- Port B enable input
WEB      => wbe_b_hi_1024(0),               -- Port B write enable input
DIB(0)   => data_write_b(7),        -- Port B data input
DOB(0)   => data_read_b_hi_1024(7),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_8_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00000648E2840112C00000418000002700500030B3132000400812082",
INIT_01 => X"100008480009004C04A100000252024840000000180800080200010040110204",
INIT_02 => X"0020042000490000004600804008000005100000000024900200000002400004",
INIT_03 => X"0A0C33400008082400000080A4004B0891000020610112000040C00000E5C000",
INIT_04 => X"18800001000000000000512080000040800150400824280110C8100000120200",
INIT_05 => X"908084A10100100200004080280008240810802206940000012C214451610800",
INIT_06 => X"81B000080860109021400008040000202048020414A0021400040200322824C1",
INIT_07 => X"000000080004408049000004860000008402001A50208000630C040800062483",
INIT_08 => X"440000428644212280800A00021004044048002124000000000021F000000244",
INIT_09 => X"00004009001001010008100414644410400102228000D20080114502006409A2",
INIT_0A => X"000051312000042200294429148A4801C80C8C81000045907118040340020832",
INIT_0B => X"4020000240404140004D0544C4AA0001150410090302500011C813428A000400",
INIT_0C => X"46501090008820240240409000240009000240009000240009000120204808A5",
INIT_0D => X"42D1A168D09A301468402480004780F00140080860280004085904309A002196",
INIT_0E => X"00783FC00044340242280000000000020000C0000442106419120004034685A3",
INIT_0F => X"8000F07F800088A80000081EA2F9EC0000064004081010001E0FF00011104040",
INIT_10 => X"0ED0FC7E00000422201080000202658FC7E0000021882020003C1FE000222080",
INIT_11 => X"018059C3F350FE0C00000002A0040500000103961FE780000110010090000800",
INIT_12 => X"FD41FF80000830200021C1CF600012200010D1CF600012121600100810000004",
INIT_13 => X"9E1FE000010A1802100004343ED8000898021000087073D80008980200800002",
INIT_14 => X"0080200000BEB07FE00002086008020000209AEE3F300000246020200000620B",
INIT_15 => X"0088881903210000440610C8000A808040000208901786E4F0FE0C0000000166",
INIT_16 => X"685A1685A769DA368DA368DA769DA36CDA121A11A141800011309284002C0810",
INIT_17 => X"95A5685A1685A5695A368DA368DA769DA368DA368DA7695A1685A1685A5695A1",
INIT_18 => X"5A1695A568DA368DA369DA768DA1685A1695A5685A168DA369DA768DA368DA16",
INIT_19 => X"A4028A0A543EBC57A10A1E75D64108080468618618630C30C30C69DA5685A168",
INIT_1A => X"9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7BF3CCD8DF5B2DB2C",
INIT_1B => X"F87D3E1F4F87D3E1F4F87D3E1F4F87D3E1F4F87C3E1F0F87C3E1F0F87C3E79E7",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000006A6D4F87D3E1F4F87D3E1F4",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"155FF00000000000000000000000000000000000000000000080000000000000",
INIT_28 => X"BFDE0055556AA005D0415555080000000087BEAA10F7803DE00FFAEBFFFF0800",
INIT_29 => X"2AA8AAA557FC0010F780154105D7FC2145005155555F780155EFAAAEA8ABAAAF",
INIT_2A => X"7FFFFF55AA80155FF087BFDF45F7AA974AAAAAA97555F784174BAF7D5555FF55",
INIT_2B => X"AAFFFDFEFAAAAAAB455D556AA00FFAE95555AAFFE8A00552EBFE00F7D17FF45F",
INIT_2C => X"A557FFDFFF5504000AAAAAAA8B55F7D140010552E821EFAAAABDF555555555EF",
INIT_2D => X"55AA8028A00A2D57FF45557BE8A00AAAE955450055421FFFFFBC0010AAD5574B",
INIT_2E => X"000557BFDFFF55003DFFFF7FBEAA00002EAAAAA082EA8A00002AA8A10F784021",
INIT_2F => X"FE10F7AEBAFFF080A175D7000000000000000000000000000000000000000000",
INIT_30 => X"175C7A2AAAAA82A2F1FAE105D556AA10410E17555080E000280071E8A00EB8E3",
INIT_31 => X"4104BAFFD1525FF492EA8AAA5571C2000FF8A17400557FC015514555757DFF8E",
INIT_32 => X"2ABDE10EBDF7AF6DE3FFF8F7DB68A105D71C7BFFF55FFA095482B6A49256DEB8",
INIT_33 => X"AA0BDF6D415B575D7AAF1FFFD7AAAAAFB7D495F6AA10E3AE90555A2FBE8A3849",
INIT_34 => X"FFFFC7010BEDF524AA5571FDFEF550E00082B6A0AFB55F7D1420104124821D7A",
INIT_35 => X"01C2EA8A00F7800017DA2842FA00B6D578F6D557FFDA00A2AE9756D145B401FF",
INIT_36 => X"00000000000000000000497BFAFFF49003AFEFEBFBEAA001C2EA8A821C2EAAA0",
INIT_37 => X"0BA08556AA00AAAABFE00F7AEAABEF082E955450000000000000000000000000",
INIT_38 => X"21555D51575EFFFAA97555A2AEA8A10AAD568A00555168A10002E9754D082E82",
INIT_39 => X"17400F780001FFAA84000AAFFD1401E7082EAAABA5D5140010F7AE974105D7BC",
INIT_3A => X"E8215DA2FFE8ABA082ABFE00AAFBEABFFAAFBEABFFF7AA80145557BFDF55F780",
INIT_3B => X"D540000000402145AA843FFFF007BD5555AAD57DF55AAAEBDFEF007BE8A10AAA",
INIT_3C => X"AAA975FF5D7BC21EFF7FBD7400F7FBC00BA55557DFF75D2E82010F7843DF45FF",
INIT_3D => X"5D2EAAA005D2AAAA185D2AAAA10F780021FFA2803DE10FFD16ABFF5D7BFDE10A",
INIT_3E => X"0000000000000000000000000000000000000007FE8BFF080028BFFAAFFEAA10",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024,               -- Port A enable input
WEA      => wbe_a_hi_1024(1),               -- Port A write enable input
DIA(0)   => data_write_a(8),        -- Port A data input
DOA(0)   => data_read_a_hi_1024(8),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024,               -- Port B enable input
WEB      => wbe_b_hi_1024(1),               -- Port B write enable input
DIB(0)   => data_write_b(8),        -- Port B data input
DOB(0)   => data_read_b_hi_1024(8),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_9_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00018248A2840112C00002C18000002300500030B3132000400812006",
INIT_01 => X"400008000000004C0020000000100248413C0A61590001D90213C10008110204",
INIT_02 => X"01A0042080010000054600C04008000004100000001020900200200002420804",
INIT_03 => X"024003400008012400000010E4004B0891000020610310000144C00000F5C000",
INIT_04 => X"1801800100E000000000510084000040010050020810200000C8900000320200",
INIT_05 => X"918004311104100000000000200008100800002000100000002C234415610820",
INIT_06 => X"81B00008080010100000980804000008800042041080001000100200322C2481",
INIT_07 => X"0000811800044080010000058600000086020002502080006000040800062C80",
INIT_08 => X"0000004001D4618008800A00061004044048002004000000000061F000000244",
INIT_09 => X"000040090802009420409004104444084001022400214A2080014400026401A2",
INIT_0A => X"04000071200000A003CA294140200800C80C8C8100004590111C040040120800",
INIT_0B => X"12210002404848502847040164880021150400080222000200C8034200000000",
INIT_0C => X"4610088010080421021040841021000841021000841021000841010800420820",
INIT_0D => X"42D0A16C529A321068500484000500D10042080040284000084900001A002196",
INIT_0E => X"00000002804000004228010410082002C000C0002400046419120410034285A1",
INIT_0F => X"A00000000500800800000800000000000002290008001080000000A010100042",
INIT_10 => X"00000000000004C2001000000240000000000000680800280000000140202000",
INIT_11 => X"0000C0000000000000000442020001000001000000000000010C800080000804",
INIT_12 => X"08000000000801A7802010000000152780102000000015000600000800000000",
INIT_13 => X"000000000101900011E0240000000009500011E0280000000009500004DD0000",
INIT_14 => X"000137400020000000000201C000136C00101000000000002340002947000240",
INIT_15 => X"0080881901210000000600C280028000419480D4000010040000000000002304",
INIT_16 => X"68DA368DA1685A1685A1685A1685A16C5A121A13A141950051309284A82C0010",
INIT_17 => X"85A1685A1685A1685A368DA368DA368DA368DA368DA368DA368DA368DA368DA3",
INIT_18 => X"5A1685A168DA368DA368DA368DA368DA368DA368DA3685A1685A1685A1685A16",
INIT_19 => X"0157344CCCF48DE68A895C38E2540A8010100000000000000000685A1685A168",
INIT_1A => X"14514514514514514514514514514514514D34D34D34D34D28E1004039248209",
INIT_1B => X"D268341A4D268341A0D069349A0D069349A0D068341A0D068341A0D068345145",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000014D490D069349A0D068341A4",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"EAABA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"03DE00FFAEBFFFF0800155FFAAFBE8B45002A974AAAA803DFFFAA843DF45FFFF",
INIT_29 => X"7BFDE00A2FBD7400F7FBFDFFFA2AEBDE00AAFBEAABA080000000087BEAA10F78",
INIT_2A => X"055401FFF7AEAAA10F780155EFAAAEA8ABAAAFBFDE0055556AA005D041555508",
INIT_2B => X"557FC0010F780154105D7FC2145005155555557BE8BEF007FFDEAAAAD1555EF0",
INIT_2C => X"AF7D5555FFF780154AA5D2AA8A10F7AA974AA082E80010A2AAAAA10552AA8AAA",
INIT_2D => X"BAF7D17FEBAA2AEBDF45002EAAABA087BFDF45F7AA974AAAAAA97555F784174B",
INIT_2E => X"000AAFFE8A00552EBFE00F7D17FF45F7FFFFF55AA80155FF080400145FFFBEAA",
INIT_2F => X"8FC7BE8A3DF7DF7F5E8A92000000000000000000000000000000000000000000",
INIT_30 => X"000280071E8A00EB8E3FE10F7AEBAFFF080A175D7BEF1E8B6D002090482B68E3",
INIT_31 => X"56AA10410E175550871FFE00A2FBD0400FFF5FDFC7B6A0BDE38B6F5E8A92080E",
INIT_32 => X"7BFAE82A2DB555C71C5B451D7FFAAA8A38FF8E175C7A2AAAAA82A2F1FAE105D5",
INIT_33 => X"2AEADA38492EA8AAA5571C2000FF8A17400557FC015514555757D5D71E8BEF14",
INIT_34 => X"B6A49256DEB84104BAFFD1525FFFF84174BA5D20AAA00E3AA904BA142A87010A",
INIT_35 => X"7000400155FFFBEDA82FFD57DEBAAAA0BFF7D0024ADA921C7BFFF55FFA095482",
INIT_36 => X"00000000000000000000A2FBE8A38492ABDE10EBDF7AF6DE3FFF8F7DB68A105D",
INIT_37 => X"BEF080402000F7AAA8B55FFAABDFEFF7D16AA000000000000000000000000000",
INIT_38 => X"FEAAFFD16AA00082E820BA08556AA00AAAABFE00F7AEAABEF082E95545F7D568",
INIT_39 => X"A8A10AAD568A00555168A10002E9754D00517DE00A2FFC2000F7D17FF55FF803",
INIT_3A => X"1575EF555568BEF5D7FE8A10AAFFD55555D7FD5555FFAAA8AAAFFAA97555A2AE",
INIT_3B => X"AE800AA552A97400A2AEBDEAA082EAAABA5D5140010F7AE974105D7BC21555D5",
INIT_3C => X"57BFDF55F78017400F780001FFAA84000AAFFD1401E7FF80174AA5D0028A00AA",
INIT_3D => X"AAFBEABFFF7AA80145080002145F7FBFFE00FFD17FEAAA2803DFEF08043FE005",
INIT_3E => X"0000000000000000000000000000000000000A2FFE8ABA082ABFE00AAFBEABFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024,               -- Port A enable input
WEA      => wbe_a_hi_1024(1),               -- Port A write enable input
DIA(0)   => data_write_a(9),        -- Port A data input
DOA(0)   => data_read_a_hi_1024(9),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024,               -- Port B enable input
WEB      => wbe_b_hi_1024(1),               -- Port B write enable input
DIB(0)   => data_write_b(9),        -- Port B data input
DOB(0)   => data_read_b_hi_1024(9),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_10_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00018248A2840112C00002C18000202300500030B3132000400992006",
INIT_01 => X"254008000000004C002000000010026840000000080000080200010008110204",
INIT_02 => X"0020042000010000004455800008000004100000000000900200000002400004",
INIT_03 => X"020001021089000021081000C400090011000000610001540104C00000F14400",
INIT_04 => X"0811800101A00002000050088554004200C840000000200080C8100000000001",
INIT_05 => X"030080001000100800009400200000000840E020201000000024024001200020",
INIT_06 => X"81B00008080012120004CC080492500280208004148000100000020020042493",
INIT_07 => X"0000000800044080010000048404081085020002502000006000040800062480",
INIT_08 => X"100202400084410808000A00021004044048000004000000000021F020408264",
INIT_09 => X"010040090002008420401004144440004040022484214A2080110108C2C00320",
INIT_0A => X"04004166A48A0001080000000000080080181881000045901118044040020800",
INIT_0B => X"1201000200484910000F0105602622291404020902005002018002400A022000",
INIT_0C => X"0440001011808020120004801120044800120004801120044800110002400884",
INIT_0D => X"008000440210100041308480800F82F00040180260A808008848000018002104",
INIT_0E => X"000000028040000002280104100820020000400020000440100204100A000100",
INIT_0F => X"040000000500800800000000000000000002280008000400000000A010100010",
INIT_10 => X"00000000000004C2001000010000000000000000680800010000000140202000",
INIT_11 => X"200000000000000000000442000001000000000000000000010C000080001000",
INIT_12 => X"00000000000801C0008000000000154000800000000015000410000800000000",
INIT_13 => X"0000000001019800180000080000000958001800000400000009580002800000",
INIT_14 => X"0000A0000000000000000201E0000A0000400000000000002360002080000800",
INIT_15 => X"0080881000000000000600C28102800060000000000800000000000000002306",
INIT_16 => X"401004010040100401004010040100441020D0030008840051309A90BA884010",
INIT_17 => X"0902409024090240900401004010040100401004010040100401004010040100",
INIT_18 => X"1004010040902409024090240902409024090240902409024090240902409024",
INIT_19 => X"F546890A940FE0D3971243555205428290100000000000000000401004010040",
INIT_1A => X"8A28A28A28A28A28A28A28A28A28A28A28A28A28A28A28A29554199854514514",
INIT_1B => X"2B95CAE532994CA6532995CAE572B94CA6532994CA6532994CA6532994CA28A2",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000002718E72B94CA6532994CA657",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"FDE1000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"03DFFFAA843DF45FFFFEAABA007FC2155F7D155545AA80001EFAAFBEAB45557F",
INIT_29 => X"042AB55FFD168B55AA8000010FFFBE8BFFF78402155AAFBE8B45002A974AAAA8",
INIT_2A => X"AD16AABA002ABDE10080000000087BEAA10F7803DE00FFAEBFFFF0800155FF00",
INIT_2B => X"A2FBD7400F7FBFDFFFA2AEBDE00AAFBEAABAA2FFD741055003DFEFF7AA801FFA",
INIT_2C => X"05D0415555007FD74105555555EFF7FBC0145F78028A00A2D142155087BFDE00",
INIT_2D => X"55AAD168ABA002A975FFF7AEBDEBAF780155EFAAAEA8ABAAAFBFDE0055556AA0",
INIT_2E => X"000557BE8BEF007FFDEAAAAD1555EF0055401FFF7AEAAA105D042ABFF5D556AB",
INIT_2F => X"71D7AAFBEFB455D71F8E00000000000000000000000000000000000000000000",
INIT_30 => X"E8B6D002090482B68E38FC7BE8A3DF7DF7F5E8A92007BC217DEBDB55555AA8E0",
INIT_31 => X"EBAFFF080A175D700042AB7DEBDB6DB55BE8E05000EBFFE8BC7E38E07145BEF1",
INIT_32 => X"0A3DFD7F7A4821D7A2D16FA82142EB8E00080E000280071E8A00EB8E3FE10F7A",
INIT_33 => X"ED1421450871FFE00A2FBD0400FFF5FDFC7B6A0BDE38B6F5E8A92B6FBD541049",
INIT_34 => X"A2F1FAE105D556AA10410E175550071D54104951555D7EBF5C5155E3842AA00B",
INIT_35 => X"8410E2ABD749516FB55BED16FA820820955EFE3AEBDEAAFF8E175C7A2AAAAA82",
INIT_36 => X"000000000000000000005D71E8BEF147BFAE82A2DB555C71C5B451D7FFAAA8A3",
INIT_37 => X"1EFA2FFD7545AAAE97555A2FBFDF455D556AA000000000000000000000000000",
INIT_38 => X"8B45AAAA95545F7D568BEF080402000F7AAA8B55FFAABDFEFF7D16AA00087FC0",
INIT_39 => X"6AA00AAAABFE00F7AEAABEF082E9554500042ABFFA2FFFFF45F7AE97400AAFFE",
INIT_3A => X"16AA00FFFBD5400082EBFF45F78400155A2D57FE00552EA8A00082E820BA0855",
INIT_3B => X"D557555A2802AA10FFD54214500517DE00A2FFC2000F7D17FF55FF803FEAAFFD",
INIT_3C => X"FAA97555A2AEA8A10AAD568A00555168A10002E9754D085155410085557555AA",
INIT_3D => X"5D7FD5555FFAAA8AAA002AAAB4508557DF55F7D17FE000804155FFAAAABDEAAF",
INIT_3E => X"0000000000000000000000000000000000000555568BEF5D7FE8A10AAFFD5555",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024,               -- Port A enable input
WEA      => wbe_a_hi_1024(1),               -- Port A write enable input
DIA(0)   => data_write_a(10),        -- Port A data input
DOA(0)   => data_read_a_hi_1024(10),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024,               -- Port B enable input
WEB      => wbe_b_hi_1024(1),               -- Port B write enable input
DIB(0)   => data_write_b(10),        -- Port B data input
DOB(0)   => data_read_b_hi_1024(10),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_11_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"A101C4B05A0034CA2840712C2D001419000002300500030B31B20084EC992002",
INIT_01 => X"90000986B83028491800E0000C26426040000000080000088200080802512224",
INIT_02 => X"1A2004205E010640024D00800008000004100000040EC090820018003241A00C",
INIT_03 => X"28639100000C5C00000045C08400C8001100000061806A001618C03001E54400",
INIT_04 => X"1A800001000009A0804059A190000040400040008058220008C8100000120D4E",
INIT_05 => X"02000E81080250010000002022000058080400000E1200000020004401000004",
INIT_06 => X"819435143F20101010001008040800B8100102041088011100022200000024B2",
INIT_07 => X"90640D280884453E01064002944180008402001295BA100022E4340800062D82",
INIT_08 => X"400000093204802200280A0012160585C1D808D004000000000323F40C102244",
INIT_09 => X"380040098010001100009204107C5950400000220080C200800900020C006827",
INIT_0A => X"80007100004016EA080801010000080D00200081000045B0511D289940103399",
INIT_0B => X"002000024040410A000D0104408810C115D9C008050042400100D04E88000002",
INIT_0C => X"00655010009264201200C7B421ED0C7B421ED0C7B431ED087B43176843DA1085",
INIT_0D => X"0401020080400A10012494881A4F80F209500BB2602881A488485C1318002000",
INIT_0E => X"6619A540124814800228010410082022C00040002020090020220C9600040802",
INIT_0F => X"ACCC334A802491600C587949B6D0141B4CC600D5761B1599865A500490B86A56",
INIT_10 => X"BAC845542056A61686EC81E3A6CB68AA2C622C9A251C352B330CB4A0092170D8",
INIT_11 => X"BCCAD0B5A81536080CC6B21A21B1FC09CB0F1076D4A200B2AD4068F4101639B5",
INIT_12 => X"4D2CC281E31AA0103AB8D5514066380804B268A2E060901204112566F10AC418",
INIT_13 => X"D551443C47281002540B2C9AAAA8662A1152B202AE3554403028115AA88201A1",
INIT_14 => X"548A20A0492A2724A0621620402A020141F172FB182A32AB6845AB6200251BC9",
INIT_15 => X"00C00A000200074044E6801832728080D00A380B753952C4877E0104DDE4D124",
INIT_16 => X"0080200802008020080200802008020480080022020081010124988800400010",
INIT_17 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_18 => X"0000000000802008020080200802008020080200802008020080200802008020",
INIT_19 => X"55062608804180C0B10A42104201400204000000000000000000000000000000",
INIT_1A => X"00000000000000000000000000000000000820820820820801C4149470000000",
INIT_1B => X"0000000000000000040200000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000007E0F0000000000000100800",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"000AA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0001EFAAFBEAB45557FFDE10082ABDF5508557DF45002ABDFFFF7803DE10AA80",
INIT_29 => X"AEBFF45FFAEBFEAA002A801FFF7FFE8A10A28000000007FC2155F7D155545AA8",
INIT_2A => X"2AABFE10082ABFFEFAAFBE8B45002A974AAAA803DFFFAA843DF45FFFFEAABAA2",
INIT_2B => X"FFD168B55AA8000010FFFBE8BFFF78402155AAD155555A28428BFF002ABDE00A",
INIT_2C => X"F0800155FF00557FF45557FC2010002A80010A2842AAAA007BFFF4500042AB55",
INIT_2D => X"FF5D00154BAF7FBE8BEFFFD540000080000000087BEAA10F7803DE00FFAEBFFF",
INIT_2E => X"000A2FFD741055003DFEFF7AA801FFAAD16AABA002ABDE10A2D168A10A284021",
INIT_2F => X"DFC7F78E3FE28B684070AA000000000000000000000000000000000000000000",
INIT_30 => X"C217DEBDB55555AA8E071D7AAFBEFB455D71F8E00002EBDF6D005B78F7D142AB",
INIT_31 => X"A3DF7DF7F5E8A92BEAEBFF7DEBA0BDEAA1C2A801C7E3FFEFA10B68407038007B",
INIT_32 => X"8A28BFF082ABAE10B6AAB8E280820B8FEFBEF1E8B6D002090482B68E38FC7BE8",
INIT_33 => X"07FF8F7D00042AB7DEBDB6DB55BE8E05000EBFFE8BC7E38E07145B6D15756DA2",
INIT_34 => X"EB8E3FE10F7AEBAFFF080A175D708517DF7D497BC5028142A87000A28A2AA920",
INIT_35 => X"0B6DB6AA28A280001FF5D0A10482FFFFEFBC7E3DF42028080E000280071E8A00",
INIT_36 => X"00000000000000000000B6FBD5410490A3DFD7F7A4821D7A2D16FA82142EB8E0",
INIT_37 => X"FEF007BE8BFF5D2ABDF55F7AABDEAAF784154BA0000000000000000000000000",
INIT_38 => X"DE00FF84154BA087FC01EFA2FFD7545AAAE97555A2FBFDF455D556AA00082EBF",
INIT_39 => X"02000F7AAA8B55FFAABDFEFF7D16AA00FFAEBFFEFAA803DEBA5D2E82155A2FBF",
INIT_3A => X"A95545F7D5555FFAAAAA8BFF002AAAA00FFAAA8AAA080028BFFF7D568BEF0804",
INIT_3B => X"2E95400A2AEA8A00007FEABFF00042ABFFA2FFFFF45F7AE97400AAFFE8B45AAA",
INIT_3C => X"82E820BA08556AA00AAAABFE00F7AEAABEF082E9554508557DFFF007BD54BA5D",
INIT_3D => X"A2D57FE00552EA8A00FFFFE8AAAAA80001FF5D2E82000F7FFFFF45AAFFC20BA0",
INIT_3E => X"0000000000000000000000000000000000000FFFBD5400082EBFF45F78400155",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024,               -- Port A enable input
WEA      => wbe_a_hi_1024(1),               -- Port A write enable input
DIA(0)   => data_write_a(11),        -- Port A data input
DOA(0)   => data_read_a_hi_1024(11),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024,               -- Port B enable input
WEB      => wbe_b_hi_1024(1),               -- Port B write enable input
DIB(0)   => data_write_b(11),        -- Port B data input
DOB(0)   => data_read_b_hi_1024(11),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_12_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50080B01BC002006940202C0DE041196A83183000000023322287E0FC000006",
INIT_01 => X"75400D849830C84C5823E0000C17424840000000080000088200002802153231",
INIT_02 => X"18A026B43ED180040147558040090000061800000C06ED9802768F4472C52005",
INIT_03 => X"2A67E34A528D0524A52850528400C8001100000171C02B550618C91A10E55440",
INIT_04 => X"1BC0000100056C8280825DE98154004300C840800850240080CA921084520A07",
INIT_05 => X"02000F832000500C0000941024000852084060202E100001002000448100000C",
INIT_06 => X"819A1D1C3FE01A1A40045408049A50BA4020C6041090001200006200000000F2",
INIT_07 => X"C26A0719CC96CC6ED18A64019695A854870300FA3968B20068FC06080106249F",
INIT_08 => X"D002024B3E040800008C0A002610240D494A06F3460409000000E3F0AD5282E5",
INIT_09 => X"27A06009200040000400120412445D78400001000410420080218029CC807A27",
INIT_0A => X"18000006848A026F000000000000080000F010C100204593F11A6CDF48003BF8",
INIT_0B => X"000000820040402B28050400400432C9349DF21A31A00ACC0000F04F80020001",
INIT_0C => X"00357804611AE45D05D0833430CD0833420CD0C33420CD0833430668619A1000",
INIT_0D => X"0000000000000A74812DF00E87E80A079F9F90FA0280E87E800C7FF3B8002000",
INIT_0E => X"3B6B0E404D26160682082002000401EA0000C40000800A006002818808000000",
INIT_0F => X"A476D61C809A4DA84272592D6246FC1B17B541F97E1B348EDA93900B2B286C56",
INIT_10 => X"30C669E622DBC325CFD881A962454CFBE5403AB99594362B1DB52720165650D9",
INIT_11 => X"F8D2D39A3745261E4A95A110A3F855000E4B1D32BAB504BB7490FCFF912A3834",
INIT_12 => X"B90E9B018C7530200AB8F8BF41F9A22006B37DC8E1F9A21A70116D4C5080651C",
INIT_13 => X"118780319CCA08AB1001ACDF34B8F1C688AB1002AE3F7B807B6289F368828C4C",
INIT_14 => X"2AF020233376A5ECC016B1A827CDA21160F051DE610A34C50427E6E220323E4A",
INIT_15 => X"0077020000000439FDC05C5806781FAB46095A0B5199B0AC55521524F1864022",
INIT_16 => X"000000000000000000000000000000000026C000002884000130921092804010",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"8020080200000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0051B946088881360A95090CB054420290100000000000000000008020080200",
INIT_1A => X"041041041041041041041041041041041049249249249249200100002D451451",
INIT_1B => X"92C964B2592C964B2592C964B2592C964B2592C86432190C86432190C8641041",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000003800F592C964B2592C964B25",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"7DE1000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"ABDFFFF7803DE10AA80000AAAA843FE0008557DFFF0800020105D557FEAA0055",
INIT_29 => X"D5420000051555FFA2AA8200000557DFFFF7AA80000082ABDF5508557DF45002",
INIT_2A => X"82AA8AAAAAFFC00BA007FC2155F7D155545AA80001EFAAFBEAB45557FFDE10AA",
INIT_2B => X"FFAEBFEAA002A801FFF7FFE8A10A28000000A2D155410F7FFFFEBA08003FE000",
INIT_2C => X"5FFFFEAABA000028A105D2ABFE10A2AABFE1055516ABEF5D517DEAAA2AEBFF45",
INIT_2D => X"55002A820AA08557DFFFF7AA82155AAFBE8B45002A974AAAA803DFFFAA843DF4",
INIT_2E => X"000AAD155555A28428BFF002ABDE00A2AABFE10082ABFFEF0855420000004175",
INIT_2F => X"5010495B7AE921C517DE10000000000000000000000000000000000000000000",
INIT_30 => X"BDF6D005B78F7D142ABDFC7F78E3FE28B684070AABE803AE38145B78FD700000",
INIT_31 => X"BEFB455D71F8E00BED547038145B505FFB6A487000005F7AFD7F7A482038002E",
INIT_32 => X"F1FDE821C003FE001C2EAAAAAB6F5C2082007BC217DEBDB55555AA8E071D7AAF",
INIT_33 => X"D517DEAABEAEBFF7DEBA0BDEAA1C2A801C7E3FFEFA10B68407038B6D550428FF",
INIT_34 => X"B68E38FC7BE8A3DF7DF7F5E8A9200002FA285D20BDE28A2A4B8E10555B68BEF5",
INIT_35 => X"F085F47038140010555142082082005F7DFD7F7A482155BEF1E8B6D002090482",
INIT_36 => X"00000000000000000000B6D15756DA28A28BFF082ABAE10B6AAB8E280820B8FE",
INIT_37 => X"ABA5D7FEAB45080015410007FEAA0055517DE000000000000000000000000000",
INIT_38 => X"AB45F780020BA082EBFFEF007BE8BFF5D2ABDF55F7AABDEAAF784154BAF7802A",
INIT_39 => X"D7545AAAE97555A2FBFDF455D556AA00F7D1554BA5D7BC01FFFF8015410007FE",
INIT_3A => X"4154BAF7D1400BAFFD57FE005D043FE10552EAAAAAFFD140000087FC01EFA2FF",
INIT_3B => X"8428A105D7FEABEF55557DEBAFFAEBFFEFAA803DEBA5D2E82155A2FBFDE00FF8",
INIT_3C => X"7D568BEF080402000F7AAA8B55FFAABDFEFF7D16AA0008003FEBA55003DEBAA2",
INIT_3D => X"FFAAA8AAA080028BFF087BD54AA550402145550000010087FFFF45F78402145F",
INIT_3E => X"0000000000000000000000000000000000000F7D5555FFAAAAA8BFF002AAAA00",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024,               -- Port A enable input
WEA      => wbe_a_hi_1024(1),               -- Port A write enable input
DIA(0)   => data_write_a(12),        -- Port A data input
DOA(0)   => data_read_a_hi_1024(12),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024,               -- Port B enable input
WEB      => wbe_b_hi_1024(1),               -- Port B write enable input
DIB(0)   => data_write_b(12),        -- Port B data input
DOB(0)   => data_read_b_hi_1024(12),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_13_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10154A0441836CA2840512822007C18000E02700500030B31B300040081A042",
INIT_01 => X"00000804A000C04800020000000002404001000008220008A200100802110204",
INIT_02 => X"02200430000104000A4700804008000004100000000420918204D3033240400D",
INIT_03 => X"AA4003400008592400000590C40009141100000C6180C0000000C00001E14000",
INIT_04 => X"0800000102400120088054019000004160004190BAA0270000C8100000600206",
INIT_05 => X"21000012040610050040000227003AA0082400E94C1200000824424005220020",
INIT_06 => X"81963B180C001010580000080400000058000004109C00138000020024142581",
INIT_07 => X"002C8008000441600106400A9600010494020002B8AAA000EF003408000E2580",
INIT_08 => X"000000E48194408000A00A001210040441C80320040210000002ABF004102244",
INIT_09 => X"2A004009640040100400940412D4C4004000022000104200802D983000480120",
INIT_0A => X"8000202020401480000000000000080C90090881000145B0111A14004015080D",
INIT_0B => X"00000002004040AA08050400404040C11444000805200A402090024000008002",
INIT_0C => X"8410000A00280020020040800020040800020000801020000800010020400000",
INIT_0D => X"84A14250A055100050100490000500D00040080040290000084E4000B800610C",
INIT_0E => X"DCD13042BEDA36820228000000000000C000400081A08BC812A2092B02850942",
INIT_0F => X"89B9A260857DB400431969CA985D480949D32804A40AB137341C10B7D6A02EC0",
INIT_10 => X"E6ACA678001CE7D0296C213A460CA4271CA2168AEC1017606E6838216FAD4055",
INIT_11 => X"84AD4961C281B20213073C5FC0058008632D30D522CE80239DCC01AB013A4D20",
INIT_12 => X"2E6B13804A4B01D83461299900F6BD583A519104A0EEBD1A141010B2A4C8E116",
INIT_13 => X"89E5E40913419151EE0E94641828F72B5151EE0D184B321037AF5158BB02D085",
INIT_14 => X"562EC0B42162D68EE0073AE1C562EC13D521921A4170300B2B458B56B01C2280",
INIT_15 => X"00888A120240034000E6DC8285028014B82372011FC1E4F5E0A00929684EAF84",
INIT_16 => X"50942509425094250942509425094254940A1421420082020120908800480030",
INIT_17 => X"0942509425094250942509425094250942509425094250942509425094250942",
INIT_18 => X"9425094250942509425094250942509425094250942509425094250942509425",
INIT_19 => X"F7EFBBEEFF3F7DF7FF3E9F7DF7E2450228000000000000000000509425094250",
INIT_1A => X"BAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBF7DFDFDDD555555",
INIT_1B => X"EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAEBAE",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000000000F7EBF5FAFD7EBF5FAFD7",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"2ABEF00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0020105D557FEAA00557DE10AAD5554BA087FFFF55557BD54AAF7FBC01FFA280",
INIT_29 => X"7BD75EF087FFFFEF557BEAB45552E80155AA802AB45AA843FE0008557DFFF080",
INIT_2A => X"FAE820AA5D5557555082ABDF5508557DF45002ABDFFFF7803DE10AA80000AA08",
INIT_2B => X"0051555FFA2AA8200000557DFFFF7AA80000AAD1420AA087BD7555FFD168AAAF",
INIT_2C => X"5557FFDE10AAAEA8BFFA2FBD7545FFD157555085140010F7AEAABFFAAD542000",
INIT_2D => X"BA557BE8A10A284154BAFFAAAAB45007FC2155F7D155545AA80001EFAAFBEAB4",
INIT_2E => X"000A2D155410F7FFFFEBA08003FE00082AA8AAAAAFFC00BA00002AAAAF7D5574",
INIT_2F => X"0492E3F1C71C7BE8A2ABD7000000000000000000000000000000000000000000",
INIT_30 => X"3AE38145B78FD7000005010495B7AE921C517DE10A2DB50482147FFAF554971D",
INIT_31 => X"E3FE28B684070AA1C71D25D7007FFAFD7497BE8B5555208217DBE8A2AB45BE80",
INIT_32 => X"7FD257DFFD568A82FFA4870BA555F5056D002EBDF6D005B78F7D142ABDFC7F78",
INIT_33 => X"FAAAFBFFBED547038145B505FFB6A487000005F7AFD7F7A482038AADF4709214",
INIT_34 => X"AA8E071D7AAFBEFB455D71F8E00A2A0ADBC7A2FFD257DE3DF52555085142000F",
INIT_35 => X"21C002AA92FFDF574824171EAA10B680124BAFFAAAFB45007BC217DEBDB55555",
INIT_36 => X"00000000000000000000B6D550428FFF1FDE821C003FE001C2EAAAAAB6F5C208",
INIT_37 => X"0105D7BE8B55085142010AAD157545F7AEA8B550000000000000000000000000",
INIT_38 => X"01EFF7AAA8B55F7802AABA5D7FEAB45080015410007FEAA0055517DE00A2FFC0",
INIT_39 => X"E8BFF5D2ABDF55F7AABDEAAF784154BA5D5140145007BE8B55087BEAB555D040",
INIT_3A => X"0020BAA2FFD54105D7FC21EFFFD16AA10FF80174AA557FC21EF082EBFFEF007B",
INIT_3B => X"FBC0155085540000FFAEBFFEFF7D1554BA5D7BC01FFFF8015410007FEAB45F78",
INIT_3C => X"87FC01EFA2FFD7545AAAE97555A2FBFDF455D556AA00A2803FF45AAFFC21EFAA",
INIT_3D => X"552EAAAAAFFD1400005D042AA00F7FBD5410085568A10FF80020AAFFAABFF550",
INIT_3E => X"0000000000000000000000000000000000000F7D1400BAFFD57FE005D043FE10",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024,               -- Port A enable input
WEA      => wbe_a_hi_1024(1),               -- Port A write enable input
DIA(0)   => data_write_a(13),        -- Port A data input
DOA(0)   => data_read_a_hi_1024(13),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024,               -- Port B enable input
WEB      => wbe_b_hi_1024(1),               -- Port B write enable input
DIB(0)   => data_write_b(13),        -- Port B data input
DOB(0)   => data_read_b_hi_1024(13),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_14_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10020A000180000284008280000281800000030000000033022000000580002",
INIT_01 => X"000008020000204D006800000030824840000000084000084200090008510200",
INIT_02 => X"0220043170010A600A4D008040080000041000000028009002000F333240800C",
INIT_03 => X"111813400008002400000000C400090011000000610200001104D83000F14000",
INIT_04 => X"0801800100A000000000540084000040000040000800200000C8100000000748",
INIT_05 => X"0100000000001000000000002000080008000000001000000024024001200020",
INIT_06 => X"819EB84028001010000000080400000000000004108000100000020020040081",
INIT_07 => X"92040608000440100102400A94810206844200021DA2A0002000340800062C80",
INIT_08 => X"000000000084400008800A001214040441481500040000000000A7F408002244",
INIT_09 => X"0A0040090002008420401004104444004000020400214A208001000002400120",
INIT_0A => X"0400002020000000000000000000080C8008088100004590111B480040120000",
INIT_0B => X"1000000200404800000504016000002114000008020000020080024000000000",
INIT_0C => X"0410000010000000000040001000000000000040000000000001000000000000",
INIT_0D => X"04810244825010004010000000000000000000000000000000080000B8002104",
INIT_0E => X"0002C38280001202020800000000001000004000000000401022000002040902",
INIT_0F => X"20000587050001404E8084341CBA3404800828805200008000E0E0A000080002",
INIT_10 => X"4D18178E012010C00224004091C3514072C000444A0400080001C1C140001000",
INIT_11 => X"51709A07424142084458476001003809D0104B01C5710044020C4006010500C5",
INIT_12 => X"C26EE3803180C18006519462A00005001460E4730000050A1011004001060049",
INIT_13 => X"01F9E00660318000000538318740000140000001B4600CE80001400000002B62",
INIT_14 => X"0000000AD89857B0E0684411800000003799EB764D000330C300000000E3554B",
INIT_15 => X"0000021002002C000024008284001A0902000422E3F5960080480A0216A07240",
INIT_16 => X"4090240902409024090240902409024090081021020080015134920800480010",
INIT_17 => X"0902409024090240902409024090240902409024090240902409024090240902",
INIT_18 => X"9024090240902409024090240902409024090240902409024090240902409024",
INIT_19 => X"F5579B4E5C8FF0F7BE9D5F7DF650400200000000000000000000409024090240",
INIT_1A => X"9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7BF7DDDDDFCF3CF3D",
INIT_1B => X"F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE79E7",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000003FFF03F9FCFE7F3F9FCFE7F3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"420BA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"BD54AAF7FBC01FFA2802ABEFA2FBE8B55A2AE80000F7D5555555D2AAAABAAAD1",
INIT_29 => X"AA801FFA28402000AAAE955455500155EF0804155EFAAD5554BA087FFFF55557",
INIT_2A => X"7AEA8B45080417400AA843FE0008557DFFF0800020105D557FEAA00557DE10A2",
INIT_2B => X"087FFFFEF557BEAB45552E80155AA802AB4500516AA00A2AE800BAFFFFC20BAF",
INIT_2C => X"0AA80000AA005568ABAA28402010A2843FEBAFFFBD7410A2D168BFF087BD75EF",
INIT_2D => X"005D7FFDF4555517DFEF00043FEAA082ABDF5508557DF45002ABDFFFF7803DE1",
INIT_2E => X"000AAD1420AA087BD7555FFD168AAAFFAE820AA5D5557555002E80155A280000",
INIT_2F => X"0555412AA8ABAAADB40092000000000000000000000000000000000000000000",
INIT_30 => X"50482147FFAF554971D0492E3F1C71C7BE8A2ABD7A2FFEDB55B6A080038E3DB5",
INIT_31 => X"B7AE921C517DE10A2AE851FFB68402038AAAA955554900105FF0800175D7A2DB",
INIT_32 => X"A0800BAE3F1C0092EBAAADB6D080A12410BE803AE38145B78FD7000005010495",
INIT_33 => X"2D568BC71C71D25D7007FFAFD7497BE8B5555208217DBE8A2AB451C556FA00A2",
INIT_34 => X"142ABDFC7F78E3FE28B684070AA00516DABAA28402038B6803DE82F7F5D5410A",
INIT_35 => X"D002A80155B680000105D7FF8F455D5F78FD7000E3FEAA002EBDF6D005B78F7D",
INIT_36 => X"00000000000000000000AADF47092147FD257DFFD568A82FFA4870BA555F5056",
INIT_37 => X"F55FF84000AAAAFBC0145002AA8AAAAAFFC20000000000000000000000000000",
INIT_38 => X"01EF080417555A2FFC00105D7BE8B55085142010AAD157545F7AEA8B55A2FBFF",
INIT_39 => X"EAB45080015410007FEAA0055517DE00A2AA955FFFF80020BAAAAA9754508000",
INIT_3A => X"AA8B555D557FE00A280020BAAAD140000A2AEBFFEF082A82010F7802AABA5D7F",
INIT_3B => X"803DE00FFD557400AAD56AB455D5140145007BE8B55087BEAB555D04001EFF7A",
INIT_3C => X"82EBFFEF007BE8BFF5D2ABDF55F7AABDEAAF784154BA08557FEAAA284000AAFF",
INIT_3D => X"FF80174AA557FC21EF082A80145F780020105D7BEAB45557BE8B45082EBFEBA0",
INIT_3E => X"0000000000000000000000000000000000000A2FFD54105D7FC21EFFFD16AA10",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024,               -- Port A enable input
WEA      => wbe_a_hi_1024(1),               -- Port A write enable input
DIA(0)   => data_write_a(14),        -- Port A data input
DOA(0)   => data_read_a_hi_1024(14),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024,               -- Port B enable input
WEB      => wbe_b_hi_1024(1),               -- Port B write enable input
DIB(0)   => data_write_b(14),        -- Port B data input
DOB(0)   => data_read_b_hi_1024(14),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_15_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000A000000000284000280000001800020030000000033022000000180002",
INIT_01 => X"8000080000000048000000000000026040000000080000080200000000110200",
INIT_02 => X"0020042004010E60004C0080000800000410000000020090020000300245E005",
INIT_03 => X"0000010000080400000000408400480111000000610008000000C00000E54400",
INIT_04 => X"980000010000000088C2550080000040000040000008A00028C8100000120000",
INIT_05 => X"020004012E025000000001322000000A28008000011000000220004D41000000",
INIT_06 => X"819588000800101000011008040000100001060418800510000A620000000092",
INIT_07 => X"0000000800044004010C20008440810284020002102220002000340800062480",
INIT_08 => X"0000000001140800002C0A001214050540C800400406180000002DF004000244",
INIT_09 => X"1E00400900000000000016041044400440000000000042008001000000000022",
INIT_0A => X"0000000000000220000000000000080C00000081000045901118000040000000",
INIT_0B => X"0000000200404000010500004000000114000009000000000000004200000000",
INIT_0C => X"0000000000000000000040001000040001000000000000000001000020000800",
INIT_0D => X"000000000000001001208000180800000000030200000180800C400030002000",
INIT_0E => X"0000000000002600020800000000001080004000000000000002000000000000",
INIT_0F => X"A400000000000000000008000000000000000000000014800000000000000052",
INIT_10 => X"0000000000000000000000010240000000000000000000290000000000000000",
INIT_11 => X"2001C05838120800000000000000000000010000000000000000000000001804",
INIT_12 => X"081004000000000000A010000000000000902000000000180010002020000000",
INIT_13 => X"6600000000000000000024080000000000000000280400000000000000000000",
INIT_14 => X"0000000000200801000000000000000000501001920000000000000000000A40",
INIT_15 => X"0000020000000000000000003000000000000000000A101C3614000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000080000120980000000010",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000400200000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"28BEF00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"5555555D2AAAABAAAD1420BAFF8000010082A954BA00003DFEF085155400F784",
INIT_29 => X"AE95555A2FBE8BEFA2843DE00AA8015400FF84001EFA2FBE8B55A2AE80000F7D",
INIT_2A => X"2FBEAB45F7D56AABAAAD5554BA087FFFF55557BD54AAF7FBC01FFA2802ABEFF7",
INIT_2B => X"A28402000AAAE955455500155EF0804155EFFFFBE8BFF0800174AA557BFDE10A",
INIT_2C => X"A00557DE10F7D1574AAA2D16AB55FFD568BEF087FE8A1055003FE00A2AA801FF",
INIT_2D => X"00AA802AA00AAAE800BA5D0015545AA843FE0008557DFFF0800020105D557FEA",
INIT_2E => X"00000516AA00A2AE800BAFFFFC20BAF7AEA8B45080417400FFFFC21450800154",
INIT_2F => X"8FD7005150438F78A2DBFF000000000000000000000000000000000000000000",
INIT_30 => X"EDB55B6A080038E3DB50555412AA8ABAAADB40092E38E070280024904AA1C043",
INIT_31 => X"1C71C7BE8A2ABD7E3AA9257DA2FFE8BC7BE8E38E10A28017400E38A051FFA2FF",
INIT_32 => X"00124AA557FFDE10A2FBEDB6DF7D16AABAA2DB50482147FFAF554971D0492E3F",
INIT_33 => X"10038E38A2AE851FFB68402038AAAA955554900105FF0800175D7E3FFEFBD700",
INIT_34 => X"000005010495B7AE921C517DE10FFDF50482A2DB6AB45FFD56DBD7087BEAA384",
INIT_35 => X"0FFF1C017D140410400BE8E28A10AAA085082550A1057DBE803AE38145B78FD7",
INIT_36 => X"000000000000000000001C556FA00A2A0800BAE3F1C0092EBAAADB6D080A1241",
INIT_37 => X"4AA0800020BA550028B550855400AAF7AEBDFEF0000000000000000000000000",
INIT_38 => X"7400AAAE975EFA2FBFFF55FF84000AAAAFBC0145002AA8AAAAAFFC2000AAAA97",
INIT_39 => X"E8B55085142010AAD157545F7AEA8B55AAAE821EFAAFBEAB55F7AAA8A00AA841",
INIT_3A => X"417555AAFFFDF450804020AA557BFFE10A2FFFFFEFF7D568ABAA2FFC00105D7B",
INIT_3B => X"D17DF45007FE8AAA08002AAAAA2AA955FFFF80020BAAAAA975450800001EF080",
INIT_3C => X"7802AABA5D7FEAB45080015410007FEAA0055517DE00FFFBC2000AAFBE8B55F7",
INIT_3D => X"A2AEBFFEF082A82010FFD5421EF5D0000010F7AAA8A10AA8017400552A801EFF",
INIT_3E => X"00000000000000000000000000000000000005D557FE00A280020BAAAD140000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024,               -- Port A enable input
WEA      => wbe_a_hi_1024(1),               -- Port A write enable input
DIA(0)   => data_write_a(15),        -- Port A data input
DOA(0)   => data_read_a_hi_1024(15),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024,               -- Port B enable input
WEB      => wbe_b_hi_1024(1),               -- Port B write enable input
DIB(0)   => data_write_b(15),        -- Port B data input
DOB(0)   => data_read_b_hi_1024(15),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_16_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"DA22C618B1000482B688B186588884862A400438255FC38381441205BA803003",
INIT_01 => X"7045A80028404C211203A952A90341080B173340412000E1005D628000820484",
INIT_02 => X"428406A4000850848330118D0AAC55001349B108818005460229044001C01784",
INIT_03 => X"092C4020000500020000500986812C405000001A48202050000A214AC0650115",
INIT_04 => X"4804A55440256F504025E003A054F46415A4E62B6FE3307943965A00001A1152",
INIT_05 => X"0000001C40A5B950ADB8EA097057ECE14C86D2B7F85AAD17F4B100000B88148C",
INIT_06 => X"415401DCDCF2C0A8030140BCB0820A200342A1C641C1E8782F508F2B00003584",
INIT_07 => X"002701881A3202080AE00480A2002840BE1480FA004342AA6F12000054004867",
INIT_08 => X"08C54828091002000002B32A8C19064E486A8001510000014140C1E2A14891E0",
INIT_09 => X"015452B103020814004088B64102680B6596594800400413CAC0208944800000",
INIT_0A => X"96AA000484094C000000000000012C9000A0000D0A80000BF8028E87C1B99270",
INIT_0B => X"014808A02004200E540480212000A448C0082024AE50064B44000000000002A2",
INIT_0C => X"0004000D5846256AAEA811150445411150445411150445411150422A088A8200",
INIT_0D => X"00000004010042A204A0C5817D00005034052E40000817D00440004004AD3240",
INIT_0E => X"632B2673FA4587978A2004102800809225545155121740000004900090000000",
INIT_0F => X"00C6564CE7F4EA4B940076D296D003030800462CBD320018CAAAACFE9164C800",
INIT_10 => X"28834ADB1440A114793A4A30A40839AA14910D08DCB2640031955559FD3AC990",
INIT_11 => X"594AB0B1A025371CA0E034E8443C097A800EB090D4AAC91208ED2FA0CE5E09B1",
INIT_12 => X"7B50446083001B94BB38C540EBE61284BB304880E3E4579EDC00992980D58033",
INIT_13 => X"5511121840E7A2CD952ECC12ABC3E6ACB3DFB12ECE315000F61FF1727A85FDBC",
INIT_14 => X"75DEB07F6F2E7084517F126F8395CB2BEFBAB8BA8AF698228CC5E2F08ECA5159",
INIT_15 => X"5580A840A8009F8B108C80A1021B080AFC0DF6422C6077F4A77F20D0C0E21084",
INIT_16 => X"0000000000000000000000000000000000044000102A0001148442A110810359",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"558D11544C690DA64C1C4F68A360400000000000000000000000000000000000",
INIT_1A => X"14D14D14D14D14D14D14D14D14D14D14D14514514514514529E5F87869E79E78",
INIT_1B => X"D1E8F47A3D1E8F47A7D3E9F4FA7D3E9F4FA7D3E9F47A7D1E9F47A7D1E9F4D14D",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000007D3E9F4FA7D3E8F47A3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"C00AA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"03DFEF085155400F78428BEF087FFFFEFF7D168B55AAD17FFFF552EBFE00007F",
INIT_29 => X"2E975EFF7D568BFFFF80175EF0004000BA552A821FFFF8000010082A954BA000",
INIT_2A => X"55540000082EAABFFA2FBE8B55A2AE80000F7D5555555D2AAAABAAAD1420BA5D",
INIT_2B => X"A2FBE8BEFA2843DE00AA8015400FF84001EF0000020AA5D00154005D043FF455",
INIT_2C => X"FA2802ABEF557BEABEF5D0415410087FD74BAAAAEBFFEF557FC00AAF7AE95555",
INIT_2D => X"FFFFAABFEAAFF84001FF002A821FFAAD5554BA087FFFF55557BD54AAF7FBC01F",
INIT_2E => X"000FFFBE8BFF0800174AA557BFDE10A2FBEAB45F7D56AABA082A97545F7D16AB",
INIT_2F => X"FFEF552AB8E38087FC2092000000000000000000000000000000000000000000",
INIT_30 => X"070280024904AA1C0438FD7005150438F78A2DBFF0871F8FC7E3D56AB6DBEDB7",
INIT_31 => X"AA8ABAAADB400924920925EFF7D16ABFFE38E175EF1400000BA412E871FFE38E",
INIT_32 => X"0A1240055003FF6D5551420101C2EAFBD7A2FFEDB55B6A080038E3DB50555412",
INIT_33 => X"57FC00BAE3AA9257DA2FFE8BC7BE8E38E10A28017400E38A051FF0804050BA41",
INIT_34 => X"4971D0492E3F1C71C7BE8A2ABD74975EDBC7550E12410087FD74AAB6AABFFC75",
INIT_35 => X"A08249756DF7D168BC7F7AABAEAAF780051C70824851D7A2DB50482147FFAF55",
INIT_36 => X"00000000000000000000E3FFEFBD70000124AA557FFDE10A2FBEDB6DF7D16AAB",
INIT_37 => X"B55A2D16ABEFFFFBFDFFF552AAAAAA007BC00000000000000000000000000000",
INIT_38 => X"20AA002A955EFAAAA974AA0800020BA550028B550855400AAF7AEBDFEF08516A",
INIT_39 => X"000AAAAFBC0145002AA8AAAAAFFC20000000021EFF7D568BFFA2AA955FF5D040",
INIT_3A => X"E975EF0800174BA002E820105D003DFEF5D51420005D2ABFF45A2FBFFF55FF84",
INIT_3B => X"7BD74AAF7AEBDF455D7BC20BAAAAE821EFAAFBEAB55F7AAA8A00AA8417400AAA",
INIT_3C => X"2FFC00105D7BE8B55085142010AAD157545F7AEA8B5500557DF45552A8200000",
INIT_3D => X"A2FFFFFEFF7D568ABA0804155FFF7D568B55FFAAAAABAFF8415545000015555A",
INIT_3E => X"0000000000000000000000000000000000000AAFFFDF450804020AA557BFFE10",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024,               -- Port A enable input
WEA      => wbe_a_hi_1024(2),               -- Port A write enable input
DIA(0)   => data_write_a(16),        -- Port A data input
DOA(0)   => data_read_a_hi_1024(16),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024,               -- Port B enable input
WEB      => wbe_b_hi_1024(2),               -- Port B write enable input
DIB(0)   => data_write_b(16),        -- Port B data input
DOB(0)   => data_read_b_hi_1024(16),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_17_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"5284CE4FB7BD2C8994A13392DBD02E14006B82AC7E800D44D3DD2FD5F9B961C0",
INIT_01 => X"2EACD01F7E03FC6793F2199B39FC233C11D93AE6F3BB92B32091DBC339B24542",
INIT_02 => X"E63CCCC00A82C08092A2AFAE667033DB50853379C10BFDC5C6F4044443C817C6",
INIT_03 => X"7FF183635AEF9E3635AEF9E18E237040404446965C0607EE6DB7854AC4DE060C",
INIT_04 => X"D78AC33FB604488B000892EF17BE6D84196482236FE100294152E294350FB697",
INIT_05 => X"081B5F9B409420D0CDB47A05403F6CE0C08A4AB7F840EDB6F48100DFC8081081",
INIT_06 => X"768465354781CBC30316367077B4BDB50646E8D87100A8201ED01C19C020F71A",
INIT_07 => X"4002A110C922480A82D0841147162C48EBB9537A0022DC67987042EE976ABEA7",
INIT_08 => X"DB931BFEF91C00002CC0E019C0C82A4E4820C15A2330E004401891181168C4D1",
INIT_09 => X"09F3A1BC11EFBC66DB65307071477FF1030C397C060B4254064302042F803A69",
INIT_0A => X"3F330802162F3B7EE3F3EC7C7DEF207000F00059D2ED56D7EED2ED3C9A867DC0",
INIT_0B => X"185C44B91BC1740B7605040BE0018CFC7429F326B9E822FFC00074D5A0AB033A",
INIT_0C => X"00367A28FC1B7F7FEFFCFBFF3EFFCFBFF3EFFCFBFF3EFFCFBFF3EFFE7DFF9E00",
INIT_0D => X"0000000008004BA78428C7AD7FC94B533F5B4FFBD2FAD7FCCA786D43FE67C218",
INIT_0E => X"BA494CEBFD4F2667ABB6F68B29760593F33FA0CF170F40006001B1A05C000000",
INIT_0F => X"7F749299D7FAEB237DFE5865B6D2BF23265CBACE542A6FEE92333AFF33E0A9BF",
INIT_10 => X"F6C24B6D18C3C9F8E2881F3F787D776B5DB94A09955054DFDD246675FE7AC153",
INIT_11 => X"BFB349E08FF9A27EDE9FA8AEFD9E7467BFCB195CFEB56A1A70D34D1706FFFA3E",
INIT_12 => X"6FE219CA80725B875EED723FF7FCB2875EDAAFEAF7FD929BFD55BBC71D79F639",
INIT_13 => X"546670D018E7A6E581D7B6AB75FDFCECA6E581D7BB5DDFC6FF0EB7D7E859FDB5",
INIT_14 => X"B978177F6D6AF5ECDB5FB76A5F5FA165B456E0FB308710C49FCFB741598B9C7E",
INIT_15 => X"CFDAAB00AC00A8BBFC8B501CF7A0FED9A540EA1952586CEB54D143ACFF9A3BA9",
INIT_16 => X"000000000000000000000000000000000026E100002F382DBD9ECFE117805F20",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"4372003009EDCC4052E917114F981800C0000000000000000000000000000000",
INIT_1A => X"BA69A69AEBA69AEBA69A69AEBA69AEBA69A69A69A69A69A68698686981D75D74",
INIT_1B => X"6A351A8D46A351A8D068341A0D068341A0D068341A0D46A341A0D46A341A69AE",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000000000046A351A8D46A351A8D4",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"7FEAA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"17FFFF552EBFE00007FC00AA087FFFFFFFFFFFFFEFF7FBEAB450804001EFAAD5",
INIT_29 => X"D168A000004020AA5D7BE8B450051401EF087FD74AA087FFFFEFF7D168B55AAD",
INIT_2A => X"D7FEAB55FF80175EFFF8000010082A954BA00003DFEF085155400F78428BEFAA",
INIT_2B => X"F7D568BFFFF80175EF0004000BA552A821FF5D00020BA552A82000552A821555",
INIT_2C => X"AAAD1420BAFFFFFDF45AAD17FFFFAAFBC01EF5D0015555557BFDEBA5D2E975EF",
INIT_2D => X"BA007FEABEF005555555A2D1554BAA2FBE8B55A2AE80000F7D5555555D2AAAAB",
INIT_2E => X"0000000020AA5D00154005D043FF45555540000082EAABFF00516AA10552E820",
INIT_2F => X"8B550000071EFB6DF7AE92000000000000000000000000000000000000000000",
INIT_30 => X"F8FC7E3D56AB6DBEDB7FFEF552AB8E38087FC2092147FFFFFFFFFBFDFC7EBF5E",
INIT_31 => X"150438F78A2DBFFBED16AA381C0A07082497FEFB6D1451471EF007BD04920871",
INIT_32 => X"2A850105D2A80155417BEFB6DEB8E175FFE38E070280024904AA1C0438FD7005",
INIT_33 => X"D7BFAEBA4920925EFF7D16ABFFE38E175EF1400000BA412E871FF550A0009249",
INIT_34 => X"E3DB50555412AA8ABAAADB40092FFF5FFF6DAADF7FFD7B6F1C71EF55001756D5",
INIT_35 => X"7145B6AA28492487082007FEDBD700515556DA2DF50492A2FFEDB55B6A080038",
INIT_36 => X"000000000000000000000804050BA410A1240055003FF6D5551420101C2EAFBD",
INIT_37 => X"FEFF7FBFFF55A2D16AB550000175EFFFFBEAA000000000000000000000000000",
INIT_38 => X"55EF087FC200008516AB55A2D16ABEFFFFBFDFFF552AAAAAA007BC0000557FFD",
INIT_39 => X"020BA550028B550855400AAF7AEBDFEFF7D568AAA5D2A97410007BFFFFF55515",
INIT_3A => X"A955EF5D2E80010002A954005D2A82155087FFFFEFAAAA975EFAAAA974AA0800",
INIT_3B => X"D1575FF5504175EF5D7FEAAAA0000021EFF7D568BFFA2AA955FF5D04020AA002",
INIT_3C => X"2FBFFF55FF84000AAAAFBC0145002AA8AAAAAFFC2000FFD57DFFFAAFFFDF55FF",
INIT_3D => X"5D51420005D2ABFF45557FE8AAA000415410007BFFF450051555EFA2FBC0000A",
INIT_3E => X"00000000000000000000000000000000000000800174BA002E820105D003DFEF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024,               -- Port A enable input
WEA      => wbe_a_hi_1024(2),               -- Port A write enable input
DIA(0)   => data_write_a(17),        -- Port A data input
DOA(0)   => data_read_a_hi_1024(17),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024,               -- Port B enable input
WEB      => wbe_b_hi_1024(2),               -- Port B write enable input
DIB(0)   => data_write_b(17),        -- Port B data input
DOB(0)   => data_read_b_hi_1024(17),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_18_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"69844019080000A21A611406840014122A641074155FC28A2024001001801003",
INIT_01 => X"7443D920034004180005E9E3C90360C0041C0181002001602025800008440084",
INIT_02 => X"E2DCCCE61D5C008103F2000781FC0FEDEAC2161B0B8FB0008620044443006010",
INIT_03 => X"884E300802006900802006995C896D605200000856E24A040000640052141103",
INIT_04 => X"480520FC026125AC0025C9122644E3E40EC8E2001001302281841A009038A86A",
INIT_05 => X"432000040089983070019400F01010004C8DB841405A80A100B586200FAC24AE",
INIT_06 => X"09044359DC7040000000002C109B0E0A00A1104641C0803804000707284600E1",
INIT_07 => X"400D10100400481D5EB08501620000007500CE801241021FE78E404860140060",
INIT_08 => X"00880C0106A0528020019307CC082A0A4A6A01ED725021400040D028000A9729",
INIT_09 => X"00117063038000282081402E4106400B6186128040600C10C1C0200950508110",
INIT_0A => X"C0C30C2E21580C874004008080003C32A10A19090C02010E1022944061688000",
INIT_0B => X"0180A8062026000DC425C0301311324AA2373088479105D044A1022000001835",
INIT_0C => X"0D89844703649000000200000000000000000000000000000000000000000010",
INIT_0D => X"0D8306C182701404C1973010802020404084001E00010802046092B5001FB365",
INIT_0E => X"528EB314068AB8B803DB00002900800400FC503F08180050942E4200020C1B06",
INIT_0F => X"40A51D66280D6032C5F96D3C51555D5D7D5AA87285820814A3CCC501C2A60820",
INIT_10 => X"8B35A3FEBF1FEDFD9C2B30E0468AAAD5D48F37E8FC1304102947998A03984C10",
INIT_11 => X"440FE1DD772D37A0A321BC6968F32658BF2D4F2A80BF8FE3F9FE3AC362080529",
INIT_12 => X"5487910D7E5A6D961A28456A1832E5161A100DD5182BC54020EA67A189C6ED36",
INIT_13 => X"AA444CAF91EDD1B725868403BE06323551B725868A100ABD119753B70964122B",
INIT_14 => X"EDC259048ACD868EE3803D65CEDC258A8F80D55E007C3F8EBB56F4C5362C978F",
INIT_15 => X"3F240014BE84370001B6922070440556B15F7FABBC0031BCF2257C41634B14D4",
INIT_16 => X"C1B06C1B06C1B06C1B06C1B06C1B06C1B0491069068000004060300A005A0118",
INIT_17 => X"1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06",
INIT_18 => X"B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C",
INIT_19 => X"B28BBECEB80EE173C2300F7DF16000000000000000000000000041B06C1B06C1",
INIT_1A => X"8A28A28AAAAAAA28A28A28AAAAAAA28A28A28A28A28A28A2910591505C104104",
INIT_1B => X"28944A25128944A25128944A25128944A25128944A2552A954AA5128944AAAA2",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000128944A25128944A251",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"9540000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"BEAB450804001EFAAD57FEAA087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974BA082E",
INIT_29 => X"7FFFFFFFFFBFDF45AAD568B55080028B55002E82000087FFFFFFFFFFFFFEFF7F",
INIT_2A => X"0043DE10AA843DE00087FFFFEFF7D168B55AAD17FFFF552EBFE00007FC00AA08",
INIT_2B => X"0004020AA5D7BE8B450051401EF087FD74AAAAFFFDF45A2D16AB55F7FFFFFFF0",
INIT_2C => X"0F78428BEFAA80000000804154BA55042ABEF5D7FD75FFAAD540145AAD168A00",
INIT_2D => X"00082E95555085168A10557FD7545FF8000010082A954BA00003DFEF08515540",
INIT_2E => X"0005D00020BA552A82000552A821555D7FEAB55FF80175EF5D00020105D2A974",
INIT_2F => X"DFFF5D2A954AA082A92428000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFBFDFC7EBF5E8B550000071EFB6DF7AE921C7FFFFFFFFFFFFFFFF7FBF",
INIT_31 => X"AB8E38087FC2092087FFDFC7E3F1FAF55A2DF6DB7D1C002AB7D002A82028147F",
INIT_32 => X"DF6DB7DE3F5FAFC708003DE28B68E38E280871F8FC7E3D56AB6DBEDB7FFEF552",
INIT_33 => X"ADF4516DBED16AA381C0A07082497FEFB6D1451471EF007BD0492B6F1F8F55AA",
INIT_34 => X"1C0438FD7005150438F78A2DBFFA28407038140410492550A2ABC7497BD25FFA",
INIT_35 => X"F5D0E05000492097428002E9557D1C516FA28417BD5545E38E070280024904AA",
INIT_36 => X"00000000000000000000550A00092492A850105D2A80155417BEFB6DEB8E175F",
INIT_37 => X"FFFFFFFFDFEFF7FBFFFEF552E974AA082A820AA0000000000000000000000000",
INIT_38 => X"ABEF002A800AA557FFDFEFF7FBFFF55A2D16AB550000175EFFFFBEAA00557FFF",
INIT_39 => X"6ABEFFFFBFDFFF552AAAAAA007BC0000087BFDF45AAD568B55AAFBFDFEF55042",
INIT_3A => X"FC2000FFD56AB45A2FFFDFFFAAD16AB4500043DEAAFFAEAAAAA08516AB55A2D1",
INIT_3B => X"2AA8B45087FC01EFA2FFD55EFF7D568AAA5D2A97410007BFFFFF5551555EF087",
INIT_3C => X"AAA974AA0800020BA550028B550855400AAF7AEBDFEFA280154BA55040000055",
INIT_3D => X"087FFFFEFAAAA975EF5D2E974000804154BA082A975EF5D517DEAA007BD5545A",
INIT_3E => X"00000000000000000000000000000000000005D2E80010002A954005D2A82155",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024,               -- Port A enable input
WEA      => wbe_a_hi_1024(2),               -- Port A write enable input
DIA(0)   => data_write_a(18),        -- Port A data input
DOA(0)   => data_read_a_hi_1024(18),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024,               -- Port B enable input
WEB      => wbe_b_hi_1024(2),               -- Port B write enable input
DIB(0)   => data_write_b(18),        -- Port B data input
DOB(0)   => data_read_b_hi_1024(18),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_19_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"042200000000000041088001001AA00000000000000000000000500802000003",
INIT_01 => X"040048000024000000000404000000000A22000800000800004A200000000001",
INIT_02 => X"200C8840085EB00480060000001C008002489E0F000405EA0004040404000000",
INIT_03 => X"24004000000000000000000900002C4050000000000069500208400002E14100",
INIT_04 => X"4800200C0000000044002000C80020E40000E200000130200188000000800100",
INIT_05 => X"000000000080181000000000701000004C8000000058800000B1000009880480",
INIT_06 => X"80500081081040000000002C100040400000004641C080380400070100000000",
INIT_07 => X"4020109801A4CE005C00048380142810010564C4100114012002402028044808",
INIT_08 => X"0070700000000000000083004C3902420062000020E0000100004082A140102B",
INIT_09 => X"001150200000000000000026400000016186100000000010C04002C000000000",
INIT_0A => X"007C00008082C0002000000000002C3000000004050001030102040000000000",
INIT_0B => X"0000000000000000000000000000010000800011000000000000000000000BC0",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"000000000000000000000000000000042000760000000000000000010004B200",
INIT_0E => X"0D74002280300F0002FB069040000060000C5003000800000000000000000000",
INIT_0F => X"C01AE8004500744C780687DBA828008080A5FC0D385598035D0008A00C015660",
INIT_10 => X"39D8140040201BF861F0E7D693E6170022408116DFE0AB3006BA0011401D02AC",
INIT_11 => X"5412E4997F5249FD005043B8680CC98F00D0F2DD0140100406FE053A98F6ECC7",
INIT_12 => X"7418663001858040E153888000010840E165D0000000285C246A181C03FE4662",
INIT_13 => X"8199830066F0020858385974000001260208583854E2200000660208D6B1423F",
INIT_14 => X"8235AC508FCE8811042040F008235AE04420C040CF00C031C80009B8F224978B",
INIT_15 => X"030004E00000C220010808C10D9A92A74CD7CF4A09051110AD5A3C9200B7F280",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000118",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"07208BBA3F0C7010C660C7441920000000000000000000000000000000000000",
INIT_1A => X"861869A61861861861869A61861861861861861861861861A8208C4C1534D34C",
INIT_1B => X"984C26130984C26130984C26130984C26130984D26930984C26130984C261861",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000984C26130984C26130",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"174BA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFDFEF5D2A974BA082E95400F7FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0004",
INIT_29 => X"FFFFFFFFFFFFFFFFF7FBFDFFF552E974BAA2FFFFE10087FFFFFFFFFFFFFFFFFF",
INIT_2A => X"004001EFAAAEA8ABA087FFFFFFFFFFFFFEFF7FBEAB450804001EFAAD57FEAAF7",
INIT_2B => X"FFFBFDF45AAD568B55080028B55002E82000F7FFFFFFFFFFFFDFEFA2D568B550",
INIT_2C => X"0007FC00AAF7FFFFFFFF7FBE8B55AAD16ABEF5D2ABFF55080402010087FFFFFF",
INIT_2D => X"55A2FFFDFEF5D2EBFE00AAFFFFEBA087FFFFEFF7D168B55AAD17FFFF552EBFE0",
INIT_2E => X"000AAFFFDF45A2D16AB55F7FFFFFFF00043DE10AA843DE00557FFDFEFA2D16AB",
INIT_2F => X"FFEF552A974AA0000104AA000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFF7FBFDFFF5D2A954AA082A92428E3FFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"0071EFB6DF7AE92EBFFFFFFFFFFFFDFEFF7F5FAFC7492A974AAB6F5F8E101C7F",
INIT_32 => X"F1F8FD7AAD16AB450000001FFBEA4A8AAA147FFFFFFFFFBFDFC7EBF5E8B55000",
INIT_33 => X"00000010087FFDFC7E3F1FAF55A2DF6DB7D1C002AB7D002A82028FFFFFFFEFF7",
INIT_34 => X"BEDB7FFEF552AB8E38087FC2092F7FBF8FC7E3F5EAB45B6DF6FBEF5D2AB8F7D0",
INIT_35 => X"84971F8FC7AAD56DB6DBEF5F8FD7412ABFE28B6F5F8E820871F8FC7E3D56AB6D",
INIT_36 => X"00000000000000000000B6F1F8F55AADF6DB7DE3F5FAFC708003DE28B68E38E2",
INIT_37 => X"FFFFFFFFFFFFFFFFFDFEF552E954AA0004000AA0000000000000000000000000",
INIT_38 => X"54AAF7D568A00557FFFFFFFFFFFDFEFF7FBFFFEF552E974AA082A820AAA2FFFF",
INIT_39 => X"FFF55A2D16AB550000175EFFFFBEAA00A2FFFFFFFF7FBFDFFFFFD568B55002A9",
INIT_3A => X"A800AAF7FBFDFEFF7D56AB45AAD56AB450004001EFFF842AAAA557FFDFEFF7FB",
INIT_3B => X"FFFFFFF552AA8BEF080402000087BFDF45AAD568B55AAFBFDFEF55042ABEF002",
INIT_3C => X"8516AB55A2D16ABEFFFFBFDFFF552AAAAAA007BC0000FFFBE8B55AAD168B55F7",
INIT_3D => X"00043DEAAFFAEAAAAA08556AB55A2D57FFFFF7D568B45002ABDEAAFFD16AA000",
INIT_3E => X"0000000000000000000000000000000000000FFD56AB45A2FFFDFFFAAD16AB45",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024,               -- Port A enable input
WEA      => wbe_a_hi_1024(2),               -- Port A write enable input
DIA(0)   => data_write_a(19),        -- Port A data input
DOA(0)   => data_read_a_hi_1024(19),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024,               -- Port B enable input
WEB      => wbe_b_hi_1024(2),               -- Port B write enable input
DIB(0)   => data_write_b(19),        -- Port B data input
DOB(0)   => data_read_b_hi_1024(19),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_20_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000003",
INIT_01 => X"F55FF80000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"E05022020800008400F655001FFCFF80018FA804400000000000004400000001",
INIT_03 => X"00000000000000000000000900002CC07000000000000000000000000000013F",
INIT_04 => X"68002FFE40900010000180000001FFEC0012EE0C001370F40780000000000000",
INIT_05 => X"0840000880FCBBF0100E204DF0F88311DD8005080679800000F3000029980580",
INIT_06 => X"001000030817C8E8840155FDF9001001050023F6C3C3D0F87FA19F7F011000E4",
INIT_07 => X"000000090492260800008000EE00000000000000002101FF2002C00000004018",
INIT_08 => X"2A040001071004000013FF7FCA302C0C0008214800002101554031F800000000",
INIT_09 => X"801F57F200000090000489FEC0000001EFBEF0040008023FDFC0000000004006",
INIT_0A => X"0000000008000000000000000000ADF000000200000008000008028300110230",
INIT_0B => X"0000000000000800080000000000000000000000000000000800800A40000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"000000040900005C848538000020000000800000080000020000800101FFB600",
INIT_0E => X"00800000003A010003000000000000600FFC53FF001800000002004080000000",
INIT_0F => X"0001000000007408040000004000000004E9000008020000200000000E800800",
INIT_10 => X"00200000000313100010002000008000000000129600040000400000001D0010",
INIT_11 => X"81C012060000000000218F7840000100800004000000000066C0000080080000",
INIT_12 => X"800000000017C000100000000001A800080000000001A8040000002840008185",
INIT_13 => X"0000000006F00000100200000000012600001004000000000066000000801040",
INIT_14 => X"0000200410100000000005F00000020080090A0000000085C800002000586000",
INIT_15 => X"FF00400000000000020020020001000040283024E4F2860400008000030ED080",
INIT_16 => X"00000000000000000000000000000004010201001003020200000000000127DB",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"A0700030038200010089120104D2040020000000000000000000000000000000",
INIT_1A => X"2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2C30C30C30C30C306982121A1E79E79",
INIT_1B => X"32190C86432190C86432190C86432190C86432190C86432190C86432190CB2CB",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000432190C86432190C864",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0201000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF552A974AA0004174BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA0804",
INIT_29 => X"7FFFFFFFFFFFFFFFFFFFFFFEF552E954AA000400000F7FFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E954BA007FC00BA087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974BA082E9540000",
INIT_2B => X"FFFFFFFFFF7FBFDFFF552E974BAA2FFFFE10FFFFFFFFFFFFFFFFFFFFFBFDFFF5",
INIT_2C => X"FAAD57FEAA007FFFFFFFFFFFFFEFF7FBFFF550800020BAAAD56AAAAF7FFFFFFF",
INIT_2D => X"EFF7D56AB450000021EFA2D57DE10087FFFFFFFFFFFFFEFF7FBEAB450804001E",
INIT_2E => X"000F7FFFFFFFFFFFFDFEFA2D568B550004001EFAAAEA8ABA5D7FFFFFFFFFFFDF",
INIT_2F => X"FFFF5D2E954AA080005000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFEF552A974AA0000104AAFFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"A954AA082A92428087FFFFFFFFFFFFFFFFFFBFDFEF5D2E974AA000A07000E3FF",
INIT_32 => X"FFFFFEFF7FBFFFFF552E974AA0071C50BA1C7FFFFFFFFFFFFFFFF7FBFDFFF5D2",
INIT_33 => X"EDF6FABAEBFFFFFFFFFFFFDFEFF7F5FAFC7492A974AAB6F5F8E10E3FFFFFFFFF",
INIT_34 => X"EBF5E8B550000071EFB6DF7AE921C7FFFFFFFFFBFDFEFE3F5F8F450004050AAB",
INIT_35 => X"A497FFFFFFF7FBF8FC7EBD168B450804021FFB6D57DE28147FFFFFFFFFBFDFC7",
INIT_36 => X"00000000000000000000FFFFFFFEFF7F1F8FD7AAD16AB450000001FFBEA4A8AA",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2A954AA0800174100000000000000000000000000",
INIT_38 => X"74AA002E95410A2FFFFFFFFFFFFFFFFFFFFFDFEF552E954AA0004000AAFFFFFF",
INIT_39 => X"FDFEFF7FBFFFEF552E974AA082A820AA087FFFFFFFFFFFFFEFF7FBFDFFF5D2A9",
INIT_3A => X"568A00AAFFFFFFFFFFBFDFEFFFFFFDFEF5D2E954AA0051554BA557FFFFFFFFFF",
INIT_3B => X"D16AB450804174AAFFFFFFEBAA2FFFFFFFF7FBFDFFFFFD568B55002A954AAF7D",
INIT_3C => X"57FFDFEFF7FBFFF55A2D16AB550000175EFFFFBEAA005D7FFFFEFF7FBFDFFFAA",
INIT_3D => X"0004001EFFF842AAAA087BFDFEFF7FFEAB45A2D568B550804001EFF7D57DEBA5",
INIT_3E => X"0000000000000000000000000000000000000F7FBFDFEFF7D56AB45AAD56AB45",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024,               -- Port A enable input
WEA      => wbe_a_hi_1024(2),               -- Port A write enable input
DIA(0)   => data_write_a(20),        -- Port A data input
DOA(0)   => data_read_a_hi_1024(20),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024,               -- Port B enable input
WEB      => wbe_b_hi_1024(2),               -- Port B write enable input
DIB(0)   => data_write_b(20),        -- Port B data input
DOB(0)   => data_read_b_hi_1024(20),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_21_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"4A302428B824900A128C090A5C1800261500213C005FE812D10420054085A202",
INIT_01 => X"001FFE3440B609703B0427F801A40B8115BC4F655300340288A40D30040E4DD8",
INIT_02 => X"E00424256888D8819801000F9FFFFFFFF149FF1FCA448046C60A0D2437C517F9",
INIT_03 => X"20030640003250640003250F06002CC1740002019824E001CD357832440001FF",
INIT_04 => X"EA2C3FFD400006E04401A8837001FFFC004AEF00080B70E08FB5789421007C5C",
INIT_05 => X"00011A0C40F9FFF80920954FF0F00809DF84A0202879800000F3000029980780",
INIT_06 => X"0805984B7A1FC0A0000101FFF0480080002281F7C3C381F87C03DFFF00009004",
INIT_07 => X"B424068086A205481A60A19000908204A855B000A08A61FF20C3D004D331D340",
INIT_08 => X"1BFA0001600802000023F7FFC08D234B40C2028253000040114200000D0226C0",
INIT_09 => X"EF1F5FF054096C6ADBA169FFC202B1C1FFBEF0440021083DFFCE22DC2880E24D",
INIT_0A => X"45FF0C004041D84862A28C54518DBFF00020004C0A6044901112A0908AA0A300",
INIT_0B => X"018C241102068006C620C03882019480E63180855A492712CC01C49C20201BFE",
INIT_0C => X"08A9464116544302C02D92236488D92236488D92236488D922366446C911B210",
INIT_0D => X"08800444021048034004001890000806002804A0822189000900D80621FFBE00",
INIT_0E => X"060580261013813A2CC396506102C4053FFD5BFF00A04A00200602CA52001100",
INIT_0F => X"080C0B004C202621A85C09411500135844C196D3606941018150098404C1A304",
INIT_10 => X"B02901013416181C96C2C9C600890A2028172192C460D1820302A0130809834A",
INIT_11 => X"9C5E803408250180AC268D185DB3F4350B811068C00049A0A4AA68F05C96A001",
INIT_12 => X"002C006560138F032B1804101244C883052208209040CC849063A747512B7678",
INIT_13 => X"41401E240665750440C9488280254530314080C2C601040420352148A00501B1",
INIT_14 => X"500811204D000700114204A70422016149916011008CAA8858850B00C32591C0",
INIT_15 => X"FFC06E60AC0496022300233104663040808E991765205000070121D41D18D098",
INIT_16 => X"40100401004010040100401004010040102090010008000001C0E010020007DF",
INIT_17 => X"0100401004010040100401004010040100401004010040100401004010040100",
INIT_18 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_19 => X"FFEF9FEEFF7FFDF7FF3E3DFDF7E0000000000000000000000000401004010040",
INIT_1A => X"BEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBFFDFDFFFCF3CF3F",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFEFF7FBFDFEFF7FBFDFEFBEF",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000FFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0001000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E954AA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0004",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA0004154BAFFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"52E974BA0804000AAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0004174BAFF",
INIT_2B => X"FFFFFFFFFFFFFFFFEF552E954AA000400000007FFFFFFFFFFFFFFFFFFFFFFEF5",
INIT_2C => X"A082E95400007FFFFFFFFFFFFFFFFFFFFDFEF5D2E974BA002E97400007FFFFFF",
INIT_2D => X"FFFFFBFDFEF5D2A954AA002E974BA087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFBFDFFF5D2E954BA007FC00BA5D7FFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA000002000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080005000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"A974AA0000104AAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974BA0000174AAFFFF",
INIT_32 => X"FFFFFFFFFFFFDFEF552E954BA080A000AAE3FFFFFFFFFFFFFFFFFFFFFFFEF552",
INIT_33 => X"02A95400087FFFFFFFFFFFFFFFFFFBFDFEF5D2E974AA000A07000007FFFFFFFF",
INIT_34 => X"F7FBFDFFF5D2A954AA082A924281C7FFFFFFFFFFFFFFFFFFBFDFEF5D2A974BA0",
INIT_35 => X"A557FFFFFFFFFFFFFFFF7FBFDFFF552E974BA0020924BA1C7FFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000E3FFFFFFFFFFFFFFEFF7FBFFFFF552E974AA0071C50B",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0000020000000000000000000000000000",
INIT_38 => X"74BA0000174BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954AA080017410FFFFFF",
INIT_39 => X"FFFFFFFFFFDFEF552E954AA0004000AAF7FFFFFFFFFFFFFFFFFFFFFFFEF552A9",
INIT_3A => X"E95410087FFFFFFFFFFFFFFFF7FBFDFEF5D2A954BA082E800AAA2FFFFFFFFFFF",
INIT_3B => X"FBFFFFF552E954BA002E97410087FFFFFFFFFFFFFEFF7FBFDFFF5D2A974AA002",
INIT_3C => X"57FFFFFFFFFFFDFEFF7FBFFFEF552E974AA082A820AA557FFFFFFFFFFFFFEFF7",
INIT_3D => X"5D2E954AA0051554BA5D7FFFFFFFFFBFDFEFF7FFFFFEF5D2A974BA0000020AA5",
INIT_3E => X"0000000000000000000000000000000000000AAFFFFFFFFFFBFDFEFFFFFFDFEF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024,               -- Port A enable input
WEA      => wbe_a_hi_1024(2),               -- Port A write enable input
DIA(0)   => data_write_a(21),        -- Port A data input
DOA(0)   => data_read_a_hi_1024(21),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024,               -- Port B enable input
WEB      => wbe_b_hi_1024(2),               -- Port B write enable input
DIB(0)   => data_write_b(21),        -- Port B data input
DOB(0)   => data_read_b_hi_1024(21),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_22_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"5290F4CDE914905A14A43D33F488243E17122300F55FEB189B343A1140548380",
INIT_01 => X"A54007B259F6A975386262000C344BA9573C6FF57B18A5FB0ABFCD3C2C5F4F0C",
INIT_02 => X"021DFF8C38B3C009D203551040030071869D0040180AA2DC53DB89BEA8204001",
INIT_03 => X"2603475A969D0475A969D0460EAA401005111011BD506954EDB40F5EF41434C0",
INIT_04 => X"922D9002100ED69E443D988B0D5400103E48003D0800011E803B06B5B9125A15",
INIT_05 => X"281B5A0C06000408F4DF9422010D8802022F2124A8022492580040440002021C",
INIT_06 => X"F780C4C052881ADA0E05440205DA50930FA182010004700083E220800440B588",
INIT_07 => X"049D028B93FB561833D8094A02F5EA92FD7247E10305C40040D136E6A023F7FC",
INIT_08 => X"00028241680A0E002A9400803A884B5B5206B7C2E53CA25144009007A64EBD64",
INIT_09 => X"41008810240240C6694008010392354010000560141801002028A83D2A08E06D",
INIT_0A => X"34000000848BCA6902A29C54539C020E11810098D4067EFF9FF284D483E2AB41",
INIT_0B => X"500001840000C80B410014088040F4A944B1AA313C0022AA0011C0DC00028001",
INIT_0C => X"80B14004D158C8CA24A1C2A870AA1C2A870AA1C2A870AA1C2A872550E1543800",
INIT_0D => X"80A14050A01509E050854498B5281A1C34E506A2C6898B52A154DAC6B6000850",
INIT_0E => X"0B03001A483A4146603050080410089180008800143D83888281A2034A850142",
INIT_0F => X"A4160600349075238473F1210006133835E92273612B3482C090068A0E84AC56",
INIT_10 => X"30060181BA1B13959DC08DA902458870201970B29602562B0581200D141D0959",
INIT_11 => X"E042021C040D0152C8058B3840F044708E7E1C20A0106EA166C13AFC14AA3804",
INIT_12 => X"080E004B0C17C1439A9838301DC1A8438EA32C009DC1A8255300650458A1D588",
INIT_13 => X"018010E186F110A908E3A8CB0026C9A610A908E6A60F0807626610E160589C4C",
INIT_14 => X"2A701667334005800B1605F043858125E0D04110408D2485CA034681E43A1E40",
INIT_15 => X"00646002304244A91102C93A2D608D2A258DF8034188200C050171A41108F084",
INIT_16 => X"110441104411044110441104411044110466C440446CA06951D4EA8010009804",
INIT_17 => X"0040100401004411044110441104411044110441104411044110441104411044",
INIT_18 => X"0401004010040100401004010040100401004010040100401004010040100401",
INIT_19 => X"F7DFBFDEFE8FF1F7DEBDDF7DF7D05122890000000003FFFFFFFF900401004010",
INIT_1A => X"9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7BFFDFD7DDDF7DF7D",
INIT_1B => X"F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE79E7",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000003F9FCFE7F3F9FCFE7F3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA000400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0800",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000002000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2A954BA000015400FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080402010FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2A954BA0004154BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A0004174BAFFFFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0800154AAFFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF552A974AA0000174BAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974A",
INIT_2E => X"000007FFFFFFFFFFFFFFFFFFFFFFEF552E974BA0804000AAA2FFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080400010000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E954AA080005000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000402010FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2A954BA000417410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"804154BAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974BA0000174AAFFFFFFFFFFF",
INIT_34 => X"FFFFFFFEF552A974AA0000104AAE3FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0",
INIT_35 => X"AA2FFFFFFFFFFFFFFFFFFFFFFFEF552E954BA000E124BAE3FFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000007FFFFFFFFFFFFFFFFFFFFDFEF552E954BA080A000A",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804000100000000000000000000000000",
INIT_38 => X"54AA000400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2A954AA080017410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"0174BAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A954BA000415400FFFFFFFFFFFFF",
INIT_3B => X"FFFDFEF552E974AA0804174AAF7FFFFFFFFFFFFFFFFFFFFFFFEF552A974BA000",
INIT_3C => X"2FFFFFFFFFFFFFFFFFFFFFDFEF552E954AA0004000AAA2FFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2A954BA082E800AAAAFFFFFFFFFFFFFFFFFFFBFDFEF5D2E954BA002A820BAA",
INIT_3E => X"0000000000000000000000000000000000000087FFFFFFFFFFFFFFFF7FBFDFEF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024,               -- Port A enable input
WEA      => wbe_a_hi_1024(2),               -- Port A write enable input
DIA(0)   => data_write_a(22),        -- Port A data input
DOA(0)   => data_read_a_hi_1024(22),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024,               -- Port B enable input
WEB      => wbe_b_hi_1024(2),               -- Port B write enable input
DIB(0)   => data_write_b(22),        -- Port B data input
DOB(0)   => data_read_b_hi_1024(22),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_23_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"EF20906D902424807BC8241BC81801B97D38AD3C0800103362A6741C80A12A02",
INIT_01 => X"001FFF8409F089003B4422000D80C80106804A7951C5B9D1C828043EA28838F9",
INIT_02 => X"E01CEE21649C82C40800000F9FFEFF8E72CA7F5FC2E22809925A0D3611C877F8",
INIT_03 => X"24000400402670400402670D48222DC1764446838624000080007460C40001BF",
INIT_04 => X"68403FFC020560E0443E21037C01FFFC0002EE00628BF0E02FAD781014085014",
INIT_05 => X"0112000202FBFFF00920017FF0F0628BFF8488890979800002F702002BB807A0",
INIT_06 => X"EF85788B681FC000000001FFF0010000000001F7CBC385F87C0BFFFF20040001",
INIT_07 => X"F6E200000000C1440E3AE408009120071070FA07A1CB23FFA403F0C4D23BF7C0",
INIT_08 => X"0BF87CA400804000003FF7FFD8880A034AC09662305AB10555421006891A1089",
INIT_09 => X"BE1F5FEA10092C0896A243FFC0008087FFBEF2000000001DFFC612C0C0400100",
INIT_0A => X"41FF0C2060501000600000000001BFFA800808189A657EF81DD0C00079CC8001",
INIT_0B => X"018C24110A860006C620C0312241C482B20400CC52492710CC80060020A81BFE",
INIT_0C => X"0C08866907048320C20C10030400C10030400C10030400C10030400608018210",
INIT_0D => X"040002000041500300100040000500C000801000C02400000952800001FFBF04",
INIT_0E => X"FC850015385380380CDB86106502C5043FFD5FFF00A04BC010A7724B10000800",
INIT_0F => X"89F90A002A70A710A51C01C05904014861433602A1CAF13F2110055614C72FC0",
INIT_10 => X"E02D02001C1E14981B43253EE50C8220180F1082E06397E07E42200AAC298E57",
INIT_11 => X"8421802400A90022B0070FAE18019214A380344920080B21A58B02AC60BACDF0",
INIT_12 => X"0A2A000C480B0704B54028101AC49C84BB4100009AC49C80857A82D20CE8CB22",
INIT_13 => X"01E00C8103416445C12ED0400027C5292445C12D500B0005A62D344CB241D095",
INIT_14 => X"132C907425604680038706A35132C94BDD011010404428886AC91B11311C8280",
INIT_15 => X"FF000470BE0692020328CA0028042054A92771C50FC070110001C1680809591D",
INIT_16 => X"00802008020080200802008020080200800800200200000000000008004807DF",
INIT_17 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_18 => X"8020080200802008020080200802008020080200802008020080200802008020",
INIT_19 => X"0000000000000000000000000000000000000000000000000000008020080200",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080002010FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974AA000400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000400010FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974AA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080000010FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E954AA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954A",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA000015400FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080002010FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974AA000400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000402010FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E954AA080005000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA080407000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA00041741",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080000010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000402010FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2A954AA080002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954AA080017410FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"552A954BA000415400F7FFFFFFFFFFFFFFFFFFFFFFFFF552A954BA080015410F",
INIT_3E => X"0000000000000000000000000000000000000F7FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024,               -- Port A enable input
WEA      => wbe_a_hi_1024(2),               -- Port A write enable input
DIA(0)   => data_write_a(23),        -- Port A data input
DOA(0)   => data_read_a_hi_1024(23),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024,               -- Port B enable input
WEB      => wbe_b_hi_1024(2),               -- Port B write enable input
DIB(0)   => data_write_b(23),        -- Port B data input
DOB(0)   => data_read_b_hi_1024(23),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_24_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100600007FFF000080108004000800020000840041000080808",
INIT_02 => X"FC5CA803400EB8209000000F9FFEFF8E7240FF1FC22409EA04018E50074017F0",
INIT_03 => X"11100400000000400000000D00002CC07400000090C080019001010A000001BF",
INIT_04 => X"68003FFC00040000000000008001FFFC0002EE00000370E007A100000000E468",
INIT_05 => X"0000000000F8BFF00920004DF0F00001DF8000000079800000F3000029980780",
INIT_06 => X"6E461803081FC000000001FFF0000000000001F7C3C380F87C019FFF00000000",
INIT_07 => X"600C2400013649609C8000980040814210254000A00B21FF2003F2A80D500000",
INIT_08 => X"0BF80000000000000003F7FFD88D2B4A02C0940062EC2804001610020408178B",
INIT_09 => X"8E1F5FE010092C0892A041FFC0000001FFBEF0000000001DFFC002C000000000",
INIT_0A => X"41FF0C0000000000600000000001BFFA0000005501AA00000CE2000009400000",
INIT_0B => X"018C0411020600048620C030020502000200000400490510CC00040020201BF4",
INIT_0C => X"0808064106040300C00C10030400C10030400C10030400C10030400608018210",
INIT_0D => X"0000000000004003000000000000001200580000000000000000000001FFBE00",
INIT_0E => X"0086C022005381380FDB96516140C6043FFD5BFF000041000000004110000000",
INIT_0F => X"80010D804400A7240C840C201D0210840043B4804012500021E0088014C04940",
INIT_10 => X"4109038041021C980200D06410C1924030008142E06024A00043C01100298092",
INIT_11 => X"587CC200002100C14428090A1D02348190814C09C010104025AA40041A0D8005",
INIT_12 => X"022E0030300B0E46177004208000D8C61D7004300000D884817B00011306B2D9",
INIT_13 => X"01E003060344710009875C018100013831000985DC000C20003C310006143B70",
INIT_14 => X"4001850EDC004780144806A64400186CBF8961104000C3807884000846EB9500",
INIT_15 => X"FF0006E08C063C0220002201490418082010A57263E0100008000290161E711C",
INIT_16 => X"00000000000000000000000000000000000000000000000000000000000007DF",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"F2D0AEEAF6E7CC1132CDB4441990000000000000000000000000000000000000",
INIT_1A => X"BEFBE79E79E79E79E79EFBEFBEFBEFBEFBEF9EF9EF9EF9EFA69861219575D75F",
INIT_1B => X"783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1EFBEF",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000783C1E0F0783C1E0F0",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0201000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A000400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA000400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000400000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402010000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"00002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080002010FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000400010FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA00040000",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020100000000000000000000000000",
INIT_38 => X"74BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"000010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA000002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974AA000402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000002010F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024,               -- Port A enable input
WEA      => wbe_a_hi_1024(3),               -- Port A write enable input
DIA(0)   => data_write_a(24),        -- Port A data input
DOA(0)   => data_read_a_hi_1024(24),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024,               -- Port B enable input
WEB      => wbe_b_hi_1024(3),               -- Port B write enable input
DIB(0)   => data_write_b(24),        -- Port B data input
DOB(0)   => data_read_b_hi_1024(24),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_25_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100200002000000080100004000000020000800041000080808",
INIT_02 => X"FC400086000000800000000F9FFEFF8E738FFF1FC204010000000111568DD7F8",
INIT_03 => X"00000400000000400000000D00002CC4740000008000000080000000000001BF",
INIT_04 => X"68003FFF64A564AC000000000001FFFE0082EF00010370E007A1000000004000",
INIT_05 => X"0A00040148F8BFF80920804DF0F00101DFC040000079C92484F30499299837C1",
INIT_06 => X"66041803081FC0E0801101FFFD000E41002299F7E3C380F87C019FFF81200096",
INIT_07 => X"000000080480AE00000080000000000000000000A00B21FF2003E00000000000",
INIT_08 => X"1BF80000400A02000003F7FFFA0008000200A0400008A0000014100200081000",
INIT_09 => X"8E1F5FFA53EFBCACB2E369FFE0010001FFBEF80C40630C7DFFEEBAF000800202",
INIT_0A => X"41FF0C0600000000600000000001BFFE00301000000000000CC020000140000C",
INIT_0B => X"01DCCC31222730A49620C030020100000200000400490D10EC00040220201BF4",
INIT_0C => X"0808064106240300C00C10030400C10030400C10030400C10030400608018210",
INIT_0D => X"0883044582114013412080000000000000000000000000000012800001FFBE00",
INIT_0E => X"00040020000180380FC386106140C6043FFD5BFF00A04B80608003CB120C1106",
INIT_0F => X"0000080040000200040400000100000000009480000240000100080000400900",
INIT_10 => X"0001000000000808000000240000020000000100006004800002001000008012",
INIT_11 => X"0001001808220000002004001900000080800008000000000022400000088000",
INIT_12 => X"0010000000000E00110000000000408009000000000040808063004000008200",
INIT_13 => X"6000000000046100000240000000001021000004400000000010210000001010",
INIT_14 => X"4000000404000800000000060400000088000001800000001084000000088000",
INIT_15 => X"FF800C608C041002000002000006100000002100000000180600000000100018",
INIT_16 => X"4110441104411044110441104411044510629041040D180400000010028047DF",
INIT_17 => X"1104411044110441104411044110441104411044110441104411044110441104",
INIT_18 => X"1044110441104411044110441104411044110441104411044110441104411044",
INIT_19 => X"FBA2894A196A8C5A2932EC15DA080800002FFFFFFFFFFFFFFFFFC11044110441",
INIT_1A => X"2492492492492492492410410410410410410492410492412000531215A69A6B",
INIT_1B => X"158AC562B158AC562B158AC562B158AC562B1588C46231188C46231188C49249",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000B158AC562B158AC562B",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080000010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000010FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08000000",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024,               -- Port A enable input
WEA      => wbe_a_hi_1024(3),               -- Port A write enable input
DIA(0)   => data_write_a(25),        -- Port A data input
DOA(0)   => data_read_a_hi_1024(25),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024,               -- Port B enable input
WEB      => wbe_b_hi_1024(3),               -- Port B write enable input
DIB(0)   => data_write_b(25),        -- Port B data input
DOB(0)   => data_read_b_hi_1024(25),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_26_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"E9264EAB20190CA3BA4997AA9002AE9C001006B0778015CFA17E0811039879C7",
INIT_01 => X"2FFFF9BB1F773C7F9BB07DFFFDD863FC5FFF3FEFFBBF9FFB22FFFBC7B9F30686",
INIT_02 => X"E06CCC62052E708180F6FFBFFFFCFFFFF9C7FF7FC24332E642090000074037F6",
INIT_03 => X"428003739CD9863739CD9869FE2B7DEAF300029E4E300DFE69A6E644E6FF473F",
INIT_04 => X"7C2FEFFFF5BA124F003DD31EAFFFFFEE9FF7EE6F4C0770FFD7DC7CA53997B2B1",
INIT_05 => X"DFFB5421C1F8BBFAFDBFFACDF0FFCC05DDDBFF3690F9EDB7F5F7AFF639BD7DE3",
INIT_06 => X"EFD044ABC817C3E3A74667FDFFB6FF5727CC3BFEF7C3FAF87FF59F7FFBFEF69F",
INIT_07 => X"00003002132462052E708180EF060C18E5BEFB051225CDFF7002C4EEDE77F6E0",
INIT_08 => X"3FFF7D5000EC75088ED3FF7FC8790E46426CE06CB1F8E041051831FA3068D77E",
INIT_09 => X"C05FD7FF9BEFBDCEFBEE59FEF44F6603EFBEFAFCC2E35E7FDFD147CCF3F583FA",
INIT_0A => X"67FF1C7FBFADEB31E35768E8ED6BFDF3EB3EBF9DDBCE7FDC1DF8A760F3EACC02",
INIT_0B => X"5BDDCC3B336F7C548667D47B7737AF3FD62601EDC25B3533DCEB07F262213FFC",
INIT_0C => X"5F9A06E19F4D93A0EA0F78C35E30D78C35E30D78C35E30D78C35E986BC61AE31",
INIT_0D => X"5FD7AFEFDFFAF59B6FF28FE1D80D73D840607307DCFE1D80EF69A004DFFFF7FF",
INIT_0E => X"0004001F8041897B2FFFC6D86D70CE04FFFFF3FF1F5F5475BD7F72E4D75EBFAF",
INIT_0F => X"F60008003F008237B0040A00010003E020023E0201F45EC0010007E01047D17B",
INIT_10 => X"00010001DC0004C81003DE050A700200001DC0006863E8BD8002000FC0208FA2",
INIT_11 => X"2200E400002801E1A00004C21C0206F60081800800007B00010F02007EC09A0E",
INIT_12 => X"0880007E000807C7C1A612001E0015C7C19C22001E0015C59DFE82011A311AA0",
INIT_13 => X"00001BC00101F60409F0670840070809760409F06984800780097604067D0010",
INIT_14 => X"81019F40042100001F800203D81019EC085614000085C80023D81009CF008A74",
INIT_15 => X"FF802FFDFFAFD082003B032FB987E04021D481D4000819060801E0D00001231D",
INIT_16 => X"EBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEFFBFBFBFBBFCFBB0FFDFEFFEF2DFFFFFB",
INIT_17 => X"BFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAF",
INIT_18 => X"FAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFE",
INIT_19 => X"475B15BCF491E166CC8553F86EDB5C88646FFFFFFFFFFFFFFFFFEBFAFEBFAFEB",
INIT_1A => X"861861861861861861861861861861861861869A69A61861AFBD54D5F871C71D",
INIT_1B => X"984C26130984C26130984C26130984C26130984C26130984C26130984C261861",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000984C26130984C26130",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040201",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024,               -- Port A enable input
WEA      => wbe_a_hi_1024(3),               -- Port A write enable input
DIA(0)   => data_write_a(26),        -- Port A data input
DOA(0)   => data_read_a_hi_1024(26),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024,               -- Port B enable input
WEB      => wbe_b_hi_1024(3),               -- Port B write enable input
DIB(0)   => data_write_b(26),        -- Port B data input
DOB(0)   => data_read_b_hi_1024(26),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_27_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"00080A40000A41248002029000050A088000008242A0004404480002000A1155",
INIT_01 => X"2FFFF1C11F781C129C107DFFFE0860941E81258CA2B71C2220EC1B86E1A00002",
INIT_02 => X"E1000000810000014400FF6FFFF0FFFFF8007F1FC21110005080200000221FF0",
INIT_03 => X"4080026318C18226318C1821302232EAE00002BE001115FE48620040840A863F",
INIT_04 => X"643D4FFC2530000F003D821C0BFFFF8E9EF79E6D440748FED70060842105B0B0",
INIT_05 => X"D6F39020D1F8A3FAFDBFBACDC8FDC405D1DB7F1490E5EDB7D5CBADB2385D79C3",
INIT_06 => X"6FE000A38007C3032646EFF1F0B6FF46A78C39F8E723F2E47FE59C7F9ADA2612",
INIT_07 => X"00002820000000810000014401060C180190310540118DFF1000C0849673F6C0",
INIT_08 => X"3FF779100062B12A8EC3F47FC80208808210880C00082050000110023068D030",
INIT_09 => X"005F07E09BFFBD07FBAC09F8E42922038F7DF8BEC2E39C5F1FD047CEF1B582D8",
INIT_0A => X"63FF5D5F9FADE911E81C09818109E1F16B16B71092CE7ED81CF403601228C402",
INIT_0B => X"1BFDCC39732F3554866AD57C37BEAF1C152201A4C05B7531D56B05B06A213FF8",
INIT_0C => X"5BCA06F18FC59380F00E34430D10C34430D10C34430D10C34430F0861A2186B5",
INIT_0D => X"5B56ADAB5FAAE58B2F628EA0C80FA3F04040510768EA0C80CC61A0044DFFC6EB",
INIT_0E => X"0004001D800188792CE79715710AE4047FFD23FF315D54358D593474955AB6AD",
INIT_0F => X"520008003B000297B0040200010003E020001F0201E44A400100076000579129",
INIT_10 => X"00010001DC00004A10035E0408300200001DC000086BC8948002000EC000AF22",
INIT_11 => X"02002400002801E1A00000C01E0202F60080800800007B00000782006EC0820A",
INIT_12 => X"0080007E000006A7C10602001E0001A7C10C02001E0001C18DE282010A311AA0",
INIT_13 => X"00001BC00000FE0401F04300400708007E0401F04180800780007E04047D0010",
INIT_14 => X"81011F40040100001F800002F81011EC080604000085C80001F810094F008034",
INIT_15 => X"FF800C6DDDAFD082001B03249887E04001D481D4000009020801E0D00001021F",
INIT_16 => X"AB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6BF1EBDABD8E270BF84A25C6ACB777E3",
INIT_17 => X"B6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6AD",
INIT_18 => X"6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADA",
INIT_19 => X"490E2168100481CA860402104A471688747FFFFFFFFFFFFFFFFFAB6ADAB6ADAB",
INIT_1A => X"000000000000000000000000000000000008200000000000200072F210000001",
INIT_1B => X"05028140A05028140A05028140A05028140A0500804020100804020100800000",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000A05028140A05028140A",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040201",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024,               -- Port A enable input
WEA      => wbe_a_hi_1024(3),               -- Port A write enable input
DIA(0)   => data_write_a(27),        -- Port A data input
DOA(0)   => data_read_a_hi_1024(27),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024,               -- Port B enable input
WEB      => wbe_b_hi_1024(3),               -- Port B write enable input
DIB(0)   => data_write_b(27),        -- Port B data input
DOB(0)   => data_read_b_hi_1024(27),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_28_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"02200AA400180030808802A900002A08001280A08A801044104A1000001818C3",
INIT_01 => X"0AA00011460214428114180000882214413D0A71592A01D92213D28005210202",
INIT_02 => X"0451110A012100884000AA30200000000C100040104112101100008888200000",
INIT_03 => X"448000318C52A20318C52A20148810200111100C211004AA00034204200A2200",
INIT_04 => X"04004001001A90110000121402AA0000003C00000500000040080421080D0080",
INIT_05 => X"4060000C8001000000002E000000050000001610300000010000802202040012",
INIT_06 => X"1000002080001111001222000425A1040026A008000000000000000009328280",
INIT_07 => X"2491008A00491201210088400122448908A20402000408001000040820000000",
INIT_08 => X"20058310402A160026500000028040101004200C840082115554000112244814",
INIT_09 => X"4140000800000060000720000102028000000490160801020002200011100010",
INIT_0A => X"020000081B34211082B694D4D294000020020381040000000200032040004400",
INIT_0B => X"4800210C19808400500010009110091500020B408810000100200020408B0000",
INIT_0C => X"01028000080118020023604858121604858121604858121604858090B0242C00",
INIT_0D => X"010000800920040804020A6058003108402043058C460580653020005A004039",
INIT_0E => X"00000002800008014004104104420A00C000200005000010040A0020CC000200",
INIT_0F => X"520000000500000010000200000000000000280000040A40000000A000001029",
INIT_10 => X"00000000000000C0000002000830000000000000480008148000000140000020",
INIT_11 => X"020024000000000000000440000000020000800000000000000C00000040020A",
INIT_12 => X"00800000000001804006020000000500400C0200000005400A90000000100000",
INIT_13 => X"0000000000018200001003004000000142000010018080000001420000200000",
INIT_14 => X"8000080000010000000000018800008000060400000000000310000008000034",
INIT_15 => X"000002040080000000110006B081400000400000000009020000000000002200",
INIT_16 => X"802008020080200802008020080200802101210810C39A66A90A85420413A820",
INIT_17 => X"0200802008020080200802008020080200802008020080200802008020080200",
INIT_18 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_19 => X"DE21102C110A00246972BD89A40A0C22E1000000000000000000002008020080",
INIT_1A => X"2082082082082082082082082082082082082082082082080D35050758C30C31",
INIT_1B => X"0582C160B0582C160B0582C160B0582C160B0580C06030180C06030180C08208",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000B0582C160B0582C160B",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024,               -- Port A enable input
WEA      => wbe_a_hi_1024(3),               -- Port A write enable input
DIA(0)   => data_write_a(28),        -- Port A data input
DOA(0)   => data_read_a_hi_1024(28),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024,               -- Port B enable input
WEB      => wbe_b_hi_1024(3),               -- Port B write enable input
DIB(0)   => data_write_b(28),        -- Port B data input
DOB(0)   => data_read_b_hi_1024(28),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_29_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"79964E4BA01DACAB9E659792D00AAE160002829C7FDFEFCEE97C2815039D70C3",
INIT_01 => X"0ABFF9AB0775343F9AB01DF80D5821FC0FFF3FEFD1AF9FF1207FFBC7B9720586",
INIT_02 => X"002CCC60050E700080F6AAA7BFFC007189C7FF2FC00330E602800000074037F6",
INIT_03 => X"468003210868A63210868A68DA017D207200021C4E200CAA6186A40042FF4300",
INIT_04 => X"7C2FE002F0900001003C5316A6ABFFE21F36E02F0D03701F47D41800109FB281",
INIT_05 => X"4979440580F9B808F49F6A4DF00F8D01DC4B97369078249370F482E62BA41462",
INIT_06 => X"B250442BC81001E1870223FC0BF7F11507C423FE33C078F803F19F00E936721D",
INIT_07 => X"00011080012460050E700080EF020408EC8CFA01122149FF700200665A35D260",
INIT_08 => X"2BFD055040A452000443FF00007906464068406C31F84000000831FA1028575A",
INIT_09 => X"805FD017102690AA694551FE30444681E0820AD40201423FC00122C493500172",
INIT_0A => X"0600002AFFBE2330815568A8AD6ABC02A02A0B0CCB463B4C0748A720B1EA4C00",
INIT_0B => X"0850400A11414C005005000B51158936D20601A98A10200308A002E240010BFC",
INIT_0C => X"05928020194918A22A2268C81A32068C81A32068C81A32068C81A99034640C00",
INIT_0D => X"058102C48970541944B20FA1580561D040406305587A158046282000DBFFF13D",
INIT_0E => X"000000028040890327DCD28928324400DFFFF0001F1F0050342D42A086040B02",
INIT_0F => X"F60000000500802010000A000000000000022A0000141EC0000000A01000507B",
INIT_10 => X"00000000000004C0000082010A700000000000006800283D80000001402000A0",
INIT_11 => X"2200E4000000000000000442040004020001800000000000010D000010401A0E",
INIT_12 => X"08800000000801C040A6120000001540409C2200000015441DAC800010100000",
INIT_13 => X"0000000001019600081027084000000956000810298480000009560002200000",
INIT_14 => X"800088000021000000000201D800088000561400000000002358000088000A74",
INIT_15 => X"00802594A282C0000033010FB181E00020400000000819060000000000002305",
INIT_16 => X"C0B02C0B02C0B02C0B02C0B02C0B02C4B12B312912831A27FCFE7FFB175B6FF8",
INIT_17 => X"0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02",
INIT_18 => X"B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C",
INIT_19 => X"BBCF9F96EE7FFDF7FE783FFDFFEA0C00602FFFFFFFFFFFFFFFFFC0B02C0B02C0",
INIT_1A => X"EFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEEBAEBAEBAEBAEBBFFDF9FBEFFFFFFE",
INIT_1B => X"BFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFBEFB",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000FBFDFEFF7FBFDFEFF7F",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024,               -- Port A enable input
WEA      => wbe_a_hi_1024(3),               -- Port A write enable input
DIA(0)   => data_write_a(29),        -- Port A data input
DOA(0)   => data_read_a_hi_1024(29),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024,               -- Port B enable input
WEB      => wbe_b_hi_1024(3),               -- Port B write enable input
DIB(0)   => data_write_b(29),        -- Port B data input
DOB(0)   => data_read_b_hi_1024(29),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_30_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"F7FFBFFEFF9FE1F7FFBFFFFDFFD0000000000000000000000000000000000000",
INIT_1A => X"9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7AFBD75F5FDF7DF7F",
INIT_1B => X"F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE79E7",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000003F9FCFE7F3F9FCFE7F3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024,               -- Port A enable input
WEA      => wbe_a_hi_1024(3),               -- Port A write enable input
DIA(0)   => data_write_a(30),        -- Port A data input
DOA(0)   => data_read_a_hi_1024(30),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024,               -- Port B enable input
WEB      => wbe_b_hi_1024(3),               -- Port B write enable input
DIB(0)   => data_write_b(30),        -- Port B data input
DOB(0)   => data_read_b_hi_1024(30),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_31_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"129000008004A00804A40000400800020000000C005FEA005800200400050100",
INIT_01 => X"255FF18019700810180065FFFC0040801E80258CA2951C2200EC0906A0804140",
INIT_02 => X"E0000000000000011000550FDFF0FFFFF0007F1FC200000044000000000817F0",
INIT_03 => X"0000024210A30024210A3001002220C06044469200040154482000408400043F",
INIT_04 => X"602D0FFC2420000E003D80080955FF8E1ECA8E2D400340FE870060842100B030",
INIT_05 => X"0213100040F8A3F8FDBF944DC0FDC001D1CB6904A061EDB6D4C30490281831C1",
INIT_06 => X"6FC000830007C202060445F1F0D25E4207A099F0E303F0E07FE19C7F80402412",
INIT_07 => X"0000200000000000000001100004081001103107000185FF0000C0849673F6C0",
INIT_08 => X"1BF27A00000000000883F47FC800080002008000000820440000100220489020",
INIT_09 => X"011F07E013EFBC06FBA009F8E00120038F3CF82C44630C5D1FC002CCE0808248",
INIT_0A => X"61FF0C06C48BC801600000000001A1F00110101092CE7ED81CF0004012288000",
INIT_0B => X"11DCCC31222730048620C4382204A608142002A440492530C401049020221BF8",
INIT_0C => X"0888066187448380E00C10030400C10030400C10030400C10030600608018210",
INIT_0D => X"080204010200418301208480800D02D00040100240A808008840800405FF8640",
INIT_0E => X"0004001D000180780CE386106100C4043FFD03FF101D40008001304018081004",
INIT_0F => X"000008003A000217A0040000010003E02000160201E040000100074000478100",
INIT_10 => X"00010001DC00000810035C0400000200001DC0000063C0800002000E80008F02",
INIT_11 => X"00000000002801E1A00000801C0202F40080000800007B00000302006E808000",
INIT_12 => X"0000007E00000607810000001E000087810000001E000081846282010A211AA0",
INIT_13 => X"00001BC00000740401E0400000070800340401E04000000780003404045D0010",
INIT_14 => X"01011740040000001F8000025010116C080000000085C80000C8100947008000",
INIT_15 => X"FF800C609C06D082000A03200806A040019481D4000000000801E0D00001001D",
INIT_16 => X"010040100401004010040100401004010060C040040C200950402090128057C3",
INIT_17 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_18 => X"0040100401004010040100401004010040100401004010040100401004010040",
INIT_19 => X"00000000000000000000000000001000802FFFFFFFFFFFFFFFFF810040100401",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024,               -- Port A enable input
WEA      => wbe_a_hi_1024(3),               -- Port A write enable input
DIA(0)   => data_write_a(31),        -- Port A data input
DOA(0)   => data_read_a_hi_1024(31),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024,               -- Port B enable input
WEB      => wbe_b_hi_1024(3),               -- Port B write enable input
DIB(0)   => data_write_b(31),        -- Port B data input
DOB(0)   => data_read_b_hi_1024(31),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_0_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"ED39BA795990D275FB4A6E96ACC4731DEA4598B0AFB54867F6EE4618C3749803",
INIT_01 => X"8AA0047D8607944AC7DA180001ECA2444042106208408208C20022E9173734B3",
INIT_02 => X"1A7DDD79F9A73E6CCA7DAAF00001000008478020113D98E382FEDF333027C80F",
INIT_03 => X"75D341110C58F31110C58F32A208921F8051500147A0E4AB3493FB3A01EBE240",
INIT_04 => X"86424001531009B100425A97B2AA0001E03501D0A39C8F0078420001106D0C4C",
INIT_05 => X"BCC8CA2EBF03400700402BB20F00239E20341699198600000B08694B16434804",
INIT_06 => X"103FB860B2800161F8432200012DA185F80F24081C3C0707800E600056881308",
INIT_07 => X"B24197ABCDA467F9A73E6CCAFDC3870EEEEC44E2BDFE220094D03022210C011C",
INIT_08 => X"240581B5695EAA80262C080032BF07C7C1FC3F8E94F65B11555EAFFC1C306758",
INIT_09 => X"7E40000BEC004170040DB60017FED1CC0001045002984202003DB931192D60A5",
INIT_0A => X"120071411A74315881A28C141118000C5A85A60444210123820B43B40804674D",
INIT_0B => X"0820008E514045BB514F0106D1D8599581D3A958BC104A89215AC14C48898403",
INIT_0C => X"C261C01C48B1584A0CA3E2687A9A1E2687A9A1E2687A9A1E26870CD061343885",
INIT_0D => X"D274E93A758FA8683AC54B287522E10A74AF4AA59C568752662F5AC218000002",
INIT_0E => X"FF83C002783A0904231C70470C7E0B92800224008AE09FAD4BD48D1FC5D3A4E9",
INIT_0F => X"5BFF078004F075885DFBF7E15C06101C55E921F1F80FAB7FE0F0009E0E903EAD",
INIT_10 => X"F12E0380231F13978FF023FAFDBD9870380230F2D6081F56FFC1E0013C1D207D",
INIT_11 => X"DE7F263C0C8700125C0F8F3C43F1F10BBF7EFC61E01804E1E6C8F8FE807F67FB",
INIT_12 => X"02BE00017C17C1007E5E2E3081C5AC007E6F0E3081C5AC44418D65FE45DEE55B",
INIT_13 => X"61E0042786F103E9F01F9BC3C120C5A703E9F01F978B8C20666703E9F8A0FFED",
INIT_14 => X"FA7E283FFB414F80005F05F10FA7E283F78F6511C048278DCA174FF038FF15B4",
INIT_15 => X"0066A20B61692F293185D8D724E15D3FCC6B7C236FE0691B0700132C1F0EF880",
INIT_16 => X"3A4E93A4E93A4E93A4E93A4E93A4E93A4F942F92E9628540AD2A91442525A000",
INIT_17 => X"A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E9",
INIT_18 => X"4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93",
INIT_19 => X"55F3898E09B56C74DAB15D1CF13501AA495000000000000000003A4E93A4E93A",
INIT_1A => X"082082082082082082082082082082082082082082082082082084E41DC71C71",
INIT_1B => X"E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F82082",
INIT_1C => X"FFFFFFFFFFFFFFF94A5294A5294A5294A5294A52800003E1F0F87C3E1F0F87C3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"3060C183060C187FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"BDEBA0000000000000000000000000000000000000000000003060C183060C18",
INIT_28 => X"168ABA002E82145085155545F7AA975EFFFAABDE00FFAEBDFFF5D2EAAAAAF7AE",
INIT_29 => X"7FFFE10005542145557FD5545FF8000155087FC0155F7D168B55007BFDF45085",
INIT_2A => X"7FFC0010080017555555568AAAFFFFD7545AA8028A00A2802AABAFF8028BEF5D",
INIT_2B => X"FF842AABAA2AE95545FFD168ABAF7AEAAAAAA2FFFDF4500043FE105D2E954BAF",
INIT_2C => X"5007FD7400550415410002E974BA5D5168A00A2D142155005142010FFAE820AA",
INIT_2D => X"FFF780000BA007FE8AAAFF803FFFF5D2A821550000000BA007FD55FF5D7FC014",
INIT_2E => X"000AAFBEAA00007BFDFFF082EBDF455D5142000082E82145FFD17DFEFFFD168B",
INIT_2F => X"DFD75D2AA8A80EA8E2FE3F000000000000000000000000000000000000000000",
INIT_30 => X"68B551475FAF6D1C556F0AA1C24AABEA495FC716F002A975FFE3AA95E00EBAEB",
INIT_31 => X"42A0070071C50BAFEF1FAE0016D56A16D557BC257D415E0216FA3F1E8FC0145B",
INIT_32 => X"8010E004924874825D7FEAA85487FD24AFE3D02DAAAE12BD5545A2803AA00005",
INIT_33 => X"120155EA568E870BAEB8A05A2AEA8B50F55A2F150005A3A438BD04AFAB8F550A",
INIT_34 => X"545E055FFBE81D0BE8EA8A3AA05A2A5504001C74BA42A1571E8028E3DB7816D0",
INIT_35 => X"A5C7E3DFFFE90B45B47ABA497A82FFAFD2A82485FD2415A105C21451ED42A002",
INIT_36 => X"00000000000000000000B55EAAA100AA1D0F6F480B6A555A2A57A002A3D5FDB6",
INIT_37 => X"5EFAAAAB5E1AF3AABFF45592E88A0AFE80A8B0A0000000000000000000000000",
INIT_38 => X"65F520EBE9EF67D7BEA1FD5D556ABEF5D557FEBA55022A3F70C6B405F4D2AE97",
INIT_39 => X"C114728007521170821CE0FDE69411A8DED57CE1055555E5F58EFFC01FE2CACB",
INIT_3A => X"42341D5DEEBEF55080034E0A592A4AD0079C75D6070CC5CBB0280C029ABAA3EB",
INIT_3B => X"7F353AAF6C77F7F20D968BF57812A95E02A2AAB5EB0F280800EFAEE9F5D18F31",
INIT_3C => X"C91565455C141E41887D58AC448B69C30E02116220415A9540AA854140A0A204",
INIT_3D => X"DE6BE93172D7D625B556EEAB157ABEBE1B4D792A4AD1183454180DD3FDCAAAB7",
INIT_3E => X"F0000001FF0000001FF0000001FF0000001FF01EABC4B8014174FF7DA80F52FE",
INIT_3F => X"FF0000001FF0000001FF0000001FF0000001FF0000001FF0000001FF0000001F")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_2,               -- Port A enable input
WEA      => wbe_a_lo_1024_2(0),               -- Port A write enable input
DIA(0)   => data_write_a(0),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_2(0),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_2,               -- Port B enable input
WEB      => wbe_b_lo_1024_2(0),               -- Port B write enable input
DIB(0)   => data_write_b(0),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_2(0),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_1_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"212C001411984004084D000508C53810A03D1450E839B003342114428A000803",
INIT_01 => X"00000019400B100A8196000000CC004400400002000000000000028001340000",
INIT_02 => X"052137AE8031800C0044009000000000061800001CD4019802AD04CCCFC20004",
INIT_03 => X"04514108C60C21008C6042108400000201440020505100000043C30E10E9F000",
INIT_04 => X"02104001011DEFE088805681920000008000004001900800004002108C280008",
INIT_05 => X"040002340105000200000000080001900010000108040000000008411600401C",
INIT_06 => X"1034001042800808201000000001000820020000102000040000000000800180",
INIT_07 => X"64BF81A15EDFDE8031800C00843060C19E030022103600000450020800040004",
INIT_08 => X"00008004691687AA840008000090248CC84E000046000311555521F183060AC5",
INIT_09 => X"0820800D08100171000DB000154440C800400500000852020011200201012021",
INIT_0A => X"02000040001000880A2A04445004000102002041000001008208001440004140",
INIT_0B => X"4820018A1140440078050040511000102000A008183000010002404400000000",
INIT_0C => X"1000C80008000C030030880C2A030A00C28030A80C2A030A00C28018D4061401",
INIT_0D => X"10040802050080200284401C0022880F009E08008205C0020118088018000000",
INIT_0E => X"0F03C00280000000420860C60C0C0B92C0000000004000010042000040102008",
INIT_0F => X"001E078005000108400005E11C0610000000288058000003C0F000A000100000",
INIT_10 => X"F10E0380000000C202300000008D187038000000480800000781E00140002000",
INIT_11 => X"806302380C870010000004400100110800007861E0180000000C400680000001",
INIT_12 => X"023E00000000018000580C308000050000610C30800005000215006800000101",
INIT_13 => X"61E0000000018100B0001843812000014100B00016030C20000141002880026D",
INIT_14 => X"400A20009B404F80000000018400A20044096111C04000000304026000501580",
INIT_15 => X"0046820040082300218450C2800010094000482141E060190700100000002200",
INIT_16 => X"020080200802008020080200802008020080008008600500A82A1100A8000000",
INIT_17 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_18 => X"0080200802008020080200802008020080200802008020080200802008020080",
INIT_19 => X"81328A46BABEFC54A0810C7452B4428A14000000000000000000020080200802",
INIT_1A => X"AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA28A28A28A28A2A8218D2C0C924925",
INIT_1B => X"E974BA5D2E974BA5D2E974BA5D2E974BA5D2E975BADD6EB75BADD6EB75BAAAAA",
INIT_1C => X"FFFFFFFFFFFFFFFD8C6318C6318C6318C6318C63000002E974BA5D2E974BA5D2",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"70E1C3870E1C387FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"5555500000000000000000000000000000000000000000000070E1C3870E1C38",
INIT_28 => X"EBDF455D2EAABEFF7FFE8BFF5D0002155557FFFFFF007FC21EFA2FFD74AAAAD5",
INIT_29 => X"AA95400552AAAABAFFD1574105D7FD75FFAAAA800AAF7AA974BAFFFBE8B45F7A",
INIT_2A => X"0517DF555D2EAAA1055000015500557DF45AAD1400BAA2AE801550051555EFF7",
INIT_2B => X"FFD540155557FD5400F78028BFFFFFBEAB55F780020AAAA80020AA082EAAB550",
INIT_2C => X"AFF842ABEF5D517DF55552A974AAF7AE820AA0851574BAA2D1574AA5D7BFDEBA",
INIT_2D => X"EFAAD1575EF557FFFE10557FFFFFFFFD56AAAAFFFFD7555AAD168B45AAAEAAAB",
INIT_2E => X"0005D7FFDF4500043FE105D2E954BAF7AE80010082A97410557FEABFFAAFBE8B",
INIT_2F => X"51C7A2FBD5490BFD1C056A000000000000000000000000000000000000000000",
INIT_30 => X"974BAF7FFEFB45FFAABDF55492AA8BC2EBDFEAF7F1F840017D4975D2FEF147FC",
INIT_31 => X"080BEF495FC71D54124924385FAAA8AAAE3D145410F7F1D55D71C002DABAEBAA",
INIT_32 => X"002D082082AB8B6DBEDB7DF7F540E2AE85028B40155145F7AF6DBED5450AA1C2",
INIT_33 => X"78E021FF1471FDEAAFFD56F16D5571D2E28E38E0216FA2D1E8E80140F45082B4",
INIT_34 => X"A2DA3FB7DAAD4AAAAF487BC70BFA97F7AF6D417E92482BF84020BA495557E3FF",
INIT_35 => X"55554ADBD7A2FFC7BEFF6FFD7FC7002FD74951D71EDFFABFD16FAAAE92BD5545",
INIT_36 => X"00000000000000000000547AB8F550A8010E00492487482FFFE82A85EBAE2FFC",
INIT_37 => X"1EF005162BEF047FD5545AAFBF7400FBF9424F70000000000000000000000000",
INIT_38 => X"714F8338AAAA1D0AE974AAF7FFFDF55F7AABFF55082CA8B4DF6C1E8F5E540002",
INIT_39 => X"EABEF75550ACBB7582225FF5843404547184164AA5D2EBEEB0A2D555410D3555",
INIT_3A => X"FEAAEB083BC1000FF8409000512AEABFFDF79DCBF755962010BDCBBC21455D7F",
INIT_3B => X"801F8BA0C57740BDAA0688E5405D57D412F7D55F5E50C7F401BAAE8403CF5A3F",
INIT_3C => X"5D16BABAA3EBC3157ABD5FFE55F2AA9FEAFDF7F431A9F7FFE81FF013A8001AFF",
INIT_3D => X"FB863550229BCABEB7DA403FFFDA2FBF7FED2C7F955445079E280A00C56145EF",
INIT_3E => X"0000000000000000000000000000000000000596EBEF55080034E0A592A4AD00",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_2,               -- Port A enable input
WEA      => wbe_a_lo_1024_2(0),               -- Port A write enable input
DIA(0)   => data_write_a(1),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_2(1),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_2,               -- Port B enable input
WEB      => wbe_b_lo_1024_2(0),               -- Port B write enable input
DIB(0)   => data_write_b(1),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_2(1),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_2_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10E006600180111284380310006289800480032283E000A34301002001A0817",
INIT_01 => X"0005A00810790848048044A54E404350404000720885800802000906E4910200",
INIT_02 => X"407004208400408044C600C50AA055254010541A110222841200000002402544",
INIT_03 => X"0600011004182401004102408C28414043101000408118000145840440F5C415",
INIT_04 => X"5035855703A2900A000CD3088400F40688C9844409060850925E58A4081A0221",
INIT_05 => X"0200840D1021A15AC50494894850890540D1E12020C6E510818500440A280090",
INIT_06 => X"113044094002801020440090A8011A1224AB9380552102442884882A20004097",
INIT_07 => X"000100880004428400408044860000008C022402102100AA40004404B5075460",
INIT_08 => X"15C23440408C862A2A12382A8A5244145048C06085008010141521F000001240",
INIT_09 => X"400582B9033AA0E7AA4110B0506744810554542450694E710A836188C2C00222",
INIT_0A => X"443518360012C2210B020414109130A28038188096A06B8C120CA440A9C00802",
INIT_0B => X"1345E53300EC68005605002964AF222A5704004D080211121C80024200821780",
INIT_0C => X"181080C1110C882202211488452213C88472213C88472213488441109A442231",
INIT_0D => X"008204440210091341208041000810C00000300220201800A908000038AD0284",
INIT_0E => X"00040002804180300E88D28D206A40000554815500481440300000C44A081100",
INIT_0F => X"000008000500828700000000010000000002380000A00000010000A010050000",
INIT_10 => X"00010000000004CA000214000000020000000000684280000002000140200500",
INIT_11 => X"000000000020000000000442100002840000000800000000010C000026000000",
INIT_12 => X"00000000000805A4800000000000152300000000000015801272000100210020",
INIT_13 => X"000000000101C00000C000000000000940000120000000000009600004050000",
INIT_14 => X"0000130000000000000002018000106000000000000000002380000141000000",
INIT_15 => X"55000190000000000002000280000000011080C0000000000000000000002310",
INIT_16 => X"40902409064190641906419024090244902A9003004800415120D4A190804241",
INIT_17 => X"0900409004090641906419064190240902409024090641906419064190240902",
INIT_18 => X"9044090040900409004190441904419044090040900409004190441904419044",
INIT_19 => X"75960040138D70C030B51C50C7D100A2052F81F81F83F03F03F0419044190441",
INIT_1A => X"0410410410410410410410410410410410410410410410410248602081659659",
INIT_1B => X"5128944A25128944A25128944A25128944A25128944A25128944A25128941041",
INIT_1C => X"FFFFFFFFFFFFFFFE1084210842108421084210843FFF825128944A25128944A2",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"7FD5FF555815607FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"2AA000000000000000000000000000000000000000000000007FD5FF55581560",
INIT_28 => X"FC21EFA2FFD75EFAA8415410AA8415555087BFFF55A2AA800BAFFAE954000800",
INIT_29 => X"84155EFA2AEBDEAAA2FBEAABA5D7FE8B555551421455D0002145552EBFEBA007",
INIT_2A => X"2AEBDF555D2E954BAA2AA974BAFFFFE8B45552EBDF45FFAEAABFFF7FFE8B55F7",
INIT_2B => X"AAAAAAAAAFFD1574105D7FFFF555D2AAAAAA5D2E820BAA2FBEAB5555557DF55A",
INIT_2C => X"50055575EFFF84021555D043DEAA5D04021EF557FC21FFAA8428BFFAAAA954AA",
INIT_2D => X"10085568A00FF80175FFA2D17DFEFF7800215500557DF55AA80001FFAA800015",
INIT_2E => X"0005D00020AAAA80020AA082EAAB5500517DF555D042AA10A284154005D00154",
INIT_2F => X"00AAFFAA9543A080038A2A000000000000000000000000000000000000000000",
INIT_30 => X"0017D5D20B8EAA007FC51C7A2FBD55D2BE800042AFE8E1557D0075D2F45BEAA8",
INIT_31 => X"AA8BC7EBDFEAFEFFD00105FFBC20BDEAAA2FBF8AAA557BE8B6D5D5FFABEF4904",
INIT_32 => X"FFEFB6D555578F7DB6A0BDF7D480E174BFA02A974BAF7F5EFB455D2ABDF55492",
INIT_33 => X"ED1FDE90E3A497492B6AAADAAAE3D155E105571D55D71C002DABA5524820BAB6",
INIT_34 => X"BE8F401D7B6A0001470155C51D0092A071555D5E3AE821D00001FF0871C016DB",
INIT_35 => X"5BE8555400550A38428007FED000E3DA3DFD5E3DFFFBD5A38A021551C5F7AF6D",
INIT_36 => X"00000000000000000000410F45082B4002D082082AB8B6D1C5B7DF7FF78E075C",
INIT_37 => X"5EF005560B55F7AA800AAF7AA954AA00042AAA20000000000000000000000000",
INIT_38 => X"ABEF057D68F5F5A00021EF55042AAAA007FD5555AAFBD7545FBB8020A3F7AE97",
INIT_39 => X"7DF55D7AABFF5428ACA8F45A6C1E8F5EFF84165EFF7802BAB0A2FFEAABA557BE",
INIT_3A => X"CA8AA80800020AAF7FBFFFEF04552ABFFFF841FFE75CA882108202E974AAF7D5",
INIT_3B => X"00151FF0C57401E5F3D1E00A1A884174A8FFAEBFEB0A2D55541051555694F002",
INIT_3C => X"2AA801455D7FE8BFFF680800FFF7AAA155F595542455512A975455D3AA8A0055",
INIT_3D => X"5D79FCAF774AE005BE7895554005D2A8A0B882FFFFE10AAAAAB755A66B6AF56A",
INIT_3E => X"00000000000000000000000000000000000000C3BC1000FF8409000512AEABFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_2,               -- Port A enable input
WEA      => wbe_a_lo_1024_2(0),               -- Port A write enable input
DIA(0)   => data_write_a(2),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_2(2),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_2,               -- Port B enable input
WEB      => wbe_b_lo_1024_2(0),               -- Port B write enable input
DIB(0)   => data_write_b(2),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_2(2),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_3_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"210C00A20020000108430020001600B8156021104940741B3530400E02B92203",
INIT_01 => X"014C9BCA58B1296D24A402C992500B69404040028804A0080A000416A8D90A08",
INIT_02 => X"C12026A484318004404405C9C66E331352180D468B8203980300204442E02B34",
INIT_03 => X"04000748D60D24648D60524C88804D0215011020D15018148040C10A70E1D58C",
INIT_04 => X"18283333240FE41244187308C9104D70944852640901083801750EB0A418C220",
INIT_05 => X"0613142D01912CC2A1B4140528348900C612A104201C689044340ED413A07649",
INIT_06 => X"119000034019881822104C5E68035250A222829710A0A02C18C01A9920842413",
INIT_07 => X"402F00AB0016CA0431800444841020509D038B021230C1990001C644C8273200",
INIT_08 => X"16905000408482088290E8E64010248C4A5AA840C2000110001521F0810A92E7",
INIT_09 => X"0003CE6581BD016342A951AB146C4480530C3B2A8088D3542651670200C1826A",
INIT_0A => X"00735D36209A8A20020894004284B660821030C8990467401218004041020002",
INIT_0B => X"512445B740457154562F957CC08B00093700080D0A4851001D8302D20A0A1530",
INIT_0C => X"00508650008008021021A40861021840869021A408610218C0869810D6043095",
INIT_0D => X"1C8508438450801043A08090380A8834207007022209038080190000999C8F84",
INIT_0E => X"000400200000C0002A48A206204C4205F3304B33004C0041006240140A1C310A",
INIT_0F => X"0000080040000083800400000100000000008400018040000100080000510100",
INIT_10 => X"0001000000000800000244040000020000000100002A0080000200100000A702",
INIT_11 => X"000000000020000000200000080002C000800008000000000022000006808000",
INIT_12 => X"0000000000000A2281000000000040A3810000000000402001400000022002A0",
INIT_13 => X"000000000004200001C0400000000010200001C0400000000010000004490010",
INIT_14 => X"0001070004000000000000060000104C08000000000000001000000903008000",
INIT_15 => X"CC004050CA0C00020220200070040000010401C4000000000000000000100008",
INIT_16 => X"4310E4310A4210A4210A4210A4210A4210A8D0830A68010001B4DA881048061C",
INIT_17 => X"21084290A4210A4210A4210A4210A4210A4210A4210E4310E4310E4310E4310E",
INIT_18 => X"90A421084290A421084390E4310C4390E4310C4390E4310C4290A421084290A4",
INIT_19 => X"015303C0C78C706428A14C586291000A044001FFE000003FFC004290A4210842",
INIT_1A => X"2492492492492492492492492492492492410410410410412821600001249249",
INIT_1B => X"51A8D46A351A8D46A351A8D46A351A8D46A351A9D4EA753A9D4EA753A9D49249",
INIT_1C => X"FFFFFFFFFFFFFFFC00000000000000000000000038F56351A8D46A351A8D46A3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"55AB02055AB0207FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"420000000000000000000000000000000000000000000000007FFFAB57FFFAB5",
INIT_28 => X"A800BAFFAE9554508002AA00AA843DF55FFAA955EFA2D168B55557BEAA000055",
INIT_29 => X"002AB55AAAA955EF005568A00087BE8BFFA2D155410AA8415555087BFFF55A2A",
INIT_2A => X"AAABFF5508003FF555D0002145552ABFEBA007FC21EF007FD75FFAA841541008",
INIT_2B => X"082EBDEAAA2FBEAABA5D7FC0155005168B455D042AB45F7FFD741000042AA10A",
INIT_2C => X"FF7FBEAB55F7AABDEBA5D7FC2010A2D1575FFF7AA975555D2E80145F78415545",
INIT_2D => X"EF5555554AA087BC01FFFFAAAAB55552A954BAFFFFE8B55552EBDE00F7AEAABF",
INIT_2E => X"000082E820BAA2FBEAB5555557DF55A2AEBDF555D2E954BA002EAAABA002A821",
INIT_2F => X"FB7D5D7FEAA3808554203A000000000000000000000000000000000000000000",
INIT_30 => X"1557D1475FAF45BEAA800AAFFAA95578080038A2AA28E3AF55E3A0BA5D7AADB6",
INIT_31 => X"BD55D7BE80004AA1E8E2AB55B6A0925D7085F6AA10087FEABD7AAD57AEBAB68E",
INIT_32 => X"F5D0438140E2FA38B6AEBFF6D1D04AAFFA41040017D5D20B8EAA007FC51C7A2F",
INIT_33 => X"D0A901FFFF801557D1C20B8EAAA2FBE80AA557BE8B6D5D5FFABEF49002FB55FF",
INIT_34 => X"5D20BDE00EBAAA8BC7EBDFEAFEFAB8ABAE925D21C7010EADB525D7FFAE975C75",
INIT_35 => X"F002EADA921420871D74971D24820875C21D5EB8AA8FFF012A954BAFFF5EFB45",
INIT_36 => X"000000000000000000001C24820BAB6FFEFB6D555578F7DB6A0BDF7DEB8E125F",
INIT_37 => X"B55A28408145AAFFFFFFF5D7FEAABA0051400A20000000000000000000000000",
INIT_38 => X"AB55FAD568AA2AFAE975EF555168B55F7AA800BAF7AA955EF00042AAA2A2AEAA",
INIT_39 => X"2AAAA007FD55558A7BD7145FBB8020A35D2ABEF55F7800015F087FEAA00007FE",
INIT_3A => X"968F575D003FF55F7D5420BA5D2ABFEAAF7AE9DFF759A82AEF70800021EF5504",
INIT_3B => X"FFD5145FBAC9755F05040255FFD84175EF55002AAB0A2FFEAABA557BEA3EF057",
INIT_3C => X"82E974AAF7D57DF45552A3FF10AA8429F45A7D5EAF5FFBAEAAA10554155400AA",
INIT_3D => X"FF843FFE77C80825BC052ABFE10550415557085540000005156155FE90A8F5C0",
INIT_3E => X"00000000000000000000000000000000000005500020AAF7FBFFFEF04552ABFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_2,               -- Port A enable input
WEA      => wbe_a_lo_1024_2(0),               -- Port A write enable input
DIA(0)   => data_write_a(3),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_2(3),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_2,               -- Port B enable input
WEB      => wbe_b_lo_1024_2(0),               -- Port B write enable input
DIB(0)   => data_write_b(3),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_2(3),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_4_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"A108400020612C80284210081034849800A00030300004833522C82D04A16002",
INIT_01 => X"2043998A1839284D1CA0650E1E504368403008418984014902030806A0D10200",
INIT_02 => X"C120042200000000044441CE01E80F00A49043118680008002000000026208E4",
INIT_03 => X"040001020019200020011209CC0164C060000000690111040144800042F5C403",
INIT_04 => X"7029AF0F81A00010CCA47700CC513CAC0D0B8E02010740E19754080108988021",
INIT_05 => X"02139405007133C0712244CD20F20105D583000020E9892201D304D42A9835E1",
INIT_06 => X"9190440300078002014405D9EE814C0284A883B6D7038AE079059B7800048092",
INIT_07 => X"000100AA0004408000000004840400008D200102503000782000C00C8025C000",
INIT_08 => X"00728A00408403220811991E02120C044058080004000001101121F220000260",
INIT_09 => X"811001E1185B38AD23C3707AD46440818F3CF80EC423CA7D01D123C80200816A",
INIT_0A => X"45810810A01B40216361056D6150F41200280001900439001FD8A00041400000",
INIT_0B => X"11FC88076266E800D605402962A820211500024808010512C40106D222223B14",
INIT_0C => X"0408804116040B02C02C500B0C02C100B0C02C100B0402C300B0401618058611",
INIT_0D => X"040200050200501301208482200D00D0A0408402C4282200A84800009B878680",
INIT_0E => X"00000020000100024AC88300300060090F0D830F00025400300204D018000804",
INIT_0F => X"8000000040000206A2000800000000000000950002E010000000080000588040",
INIT_10 => X"0000000000000808000554000200000000000100006D0020000000100000BB00",
INIT_11 => X"0000400000000000002000001A0002504001000000000000002280000D800800",
INIT_12 => X"0800000000000E2C802000000000408D801000000000408012440000200110A0",
INIT_13 => X"000000000004680003A0040000000010280003800800000000102800000B0000",
INIT_14 => X"000005C0002000000000000620000158000010000000000010A0000B00000200",
INIT_15 => X"C30146200400104002602600400000000294004000000004000000000010001A",
INIT_16 => X"0080200000008020000000802000000080080000004090014134DA101288C6DB",
INIT_17 => X"0802000000000401806010040180601004018060100000802000000080200000",
INIT_18 => X"8060180601004010040080200802000000000000802008020000000000008020",
INIT_19 => X"C0A28A063807E0500014063450404882846FFE000003FFC00000010040100401",
INIT_1A => X"AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA28A28A28A28A2934C8D0CCD145144",
INIT_1B => X"68341A0D068341A0D068341A0D068341A0D068351A8D46A351A8D46A351AAAAA",
INIT_1C => X"FFFFFFFFFFFFFFFC0000000000000000000000001FE32068341A0D068341A0D0",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"408102040810207FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"800AA00000000000000000000000000000000000000000000040810204081020",
INIT_28 => X"168B55557BEAB4500554200000557FE10FFFBEAA10007FD7410FFAA97555082A",
INIT_29 => X"55574105D2A800AA00043FEBA5D7FEAA00007BE8AAAAA843DF55FFAA955EFA2D",
INIT_2A => X"57BC00AAA2FFEAAAAAA8415555087BFFF55A2AA800BAFFAE9555508002AA0000",
INIT_2B => X"A2AA955EF005568A00087BE8BFFA2D17DE1000517FE10AAAAA8AAA002E975455",
INIT_2C => X"FAA8417410A2D140000F7FBC2010A2D157400AAAE974AAAAAA974BA08002AB55",
INIT_2D => X"EFA2AABDEAA087BEAAAAA2FBD54BA080002145552ABFEAA007FC21EF007FD75F",
INIT_2E => X"00055042AB45F7FFD741000042AA10AAAABFF5508003FF55F7D568A00552EA8B",
INIT_2F => X"5400F7A49057D0824850B8000000000000000000000000000000000000000000",
INIT_30 => X"3AF55F7A0925D7AADB6FB7D5D7FEAB7808554203A145178E00FFFBE8A101475D",
INIT_31 => X"A9557D080038AAA145157428492E8008200043FE925571EFA380871C7028A28E",
INIT_32 => X"AEA8A9200249056D4175C5092AAF5FDA38BE8E1557D1475FAF45BEAA800AAFFA",
INIT_33 => X"AA4954281C0E2FB55B6A0925D7085F6AA10087FEABD7AAD57AEBA08517DE00AA",
INIT_34 => X"007FC51C7007BD55D7BE80004AAFEDB42028EBFBC2028BED152438AAA092492A",
INIT_35 => X"AF7DF6AA00412EAABFFAA803DEBA0875EDA80BEF1C743840040017D5520B8EAA",
INIT_36 => X"0000000000000000000041002FB55FFF5D0438140E2FA38B6AEBFF6DBE84AAEB",
INIT_37 => X"A00FFFFEAA105D5155410FF84021EF0800154B20000000000000000000000000",
INIT_38 => X"DEBA0851574B2AAAEAAB55F78400145AAFFFFFEF5D7FEABFF0051400A25D5568",
INIT_39 => X"68B55F7AA800BAF7AA955EF00042AAA25555410BA082E8201000043FE005D517",
INIT_3A => X"568AA200557DE00AAAAAAA000804001FF005575408AA557FEB2FFAE975EF5551",
INIT_3B => X"D1550AAAA8002010F2AC154B25F2ABFF55F7800015F087FEAA00007FEAB55FAD",
INIT_3C => X"800021EF55042AAAA007FD5555087BD6145FAAC000A2A6FBC00BAAAFBC00BAF7",
INIT_3D => X"F7AEBDFF779A82AA43F7FBE8A00082EA8BFFAA843FEBA08517DE00F3F9574B30",
INIT_3E => X"000000000000000000000000000000000000008003FF55F7D5420BA5D2ABFEAA",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_2,               -- Port A enable input
WEA      => wbe_a_lo_1024_2(0),               -- Port A write enable input
DIA(0)   => data_write_a(4),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_2(4),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_2,               -- Port B enable input
WEB      => wbe_b_lo_1024_2(0),               -- Port B write enable input
DIB(0)   => data_write_b(4),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_2(4),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_5_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50DF4A0791B3FCB694379283C81FD996A091832102004A336A20E03C040C002",
INIT_01 => X"805FBDC69830A84D5C6A60000C34C26841280A00084000C8C212892EEAD53235",
INIT_02 => X"3B2026B578918E640A4F01CF8011FF0002080000082CA9998276DF7772C7C80D",
INIT_03 => X"37134108420D700084205702A4008A1D9100002171C0E0051554D93A11F5D140",
INIT_04 => X"8A41A0FC03A56DA000425A819410E3816C086198A388B702A8CA1210844A0C4C",
INIT_05 => X"B1808A062E8BC835F5E84532D708238A282F00A9291224800A2861490343082C",
INIT_06 => X"903FB8483A90581859050424100940825C6184401CDC451B860A6507160C4100",
INIT_07 => X"D26F068BCC96CDF8918E640E96D1A3469D6300E2FFEA27F8E4D23248130E259C",
INIT_08 => X"0BFA82E568442B2A082C0A7E3014250D49DA37A2420619000002AFF48D1222E5",
INIT_09 => X"3F005001E40969289429360416DCD1C46083030604B1CA20C03DF83B0A2C60A5",
INIT_0A => X"14613C71005A10492B888120288F480D58858449026145B3830F449449062B4F",
INIT_0B => X"11AC04934AC648BFD727C031E64170A137D5AA5C3E4B0F8A3C58C34C002290E3",
INIT_0C => X"CA29C6CC50384B6AC6AC86AB31AACA6AB39AAC86AB39AACA6AB3055643559C31",
INIT_0D => X"C673E33CF28F38603855401985228A0614BD30A0A2819852011E5AC2B87F9182",
INIT_0E => X"FF87C002F87A803E460B2516510CA594FF0044FFA4B08BAC4BB2CD0F09CF84E3",
INIT_0F => X"0DFF0F8005F0F5100DFFF5E15D06101C55EB29F1E00BE53FE1F000BE1E802F94",
INIT_10 => X"F12F0380231F17D78FC029FFF58D9A70380230F2FE0017C37FC3E0017C3D005F",
INIT_11 => X"FC7F023C0CA700125C0F8F7E43F1F001BFFE7C69E01804E1E7CCF8FC003FF5F1",
INIT_12 => X"023E00017C1FC1A4BFD82C3081C5BD27BFE30C3081C5BD00C02365D645CEEF5B",
INIT_13 => X"61E0042787F181E9C1EFD8CB8120C5AF41E9C18FD60F0C20666F41E9F009FFFD",
INIT_14 => X"7A7C077FFF404F80005F07F187A7D14BFFC96111C048278DEB074F9930FF9D80",
INIT_15 => X"C064014B8B652E2B3120C81284641D3E8DBF7D636FE860190700132C1F0EFB80",
INIT_16 => X"38CE1384E3384E338CE138CE1384E33C4E3ECE32E128882551349A1CBAA44103",
INIT_17 => X"84E3384E3384E3384E338CE138CE1384E3384E338CE138CE1384E3384E338CE1",
INIT_18 => X"CE138CE138CE138CE1384E3384E3384E3384E338CE138CE138CE138CE1384E33",
INIT_19 => X"F5E5BB4E7F7B9DB7FF3A1B6DB7E8410A8C000000000000000000384E3384E338",
INIT_1A => X"BEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEF9F7CFDFDDCF3CF3D",
INIT_1B => X"BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEFBEF",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000001711C7BBDDEEF77BBDDEEF77",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"FDFFF00000000000000000000000000000000000000000000080000000000000",
INIT_28 => X"FD7410FFAA97410082A800AAAAAE955450055421FFFFFBC0010AAD5574BA557F",
INIT_29 => X"7FD74000055574BA5D7FD7555A2D5575EF55517FF5500557FE10FFFBEAA10007",
INIT_2A => X"0002AABA5D2ABFFFFAA843DF55FFAA955EFA2D168B55557BEAB5500554200000",
INIT_2B => X"5D2A800AA00043FEBA5D7FEAA00007BC00AAAAAEBDF45A28428B45FFD168BFF0",
INIT_2C => X"5080028A00A2FFFDE00F7D57FEBAFF80174BAAAD1555EF555555555005557410",
INIT_2D => X"BA5D2E821FFA2D5554BA557BD75FFAA8415555087BFFF55A2AA800BAFFAE9555",
INIT_2E => X"00000517FE10AAAAA8AAA002E97545557BC00AAA2FFEAAAA082A97545F7D5420",
INIT_2F => X"7010BEDF524AA5571FDFEF000000000000000000000000000000000000000000",
INIT_30 => X"78E00EBFBE8A101475D5400F7A49043D0824850B8A2AE9756D145B401FFFFFFC",
INIT_31 => X"FEAB7D0855420BA1471D74380851524BA5571D757DB6D5525EF555178F6D1451",
INIT_32 => X"8A28B6DEBDF6DBEF1C0A28AAA5524BFFFFA28E3AF55F7A0925D7AADB6FB7D5D7",
INIT_33 => X"5555057D145152428492E8008200043FE925571EFA380871C7028B6AEBDF45B6",
INIT_34 => X"BEAA800AAFFAA9557D080038AAAA2FBF8E10EBD578EAAFF8415482BED1555EF5",
INIT_35 => X"81C209256DFFDF420BA552A821FFB6DF574A85575C55EFBE8E1557D1475FAF45",
INIT_36 => X"0000000000000000000008517DE00AAAEA8A9200249056D4175C50920875FDA3",
INIT_37 => X"5FF5D7BC21EFF7FBD7400F7FBC00BA55557DFF70000000000000000000000000",
INIT_38 => X"01FF5D5568BE7555568A00AAFFEAA105D5155410FF84020AA0800154B2AAAA97",
INIT_39 => X"00145AAFFFFFEF5D7FEABFF0051400A25551554BA0051400BA5551575EFF7D14",
INIT_3A => X"1574B2FFAABFF45FFAAAABFFAAFFFDFFF552EA8AAA55043DFF7AAAEAAB55F784",
INIT_3B => X"8002410FFD5575EF5555421E75555400BA082E8201000043FE005D517DEBA085",
INIT_3C => X"FAE975EF555168B55F7AA800BAF7AA955EF00002AAA2A2FBE8A00A2D16AAAAFF",
INIT_3D => X"0055554088A557FEB25D00021FFFFFFC00BA552A821EFFFFFD74BA5D51575F7F",
INIT_3E => X"000000000000000000000000000000000000000557DE00AAAAAAA000804001FF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_2,               -- Port A enable input
WEA      => wbe_a_lo_1024_2(0),               -- Port A write enable input
DIA(0)   => data_write_a(5),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_2(5),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_2,               -- Port B enable input
WEB      => wbe_b_lo_1024_2(0),               -- Port B write enable input
DIB(0)   => data_write_b(5),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_2(5),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_6_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10800B0061A01002840002C03002818000402322520070B313301C4389B2082",
INIT_01 => X"250041CA3839684D18A160000C52426841000000090800090210080008110200",
INIT_02 => X"0020042080010000044654C0000C008010000000001020900200200002620814",
INIT_03 => X"060881021088200021080200E4000A0891000020610111500104C00000F14400",
INIT_04 => X"0880000100000002000052288144004281C050400100280000C8100000080001",
INIT_05 => X"928080840001100A08009000280201000850E022401400002028214043410820",
INIT_06 => X"10100518090012122100C808049310002040000410A0001400000200120840D2",
INIT_07 => X"000100800004400001000000860408108C22000A502010074120044800040001",
INIT_08 => X"50000040D0C4E2088003FD01C01004044058082004000000000121F020408244",
INIT_09 => X"00BF17E9001205A5204911F814444080400100020000D200DFD16400C2A40AA0",
INIT_0A => X"04611C17849000022862A1596C8B5DF04834948900000100220C244840000880",
INIT_0B => X"03AD0413424E4044D665C070C22602291504400D084915020448114080201000",
INIT_0C => X"5E08864011088B22D22C008B0022C408B1022C208B0822C608B1111600458010",
INIT_0D => X"4251A12CD28A300429688001000800000020280204001000A00804309A002182",
INIT_0E => X"0000000280402400420800000000006200FC10002442042429324294014E8CA7",
INIT_0F => X"A40000000500800840000800000000000002280018001480000000A010100052",
INIT_10 => X"00000000000004C2003000010240000000000000680800290000000140202000",
INIT_11 => X"2000C0000000000000000442000001080001000000000000010C000280001804",
INIT_12 => X"08000000000801C300A010000000156000902000000015101200002800000000",
INIT_13 => X"000000000101800038002408000000094000386028040000000940000ED40000",
INIT_14 => X"0003B000002000000000020180002A24005010000000000023000060C7000A40",
INIT_15 => X"3F0280090321000040A410C28108000160008094000810040000000000002300",
INIT_16 => X"284A5284A728CA5284A528CA728CA52C4A5A0A32A300940101349A0408240818",
INIT_17 => X"9CA1294A329CA5284A728CA7284A5284A728CA5284A528CA728CA5284A728CA7",
INIT_18 => X"CA3294A129CA3294A129CA1294A329CA1294A3294A129CA3294A129CA3294A32",
INIT_19 => X"F5F78BCE7F8FF0F4FA955F7CF7F40A80145D55555556AAAAAAAAA94A329CA129",
INIT_1A => X"8E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E39B6CEDECDDF7DF7D",
INIT_1B => X"F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE38E3",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000001A1A33F9FCFE7F3F9FCFE7F3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"555FF00000000000000000000000000000000000000000000080000000000000",
INIT_28 => X"BC0010AAD5574BA557FFDFFF087BFDF45F7AA974AAAAAA97555F784174BAF7D5",
INIT_29 => X"515555508043FE00F7AA97555A2FBD7410AA8428AAAAAAE955450055421FFFFF",
INIT_2A => X"7D1575EFFFAA9555500557FE10FFFBEAA10007FD7410FFAA97400082A800AA08",
INIT_2B => X"0055574BA5D7FD7555A2D5575EF55517FF55A2AA97400552AAAB45082E80155F",
INIT_2C => X"500554200000003DE10FFD5401FFF7AAA8A10082EAAB45A2FFC2000007FD7400",
INIT_2D => X"10AA803FE105D516AABAFF843FFFFAA843DF55FFAA955EFA2D168B55557BEAB5",
INIT_2E => X"000AAAEBDF45A28428B45FFD168BFF00002AABA5D2ABFFFF087BD5545007BFDE",
INIT_2F => X"256DEB84104BAFFD1525FF000000000000000000000000000000000000000000",
INIT_30 => X"9756D145B401FFFFFFC7010BEDF524AA5571FDFEF1C7BFFF55FFA095482B6A49",
INIT_31 => X"4904380824850381C5B5057D1C003DE28F7A49057DAAF5D2428A2842AAAAA2AE",
INIT_32 => X"2AAFB451C2A8017DE3DF525FFFFA49756D145178E00EBFBE8A101475D5400F7A",
INIT_33 => X"2F1C50381471D74380851524BA5571D757DB6D5525EF555178F6DAAA49542841",
INIT_34 => X"AADB6FB7D5D7FEAB7D0855420BA1C0E3FE00E3DB471EFE3AAAAA00082EA8B6DA",
INIT_35 => X"F1C7BD057D1C71FFE10A28038E1049516AAB8FF8428FEFA28E3AF55F7A0925D7",
INIT_36 => X"00000000000000000000B6AEBDF45B68A28B6DEBDF6DBEF1C0A28AAA5524BFFF",
INIT_37 => X"F55F78017400F780001FFAA84000AAFFD1401E70000000000000000000000000",
INIT_38 => X"20BAAA8428AA2AAAA975FF5D7BC21EFF7FBD7400F7FBC00BA55557DFF7557BFD",
INIT_39 => X"EAA105D5155410FF84020AA0800154B2557FC01EF55043FEAAFF80021EFA2D14",
INIT_3A => X"568BE7AA80174AA082ABDF555D2A821EFAAFBC01FFF780155F7555568A00AAFF",
INIT_3B => X"AEA8A10082EA8BEFAAD5554B25551554BA0051400BA5551575EFF7D1401FF5D5",
INIT_3C => X"AAEAAB55F78400145AAFFFFFEF5D7FEABFF0051400A25D2EBFE10AAFFD55EFA2",
INIT_3D => X"552EA8AAA55043DFF7557BC01EF55557DE00AA842AA0000516AABAFF8428BE7A",
INIT_3E => X"0000000000000000000000000000000000000FFAABFF45FFAAAABFFAAFFFDFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_2,               -- Port A enable input
WEA      => wbe_a_lo_1024_2(0),               -- Port A write enable input
DIA(0)   => data_write_a(6),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_2(6),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_2,               -- Port B enable input
WEB      => wbe_b_lo_1024_2(0),               -- Port B write enable input
DIB(0)   => data_write_b(6),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_2(6),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_7_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10844B00482258A2842112C02450418800002300500030B313300C418992002",
INIT_01 => X"000009CA3839684D1CA0E0000E51424840000000080000080200080008510204",
INIT_02 => X"0120042086010000044600C00008000004100000000260900200000002402004",
INIT_03 => X"8628A10000082400000002408400080011000000610008000208C00000E14400",
INIT_04 => X"0911800100A000000000524084000040000050001140200100C8100000080102",
INIT_05 => X"0300812401011000000000002000114008008060441000000020024093000000",
INIT_06 => X"9190431C0D4010100000880804010010800000041080081000000200010424B2",
INIT_07 => X"000100AA0004408601000004860000008C02000A103010006928040800062481",
INIT_08 => X"84000048D484C20888000A0002120484C048007004000000000021F000000244",
INIT_09 => X"00A06009881201A520491004106C48A04040002400A15A208001650004001020",
INIT_0A => X"C99E1060201002044809C1040140A001004808810000459033189C0A400118A0",
INIT_0B => X"102000024040484050050041648A0041140C500B08821054C000264120000400",
INIT_0C => X"0404A083260E0832132011880462011880462051881462051881D31018C40620",
INIT_0D => X"0001000080001000813094801A8F80F00A600B52602801A88848011118003700",
INIT_0E => X"000003C007C002808228010410082042C000C000000004001002000400040002",
INIT_0F => X"A4000007800F80C840000800009864038A1200081C0014800000F001F0200052",
INIT_10 => X"00002C0E00E0E4004038000102400002C0E00E0D20100029000001E003E04000",
INIT_11 => X"2000C04031100E0403D0700300080908000100000661801E1900040380001804",
INIT_12 => X"0840878083E8003780A01043203A101780902043203A10082410082880000000",
INIT_13 => X"0601E0187900181035E0240806483248181035E0280410C8198818100DDD0000",
INIT_14 => X"0403774000201021E020FA006040376C00501022131210722060806D47000A40",
INIT_15 => X"00928A0002000110888600C032128201519480D40009902430160403E0E00506",
INIT_16 => X"01000000020080601802000000000405000A0020020081014134928820480010",
INIT_17 => X"0802018040000000006018020080200804010000000000806018020080000004",
INIT_18 => X"0000000001806008020000001006008020080001004008020080201004000020",
INIT_19 => X"0000000000000000000000000000400A004618618618C30C30C3000020180600",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000000B0840000000000000000000",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"1555500000000000000000000000000000000000000000000080000000000000",
INIT_28 => X"A97555F784174BAF7D5555FFF780155EFAAAEA8ABAAAFBFDE0055556AA005D04",
INIT_29 => X"55555EFAAFFFDFEFAAAAAAB455D556AA00FFAE95555087BFDF45F7AA974AAAAA",
INIT_2A => X"02EAAAAA082EA8A00AAAE955450055421FFFFFBC0010AAD5574BA557FFDFFF55",
INIT_2B => X"08043FE00F7AA97555A2FBD7410AA8428AAA557BFDFFF55003DFFFF7FBEAA000",
INIT_2C => X"0082A800AAF7AE975FFA28000010552EBDE00007BEAAAAA2D140000085155555",
INIT_2D => X"45087FEAB455D516AB55557BD55FF00557FE10FFFBEAA10007FD7410FFAA9740",
INIT_2E => X"000A2AA97400552AAAB45082E80155F7D1575EFFFAA955555D51574AAAAFFD55",
INIT_2F => X"AE105D556AA10410E17555000000000000000000000000000000000000000000",
INIT_30 => X"FFF55FFA095482B6A49256DEB84104BAFFD1525FFFF8E175C7A2AAAAA82A2F1F",
INIT_31 => X"F524AA5571FDFEF415B575D7AAF1FFFD7AAAAAFB7D495F6AA10E3AE905551C7B",
INIT_32 => X"003AFEFEBFBEAA001C2EA8A821C2EAAA00A2AE9756D145B401FFFFFFC7010BED",
INIT_33 => X"EDB470101C5B5057D1C003DE28F7A49057DAAF5D2428A2842AAAA497BFAFFF49",
INIT_34 => X"1475D5400F7A490438082485038F7A4905C7A28A070384120BDE100075EAA82B",
INIT_35 => X"D495150492BEF1D2555087BE8B7D555F6AB57417BC05D7145178E00EBFBE8A10",
INIT_36 => X"00000000000000000000AAA495428412AAFB451C2A8017DE3DF525FFFFA49756",
INIT_37 => X"555A2AEA8A10AAD568A00555168A10002E9754D0000000000000000000000000",
INIT_38 => X"8A10AAAE8215D557BFDF55F78017400F780001FFAA84000AAFFD1401E7FFAA97",
INIT_39 => X"C21EFF7FBD7400F7FBC00BA55557DFF7007BD5555AAD57DF55AAAEBDFEF007BE",
INIT_3A => X"428AA2007FE8BFF080028BFFAAFFEAA105D2EAAA005D2AAAA18AAAA975FF5D7B",
INIT_3B => X"043DE0000516AA10F7FBD7408557FC01EF55043FEAAFF80021EFA2D1420BAAA8",
INIT_3C => X"55568A00AAFFEAA105D5155410FF84020AA0800154B2FF8402145A2AA954AA00",
INIT_3D => X"AAFBC01FFF780155F7005140000FFD140145007FE8BEF557BEAB55087FC215D5",
INIT_3E => X"0000000000000000000000000000000000000AA80174AA082ABDF555D2A821EF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_2,               -- Port A enable input
WEA      => wbe_a_lo_1024_2(0),               -- Port A write enable input
DIA(0)   => data_write_a(7),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_2(7),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_2,               -- Port B enable input
WEB      => wbe_b_lo_1024_2(0),               -- Port B write enable input
DIB(0)   => data_write_b(7),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_2(7),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_8_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00000648E2840112C00000418000002700500030B3132000400812082",
INIT_01 => X"100008480009004C04A100000252024840000000180800080200010040110204",
INIT_02 => X"0020042000490000004600804008000005100000000024900200000002400004",
INIT_03 => X"0A0C33400008082400000080A4004B0891000020610112000040C00000E5C000",
INIT_04 => X"18800001000000000000512080000040800150400824280110C8100000120200",
INIT_05 => X"908084A10100100200004080280008240810802206940000012C214451610800",
INIT_06 => X"81B000080860109021400008040000202048020414A0021400040200322824C1",
INIT_07 => X"000000080004408049000004860000008402001A50208000630C040800062483",
INIT_08 => X"440000428644212280800A00021004044048002124000000000021F000000244",
INIT_09 => X"00004009001001010008100414644410400102228000D20080114502006409A2",
INIT_0A => X"000051312000042200294429148A4801C80C8C81000045907118040340020832",
INIT_0B => X"4020000240404140004D0544C4AA0001150410090302500011C813428A000400",
INIT_0C => X"46501090008820240240409000240009000240009000240009000120204808A5",
INIT_0D => X"42D1A168D09A301468402480004780F00140080860280004085904309A002196",
INIT_0E => X"00783FC00044340242280000000000020000C0000442106419120004034685A3",
INIT_0F => X"8000F07F800088A80000081EA2F9EC0000064004081010001E0FF00011104040",
INIT_10 => X"0ED0FC7E00000422201080000202658FC7E0000021882020003C1FE000222080",
INIT_11 => X"018059C3F350FE0C00000002A0040500000103961FE780000110010090000800",
INIT_12 => X"FD41FF80000830200021C1CF600012200010D1CF600012121600100810000004",
INIT_13 => X"9E1FE000010A1802100004343ED8000898021000087073D80008980200800002",
INIT_14 => X"0080200000BEB07FE00002086008020000209AEE3F300000246020200000620B",
INIT_15 => X"0088881903210000440610C8000A808040000208901786E4F0FE0C0000000166",
INIT_16 => X"685A1685A769DA368DA368DA769DA36CDA121A11A141800011309284002C0810",
INIT_17 => X"95A5685A1685A5695A368DA368DA769DA368DA368DA7695A1685A1685A5695A1",
INIT_18 => X"5A1695A568DA368DA369DA768DA1685A1695A5685A168DA369DA768DA368DA16",
INIT_19 => X"A4028A0A543EBC57A10A1E75D64108080468618618630C30C30C69DA5685A168",
INIT_1A => X"9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7BF3CCD8DF5B2DB2C",
INIT_1B => X"F87D3E1F4F87D3E1F4F87D3E1F4F87D3E1F4F87C3E1F0F87C3E1F0F87C3E79E7",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000006A6D4F87D3E1F4F87D3E1F4",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"155FF00000000000000000000000000000000000000000000080000000000000",
INIT_28 => X"BFDE0055556AA005D0415555080000000087BEAA10F7803DE00FFAEBFFFF0800",
INIT_29 => X"2AA8AAA557FC0010F780154105D7FC2145005155555F780155EFAAAEA8ABAAAF",
INIT_2A => X"7FFFFF55AA80155FF087BFDF45F7AA974AAAAAA97555F784174BAF7D5555FF55",
INIT_2B => X"AAFFFDFEFAAAAAAB455D556AA00FFAE95555AAFFE8A00552EBFE00F7D17FF45F",
INIT_2C => X"A557FFDFFF5504000AAAAAAA8B55F7D140010552E821EFAAAABDF555555555EF",
INIT_2D => X"55AA8028A00A2D57FF45557BE8A00AAAE955450055421FFFFFBC0010AAD5574B",
INIT_2E => X"000557BFDFFF55003DFFFF7FBEAA00002EAAAAA082EA8A00002AA8A10F784021",
INIT_2F => X"FE10F7AEBAFFF080A175D7000000000000000000000000000000000000000000",
INIT_30 => X"175C7A2AAAAA82A2F1FAE105D556AA10410E17555080E000280071E8A00EB8E3",
INIT_31 => X"4104BAFFD1525FF492EA8AAA5571C2000FF8A17400557FC015514555757DFF8E",
INIT_32 => X"2ABDE10EBDF7AF6DE3FFF8F7DB68A105D71C7BFFF55FFA095482B6A49256DEB8",
INIT_33 => X"AA0BDF6D415B575D7AAF1FFFD7AAAAAFB7D495F6AA10E3AE90555A2FBE8A3849",
INIT_34 => X"FFFFC7010BEDF524AA5571FDFEF550E00082B6A0AFB55F7D1420104124821D7A",
INIT_35 => X"01C2EA8A00F7800017DA2842FA00B6D578F6D557FFDA00A2AE9756D145B401FF",
INIT_36 => X"00000000000000000000497BFAFFF49003AFEFEBFBEAA001C2EA8A821C2EAAA0",
INIT_37 => X"0BA08556AA00AAAABFE00F7AEAABEF082E955450000000000000000000000000",
INIT_38 => X"21555D51575EFFFAA97555A2AEA8A10AAD568A00555168A10002E9754D082E82",
INIT_39 => X"17400F780001FFAA84000AAFFD1401E7082EAAABA5D5140010F7AE974105D7BC",
INIT_3A => X"E8215DA2FFE8ABA082ABFE00AAFBEABFFAAFBEABFFF7AA80145557BFDF55F780",
INIT_3B => X"D540000000402145AA843FFFF007BD5555AAD57DF55AAAEBDFEF007BE8A10AAA",
INIT_3C => X"AAA975FF5D7BC21EFF7FBD7400F7FBC00BA55557DFF75D2E82010F7843DF45FF",
INIT_3D => X"5D2EAAA005D2AAAA185D2AAAA10F780021FFA2803DE10FFD16ABFF5D7BFDE10A",
INIT_3E => X"0000000000000000000000000000000000000007FE8BFF080028BFFAAFFEAA10",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_2,               -- Port A enable input
WEA      => wbe_a_lo_1024_2(1),               -- Port A write enable input
DIA(0)   => data_write_a(8),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_2(8),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_2,               -- Port B enable input
WEB      => wbe_b_lo_1024_2(1),               -- Port B write enable input
DIB(0)   => data_write_b(8),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_2(8),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_9_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00018248A2840112C00002C18000002300500030B3132000400812006",
INIT_01 => X"400008000000004C0020000000100248413C0A61590001D90213C10008110204",
INIT_02 => X"01A0042080010000054600C04008000004100000001020900200200002420804",
INIT_03 => X"024003400008012400000010E4004B0891000020610310000144C00000F5C000",
INIT_04 => X"1801800100E000000000510084000040010050020810200000C8900000320200",
INIT_05 => X"918004311104100000000000200008100800002000100000002C234415610820",
INIT_06 => X"81B00008080010100000980804000008800042041080001000100200322C2481",
INIT_07 => X"0000811800044080010000058600000086020002502080006000040800062C80",
INIT_08 => X"0000004001D4618008800A00061004044048002004000000000061F000000244",
INIT_09 => X"000040090802009420409004104444084001022400214A2080014400026401A2",
INIT_0A => X"04000071200000A003CA294140200800C80C8C8100004590111C040040120800",
INIT_0B => X"12210002404848502847040164880021150400080222000200C8034200000000",
INIT_0C => X"4610088010080421021040841021000841021000841021000841010800420820",
INIT_0D => X"42D0A16C529A321068500484000500D10042080040284000084900001A002196",
INIT_0E => X"00000002804000004228010410082002C000C0002400046419120410034285A1",
INIT_0F => X"A00000000500800800000800000000000002290008001080000000A010100042",
INIT_10 => X"00000000000004C2001000000240000000000000680800280000000140202000",
INIT_11 => X"0000C0000000000000000442020001000001000000000000010C800080000804",
INIT_12 => X"08000000000801A7802010000000152780102000000015000600000800000000",
INIT_13 => X"000000000101900011E0240000000009500011E0280000000009500004DD0000",
INIT_14 => X"000137400020000000000201C000136C00101000000000002340002947000240",
INIT_15 => X"0080881901210000000600C280028000419480D4000010040000000000002304",
INIT_16 => X"68DA368DA1685A1685A1685A1685A16C5A121A13A141950051309284A82C0010",
INIT_17 => X"85A1685A1685A1685A368DA368DA368DA368DA368DA368DA368DA368DA368DA3",
INIT_18 => X"5A1685A168DA368DA368DA368DA368DA368DA368DA3685A1685A1685A1685A16",
INIT_19 => X"0157344CCCF48DE68A895C38E2540A8010100000000000000000685A1685A168",
INIT_1A => X"14514514514514514514514514514514514D34D34D34D34D28E1004039248209",
INIT_1B => X"D268341A4D268341A0D069349A0D069349A0D068341A0D068341A0D068345145",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000014D490D069349A0D068341A4",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"EAABA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"03DE00FFAEBFFFF0800155FFAAFBE8B45002A974AAAA803DFFFAA843DF45FFFF",
INIT_29 => X"7BFDE00A2FBD7400F7FBFDFFFA2AEBDE00AAFBEAABA080000000087BEAA10F78",
INIT_2A => X"055401FFF7AEAAA10F780155EFAAAEA8ABAAAFBFDE0055556AA005D041555508",
INIT_2B => X"557FC0010F780154105D7FC2145005155555557BE8BEF007FFDEAAAAD1555EF0",
INIT_2C => X"AF7D5555FFF780154AA5D2AA8A10F7AA974AA082E80010A2AAAAA10552AA8AAA",
INIT_2D => X"BAF7D17FEBAA2AEBDF45002EAAABA087BFDF45F7AA974AAAAAA97555F784174B",
INIT_2E => X"000AAFFE8A00552EBFE00F7D17FF45F7FFFFF55AA80155FF080400145FFFBEAA",
INIT_2F => X"8FC7BE8A3DF7DF7F5E8A92000000000000000000000000000000000000000000",
INIT_30 => X"000280071E8A00EB8E3FE10F7AEBAFFF080A175D7BEF1E8B6D002090482B68E3",
INIT_31 => X"56AA10410E175550871FFE00A2FBD0400FFF5FDFC7B6A0BDE38B6F5E8A92080E",
INIT_32 => X"7BFAE82A2DB555C71C5B451D7FFAAA8A38FF8E175C7A2AAAAA82A2F1FAE105D5",
INIT_33 => X"2AEADA38492EA8AAA5571C2000FF8A17400557FC015514555757D5D71E8BEF14",
INIT_34 => X"B6A49256DEB84104BAFFD1525FFFF84174BA5D20AAA00E3AA904BA142A87010A",
INIT_35 => X"7000400155FFFBEDA82FFD57DEBAAAA0BFF7D0024ADA921C7BFFF55FFA095482",
INIT_36 => X"00000000000000000000A2FBE8A38492ABDE10EBDF7AF6DE3FFF8F7DB68A105D",
INIT_37 => X"BEF080402000F7AAA8B55FFAABDFEFF7D16AA000000000000000000000000000",
INIT_38 => X"FEAAFFD16AA00082E820BA08556AA00AAAABFE00F7AEAABEF082E95545F7D568",
INIT_39 => X"A8A10AAD568A00555168A10002E9754D00517DE00A2FFC2000F7D17FF55FF803",
INIT_3A => X"1575EF555568BEF5D7FE8A10AAFFD55555D7FD5555FFAAA8AAAFFAA97555A2AE",
INIT_3B => X"AE800AA552A97400A2AEBDEAA082EAAABA5D5140010F7AE974105D7BC21555D5",
INIT_3C => X"57BFDF55F78017400F780001FFAA84000AAFFD1401E7FF80174AA5D0028A00AA",
INIT_3D => X"AAFBEABFFF7AA80145080002145F7FBFFE00FFD17FEAAA2803DFEF08043FE005",
INIT_3E => X"0000000000000000000000000000000000000A2FFE8ABA082ABFE00AAFBEABFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_2,               -- Port A enable input
WEA      => wbe_a_lo_1024_2(1),               -- Port A write enable input
DIA(0)   => data_write_a(9),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_2(9),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_2,               -- Port B enable input
WEB      => wbe_b_lo_1024_2(1),               -- Port B write enable input
DIB(0)   => data_write_b(9),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_2(9),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_10_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00018248A2840112C00002C18000202300500030B3132000400992006",
INIT_01 => X"254008000000004C002000000010026840000000080000080200010008110204",
INIT_02 => X"0020042000010000004455800008000004100000000000900200000002400004",
INIT_03 => X"020001021089000021081000C400090011000000610001540104C00000F14400",
INIT_04 => X"0811800101A00002000050088554004200C840000000200080C8100000000001",
INIT_05 => X"030080001000100800009400200000000840E020201000000024024001200020",
INIT_06 => X"81B00008080012120004CC080492500280208004148000100000020020042493",
INIT_07 => X"0000000800044080010000048404081085020002502000006000040800062480",
INIT_08 => X"100202400084410808000A00021004044048000004000000000021F020408264",
INIT_09 => X"010040090002008420401004144440004040022484214A2080110108C2C00320",
INIT_0A => X"04004166A48A0001080000000000080080181881000045901118044040020800",
INIT_0B => X"1201000200484910000F0105602622291404020902005002018002400A022000",
INIT_0C => X"0440001011808020120004801120044800120004801120044800110002400884",
INIT_0D => X"008000440210100041308480800F82F00040180260A808008848000018002104",
INIT_0E => X"000000028040000002280104100820020000400020000440100204100A000100",
INIT_0F => X"040000000500800800000000000000000002280008000400000000A010100010",
INIT_10 => X"00000000000004C2001000010000000000000000680800010000000140202000",
INIT_11 => X"200000000000000000000442000001000000000000000000010C000080001000",
INIT_12 => X"00000000000801C0008000000000154000800000000015000410000800000000",
INIT_13 => X"0000000001019800180000080000000958001800000400000009580002800000",
INIT_14 => X"0000A0000000000000000201E0000A0000400000000000002360002080000800",
INIT_15 => X"0080881000000000000600C28102800060000000000800000000000000002306",
INIT_16 => X"401004010040100401004010040100441020D0030008840051309A90BA884010",
INIT_17 => X"0902409024090240900401004010040100401004010040100401004010040100",
INIT_18 => X"1004010040902409024090240902409024090240902409024090240902409024",
INIT_19 => X"F546890A940FE0D3971243555205428290100000000000000000401004010040",
INIT_1A => X"8A28A28A28A28A28A28A28A28A28A28A28A28A28A28A28A29554199854514514",
INIT_1B => X"2B95CAE532994CA6532995CAE572B94CA6532994CA6532994CA6532994CA28A2",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000002718E72B94CA6532994CA657",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"FDE1000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"03DFFFAA843DF45FFFFEAABA007FC2155F7D155545AA80001EFAAFBEAB45557F",
INIT_29 => X"042AB55FFD168B55AA8000010FFFBE8BFFF78402155AAFBE8B45002A974AAAA8",
INIT_2A => X"AD16AABA002ABDE10080000000087BEAA10F7803DE00FFAEBFFFF0800155FF00",
INIT_2B => X"A2FBD7400F7FBFDFFFA2AEBDE00AAFBEAABAA2FFD741055003DFEFF7AA801FFA",
INIT_2C => X"05D0415555007FD74105555555EFF7FBC0145F78028A00A2D142155087BFDE00",
INIT_2D => X"55AAD168ABA002A975FFF7AEBDEBAF780155EFAAAEA8ABAAAFBFDE0055556AA0",
INIT_2E => X"000557BE8BEF007FFDEAAAAD1555EF0055401FFF7AEAAA105D042ABFF5D556AB",
INIT_2F => X"71D7AAFBEFB455D71F8E00000000000000000000000000000000000000000000",
INIT_30 => X"E8B6D002090482B68E38FC7BE8A3DF7DF7F5E8A92007BC217DEBDB55555AA8E0",
INIT_31 => X"EBAFFF080A175D700042AB7DEBDB6DB55BE8E05000EBFFE8BC7E38E07145BEF1",
INIT_32 => X"0A3DFD7F7A4821D7A2D16FA82142EB8E00080E000280071E8A00EB8E3FE10F7A",
INIT_33 => X"ED1421450871FFE00A2FBD0400FFF5FDFC7B6A0BDE38B6F5E8A92B6FBD541049",
INIT_34 => X"A2F1FAE105D556AA10410E175550071D54104951555D7EBF5C5155E3842AA00B",
INIT_35 => X"8410E2ABD749516FB55BED16FA820820955EFE3AEBDEAAFF8E175C7A2AAAAA82",
INIT_36 => X"000000000000000000005D71E8BEF147BFAE82A2DB555C71C5B451D7FFAAA8A3",
INIT_37 => X"1EFA2FFD7545AAAE97555A2FBFDF455D556AA000000000000000000000000000",
INIT_38 => X"8B45AAAA95545F7D568BEF080402000F7AAA8B55FFAABDFEFF7D16AA00087FC0",
INIT_39 => X"6AA00AAAABFE00F7AEAABEF082E9554500042ABFFA2FFFFF45F7AE97400AAFFE",
INIT_3A => X"16AA00FFFBD5400082EBFF45F78400155A2D57FE00552EA8A00082E820BA0855",
INIT_3B => X"D557555A2802AA10FFD54214500517DE00A2FFC2000F7D17FF55FF803FEAAFFD",
INIT_3C => X"FAA97555A2AEA8A10AAD568A00555168A10002E9754D085155410085557555AA",
INIT_3D => X"5D7FD5555FFAAA8AAA002AAAB4508557DF55F7D17FE000804155FFAAAABDEAAF",
INIT_3E => X"0000000000000000000000000000000000000555568BEF5D7FE8A10AAFFD5555",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_2,               -- Port A enable input
WEA      => wbe_a_lo_1024_2(1),               -- Port A write enable input
DIA(0)   => data_write_a(10),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_2(10),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_2,               -- Port B enable input
WEB      => wbe_b_lo_1024_2(1),               -- Port B write enable input
DIB(0)   => data_write_b(10),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_2(10),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_11_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"A101C4B05A0034CA2840712C2D001419000002300500030B31B20084EC992002",
INIT_01 => X"90000986B83028491800E0000C26426040000000080000088200080802512224",
INIT_02 => X"1A2004205E010640024D00800008000004100000040EC090820018003241A00C",
INIT_03 => X"28639100000C5C00000045C08400C8001100000061806A001618C03001E54400",
INIT_04 => X"1A800001000009A0804059A190000040400040008058220008C8100000120D4E",
INIT_05 => X"02000E81080250010000002022000058080400000E1200000020004401000004",
INIT_06 => X"819435143F20101010001008040800B8100102041088011100022200000024B2",
INIT_07 => X"90640D280884453E01064002944180008402001295BA100022E4340800062D82",
INIT_08 => X"400000093204802200280A0012160585C1D808D004000000000323F40C102244",
INIT_09 => X"380040098010001100009204107C5950400000220080C200800900020C006827",
INIT_0A => X"80007100004016EA080801010000080D00200081000045B0511D289940103399",
INIT_0B => X"002000024040410A000D0104408810C115D9C008050042400100D04E88000002",
INIT_0C => X"00655010009264201200C7B421ED0C7B421ED0C7B431ED087B43176843DA1085",
INIT_0D => X"0401020080400A10012494881A4F80F209500BB2602881A488485C1318002000",
INIT_0E => X"6619A540124814800228010410082022C00040002020090020220C9600040802",
INIT_0F => X"ACCC334A802491600C587949B6D0141B4CC600D5761B1599865A500490B86A56",
INIT_10 => X"BAC845542056A61686EC81E3A6CB68AA2C622C9A251C352B330CB4A0092170D8",
INIT_11 => X"BCCAD0B5A81536080CC6B21A21B1FC09CB0F1076D4A200B2AD4068F4101639B5",
INIT_12 => X"4D2CC281E31AA0103AB8D5514066380804B268A2E060901204112566F10AC418",
INIT_13 => X"D551443C47281002540B2C9AAAA8662A1152B202AE3554403028115AA88201A1",
INIT_14 => X"548A20A0492A2724A0621620402A020141F172FB182A32AB6845AB6200251BC9",
INIT_15 => X"00C00A000200074044E6801832728080D00A380B753952C4877E0104DDE4D124",
INIT_16 => X"0080200802008020080200802008020480080022020081010124988800400010",
INIT_17 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_18 => X"0000000000802008020080200802008020080200802008020080200802008020",
INIT_19 => X"55062608804180C0B10A42104201400204000000000000000000000000000000",
INIT_1A => X"00000000000000000000000000000000000820820820820801C4149470000000",
INIT_1B => X"0000000000000000040200000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000007E0F0000000000000100800",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"000AA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0001EFAAFBEAB45557FFDE10082ABDF5508557DF45002ABDFFFF7803DE10AA80",
INIT_29 => X"AEBFF45FFAEBFEAA002A801FFF7FFE8A10A28000000007FC2155F7D155545AA8",
INIT_2A => X"2AABFE10082ABFFEFAAFBE8B45002A974AAAA803DFFFAA843DF45FFFFEAABAA2",
INIT_2B => X"FFD168B55AA8000010FFFBE8BFFF78402155AAD155555A28428BFF002ABDE00A",
INIT_2C => X"F0800155FF00557FF45557FC2010002A80010A2842AAAA007BFFF4500042AB55",
INIT_2D => X"FF5D00154BAF7FBE8BEFFFD540000080000000087BEAA10F7803DE00FFAEBFFF",
INIT_2E => X"000A2FFD741055003DFEFF7AA801FFAAD16AABA002ABDE10A2D168A10A284021",
INIT_2F => X"DFC7F78E3FE28B684070AA000000000000000000000000000000000000000000",
INIT_30 => X"C217DEBDB55555AA8E071D7AAFBEFB455D71F8E00002EBDF6D005B78F7D142AB",
INIT_31 => X"A3DF7DF7F5E8A92BEAEBFF7DEBA0BDEAA1C2A801C7E3FFEFA10B68407038007B",
INIT_32 => X"8A28BFF082ABAE10B6AAB8E280820B8FEFBEF1E8B6D002090482B68E38FC7BE8",
INIT_33 => X"07FF8F7D00042AB7DEBDB6DB55BE8E05000EBFFE8BC7E38E07145B6D15756DA2",
INIT_34 => X"EB8E3FE10F7AEBAFFF080A175D708517DF7D497BC5028142A87000A28A2AA920",
INIT_35 => X"0B6DB6AA28A280001FF5D0A10482FFFFEFBC7E3DF42028080E000280071E8A00",
INIT_36 => X"00000000000000000000B6FBD5410490A3DFD7F7A4821D7A2D16FA82142EB8E0",
INIT_37 => X"FEF007BE8BFF5D2ABDF55F7AABDEAAF784154BA0000000000000000000000000",
INIT_38 => X"DE00FF84154BA087FC01EFA2FFD7545AAAE97555A2FBFDF455D556AA00082EBF",
INIT_39 => X"02000F7AAA8B55FFAABDFEFF7D16AA00FFAEBFFEFAA803DEBA5D2E82155A2FBF",
INIT_3A => X"A95545F7D5555FFAAAAA8BFF002AAAA00FFAAA8AAA080028BFFF7D568BEF0804",
INIT_3B => X"2E95400A2AEA8A00007FEABFF00042ABFFA2FFFFF45F7AE97400AAFFE8B45AAA",
INIT_3C => X"82E820BA08556AA00AAAABFE00F7AEAABEF082E9554508557DFFF007BD54BA5D",
INIT_3D => X"A2D57FE00552EA8A00FFFFE8AAAAA80001FF5D2E82000F7FFFFF45AAFFC20BA0",
INIT_3E => X"0000000000000000000000000000000000000FFFBD5400082EBFF45F78400155",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_2,               -- Port A enable input
WEA      => wbe_a_lo_1024_2(1),               -- Port A write enable input
DIA(0)   => data_write_a(11),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_2(11),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_2,               -- Port B enable input
WEB      => wbe_b_lo_1024_2(1),               -- Port B write enable input
DIB(0)   => data_write_b(11),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_2(11),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_12_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50080B01BC002006940202C0DE041196A83183000000023322287E0FC000006",
INIT_01 => X"75400D849830C84C5823E0000C17424840000000080000088200002802153231",
INIT_02 => X"18A026B43ED180040147558040090000061800000C06ED9802768F4472C52005",
INIT_03 => X"2A67E34A528D0524A52850528400C8001100000171C02B550618C91A10E55440",
INIT_04 => X"1BC0000100056C8280825DE98154004300C840800850240080CA921084520A07",
INIT_05 => X"02000F832000500C0000941024000852084060202E100001002000448100000C",
INIT_06 => X"819A1D1C3FE01A1A40045408049A50BA4020C6041090001200006200000000F2",
INIT_07 => X"C26A0719CC96CC6ED18A64019695A854870300FA3968B20068FC06080106249F",
INIT_08 => X"D002024B3E040800008C0A002610240D494A06F3460409000000E3F0AD5282E5",
INIT_09 => X"27A06009200040000400120412445D78400001000410420080218029CC807A27",
INIT_0A => X"18000006848A026F000000000000080000F010C100204593F11A6CDF48003BF8",
INIT_0B => X"000000820040402B28050400400432C9349DF21A31A00ACC0000F04F80020001",
INIT_0C => X"00357804611AE45D05D0833430CD0833420CD0C33420CD0833430668619A1000",
INIT_0D => X"0000000000000A74812DF00E87E80A079F9F90FA0280E87E800C7FF3B8002000",
INIT_0E => X"3B6B0E404D26160682082002000401EA0000C40000800A006002818808000000",
INIT_0F => X"A476D61C809A4DA84272592D6246FC1B17B541F97E1B348EDA93900B2B286C56",
INIT_10 => X"30C669E622DBC325CFD881A962454CFBE5403AB99594362B1DB52720165650D9",
INIT_11 => X"F8D2D39A3745261E4A95A110A3F855000E4B1D32BAB504BB7490FCFF912A3834",
INIT_12 => X"B90E9B018C7530200AB8F8BF41F9A22006B37DC8E1F9A21A70116D4C5080651C",
INIT_13 => X"118780319CCA08AB1001ACDF34B8F1C688AB1002AE3F7B807B6289F368828C4C",
INIT_14 => X"2AF020233376A5ECC016B1A827CDA21160F051DE610A34C50427E6E220323E4A",
INIT_15 => X"0077020000000439FDC05C5806781FAB46095A0B5199B0AC55521524F1864022",
INIT_16 => X"000000000000000000000000000000000026C000002884000130921092804010",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"8020080200000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0051B946088881360A95090CB054420290100000000000000000008020080200",
INIT_1A => X"041041041041041041041041041041041049249249249249200100002D451451",
INIT_1B => X"92C964B2592C964B2592C964B2592C964B2592C86432190C86432190C8641041",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000003800F592C964B2592C964B25",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"7DE1000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"ABDFFFF7803DE10AA80000AAAA843FE0008557DFFF0800020105D557FEAA0055",
INIT_29 => X"D5420000051555FFA2AA8200000557DFFFF7AA80000082ABDF5508557DF45002",
INIT_2A => X"82AA8AAAAAFFC00BA007FC2155F7D155545AA80001EFAAFBEAB45557FFDE10AA",
INIT_2B => X"FFAEBFEAA002A801FFF7FFE8A10A28000000A2D155410F7FFFFEBA08003FE000",
INIT_2C => X"5FFFFEAABA000028A105D2ABFE10A2AABFE1055516ABEF5D517DEAAA2AEBFF45",
INIT_2D => X"55002A820AA08557DFFFF7AA82155AAFBE8B45002A974AAAA803DFFFAA843DF4",
INIT_2E => X"000AAD155555A28428BFF002ABDE00A2AABFE10082ABFFEF0855420000004175",
INIT_2F => X"5010495B7AE921C517DE10000000000000000000000000000000000000000000",
INIT_30 => X"BDF6D005B78F7D142ABDFC7F78E3FE28B684070AABE803AE38145B78FD700000",
INIT_31 => X"BEFB455D71F8E00BED547038145B505FFB6A487000005F7AFD7F7A482038002E",
INIT_32 => X"F1FDE821C003FE001C2EAAAAAB6F5C2082007BC217DEBDB55555AA8E071D7AAF",
INIT_33 => X"D517DEAABEAEBFF7DEBA0BDEAA1C2A801C7E3FFEFA10B68407038B6D550428FF",
INIT_34 => X"B68E38FC7BE8A3DF7DF7F5E8A9200002FA285D20BDE28A2A4B8E10555B68BEF5",
INIT_35 => X"F085F47038140010555142082082005F7DFD7F7A482155BEF1E8B6D002090482",
INIT_36 => X"00000000000000000000B6D15756DA28A28BFF082ABAE10B6AAB8E280820B8FE",
INIT_37 => X"ABA5D7FEAB45080015410007FEAA0055517DE000000000000000000000000000",
INIT_38 => X"AB45F780020BA082EBFFEF007BE8BFF5D2ABDF55F7AABDEAAF784154BAF7802A",
INIT_39 => X"D7545AAAE97555A2FBFDF455D556AA00F7D1554BA5D7BC01FFFF8015410007FE",
INIT_3A => X"4154BAF7D1400BAFFD57FE005D043FE10552EAAAAAFFD140000087FC01EFA2FF",
INIT_3B => X"8428A105D7FEABEF55557DEBAFFAEBFFEFAA803DEBA5D2E82155A2FBFDE00FF8",
INIT_3C => X"7D568BEF080402000F7AAA8B55FFAABDFEFF7D16AA0008003FEBA55003DEBAA2",
INIT_3D => X"FFAAA8AAA080028BFF087BD54AA550402145550000010087FFFF45F78402145F",
INIT_3E => X"0000000000000000000000000000000000000F7D5555FFAAAAA8BFF002AAAA00",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_2,               -- Port A enable input
WEA      => wbe_a_lo_1024_2(1),               -- Port A write enable input
DIA(0)   => data_write_a(12),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_2(12),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_2,               -- Port B enable input
WEB      => wbe_b_lo_1024_2(1),               -- Port B write enable input
DIB(0)   => data_write_b(12),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_2(12),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_13_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10154A0441836CA2840512822007C18000E02700500030B31B300040081A042",
INIT_01 => X"00000804A000C04800020000000002404001000008220008A200100802110204",
INIT_02 => X"02200430000104000A4700804008000004100000000420918204D3033240400D",
INIT_03 => X"AA4003400008592400000590C40009141100000C6180C0000000C00001E14000",
INIT_04 => X"0800000102400120088054019000004160004190BAA0270000C8100000600206",
INIT_05 => X"21000012040610050040000227003AA0082400E94C1200000824424005220020",
INIT_06 => X"81963B180C001010580000080400000058000004109C00138000020024142581",
INIT_07 => X"002C8008000441600106400A9600010494020002B8AAA000EF003408000E2580",
INIT_08 => X"000000E48194408000A00A001210040441C80320040210000002ABF004102244",
INIT_09 => X"2A004009640040100400940412D4C4004000022000104200802D983000480120",
INIT_0A => X"8000202020401480000000000000080C90090881000145B0111A14004015080D",
INIT_0B => X"00000002004040AA08050400404040C11444000805200A402090024000008002",
INIT_0C => X"8410000A00280020020040800020040800020000801020000800010020400000",
INIT_0D => X"84A14250A055100050100490000500D00040080040290000084E4000B800610C",
INIT_0E => X"DCD13042BEDA36820228000000000000C000400081A08BC812A2092B02850942",
INIT_0F => X"89B9A260857DB400431969CA985D480949D32804A40AB137341C10B7D6A02EC0",
INIT_10 => X"E6ACA678001CE7D0296C213A460CA4271CA2168AEC1017606E6838216FAD4055",
INIT_11 => X"84AD4961C281B20213073C5FC0058008632D30D522CE80239DCC01AB013A4D20",
INIT_12 => X"2E6B13804A4B01D83461299900F6BD583A519104A0EEBD1A141010B2A4C8E116",
INIT_13 => X"89E5E40913419151EE0E94641828F72B5151EE0D184B321037AF5158BB02D085",
INIT_14 => X"562EC0B42162D68EE0073AE1C562EC13D521921A4170300B2B458B56B01C2280",
INIT_15 => X"00888A120240034000E6DC8285028014B82372011FC1E4F5E0A00929684EAF84",
INIT_16 => X"50942509425094250942509425094254940A1421420082020120908800480030",
INIT_17 => X"0942509425094250942509425094250942509425094250942509425094250942",
INIT_18 => X"9425094250942509425094250942509425094250942509425094250942509425",
INIT_19 => X"F7EFBBEEFF3F7DF7FF3E9F7DF7E2450228000000000000000000509425094250",
INIT_1A => X"BAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBF7DFDFDDD555555",
INIT_1B => X"EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAEBAE",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000000000F7EBF5FAFD7EBF5FAFD7",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"2ABEF00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0020105D557FEAA00557DE10AAD5554BA087FFFF55557BD54AAF7FBC01FFA280",
INIT_29 => X"7BD75EF087FFFFEF557BEAB45552E80155AA802AB45AA843FE0008557DFFF080",
INIT_2A => X"FAE820AA5D5557555082ABDF5508557DF45002ABDFFFF7803DE10AA80000AA08",
INIT_2B => X"0051555FFA2AA8200000557DFFFF7AA80000AAD1420AA087BD7555FFD168AAAF",
INIT_2C => X"5557FFDE10AAAEA8BFFA2FBD7545FFD157555085140010F7AEAABFFAAD542000",
INIT_2D => X"BA557BE8A10A284154BAFFAAAAB45007FC2155F7D155545AA80001EFAAFBEAB4",
INIT_2E => X"000A2D155410F7FFFFEBA08003FE00082AA8AAAAAFFC00BA00002AAAAF7D5574",
INIT_2F => X"0492E3F1C71C7BE8A2ABD7000000000000000000000000000000000000000000",
INIT_30 => X"3AE38145B78FD7000005010495B7AE921C517DE10A2DB50482147FFAF554971D",
INIT_31 => X"E3FE28B684070AA1C71D25D7007FFAFD7497BE8B5555208217DBE8A2AB45BE80",
INIT_32 => X"7FD257DFFD568A82FFA4870BA555F5056D002EBDF6D005B78F7D142ABDFC7F78",
INIT_33 => X"FAAAFBFFBED547038145B505FFB6A487000005F7AFD7F7A482038AADF4709214",
INIT_34 => X"AA8E071D7AAFBEFB455D71F8E00A2A0ADBC7A2FFD257DE3DF52555085142000F",
INIT_35 => X"21C002AA92FFDF574824171EAA10B680124BAFFAAAFB45007BC217DEBDB55555",
INIT_36 => X"00000000000000000000B6D550428FFF1FDE821C003FE001C2EAAAAAB6F5C208",
INIT_37 => X"0105D7BE8B55085142010AAD157545F7AEA8B550000000000000000000000000",
INIT_38 => X"01EFF7AAA8B55F7802AABA5D7FEAB45080015410007FEAA0055517DE00A2FFC0",
INIT_39 => X"E8BFF5D2ABDF55F7AABDEAAF784154BA5D5140145007BE8B55087BEAB555D040",
INIT_3A => X"0020BAA2FFD54105D7FC21EFFFD16AA10FF80174AA557FC21EF082EBFFEF007B",
INIT_3B => X"FBC0155085540000FFAEBFFEFF7D1554BA5D7BC01FFFF8015410007FEAB45F78",
INIT_3C => X"87FC01EFA2FFD7545AAAE97555A2FBFDF455D556AA00A2803FF45AAFFC21EFAA",
INIT_3D => X"552EAAAAAFFD1400005D042AA00F7FBD5410085568A10FF80020AAFFAABFF550",
INIT_3E => X"0000000000000000000000000000000000000F7D1400BAFFD57FE005D043FE10",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_2,               -- Port A enable input
WEA      => wbe_a_lo_1024_2(1),               -- Port A write enable input
DIA(0)   => data_write_a(13),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_2(13),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_2,               -- Port B enable input
WEB      => wbe_b_lo_1024_2(1),               -- Port B write enable input
DIB(0)   => data_write_b(13),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_2(13),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_14_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10020A000180000284008280000281800000030000000033022000000580002",
INIT_01 => X"000008020000204D006800000030824840000000084000084200090008510200",
INIT_02 => X"0220043170010A600A4D008040080000041000000028009002000F333240800C",
INIT_03 => X"111813400008002400000000C400090011000000610200001104D83000F14000",
INIT_04 => X"0801800100A000000000540084000040000040000800200000C8100000000748",
INIT_05 => X"0100000000001000000000002000080008000000001000000024024001200020",
INIT_06 => X"819EB84028001010000000080400000000000004108000100000020020040081",
INIT_07 => X"92040608000440100102400A94810206844200021DA2A0002000340800062C80",
INIT_08 => X"000000000084400008800A001214040441481500040000000000A7F408002244",
INIT_09 => X"0A0040090002008420401004104444004000020400214A208001000002400120",
INIT_0A => X"0400002020000000000000000000080C8008088100004590111B480040120000",
INIT_0B => X"1000000200404800000504016000002114000008020000020080024000000000",
INIT_0C => X"0410000010000000000040001000000000000040000000000001000000000000",
INIT_0D => X"04810244825010004010000000000000000000000000000000080000B8002104",
INIT_0E => X"0002C38280001202020800000000001000004000000000401022000002040902",
INIT_0F => X"20000587050001404E8084341CBA3404800828805200008000E0E0A000080002",
INIT_10 => X"4D18178E012010C00224004091C3514072C000444A0400080001C1C140001000",
INIT_11 => X"51709A07424142084458476001003809D0104B01C5710044020C4006010500C5",
INIT_12 => X"C26EE3803180C18006519462A00005001460E4730000050A1011004001060049",
INIT_13 => X"01F9E00660318000000538318740000140000001B4600CE80001400000002B62",
INIT_14 => X"0000000AD89857B0E0684411800000003799EB764D000330C300000000E3554B",
INIT_15 => X"0000021002002C000024008284001A0902000422E3F5960080480A0216A07240",
INIT_16 => X"4090240902409024090240902409024090081021020080015134920800480010",
INIT_17 => X"0902409024090240902409024090240902409024090240902409024090240902",
INIT_18 => X"9024090240902409024090240902409024090240902409024090240902409024",
INIT_19 => X"F5579B4E5C8FF0F7BE9D5F7DF650400200000000000000000000409024090240",
INIT_1A => X"9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7BF7DDDDDFCF3CF3D",
INIT_1B => X"F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE79E7",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000003FFF03F9FCFE7F3F9FCFE7F3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"420BA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"BD54AAF7FBC01FFA2802ABEFA2FBE8B55A2AE80000F7D5555555D2AAAABAAAD1",
INIT_29 => X"AA801FFA28402000AAAE955455500155EF0804155EFAAD5554BA087FFFF55557",
INIT_2A => X"7AEA8B45080417400AA843FE0008557DFFF0800020105D557FEAA00557DE10A2",
INIT_2B => X"087FFFFEF557BEAB45552E80155AA802AB4500516AA00A2AE800BAFFFFC20BAF",
INIT_2C => X"0AA80000AA005568ABAA28402010A2843FEBAFFFBD7410A2D168BFF087BD75EF",
INIT_2D => X"005D7FFDF4555517DFEF00043FEAA082ABDF5508557DF45002ABDFFFF7803DE1",
INIT_2E => X"000AAD1420AA087BD7555FFD168AAAFFAE820AA5D5557555002E80155A280000",
INIT_2F => X"0555412AA8ABAAADB40092000000000000000000000000000000000000000000",
INIT_30 => X"50482147FFAF554971D0492E3F1C71C7BE8A2ABD7A2FFEDB55B6A080038E3DB5",
INIT_31 => X"B7AE921C517DE10A2AE851FFB68402038AAAA955554900105FF0800175D7A2DB",
INIT_32 => X"A0800BAE3F1C0092EBAAADB6D080A12410BE803AE38145B78FD7000005010495",
INIT_33 => X"2D568BC71C71D25D7007FFAFD7497BE8B5555208217DBE8A2AB451C556FA00A2",
INIT_34 => X"142ABDFC7F78E3FE28B684070AA00516DABAA28402038B6803DE82F7F5D5410A",
INIT_35 => X"D002A80155B680000105D7FF8F455D5F78FD7000E3FEAA002EBDF6D005B78F7D",
INIT_36 => X"00000000000000000000AADF47092147FD257DFFD568A82FFA4870BA555F5056",
INIT_37 => X"F55FF84000AAAAFBC0145002AA8AAAAAFFC20000000000000000000000000000",
INIT_38 => X"01EF080417555A2FFC00105D7BE8B55085142010AAD157545F7AEA8B55A2FBFF",
INIT_39 => X"EAB45080015410007FEAA0055517DE00A2AA955FFFF80020BAAAAA9754508000",
INIT_3A => X"AA8B555D557FE00A280020BAAAD140000A2AEBFFEF082A82010F7802AABA5D7F",
INIT_3B => X"803DE00FFD557400AAD56AB455D5140145007BE8B55087BEAB555D04001EFF7A",
INIT_3C => X"82EBFFEF007BE8BFF5D2ABDF55F7AABDEAAF784154BA08557FEAAA284000AAFF",
INIT_3D => X"FF80174AA557FC21EF082A80145F780020105D7BEAB45557BE8B45082EBFEBA0",
INIT_3E => X"0000000000000000000000000000000000000A2FFD54105D7FC21EFFFD16AA10",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_2,               -- Port A enable input
WEA      => wbe_a_lo_1024_2(1),               -- Port A write enable input
DIA(0)   => data_write_a(14),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_2(14),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_2,               -- Port B enable input
WEB      => wbe_b_lo_1024_2(1),               -- Port B write enable input
DIB(0)   => data_write_b(14),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_2(14),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_15_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000A000000000284000280000001800020030000000033022000000180002",
INIT_01 => X"8000080000000048000000000000026040000000080000080200000000110200",
INIT_02 => X"0020042004010E60004C0080000800000410000000020090020000300245E005",
INIT_03 => X"0000010000080400000000408400480111000000610008000000C00000E54400",
INIT_04 => X"980000010000000088C2550080000040000040000008A00028C8100000120000",
INIT_05 => X"020004012E025000000001322000000A28008000011000000220004D41000000",
INIT_06 => X"819588000800101000011008040000100001060418800510000A620000000092",
INIT_07 => X"0000000800044004010C20008440810284020002102220002000340800062480",
INIT_08 => X"0000000001140800002C0A001214050540C800400406180000002DF004000244",
INIT_09 => X"1E00400900000000000016041044400440000000000042008001000000000022",
INIT_0A => X"0000000000000220000000000000080C00000081000045901118000040000000",
INIT_0B => X"0000000200404000010500004000000114000009000000000000004200000000",
INIT_0C => X"0000000000000000000040001000040001000000000000000001000020000800",
INIT_0D => X"000000000000001001208000180800000000030200000180800C400030002000",
INIT_0E => X"0000000000002600020800000000001080004000000000000002000000000000",
INIT_0F => X"A400000000000000000008000000000000000000000014800000000000000052",
INIT_10 => X"0000000000000000000000010240000000000000000000290000000000000000",
INIT_11 => X"2001C05838120800000000000000000000010000000000000000000000001804",
INIT_12 => X"081004000000000000A010000000000000902000000000180010002020000000",
INIT_13 => X"6600000000000000000024080000000000000000280400000000000000000000",
INIT_14 => X"0000000000200801000000000000000000501001920000000000000000000A40",
INIT_15 => X"0000020000000000000000003000000000000000000A101C3614000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000080000120980000000010",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000400200000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"28BEF00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"5555555D2AAAABAAAD1420BAFF8000010082A954BA00003DFEF085155400F784",
INIT_29 => X"AE95555A2FBE8BEFA2843DE00AA8015400FF84001EFA2FBE8B55A2AE80000F7D",
INIT_2A => X"2FBEAB45F7D56AABAAAD5554BA087FFFF55557BD54AAF7FBC01FFA2802ABEFF7",
INIT_2B => X"A28402000AAAE955455500155EF0804155EFFFFBE8BFF0800174AA557BFDE10A",
INIT_2C => X"A00557DE10F7D1574AAA2D16AB55FFD568BEF087FE8A1055003FE00A2AA801FF",
INIT_2D => X"00AA802AA00AAAE800BA5D0015545AA843FE0008557DFFF0800020105D557FEA",
INIT_2E => X"00000516AA00A2AE800BAFFFFC20BAF7AEA8B45080417400FFFFC21450800154",
INIT_2F => X"8FD7005150438F78A2DBFF000000000000000000000000000000000000000000",
INIT_30 => X"EDB55B6A080038E3DB50555412AA8ABAAADB40092E38E070280024904AA1C043",
INIT_31 => X"1C71C7BE8A2ABD7E3AA9257DA2FFE8BC7BE8E38E10A28017400E38A051FFA2FF",
INIT_32 => X"00124AA557FFDE10A2FBEDB6DF7D16AABAA2DB50482147FFAF554971D0492E3F",
INIT_33 => X"10038E38A2AE851FFB68402038AAAA955554900105FF0800175D7E3FFEFBD700",
INIT_34 => X"000005010495B7AE921C517DE10FFDF50482A2DB6AB45FFD56DBD7087BEAA384",
INIT_35 => X"0FFF1C017D140410400BE8E28A10AAA085082550A1057DBE803AE38145B78FD7",
INIT_36 => X"000000000000000000001C556FA00A2A0800BAE3F1C0092EBAAADB6D080A1241",
INIT_37 => X"4AA0800020BA550028B550855400AAF7AEBDFEF0000000000000000000000000",
INIT_38 => X"7400AAAE975EFA2FBFFF55FF84000AAAAFBC0145002AA8AAAAAFFC2000AAAA97",
INIT_39 => X"E8B55085142010AAD157545F7AEA8B55AAAE821EFAAFBEAB55F7AAA8A00AA841",
INIT_3A => X"417555AAFFFDF450804020AA557BFFE10A2FFFFFEFF7D568ABAA2FFC00105D7B",
INIT_3B => X"D17DF45007FE8AAA08002AAAAA2AA955FFFF80020BAAAAA975450800001EF080",
INIT_3C => X"7802AABA5D7FEAB45080015410007FEAA0055517DE00FFFBC2000AAFBE8B55F7",
INIT_3D => X"A2AEBFFEF082A82010FFD5421EF5D0000010F7AAA8A10AA8017400552A801EFF",
INIT_3E => X"00000000000000000000000000000000000005D557FE00A280020BAAAD140000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_2,               -- Port A enable input
WEA      => wbe_a_lo_1024_2(1),               -- Port A write enable input
DIA(0)   => data_write_a(15),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_2(15),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_2,               -- Port B enable input
WEB      => wbe_b_lo_1024_2(1),               -- Port B write enable input
DIB(0)   => data_write_b(15),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_2(15),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_16_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"DA22C618B1000482B688B186588884862A400438255FC38381441205BA803003",
INIT_01 => X"7045A80028404C211203A952A90341080B173340412000E1005D628000820484",
INIT_02 => X"428406A4000850848330118D0AAC55001349B108818005460229044001C01784",
INIT_03 => X"092C4020000500020000500986812C405000001A48202050000A214AC0650115",
INIT_04 => X"4804A55440256F504025E003A054F46415A4E62B6FE3307943965A00001A1152",
INIT_05 => X"0000001C40A5B950ADB8EA097057ECE14C86D2B7F85AAD17F4B100000B88148C",
INIT_06 => X"415401DCDCF2C0A8030140BCB0820A200342A1C641C1E8782F508F2B00003584",
INIT_07 => X"002701881A3202080AE00480A2002840BE1480FA004342AA6F12000054004867",
INIT_08 => X"08C54828091002000002B32A8C19064E486A8001510000014140C1E2A14891E0",
INIT_09 => X"015452B103020814004088B64102680B6596594800400413CAC0208944800000",
INIT_0A => X"96AA000484094C000000000000012C9000A0000D0A80000BF8028E87C1B99270",
INIT_0B => X"014808A02004200E540480212000A448C0082024AE50064B44000000000002A2",
INIT_0C => X"0004000D5846256AAEA811150445411150445411150445411150422A088A8200",
INIT_0D => X"00000004010042A204A0C5817D00005034052E40000817D00440004004AD3240",
INIT_0E => X"632B2673FA4587978A2004102800809225545155121740000004900090000000",
INIT_0F => X"00C6564CE7F4EA4B940076D296D003030800462CBD320018CAAAACFE9164C800",
INIT_10 => X"28834ADB1440A114793A4A30A40839AA14910D08DCB2640031955559FD3AC990",
INIT_11 => X"594AB0B1A025371CA0E034E8443C097A800EB090D4AAC91208ED2FA0CE5E09B1",
INIT_12 => X"7B50446083001B94BB38C540EBE61284BB304880E3E4579EDC00992980D58033",
INIT_13 => X"5511121840E7A2CD952ECC12ABC3E6ACB3DFB12ECE315000F61FF1727A85FDBC",
INIT_14 => X"75DEB07F6F2E7084517F126F8395CB2BEFBAB8BA8AF698228CC5E2F08ECA5159",
INIT_15 => X"5580A840A8009F8B108C80A1021B080AFC0DF6422C6077F4A77F20D0C0E21084",
INIT_16 => X"0000000000000000000000000000000000044000102A0001148442A110810359",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"558D11544C690DA64C1C4F68A360400000000000000000000000000000000000",
INIT_1A => X"14D14D14D14D14D14D14D14D14D14D14D14514514514514529E5F87869E79E78",
INIT_1B => X"D1E8F47A3D1E8F47A7D3E9F4FA7D3E9F4FA7D3E9F47A7D1E9F47A7D1E9F4D14D",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000007D3E9F4FA7D3E8F47A3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"C00AA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"03DFEF085155400F78428BEF087FFFFEFF7D168B55AAD17FFFF552EBFE00007F",
INIT_29 => X"2E975EFF7D568BFFFF80175EF0004000BA552A821FFFF8000010082A954BA000",
INIT_2A => X"55540000082EAABFFA2FBE8B55A2AE80000F7D5555555D2AAAABAAAD1420BA5D",
INIT_2B => X"A2FBE8BEFA2843DE00AA8015400FF84001EF0000020AA5D00154005D043FF455",
INIT_2C => X"FA2802ABEF557BEABEF5D0415410087FD74BAAAAEBFFEF557FC00AAF7AE95555",
INIT_2D => X"FFFFAABFEAAFF84001FF002A821FFAAD5554BA087FFFF55557BD54AAF7FBC01F",
INIT_2E => X"000FFFBE8BFF0800174AA557BFDE10A2FBEAB45F7D56AABA082A97545F7D16AB",
INIT_2F => X"FFEF552AB8E38087FC2092000000000000000000000000000000000000000000",
INIT_30 => X"070280024904AA1C0438FD7005150438F78A2DBFF0871F8FC7E3D56AB6DBEDB7",
INIT_31 => X"AA8ABAAADB400924920925EFF7D16ABFFE38E175EF1400000BA412E871FFE38E",
INIT_32 => X"0A1240055003FF6D5551420101C2EAFBD7A2FFEDB55B6A080038E3DB50555412",
INIT_33 => X"57FC00BAE3AA9257DA2FFE8BC7BE8E38E10A28017400E38A051FF0804050BA41",
INIT_34 => X"4971D0492E3F1C71C7BE8A2ABD74975EDBC7550E12410087FD74AAB6AABFFC75",
INIT_35 => X"A08249756DF7D168BC7F7AABAEAAF780051C70824851D7A2DB50482147FFAF55",
INIT_36 => X"00000000000000000000E3FFEFBD70000124AA557FFDE10A2FBEDB6DF7D16AAB",
INIT_37 => X"B55A2D16ABEFFFFBFDFFF552AAAAAA007BC00000000000000000000000000000",
INIT_38 => X"20AA002A955EFAAAA974AA0800020BA550028B550855400AAF7AEBDFEF08516A",
INIT_39 => X"000AAAAFBC0145002AA8AAAAAFFC20000000021EFF7D568BFFA2AA955FF5D040",
INIT_3A => X"E975EF0800174BA002E820105D003DFEF5D51420005D2ABFF45A2FBFFF55FF84",
INIT_3B => X"7BD74AAF7AEBDF455D7BC20BAAAAE821EFAAFBEAB55F7AAA8A00AA8417400AAA",
INIT_3C => X"2FFC00105D7BE8B55085142010AAD157545F7AEA8B5500557DF45552A8200000",
INIT_3D => X"A2FFFFFEFF7D568ABA0804155FFF7D568B55FFAAAAABAFF8415545000015555A",
INIT_3E => X"0000000000000000000000000000000000000AAFFFDF450804020AA557BFFE10",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_2,               -- Port A enable input
WEA      => wbe_a_lo_1024_2(2),               -- Port A write enable input
DIA(0)   => data_write_a(16),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_2(16),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_2,               -- Port B enable input
WEB      => wbe_b_lo_1024_2(2),               -- Port B write enable input
DIB(0)   => data_write_b(16),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_2(16),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_17_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"5284CE4FB7BD2C8994A13392DBD02E14006B82AC7E800D44D3DD2FD5F9B961C0",
INIT_01 => X"2EACD01F7E03FC6793F2199B39FC233C11D93AE6F3BB92B32091DBC339B24542",
INIT_02 => X"E63CCCC00A82C08092A2AFAE667033DB50853379C10BFDC5C6F4044443C817C6",
INIT_03 => X"7FF183635AEF9E3635AEF9E18E237040404446965C0607EE6DB7854AC4DE060C",
INIT_04 => X"D78AC33FB604488B000892EF17BE6D84196482236FE100294152E294350FB697",
INIT_05 => X"081B5F9B409420D0CDB47A05403F6CE0C08A4AB7F840EDB6F48100DFC8081081",
INIT_06 => X"768465354781CBC30316367077B4BDB50646E8D87100A8201ED01C19C020F71A",
INIT_07 => X"4002A110C922480A82D0841147162C48EBB9537A0022DC67987042EE976ABEA7",
INIT_08 => X"DB931BFEF91C00002CC0E019C0C82A4E4820C15A2330E004401891181168C4D1",
INIT_09 => X"09F3A1BC11EFBC66DB65307071477FF1030C397C060B4254064302042F803A69",
INIT_0A => X"3F330802162F3B7EE3F3EC7C7DEF207000F00059D2ED56D7EED2ED3C9A867DC0",
INIT_0B => X"185C44B91BC1740B7605040BE0018CFC7429F326B9E822FFC00074D5A0AB033A",
INIT_0C => X"00367A28FC1B7F7FEFFCFBFF3EFFCFBFF3EFFCFBFF3EFFCFBFF3EFFE7DFF9E00",
INIT_0D => X"0000000008004BA78428C7AD7FC94B533F5B4FFBD2FAD7FCCA786D43FE67C218",
INIT_0E => X"BA494CEBFD4F2667ABB6F68B29760593F33FA0CF170F40006001B1A05C000000",
INIT_0F => X"7F749299D7FAEB237DFE5865B6D2BF23265CBACE542A6FEE92333AFF33E0A9BF",
INIT_10 => X"F6C24B6D18C3C9F8E2881F3F787D776B5DB94A09955054DFDD246675FE7AC153",
INIT_11 => X"BFB349E08FF9A27EDE9FA8AEFD9E7467BFCB195CFEB56A1A70D34D1706FFFA3E",
INIT_12 => X"6FE219CA80725B875EED723FF7FCB2875EDAAFEAF7FD929BFD55BBC71D79F639",
INIT_13 => X"546670D018E7A6E581D7B6AB75FDFCECA6E581D7BB5DDFC6FF0EB7D7E859FDB5",
INIT_14 => X"B978177F6D6AF5ECDB5FB76A5F5FA165B456E0FB308710C49FCFB741598B9C7E",
INIT_15 => X"CFDAAB00AC00A8BBFC8B501CF7A0FED9A540EA1952586CEB54D143ACFF9A3BA9",
INIT_16 => X"000000000000000000000000000000000026E100002F382DBD9ECFE117805F20",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"4372003009EDCC4052E917114F981800C0000000000000000000000000000000",
INIT_1A => X"BA69A69AEBA69AEBA69A69AEBA69AEBA69A69A69A69A69A68698686981D75D74",
INIT_1B => X"6A351A8D46A351A8D068341A0D068341A0D068341A0D46A341A0D46A341A69AE",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000000000046A351A8D46A351A8D4",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"7FEAA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"17FFFF552EBFE00007FC00AA087FFFFFFFFFFFFFEFF7FBEAB450804001EFAAD5",
INIT_29 => X"D168A000004020AA5D7BE8B450051401EF087FD74AA087FFFFEFF7D168B55AAD",
INIT_2A => X"D7FEAB55FF80175EFFF8000010082A954BA00003DFEF085155400F78428BEFAA",
INIT_2B => X"F7D568BFFFF80175EF0004000BA552A821FF5D00020BA552A82000552A821555",
INIT_2C => X"AAAD1420BAFFFFFDF45AAD17FFFFAAFBC01EF5D0015555557BFDEBA5D2E975EF",
INIT_2D => X"BA007FEABEF005555555A2D1554BAA2FBE8B55A2AE80000F7D5555555D2AAAAB",
INIT_2E => X"0000000020AA5D00154005D043FF45555540000082EAABFF00516AA10552E820",
INIT_2F => X"8B550000071EFB6DF7AE92000000000000000000000000000000000000000000",
INIT_30 => X"F8FC7E3D56AB6DBEDB7FFEF552AB8E38087FC2092147FFFFFFFFFBFDFC7EBF5E",
INIT_31 => X"150438F78A2DBFFBED16AA381C0A07082497FEFB6D1451471EF007BD04920871",
INIT_32 => X"2A850105D2A80155417BEFB6DEB8E175FFE38E070280024904AA1C0438FD7005",
INIT_33 => X"D7BFAEBA4920925EFF7D16ABFFE38E175EF1400000BA412E871FF550A0009249",
INIT_34 => X"E3DB50555412AA8ABAAADB40092FFF5FFF6DAADF7FFD7B6F1C71EF55001756D5",
INIT_35 => X"7145B6AA28492487082007FEDBD700515556DA2DF50492A2FFEDB55B6A080038",
INIT_36 => X"000000000000000000000804050BA410A1240055003FF6D5551420101C2EAFBD",
INIT_37 => X"FEFF7FBFFF55A2D16AB550000175EFFFFBEAA000000000000000000000000000",
INIT_38 => X"55EF087FC200008516AB55A2D16ABEFFFFBFDFFF552AAAAAA007BC0000557FFD",
INIT_39 => X"020BA550028B550855400AAF7AEBDFEFF7D568AAA5D2A97410007BFFFFF55515",
INIT_3A => X"A955EF5D2E80010002A954005D2A82155087FFFFEFAAAA975EFAAAA974AA0800",
INIT_3B => X"D1575FF5504175EF5D7FEAAAA0000021EFF7D568BFFA2AA955FF5D04020AA002",
INIT_3C => X"2FBFFF55FF84000AAAAFBC0145002AA8AAAAAFFC2000FFD57DFFFAAFFFDF55FF",
INIT_3D => X"5D51420005D2ABFF45557FE8AAA000415410007BFFF450051555EFA2FBC0000A",
INIT_3E => X"00000000000000000000000000000000000000800174BA002E820105D003DFEF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_2,               -- Port A enable input
WEA      => wbe_a_lo_1024_2(2),               -- Port A write enable input
DIA(0)   => data_write_a(17),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_2(17),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_2,               -- Port B enable input
WEB      => wbe_b_lo_1024_2(2),               -- Port B write enable input
DIB(0)   => data_write_b(17),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_2(17),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_18_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"69844019080000A21A611406840014122A641074155FC28A2024001001801003",
INIT_01 => X"7443D920034004180005E9E3C90360C0041C0181002001602025800008440084",
INIT_02 => X"E2DCCCE61D5C008103F2000781FC0FEDEAC2161B0B8FB0008620044443006010",
INIT_03 => X"884E300802006900802006995C896D605200000856E24A040000640052141103",
INIT_04 => X"480520FC026125AC0025C9122644E3E40EC8E2001001302281841A009038A86A",
INIT_05 => X"432000040089983070019400F01010004C8DB841405A80A100B586200FAC24AE",
INIT_06 => X"09044359DC7040000000002C109B0E0A00A1104641C0803804000707284600E1",
INIT_07 => X"400D10100400481D5EB08501620000007500CE801241021FE78E404860140060",
INIT_08 => X"00880C0106A0528020019307CC082A0A4A6A01ED725021400040D028000A9729",
INIT_09 => X"00117063038000282081402E4106400B6186128040600C10C1C0200950508110",
INIT_0A => X"C0C30C2E21580C874004008080003C32A10A19090C02010E1022944061688000",
INIT_0B => X"0180A8062026000DC425C0301311324AA2373088479105D044A1022000001835",
INIT_0C => X"0D89844703649000000200000000000000000000000000000000000000000010",
INIT_0D => X"0D8306C182701404C1973010802020404084001E00010802046092B5001FB365",
INIT_0E => X"528EB314068AB8B803DB00002900800400FC503F08180050942E4200020C1B06",
INIT_0F => X"40A51D66280D6032C5F96D3C51555D5D7D5AA87285820814A3CCC501C2A60820",
INIT_10 => X"8B35A3FEBF1FEDFD9C2B30E0468AAAD5D48F37E8FC1304102947998A03984C10",
INIT_11 => X"440FE1DD772D37A0A321BC6968F32658BF2D4F2A80BF8FE3F9FE3AC362080529",
INIT_12 => X"5487910D7E5A6D961A28456A1832E5161A100DD5182BC54020EA67A189C6ED36",
INIT_13 => X"AA444CAF91EDD1B725868403BE06323551B725868A100ABD119753B70964122B",
INIT_14 => X"EDC259048ACD868EE3803D65CEDC258A8F80D55E007C3F8EBB56F4C5362C978F",
INIT_15 => X"3F240014BE84370001B6922070440556B15F7FABBC0031BCF2257C41634B14D4",
INIT_16 => X"C1B06C1B06C1B06C1B06C1B06C1B06C1B0491069068000004060300A005A0118",
INIT_17 => X"1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06",
INIT_18 => X"B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C",
INIT_19 => X"B28BBECEB80EE173C2300F7DF16000000000000000000000000041B06C1B06C1",
INIT_1A => X"8A28A28AAAAAAA28A28A28AAAAAAA28A28A28A28A28A28A2910591505C104104",
INIT_1B => X"28944A25128944A25128944A25128944A25128944A2552A954AA5128944AAAA2",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000128944A25128944A251",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"9540000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"BEAB450804001EFAAD57FEAA087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974BA082E",
INIT_29 => X"7FFFFFFFFFBFDF45AAD568B55080028B55002E82000087FFFFFFFFFFFFFEFF7F",
INIT_2A => X"0043DE10AA843DE00087FFFFEFF7D168B55AAD17FFFF552EBFE00007FC00AA08",
INIT_2B => X"0004020AA5D7BE8B450051401EF087FD74AAAAFFFDF45A2D16AB55F7FFFFFFF0",
INIT_2C => X"0F78428BEFAA80000000804154BA55042ABEF5D7FD75FFAAD540145AAD168A00",
INIT_2D => X"00082E95555085168A10557FD7545FF8000010082A954BA00003DFEF08515540",
INIT_2E => X"0005D00020BA552A82000552A821555D7FEAB55FF80175EF5D00020105D2A974",
INIT_2F => X"DFFF5D2A954AA082A92428000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFBFDFC7EBF5E8B550000071EFB6DF7AE921C7FFFFFFFFFFFFFFFF7FBF",
INIT_31 => X"AB8E38087FC2092087FFDFC7E3F1FAF55A2DF6DB7D1C002AB7D002A82028147F",
INIT_32 => X"DF6DB7DE3F5FAFC708003DE28B68E38E280871F8FC7E3D56AB6DBEDB7FFEF552",
INIT_33 => X"ADF4516DBED16AA381C0A07082497FEFB6D1451471EF007BD0492B6F1F8F55AA",
INIT_34 => X"1C0438FD7005150438F78A2DBFFA28407038140410492550A2ABC7497BD25FFA",
INIT_35 => X"F5D0E05000492097428002E9557D1C516FA28417BD5545E38E070280024904AA",
INIT_36 => X"00000000000000000000550A00092492A850105D2A80155417BEFB6DEB8E175F",
INIT_37 => X"FFFFFFFFDFEFF7FBFFFEF552E974AA082A820AA0000000000000000000000000",
INIT_38 => X"ABEF002A800AA557FFDFEFF7FBFFF55A2D16AB550000175EFFFFBEAA00557FFF",
INIT_39 => X"6ABEFFFFBFDFFF552AAAAAA007BC0000087BFDF45AAD568B55AAFBFDFEF55042",
INIT_3A => X"FC2000FFD56AB45A2FFFDFFFAAD16AB4500043DEAAFFAEAAAAA08516AB55A2D1",
INIT_3B => X"2AA8B45087FC01EFA2FFD55EFF7D568AAA5D2A97410007BFFFFF5551555EF087",
INIT_3C => X"AAA974AA0800020BA550028B550855400AAF7AEBDFEFA280154BA55040000055",
INIT_3D => X"087FFFFEFAAAA975EF5D2E974000804154BA082A975EF5D517DEAA007BD5545A",
INIT_3E => X"00000000000000000000000000000000000005D2E80010002A954005D2A82155",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_2,               -- Port A enable input
WEA      => wbe_a_lo_1024_2(2),               -- Port A write enable input
DIA(0)   => data_write_a(18),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_2(18),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_2,               -- Port B enable input
WEB      => wbe_b_lo_1024_2(2),               -- Port B write enable input
DIB(0)   => data_write_b(18),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_2(18),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_19_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"042200000000000041088001001AA00000000000000000000000500802000003",
INIT_01 => X"040048000024000000000404000000000A22000800000800004A200000000001",
INIT_02 => X"200C8840085EB00480060000001C008002489E0F000405EA0004040404000000",
INIT_03 => X"24004000000000000000000900002C4050000000000069500208400002E14100",
INIT_04 => X"4800200C0000000044002000C80020E40000E200000130200188000000800100",
INIT_05 => X"000000000080181000000000701000004C8000000058800000B1000009880480",
INIT_06 => X"80500081081040000000002C100040400000004641C080380400070100000000",
INIT_07 => X"4020109801A4CE005C00048380142810010564C4100114012002402028044808",
INIT_08 => X"0070700000000000000083004C3902420062000020E0000100004082A140102B",
INIT_09 => X"001150200000000000000026400000016186100000000010C04002C000000000",
INIT_0A => X"007C00008082C0002000000000002C3000000004050001030102040000000000",
INIT_0B => X"0000000000000000000000000000010000800011000000000000000000000BC0",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"000000000000000000000000000000042000760000000000000000010004B200",
INIT_0E => X"0D74002280300F0002FB069040000060000C5003000800000000000000000000",
INIT_0F => X"C01AE8004500744C780687DBA828008080A5FC0D385598035D0008A00C015660",
INIT_10 => X"39D8140040201BF861F0E7D693E6170022408116DFE0AB3006BA0011401D02AC",
INIT_11 => X"5412E4997F5249FD005043B8680CC98F00D0F2DD0140100406FE053A98F6ECC7",
INIT_12 => X"7418663001858040E153888000010840E165D0000000285C246A181C03FE4662",
INIT_13 => X"8199830066F0020858385974000001260208583854E2200000660208D6B1423F",
INIT_14 => X"8235AC508FCE8811042040F008235AE04420C040CF00C031C80009B8F224978B",
INIT_15 => X"030004E00000C220010808C10D9A92A74CD7CF4A09051110AD5A3C9200B7F280",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000118",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"07208BBA3F0C7010C660C7441920000000000000000000000000000000000000",
INIT_1A => X"861869A61861861861869A61861861861861861861861861A8208C4C1534D34C",
INIT_1B => X"984C26130984C26130984C26130984C26130984D26930984C26130984C261861",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000984C26130984C26130",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"174BA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFDFEF5D2A974BA082E95400F7FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0004",
INIT_29 => X"FFFFFFFFFFFFFFFFF7FBFDFFF552E974BAA2FFFFE10087FFFFFFFFFFFFFFFFFF",
INIT_2A => X"004001EFAAAEA8ABA087FFFFFFFFFFFFFEFF7FBEAB450804001EFAAD57FEAAF7",
INIT_2B => X"FFFBFDF45AAD568B55080028B55002E82000F7FFFFFFFFFFFFDFEFA2D568B550",
INIT_2C => X"0007FC00AAF7FFFFFFFF7FBE8B55AAD16ABEF5D2ABFF55080402010087FFFFFF",
INIT_2D => X"55A2FFFDFEF5D2EBFE00AAFFFFEBA087FFFFEFF7D168B55AAD17FFFF552EBFE0",
INIT_2E => X"000AAFFFDF45A2D16AB55F7FFFFFFF00043DE10AA843DE00557FFDFEFA2D16AB",
INIT_2F => X"FFEF552A974AA0000104AA000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFF7FBFDFFF5D2A954AA082A92428E3FFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"0071EFB6DF7AE92EBFFFFFFFFFFFFDFEFF7F5FAFC7492A974AAB6F5F8E101C7F",
INIT_32 => X"F1F8FD7AAD16AB450000001FFBEA4A8AAA147FFFFFFFFFBFDFC7EBF5E8B55000",
INIT_33 => X"00000010087FFDFC7E3F1FAF55A2DF6DB7D1C002AB7D002A82028FFFFFFFEFF7",
INIT_34 => X"BEDB7FFEF552AB8E38087FC2092F7FBF8FC7E3F5EAB45B6DF6FBEF5D2AB8F7D0",
INIT_35 => X"84971F8FC7AAD56DB6DBEF5F8FD7412ABFE28B6F5F8E820871F8FC7E3D56AB6D",
INIT_36 => X"00000000000000000000B6F1F8F55AADF6DB7DE3F5FAFC708003DE28B68E38E2",
INIT_37 => X"FFFFFFFFFFFFFFFFFDFEF552E954AA0004000AA0000000000000000000000000",
INIT_38 => X"54AAF7D568A00557FFFFFFFFFFFDFEFF7FBFFFEF552E974AA082A820AAA2FFFF",
INIT_39 => X"FFF55A2D16AB550000175EFFFFBEAA00A2FFFFFFFF7FBFDFFFFFD568B55002A9",
INIT_3A => X"A800AAF7FBFDFEFF7D56AB45AAD56AB450004001EFFF842AAAA557FFDFEFF7FB",
INIT_3B => X"FFFFFFF552AA8BEF080402000087BFDF45AAD568B55AAFBFDFEF55042ABEF002",
INIT_3C => X"8516AB55A2D16ABEFFFFBFDFFF552AAAAAA007BC0000FFFBE8B55AAD168B55F7",
INIT_3D => X"00043DEAAFFAEAAAAA08556AB55A2D57FFFFF7D568B45002ABDEAAFFD16AA000",
INIT_3E => X"0000000000000000000000000000000000000FFD56AB45A2FFFDFFFAAD16AB45",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_2,               -- Port A enable input
WEA      => wbe_a_lo_1024_2(2),               -- Port A write enable input
DIA(0)   => data_write_a(19),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_2(19),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_2,               -- Port B enable input
WEB      => wbe_b_lo_1024_2(2),               -- Port B write enable input
DIB(0)   => data_write_b(19),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_2(19),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_20_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000003",
INIT_01 => X"F55FF80000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"E05022020800008400F655001FFCFF80018FA804400000000000004400000001",
INIT_03 => X"00000000000000000000000900002CC07000000000000000000000000000013F",
INIT_04 => X"68002FFE40900010000180000001FFEC0012EE0C001370F40780000000000000",
INIT_05 => X"0840000880FCBBF0100E204DF0F88311DD8005080679800000F3000029980580",
INIT_06 => X"001000030817C8E8840155FDF9001001050023F6C3C3D0F87FA19F7F011000E4",
INIT_07 => X"000000090492260800008000EE00000000000000002101FF2002C00000004018",
INIT_08 => X"2A040001071004000013FF7FCA302C0C0008214800002101554031F800000000",
INIT_09 => X"801F57F200000090000489FEC0000001EFBEF0040008023FDFC0000000004006",
INIT_0A => X"0000000008000000000000000000ADF000000200000008000008028300110230",
INIT_0B => X"0000000000000800080000000000000000000000000000000800800A40000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"000000040900005C848538000020000000800000080000020000800101FFB600",
INIT_0E => X"00800000003A010003000000000000600FFC53FF001800000002004080000000",
INIT_0F => X"0001000000007408040000004000000004E9000008020000200000000E800800",
INIT_10 => X"00200000000313100010002000008000000000129600040000400000001D0010",
INIT_11 => X"81C012060000000000218F7840000100800004000000000066C0000080080000",
INIT_12 => X"800000000017C000100000000001A800080000000001A8040000002840008185",
INIT_13 => X"0000000006F00000100200000000012600001004000000000066000000801040",
INIT_14 => X"0000200410100000000005F00000020080090A0000000085C800002000586000",
INIT_15 => X"FF00400000000000020020020001000040283024E4F2860400008000030ED080",
INIT_16 => X"00000000000000000000000000000004010201001003020200000000000127DB",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"A0700030038200010089120104D2040020000000000000000000000000000000",
INIT_1A => X"2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2C30C30C30C30C306982121A1E79E79",
INIT_1B => X"32190C86432190C86432190C86432190C86432190C86432190C86432190CB2CB",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000432190C86432190C864",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0201000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF552A974AA0004174BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA0804",
INIT_29 => X"7FFFFFFFFFFFFFFFFFFFFFFEF552E954AA000400000F7FFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E954BA007FC00BA087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974BA082E9540000",
INIT_2B => X"FFFFFFFFFF7FBFDFFF552E974BAA2FFFFE10FFFFFFFFFFFFFFFFFFFFFBFDFFF5",
INIT_2C => X"FAAD57FEAA007FFFFFFFFFFFFFEFF7FBFFF550800020BAAAD56AAAAF7FFFFFFF",
INIT_2D => X"EFF7D56AB450000021EFA2D57DE10087FFFFFFFFFFFFFEFF7FBEAB450804001E",
INIT_2E => X"000F7FFFFFFFFFFFFDFEFA2D568B550004001EFAAAEA8ABA5D7FFFFFFFFFFFDF",
INIT_2F => X"FFFF5D2E954AA080005000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFEF552A974AA0000104AAFFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"A954AA082A92428087FFFFFFFFFFFFFFFFFFBFDFEF5D2E974AA000A07000E3FF",
INIT_32 => X"FFFFFEFF7FBFFFFF552E974AA0071C50BA1C7FFFFFFFFFFFFFFFF7FBFDFFF5D2",
INIT_33 => X"EDF6FABAEBFFFFFFFFFFFFDFEFF7F5FAFC7492A974AAB6F5F8E10E3FFFFFFFFF",
INIT_34 => X"EBF5E8B550000071EFB6DF7AE921C7FFFFFFFFFBFDFEFE3F5F8F450004050AAB",
INIT_35 => X"A497FFFFFFF7FBF8FC7EBD168B450804021FFB6D57DE28147FFFFFFFFFBFDFC7",
INIT_36 => X"00000000000000000000FFFFFFFEFF7F1F8FD7AAD16AB450000001FFBEA4A8AA",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2A954AA0800174100000000000000000000000000",
INIT_38 => X"74AA002E95410A2FFFFFFFFFFFFFFFFFFFFFDFEF552E954AA0004000AAFFFFFF",
INIT_39 => X"FDFEFF7FBFFFEF552E974AA082A820AA087FFFFFFFFFFFFFEFF7FBFDFFF5D2A9",
INIT_3A => X"568A00AAFFFFFFFFFFBFDFEFFFFFFDFEF5D2E954AA0051554BA557FFFFFFFFFF",
INIT_3B => X"D16AB450804174AAFFFFFFEBAA2FFFFFFFF7FBFDFFFFFD568B55002A954AAF7D",
INIT_3C => X"57FFDFEFF7FBFFF55A2D16AB550000175EFFFFBEAA005D7FFFFEFF7FBFDFFFAA",
INIT_3D => X"0004001EFFF842AAAA087BFDFEFF7FFEAB45A2D568B550804001EFF7D57DEBA5",
INIT_3E => X"0000000000000000000000000000000000000F7FBFDFEFF7D56AB45AAD56AB45",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_2,               -- Port A enable input
WEA      => wbe_a_lo_1024_2(2),               -- Port A write enable input
DIA(0)   => data_write_a(20),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_2(20),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_2,               -- Port B enable input
WEB      => wbe_b_lo_1024_2(2),               -- Port B write enable input
DIB(0)   => data_write_b(20),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_2(20),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_21_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"4A302428B824900A128C090A5C1800261500213C005FE812D10420054085A202",
INIT_01 => X"001FFE3440B609703B0427F801A40B8115BC4F655300340288A40D30040E4DD8",
INIT_02 => X"E00424256888D8819801000F9FFFFFFFF149FF1FCA448046C60A0D2437C517F9",
INIT_03 => X"20030640003250640003250F06002CC1740002019824E001CD357832440001FF",
INIT_04 => X"EA2C3FFD400006E04401A8837001FFFC004AEF00080B70E08FB5789421007C5C",
INIT_05 => X"00011A0C40F9FFF80920954FF0F00809DF84A0202879800000F3000029980780",
INIT_06 => X"0805984B7A1FC0A0000101FFF0480080002281F7C3C381F87C03DFFF00009004",
INIT_07 => X"B424068086A205481A60A19000908204A855B000A08A61FF20C3D004D331D340",
INIT_08 => X"1BFA0001600802000023F7FFC08D234B40C2028253000040114200000D0226C0",
INIT_09 => X"EF1F5FF054096C6ADBA169FFC202B1C1FFBEF0440021083DFFCE22DC2880E24D",
INIT_0A => X"45FF0C004041D84862A28C54518DBFF00020004C0A6044901112A0908AA0A300",
INIT_0B => X"018C241102068006C620C03882019480E63180855A492712CC01C49C20201BFE",
INIT_0C => X"08A9464116544302C02D92236488D92236488D92236488D922366446C911B210",
INIT_0D => X"08800444021048034004001890000806002804A0822189000900D80621FFBE00",
INIT_0E => X"060580261013813A2CC396506102C4053FFD5BFF00A04A00200602CA52001100",
INIT_0F => X"080C0B004C202621A85C09411500135844C196D3606941018150098404C1A304",
INIT_10 => X"B02901013416181C96C2C9C600890A2028172192C460D1820302A0130809834A",
INIT_11 => X"9C5E803408250180AC268D185DB3F4350B811068C00049A0A4AA68F05C96A001",
INIT_12 => X"002C006560138F032B1804101244C883052208209040CC849063A747512B7678",
INIT_13 => X"41401E240665750440C9488280254530314080C2C601040420352148A00501B1",
INIT_14 => X"500811204D000700114204A70422016149916011008CAA8858850B00C32591C0",
INIT_15 => X"FFC06E60AC0496022300233104663040808E991765205000070121D41D18D098",
INIT_16 => X"40100401004010040100401004010040102090010008000001C0E010020007DF",
INIT_17 => X"0100401004010040100401004010040100401004010040100401004010040100",
INIT_18 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_19 => X"FFEF9FEEFF7FFDF7FF3E3DFDF7E0000000000000000000000000401004010040",
INIT_1A => X"BEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBFFDFDFFFCF3CF3F",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFEFF7FBFDFEFF7FBFDFEFBEF",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000FFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0001000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E954AA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0004",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA0004154BAFFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"52E974BA0804000AAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0004174BAFF",
INIT_2B => X"FFFFFFFFFFFFFFFFEF552E954AA000400000007FFFFFFFFFFFFFFFFFFFFFFEF5",
INIT_2C => X"A082E95400007FFFFFFFFFFFFFFFFFFFFDFEF5D2E974BA002E97400007FFFFFF",
INIT_2D => X"FFFFFBFDFEF5D2A954AA002E974BA087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFBFDFFF5D2E954BA007FC00BA5D7FFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA000002000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080005000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"A974AA0000104AAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974BA0000174AAFFFF",
INIT_32 => X"FFFFFFFFFFFFDFEF552E954BA080A000AAE3FFFFFFFFFFFFFFFFFFFFFFFEF552",
INIT_33 => X"02A95400087FFFFFFFFFFFFFFFFFFBFDFEF5D2E974AA000A07000007FFFFFFFF",
INIT_34 => X"F7FBFDFFF5D2A954AA082A924281C7FFFFFFFFFFFFFFFFFFBFDFEF5D2A974BA0",
INIT_35 => X"A557FFFFFFFFFFFFFFFF7FBFDFFF552E974BA0020924BA1C7FFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000E3FFFFFFFFFFFFFFEFF7FBFFFFF552E974AA0071C50B",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0000020000000000000000000000000000",
INIT_38 => X"74BA0000174BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954AA080017410FFFFFF",
INIT_39 => X"FFFFFFFFFFDFEF552E954AA0004000AAF7FFFFFFFFFFFFFFFFFFFFFFFEF552A9",
INIT_3A => X"E95410087FFFFFFFFFFFFFFFF7FBFDFEF5D2A954BA082E800AAA2FFFFFFFFFFF",
INIT_3B => X"FBFFFFF552E954BA002E97410087FFFFFFFFFFFFFEFF7FBFDFFF5D2A974AA002",
INIT_3C => X"57FFFFFFFFFFFDFEFF7FBFFFEF552E974AA082A820AA557FFFFFFFFFFFFFEFF7",
INIT_3D => X"5D2E954AA0051554BA5D7FFFFFFFFFBFDFEFF7FFFFFEF5D2A974BA0000020AA5",
INIT_3E => X"0000000000000000000000000000000000000AAFFFFFFFFFFBFDFEFFFFFFDFEF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_2,               -- Port A enable input
WEA      => wbe_a_lo_1024_2(2),               -- Port A write enable input
DIA(0)   => data_write_a(21),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_2(21),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_2,               -- Port B enable input
WEB      => wbe_b_lo_1024_2(2),               -- Port B write enable input
DIB(0)   => data_write_b(21),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_2(21),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_22_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"5290F4CDE914905A14A43D33F488243E17122300F55FEB189B343A1140548380",
INIT_01 => X"A54007B259F6A975386262000C344BA9573C6FF57B18A5FB0ABFCD3C2C5F4F0C",
INIT_02 => X"021DFF8C38B3C009D203551040030071869D0040180AA2DC53DB89BEA8204001",
INIT_03 => X"2603475A969D0475A969D0460EAA401005111011BD506954EDB40F5EF41434C0",
INIT_04 => X"922D9002100ED69E443D988B0D5400103E48003D0800011E803B06B5B9125A15",
INIT_05 => X"281B5A0C06000408F4DF9422010D8802022F2124A8022492580040440002021C",
INIT_06 => X"F780C4C052881ADA0E05440205DA50930FA182010004700083E220800440B588",
INIT_07 => X"049D028B93FB561833D8094A02F5EA92FD7247E10305C40040D136E6A023F7FC",
INIT_08 => X"00028241680A0E002A9400803A884B5B5206B7C2E53CA25144009007A64EBD64",
INIT_09 => X"41008810240240C6694008010392354010000560141801002028A83D2A08E06D",
INIT_0A => X"34000000848BCA6902A29C54539C020E11810098D4067EFF9FF284D483E2AB41",
INIT_0B => X"500001840000C80B410014088040F4A944B1AA313C0022AA0011C0DC00028001",
INIT_0C => X"80B14004D158C8CA24A1C2A870AA1C2A870AA1C2A870AA1C2A872550E1543800",
INIT_0D => X"80A14050A01509E050854498B5281A1C34E506A2C6898B52A154DAC6B6000850",
INIT_0E => X"0B03001A483A4146603050080410089180008800143D83888281A2034A850142",
INIT_0F => X"A4160600349075238473F1210006133835E92273612B3482C090068A0E84AC56",
INIT_10 => X"30060181BA1B13959DC08DA902458870201970B29602562B0581200D141D0959",
INIT_11 => X"E042021C040D0152C8058B3840F044708E7E1C20A0106EA166C13AFC14AA3804",
INIT_12 => X"080E004B0C17C1439A9838301DC1A8438EA32C009DC1A8255300650458A1D588",
INIT_13 => X"018010E186F110A908E3A8CB0026C9A610A908E6A60F0807626610E160589C4C",
INIT_14 => X"2A701667334005800B1605F043858125E0D04110408D2485CA034681E43A1E40",
INIT_15 => X"00646002304244A91102C93A2D608D2A258DF8034188200C050171A41108F084",
INIT_16 => X"110441104411044110441104411044110466C440446CA06951D4EA8010009804",
INIT_17 => X"0040100401004411044110441104411044110441104411044110441104411044",
INIT_18 => X"0401004010040100401004010040100401004010040100401004010040100401",
INIT_19 => X"F7DFBFDEFE8FF1F7DEBDDF7DF7D05122890000000003FFFFFFFF900401004010",
INIT_1A => X"9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7BFFDFD7DDDF7DF7D",
INIT_1B => X"F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE79E7",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000003F9FCFE7F3F9FCFE7F3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA000400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0800",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000002000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2A954BA000015400FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080402010FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2A954BA0004154BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A0004174BAFFFFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0800154AAFFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF552A974AA0000174BAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974A",
INIT_2E => X"000007FFFFFFFFFFFFFFFFFFFFFFEF552E974BA0804000AAA2FFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080400010000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E954AA080005000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000402010FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2A954BA000417410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"804154BAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974BA0000174AAFFFFFFFFFFF",
INIT_34 => X"FFFFFFFEF552A974AA0000104AAE3FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0",
INIT_35 => X"AA2FFFFFFFFFFFFFFFFFFFFFFFEF552E954BA000E124BAE3FFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000007FFFFFFFFFFFFFFFFFFFFDFEF552E954BA080A000A",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804000100000000000000000000000000",
INIT_38 => X"54AA000400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2A954AA080017410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"0174BAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A954BA000415400FFFFFFFFFFFFF",
INIT_3B => X"FFFDFEF552E974AA0804174AAF7FFFFFFFFFFFFFFFFFFFFFFFEF552A974BA000",
INIT_3C => X"2FFFFFFFFFFFFFFFFFFFFFDFEF552E954AA0004000AAA2FFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2A954BA082E800AAAAFFFFFFFFFFFFFFFFFFFBFDFEF5D2E954BA002A820BAA",
INIT_3E => X"0000000000000000000000000000000000000087FFFFFFFFFFFFFFFF7FBFDFEF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_2,               -- Port A enable input
WEA      => wbe_a_lo_1024_2(2),               -- Port A write enable input
DIA(0)   => data_write_a(22),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_2(22),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_2,               -- Port B enable input
WEB      => wbe_b_lo_1024_2(2),               -- Port B write enable input
DIB(0)   => data_write_b(22),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_2(22),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_23_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"EF20906D902424807BC8241BC81801B97D38AD3C0800103362A6741C80A12A02",
INIT_01 => X"001FFF8409F089003B4422000D80C80106804A7951C5B9D1C828043EA28838F9",
INIT_02 => X"E01CEE21649C82C40800000F9FFEFF8E72CA7F5FC2E22809925A0D3611C877F8",
INIT_03 => X"24000400402670400402670D48222DC1764446838624000080007460C40001BF",
INIT_04 => X"68403FFC020560E0443E21037C01FFFC0002EE00628BF0E02FAD781014085014",
INIT_05 => X"0112000202FBFFF00920017FF0F0628BFF8488890979800002F702002BB807A0",
INIT_06 => X"EF85788B681FC000000001FFF0010000000001F7CBC385F87C0BFFFF20040001",
INIT_07 => X"F6E200000000C1440E3AE408009120071070FA07A1CB23FFA403F0C4D23BF7C0",
INIT_08 => X"0BF87CA400804000003FF7FFD8880A034AC09662305AB10555421006891A1089",
INIT_09 => X"BE1F5FEA10092C0896A243FFC0008087FFBEF2000000001DFFC612C0C0400100",
INIT_0A => X"41FF0C2060501000600000000001BFFA800808189A657EF81DD0C00079CC8001",
INIT_0B => X"018C24110A860006C620C0312241C482B20400CC52492710CC80060020A81BFE",
INIT_0C => X"0C08866907048320C20C10030400C10030400C10030400C10030400608018210",
INIT_0D => X"040002000041500300100040000500C000801000C02400000952800001FFBF04",
INIT_0E => X"FC850015385380380CDB86106502C5043FFD5FFF00A04BC010A7724B10000800",
INIT_0F => X"89F90A002A70A710A51C01C05904014861433602A1CAF13F2110055614C72FC0",
INIT_10 => X"E02D02001C1E14981B43253EE50C8220180F1082E06397E07E42200AAC298E57",
INIT_11 => X"8421802400A90022B0070FAE18019214A380344920080B21A58B02AC60BACDF0",
INIT_12 => X"0A2A000C480B0704B54028101AC49C84BB4100009AC49C80857A82D20CE8CB22",
INIT_13 => X"01E00C8103416445C12ED0400027C5292445C12D500B0005A62D344CB241D095",
INIT_14 => X"132C907425604680038706A35132C94BDD011010404428886AC91B11311C8280",
INIT_15 => X"FF000470BE0692020328CA0028042054A92771C50FC070110001C1680809591D",
INIT_16 => X"00802008020080200802008020080200800800200200000000000008004807DF",
INIT_17 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_18 => X"8020080200802008020080200802008020080200802008020080200802008020",
INIT_19 => X"0000000000000000000000000000000000000000000000000000008020080200",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080002010FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974AA000400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000400010FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974AA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080000010FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E954AA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954A",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA000015400FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080002010FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974AA000400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000402010FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E954AA080005000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA080407000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA00041741",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080000010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000402010FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2A954AA080002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954AA080017410FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"552A954BA000415400F7FFFFFFFFFFFFFFFFFFFFFFFFF552A954BA080015410F",
INIT_3E => X"0000000000000000000000000000000000000F7FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_2,               -- Port A enable input
WEA      => wbe_a_lo_1024_2(2),               -- Port A write enable input
DIA(0)   => data_write_a(23),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_2(23),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_2,               -- Port B enable input
WEB      => wbe_b_lo_1024_2(2),               -- Port B write enable input
DIB(0)   => data_write_b(23),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_2(23),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_24_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100600007FFF000080108004000800020000840041000080808",
INIT_02 => X"FC5CA803400EB8209000000F9FFEFF8E7240FF1FC22409EA04018E50074017F0",
INIT_03 => X"11100400000000400000000D00002CC07400000090C080019001010A000001BF",
INIT_04 => X"68003FFC00040000000000008001FFFC0002EE00000370E007A100000000E468",
INIT_05 => X"0000000000F8BFF00920004DF0F00001DF8000000079800000F3000029980780",
INIT_06 => X"6E461803081FC000000001FFF0000000000001F7C3C380F87C019FFF00000000",
INIT_07 => X"600C2400013649609C8000980040814210254000A00B21FF2003F2A80D500000",
INIT_08 => X"0BF80000000000000003F7FFD88D2B4A02C0940062EC2804001610020408178B",
INIT_09 => X"8E1F5FE010092C0892A041FFC0000001FFBEF0000000001DFFC002C000000000",
INIT_0A => X"41FF0C0000000000600000000001BFFA0000005501AA00000CE2000009400000",
INIT_0B => X"018C0411020600048620C030020502000200000400490510CC00040020201BF4",
INIT_0C => X"0808064106040300C00C10030400C10030400C10030400C10030400608018210",
INIT_0D => X"0000000000004003000000000000001200580000000000000000000001FFBE00",
INIT_0E => X"0086C022005381380FDB96516140C6043FFD5BFF000041000000004110000000",
INIT_0F => X"80010D804400A7240C840C201D0210840043B4804012500021E0088014C04940",
INIT_10 => X"4109038041021C980200D06410C1924030008142E06024A00043C01100298092",
INIT_11 => X"587CC200002100C14428090A1D02348190814C09C010104025AA40041A0D8005",
INIT_12 => X"022E0030300B0E46177004208000D8C61D7004300000D884817B00011306B2D9",
INIT_13 => X"01E003060344710009875C018100013831000985DC000C20003C310006143B70",
INIT_14 => X"4001850EDC004780144806A64400186CBF8961104000C3807884000846EB9500",
INIT_15 => X"FF0006E08C063C0220002201490418082010A57263E0100008000290161E711C",
INIT_16 => X"00000000000000000000000000000000000000000000000000000000000007DF",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"F2D0AEEAF6E7CC1132CDB4441990000000000000000000000000000000000000",
INIT_1A => X"BEFBE79E79E79E79E79EFBEFBEFBEFBEFBEF9EF9EF9EF9EFA69861219575D75F",
INIT_1B => X"783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1EFBEF",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000783C1E0F0783C1E0F0",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0201000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A000400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA000400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000400000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402010000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"00002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080002010FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000400010FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA00040000",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020100000000000000000000000000",
INIT_38 => X"74BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"000010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA000002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974AA000402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000002010F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_2,               -- Port A enable input
WEA      => wbe_a_lo_1024_2(3),               -- Port A write enable input
DIA(0)   => data_write_a(24),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_2(24),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_2,               -- Port B enable input
WEB      => wbe_b_lo_1024_2(3),               -- Port B write enable input
DIB(0)   => data_write_b(24),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_2(24),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_25_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100200002000000080100004000000020000800041000080808",
INIT_02 => X"FC400086000000800000000F9FFEFF8E738FFF1FC204010000000111568DD7F8",
INIT_03 => X"00000400000000400000000D00002CC4740000008000000080000000000001BF",
INIT_04 => X"68003FFF64A564AC000000000001FFFE0082EF00010370E007A1000000004000",
INIT_05 => X"0A00040148F8BFF80920804DF0F00101DFC040000079C92484F30499299837C1",
INIT_06 => X"66041803081FC0E0801101FFFD000E41002299F7E3C380F87C019FFF81200096",
INIT_07 => X"000000080480AE00000080000000000000000000A00B21FF2003E00000000000",
INIT_08 => X"1BF80000400A02000003F7FFFA0008000200A0400008A0000014100200081000",
INIT_09 => X"8E1F5FFA53EFBCACB2E369FFE0010001FFBEF80C40630C7DFFEEBAF000800202",
INIT_0A => X"41FF0C0600000000600000000001BFFE00301000000000000CC020000140000C",
INIT_0B => X"01DCCC31222730A49620C030020100000200000400490D10EC00040220201BF4",
INIT_0C => X"0808064106240300C00C10030400C10030400C10030400C10030400608018210",
INIT_0D => X"0883044582114013412080000000000000000000000000000012800001FFBE00",
INIT_0E => X"00040020000180380FC386106140C6043FFD5BFF00A04B80608003CB120C1106",
INIT_0F => X"0000080040000200040400000100000000009480000240000100080000400900",
INIT_10 => X"0001000000000808000000240000020000000100006004800002001000008012",
INIT_11 => X"0001001808220000002004001900000080800008000000000022400000088000",
INIT_12 => X"0010000000000E00110000000000408009000000000040808063004000008200",
INIT_13 => X"6000000000046100000240000000001021000004400000000010210000001010",
INIT_14 => X"4000000404000800000000060400000088000001800000001084000000088000",
INIT_15 => X"FF800C608C041002000002000006100000002100000000180600000000100018",
INIT_16 => X"4110441104411044110441104411044510629041040D180400000010028047DF",
INIT_17 => X"1104411044110441104411044110441104411044110441104411044110441104",
INIT_18 => X"1044110441104411044110441104411044110441104411044110441104411044",
INIT_19 => X"FBA2894A196A8C5A2932EC15DA080800002FFFFFFFFFFFFFFFFFC11044110441",
INIT_1A => X"2492492492492492492410410410410410410492410492412000531215A69A6B",
INIT_1B => X"158AC562B158AC562B158AC562B158AC562B1588C46231188C46231188C49249",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000B158AC562B158AC562B",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080000010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000010FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08000000",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_2,               -- Port A enable input
WEA      => wbe_a_lo_1024_2(3),               -- Port A write enable input
DIA(0)   => data_write_a(25),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_2(25),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_2,               -- Port B enable input
WEB      => wbe_b_lo_1024_2(3),               -- Port B write enable input
DIB(0)   => data_write_b(25),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_2(25),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_26_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"E9264EAB20190CA3BA4997AA9002AE9C001006B0778015CFA17E0811039879C7",
INIT_01 => X"2FFFF9BB1F773C7F9BB07DFFFDD863FC5FFF3FEFFBBF9FFB22FFFBC7B9F30686",
INIT_02 => X"E06CCC62052E708180F6FFBFFFFCFFFFF9C7FF7FC24332E642090000074037F6",
INIT_03 => X"428003739CD9863739CD9869FE2B7DEAF300029E4E300DFE69A6E644E6FF473F",
INIT_04 => X"7C2FEFFFF5BA124F003DD31EAFFFFFEE9FF7EE6F4C0770FFD7DC7CA53997B2B1",
INIT_05 => X"DFFB5421C1F8BBFAFDBFFACDF0FFCC05DDDBFF3690F9EDB7F5F7AFF639BD7DE3",
INIT_06 => X"EFD044ABC817C3E3A74667FDFFB6FF5727CC3BFEF7C3FAF87FF59F7FFBFEF69F",
INIT_07 => X"00003002132462052E708180EF060C18E5BEFB051225CDFF7002C4EEDE77F6E0",
INIT_08 => X"3FFF7D5000EC75088ED3FF7FC8790E46426CE06CB1F8E041051831FA3068D77E",
INIT_09 => X"C05FD7FF9BEFBDCEFBEE59FEF44F6603EFBEFAFCC2E35E7FDFD147CCF3F583FA",
INIT_0A => X"67FF1C7FBFADEB31E35768E8ED6BFDF3EB3EBF9DDBCE7FDC1DF8A760F3EACC02",
INIT_0B => X"5BDDCC3B336F7C548667D47B7737AF3FD62601EDC25B3533DCEB07F262213FFC",
INIT_0C => X"5F9A06E19F4D93A0EA0F78C35E30D78C35E30D78C35E30D78C35E986BC61AE31",
INIT_0D => X"5FD7AFEFDFFAF59B6FF28FE1D80D73D840607307DCFE1D80EF69A004DFFFF7FF",
INIT_0E => X"0004001F8041897B2FFFC6D86D70CE04FFFFF3FF1F5F5475BD7F72E4D75EBFAF",
INIT_0F => X"F60008003F008237B0040A00010003E020023E0201F45EC0010007E01047D17B",
INIT_10 => X"00010001DC0004C81003DE050A700200001DC0006863E8BD8002000FC0208FA2",
INIT_11 => X"2200E400002801E1A00004C21C0206F60081800800007B00010F02007EC09A0E",
INIT_12 => X"0880007E000807C7C1A612001E0015C7C19C22001E0015C59DFE82011A311AA0",
INIT_13 => X"00001BC00101F60409F0670840070809760409F06984800780097604067D0010",
INIT_14 => X"81019F40042100001F800203D81019EC085614000085C80023D81009CF008A74",
INIT_15 => X"FF802FFDFFAFD082003B032FB987E04021D481D4000819060801E0D00001231D",
INIT_16 => X"EBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEFFBFBFBFBBFCFBB0FFDFEFFEF2DFFFFFB",
INIT_17 => X"BFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAF",
INIT_18 => X"FAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFE",
INIT_19 => X"475B15BCF491E166CC8553F86EDB5C88646FFFFFFFFFFFFFFFFFEBFAFEBFAFEB",
INIT_1A => X"861861861861861861861861861861861861869A69A61861AFBD54D5F871C71D",
INIT_1B => X"984C26130984C26130984C26130984C26130984C26130984C26130984C261861",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000984C26130984C26130",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040201",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_2,               -- Port A enable input
WEA      => wbe_a_lo_1024_2(3),               -- Port A write enable input
DIA(0)   => data_write_a(26),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_2(26),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_2,               -- Port B enable input
WEB      => wbe_b_lo_1024_2(3),               -- Port B write enable input
DIB(0)   => data_write_b(26),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_2(26),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_27_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"00080A40000A41248002029000050A088000008242A0004404480002000A1155",
INIT_01 => X"2FFFF1C11F781C129C107DFFFE0860941E81258CA2B71C2220EC1B86E1A00002",
INIT_02 => X"E1000000810000014400FF6FFFF0FFFFF8007F1FC21110005080200000221FF0",
INIT_03 => X"4080026318C18226318C1821302232EAE00002BE001115FE48620040840A863F",
INIT_04 => X"643D4FFC2530000F003D821C0BFFFF8E9EF79E6D440748FED70060842105B0B0",
INIT_05 => X"D6F39020D1F8A3FAFDBFBACDC8FDC405D1DB7F1490E5EDB7D5CBADB2385D79C3",
INIT_06 => X"6FE000A38007C3032646EFF1F0B6FF46A78C39F8E723F2E47FE59C7F9ADA2612",
INIT_07 => X"00002820000000810000014401060C180190310540118DFF1000C0849673F6C0",
INIT_08 => X"3FF779100062B12A8EC3F47FC80208808210880C00082050000110023068D030",
INIT_09 => X"005F07E09BFFBD07FBAC09F8E42922038F7DF8BEC2E39C5F1FD047CEF1B582D8",
INIT_0A => X"63FF5D5F9FADE911E81C09818109E1F16B16B71092CE7ED81CF403601228C402",
INIT_0B => X"1BFDCC39732F3554866AD57C37BEAF1C152201A4C05B7531D56B05B06A213FF8",
INIT_0C => X"5BCA06F18FC59380F00E34430D10C34430D10C34430D10C34430F0861A2186B5",
INIT_0D => X"5B56ADAB5FAAE58B2F628EA0C80FA3F04040510768EA0C80CC61A0044DFFC6EB",
INIT_0E => X"0004001D800188792CE79715710AE4047FFD23FF315D54358D593474955AB6AD",
INIT_0F => X"520008003B000297B0040200010003E020001F0201E44A400100076000579129",
INIT_10 => X"00010001DC00004A10035E0408300200001DC000086BC8948002000EC000AF22",
INIT_11 => X"02002400002801E1A00000C01E0202F60080800800007B00000782006EC0820A",
INIT_12 => X"0080007E000006A7C10602001E0001A7C10C02001E0001C18DE282010A311AA0",
INIT_13 => X"00001BC00000FE0401F04300400708007E0401F04180800780007E04047D0010",
INIT_14 => X"81011F40040100001F800002F81011EC080604000085C80001F810094F008034",
INIT_15 => X"FF800C6DDDAFD082001B03249887E04001D481D4000009020801E0D00001021F",
INIT_16 => X"AB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6BF1EBDABD8E270BF84A25C6ACB777E3",
INIT_17 => X"B6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6AD",
INIT_18 => X"6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADA",
INIT_19 => X"490E2168100481CA860402104A471688747FFFFFFFFFFFFFFFFFAB6ADAB6ADAB",
INIT_1A => X"000000000000000000000000000000000008200000000000200072F210000001",
INIT_1B => X"05028140A05028140A05028140A05028140A0500804020100804020100800000",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000A05028140A05028140A",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040201",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_2,               -- Port A enable input
WEA      => wbe_a_lo_1024_2(3),               -- Port A write enable input
DIA(0)   => data_write_a(27),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_2(27),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_2,               -- Port B enable input
WEB      => wbe_b_lo_1024_2(3),               -- Port B write enable input
DIB(0)   => data_write_b(27),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_2(27),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_28_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"02200AA400180030808802A900002A08001280A08A801044104A1000001818C3",
INIT_01 => X"0AA00011460214428114180000882214413D0A71592A01D92213D28005210202",
INIT_02 => X"0451110A012100884000AA30200000000C100040104112101100008888200000",
INIT_03 => X"448000318C52A20318C52A20148810200111100C211004AA00034204200A2200",
INIT_04 => X"04004001001A90110000121402AA0000003C00000500000040080421080D0080",
INIT_05 => X"4060000C8001000000002E000000050000001610300000010000802202040012",
INIT_06 => X"1000002080001111001222000425A1040026A008000000000000000009328280",
INIT_07 => X"2491008A00491201210088400122448908A20402000408001000040820000000",
INIT_08 => X"20058310402A160026500000028040101004200C840082115554000112244814",
INIT_09 => X"4140000800000060000720000102028000000490160801020002200011100010",
INIT_0A => X"020000081B34211082B694D4D294000020020381040000000200032040004400",
INIT_0B => X"4800210C19808400500010009110091500020B408810000100200020408B0000",
INIT_0C => X"01028000080118020023604858121604858121604858121604858090B0242C00",
INIT_0D => X"010000800920040804020A6058003108402043058C460580653020005A004039",
INIT_0E => X"00000002800008014004104104420A00C000200005000010040A0020CC000200",
INIT_0F => X"520000000500000010000200000000000000280000040A40000000A000001029",
INIT_10 => X"00000000000000C0000002000830000000000000480008148000000140000020",
INIT_11 => X"020024000000000000000440000000020000800000000000000C00000040020A",
INIT_12 => X"00800000000001804006020000000500400C0200000005400A90000000100000",
INIT_13 => X"0000000000018200001003004000000142000010018080000001420000200000",
INIT_14 => X"8000080000010000000000018800008000060400000000000310000008000034",
INIT_15 => X"000002040080000000110006B081400000400000000009020000000000002200",
INIT_16 => X"802008020080200802008020080200802101210810C39A66A90A85420413A820",
INIT_17 => X"0200802008020080200802008020080200802008020080200802008020080200",
INIT_18 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_19 => X"DE21102C110A00246972BD89A40A0C22E1000000000000000000002008020080",
INIT_1A => X"2082082082082082082082082082082082082082082082080D35050758C30C31",
INIT_1B => X"0582C160B0582C160B0582C160B0582C160B0580C06030180C06030180C08208",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000B0582C160B0582C160B",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_2,               -- Port A enable input
WEA      => wbe_a_lo_1024_2(3),               -- Port A write enable input
DIA(0)   => data_write_a(28),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_2(28),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_2,               -- Port B enable input
WEB      => wbe_b_lo_1024_2(3),               -- Port B write enable input
DIB(0)   => data_write_b(28),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_2(28),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_29_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"79964E4BA01DACAB9E659792D00AAE160002829C7FDFEFCEE97C2815039D70C3",
INIT_01 => X"0ABFF9AB0775343F9AB01DF80D5821FC0FFF3FEFD1AF9FF1207FFBC7B9720586",
INIT_02 => X"002CCC60050E700080F6AAA7BFFC007189C7FF2FC00330E602800000074037F6",
INIT_03 => X"468003210868A63210868A68DA017D207200021C4E200CAA6186A40042FF4300",
INIT_04 => X"7C2FE002F0900001003C5316A6ABFFE21F36E02F0D03701F47D41800109FB281",
INIT_05 => X"4979440580F9B808F49F6A4DF00F8D01DC4B97369078249370F482E62BA41462",
INIT_06 => X"B250442BC81001E1870223FC0BF7F11507C423FE33C078F803F19F00E936721D",
INIT_07 => X"00011080012460050E700080EF020408EC8CFA01122149FF700200665A35D260",
INIT_08 => X"2BFD055040A452000443FF00007906464068406C31F84000000831FA1028575A",
INIT_09 => X"805FD017102690AA694551FE30444681E0820AD40201423FC00122C493500172",
INIT_0A => X"0600002AFFBE2330815568A8AD6ABC02A02A0B0CCB463B4C0748A720B1EA4C00",
INIT_0B => X"0850400A11414C005005000B51158936D20601A98A10200308A002E240010BFC",
INIT_0C => X"05928020194918A22A2268C81A32068C81A32068C81A32068C81A99034640C00",
INIT_0D => X"058102C48970541944B20FA1580561D040406305587A158046282000DBFFF13D",
INIT_0E => X"000000028040890327DCD28928324400DFFFF0001F1F0050342D42A086040B02",
INIT_0F => X"F60000000500802010000A000000000000022A0000141EC0000000A01000507B",
INIT_10 => X"00000000000004C0000082010A700000000000006800283D80000001402000A0",
INIT_11 => X"2200E4000000000000000442040004020001800000000000010D000010401A0E",
INIT_12 => X"08800000000801C040A6120000001540409C2200000015441DAC800010100000",
INIT_13 => X"0000000001019600081027084000000956000810298480000009560002200000",
INIT_14 => X"800088000021000000000201D800088000561400000000002358000088000A74",
INIT_15 => X"00802594A282C0000033010FB181E00020400000000819060000000000002305",
INIT_16 => X"C0B02C0B02C0B02C0B02C0B02C0B02C4B12B312912831A27FCFE7FFB175B6FF8",
INIT_17 => X"0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02",
INIT_18 => X"B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C",
INIT_19 => X"BBCF9F96EE7FFDF7FE783FFDFFEA0C00602FFFFFFFFFFFFFFFFFC0B02C0B02C0",
INIT_1A => X"EFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEEBAEBAEBAEBAEBBFFDF9FBEFFFFFFE",
INIT_1B => X"BFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFBEFB",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000FBFDFEFF7FBFDFEFF7F",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_2,               -- Port A enable input
WEA      => wbe_a_lo_1024_2(3),               -- Port A write enable input
DIA(0)   => data_write_a(29),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_2(29),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_2,               -- Port B enable input
WEB      => wbe_b_lo_1024_2(3),               -- Port B write enable input
DIB(0)   => data_write_b(29),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_2(29),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_30_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"F7FFBFFEFF9FE1F7FFBFFFFDFFD0000000000000000000000000000000000000",
INIT_1A => X"9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7AFBD75F5FDF7DF7F",
INIT_1B => X"F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE79E7",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000003F9FCFE7F3F9FCFE7F3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_2,               -- Port A enable input
WEA      => wbe_a_lo_1024_2(3),               -- Port A write enable input
DIA(0)   => data_write_a(30),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_2(30),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_2,               -- Port B enable input
WEB      => wbe_b_lo_1024_2(3),               -- Port B write enable input
DIB(0)   => data_write_b(30),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_2(30),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_31_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"129000008004A00804A40000400800020000000C005FEA005800200400050100",
INIT_01 => X"255FF18019700810180065FFFC0040801E80258CA2951C2200EC0906A0804140",
INIT_02 => X"E0000000000000011000550FDFF0FFFFF0007F1FC200000044000000000817F0",
INIT_03 => X"0000024210A30024210A3001002220C06044469200040154482000408400043F",
INIT_04 => X"602D0FFC2420000E003D80080955FF8E1ECA8E2D400340FE870060842100B030",
INIT_05 => X"0213100040F8A3F8FDBF944DC0FDC001D1CB6904A061EDB6D4C30490281831C1",
INIT_06 => X"6FC000830007C202060445F1F0D25E4207A099F0E303F0E07FE19C7F80402412",
INIT_07 => X"0000200000000000000001100004081001103107000185FF0000C0849673F6C0",
INIT_08 => X"1BF27A00000000000883F47FC800080002008000000820440000100220489020",
INIT_09 => X"011F07E013EFBC06FBA009F8E00120038F3CF82C44630C5D1FC002CCE0808248",
INIT_0A => X"61FF0C06C48BC801600000000001A1F00110101092CE7ED81CF0004012288000",
INIT_0B => X"11DCCC31222730048620C4382204A608142002A440492530C401049020221BF8",
INIT_0C => X"0888066187448380E00C10030400C10030400C10030400C10030600608018210",
INIT_0D => X"080204010200418301208480800D02D00040100240A808008840800405FF8640",
INIT_0E => X"0004001D000180780CE386106100C4043FFD03FF101D40008001304018081004",
INIT_0F => X"000008003A000217A0040000010003E02000160201E040000100074000478100",
INIT_10 => X"00010001DC00000810035C0400000200001DC0000063C0800002000E80008F02",
INIT_11 => X"00000000002801E1A00000801C0202F40080000800007B00000302006E808000",
INIT_12 => X"0000007E00000607810000001E000087810000001E000081846282010A211AA0",
INIT_13 => X"00001BC00000740401E0400000070800340401E04000000780003404045D0010",
INIT_14 => X"01011740040000001F8000025010116C080000000085C80000C8100947008000",
INIT_15 => X"FF800C609C06D082000A03200806A040019481D4000000000801E0D00001001D",
INIT_16 => X"010040100401004010040100401004010060C040040C200950402090128057C3",
INIT_17 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_18 => X"0040100401004010040100401004010040100401004010040100401004010040",
INIT_19 => X"00000000000000000000000000001000802FFFFFFFFFFFFFFFFF810040100401",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_2,               -- Port A enable input
WEA      => wbe_a_lo_1024_2(3),               -- Port A write enable input
DIA(0)   => data_write_a(31),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_2(31),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_2,               -- Port B enable input
WEB      => wbe_b_lo_1024_2(3),               -- Port B write enable input
DIB(0)   => data_write_b(31),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_2(31),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_0_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"ED39BA795990D275FB4A6E96ACC4731DEA4598B0AFB54867F6EE4618C3749803",
INIT_01 => X"8AA0047D8607944AC7DA180001ECA2444042106208408208C20022E9173734B3",
INIT_02 => X"1A7DDD79F9A73E6CCA7DAAF00001000008478020113D98E382FEDF333027C80F",
INIT_03 => X"75D341110C58F31110C58F32A208921F8051500147A0E4AB3493FB3A01EBE240",
INIT_04 => X"86424001531009B100425A97B2AA0001E03501D0A39C8F0078420001106D0C4C",
INIT_05 => X"BCC8CA2EBF03400700402BB20F00239E20341699198600000B08694B16434804",
INIT_06 => X"103FB860B2800161F8432200012DA185F80F24081C3C0707800E600056881308",
INIT_07 => X"B24197ABCDA467F9A73E6CCAFDC3870EEEEC44E2BDFE220094D03022210C011C",
INIT_08 => X"240581B5695EAA80262C080032BF07C7C1FC3F8E94F65B11555EAFFC1C306758",
INIT_09 => X"7E40000BEC004170040DB60017FED1CC0001045002984202003DB931192D60A5",
INIT_0A => X"120071411A74315881A28C141118000C5A85A60444210123820B43B40804674D",
INIT_0B => X"0820008E514045BB514F0106D1D8599581D3A958BC104A89215AC14C48898403",
INIT_0C => X"C261C01C48B1584A0CA3E2687A9A1E2687A9A1E2687A9A1E26870CD061343885",
INIT_0D => X"D274E93A758FA8683AC54B287522E10A74AF4AA59C568752662F5AC218000002",
INIT_0E => X"FF83C002783A0904231C70470C7E0B92800224008AE09FAD4BD48D1FC5D3A4E9",
INIT_0F => X"5BFF078004F075885DFBF7E15C06101C55E921F1F80FAB7FE0F0009E0E903EAD",
INIT_10 => X"F12E0380231F13978FF023FAFDBD9870380230F2D6081F56FFC1E0013C1D207D",
INIT_11 => X"DE7F263C0C8700125C0F8F3C43F1F10BBF7EFC61E01804E1E6C8F8FE807F67FB",
INIT_12 => X"02BE00017C17C1007E5E2E3081C5AC007E6F0E3081C5AC44418D65FE45DEE55B",
INIT_13 => X"61E0042786F103E9F01F9BC3C120C5A703E9F01F978B8C20666703E9F8A0FFED",
INIT_14 => X"FA7E283FFB414F80005F05F10FA7E283F78F6511C048278DCA174FF038FF15B4",
INIT_15 => X"0066A20B61692F293185D8D724E15D3FCC6B7C236FE0691B0700132C1F0EF880",
INIT_16 => X"3A4E93A4E93A4E93A4E93A4E93A4E93A4F942F92E9628540AD2A91442525A000",
INIT_17 => X"A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E9",
INIT_18 => X"4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93",
INIT_19 => X"55F3898E09B56C74DAB15D1CF13501AA495000000000000000003A4E93A4E93A",
INIT_1A => X"082082082082082082082082082082082082082082082082082084E41DC71C71",
INIT_1B => X"E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F82082",
INIT_1C => X"FFFFFFFFFFFFFFF94A5294A5294A5294A5294A52800003E1F0F87C3E1F0F87C3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"3060C183060C187FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"BDEBA0000000000000000000000000000000000000000000003060C183060C18",
INIT_28 => X"168ABA002E82145085155545F7AA975EFFFAABDE00FFAEBDFFF5D2EAAAAAF7AE",
INIT_29 => X"7FFFE10005542145557FD5545FF8000155087FC0155F7D168B55007BFDF45085",
INIT_2A => X"7FFC0010080017555555568AAAFFFFD7545AA8028A00A2802AABAFF8028BEF5D",
INIT_2B => X"FF842AABAA2AE95545FFD168ABAF7AEAAAAAA2FFFDF4500043FE105D2E954BAF",
INIT_2C => X"5007FD7400550415410002E974BA5D5168A00A2D142155005142010FFAE820AA",
INIT_2D => X"FFF780000BA007FE8AAAFF803FFFF5D2A821550000000BA007FD55FF5D7FC014",
INIT_2E => X"000AAFBEAA00007BFDFFF082EBDF455D5142000082E82145FFD17DFEFFFD168B",
INIT_2F => X"DFD75D2AA8A80EA8E2FE3F000000000000000000000000000000000000000000",
INIT_30 => X"68B551475FAF6D1C556F0AA1C24AABEA495FC716F002A975FFE3AA95E00EBAEB",
INIT_31 => X"42A0070071C50BAFEF1FAE0016D56A16D557BC257D415E0216FA3F1E8FC0145B",
INIT_32 => X"8010E004924874825D7FEAA85487FD24AFE3D02DAAAE12BD5545A2803AA00005",
INIT_33 => X"120155EA568E870BAEB8A05A2AEA8B50F55A2F150005A3A438BD04AFAB8F550A",
INIT_34 => X"545E055FFBE81D0BE8EA8A3AA05A2A5504001C74BA42A1571E8028E3DB7816D0",
INIT_35 => X"A5C7E3DFFFE90B45B47ABA497A82FFAFD2A82485FD2415A105C21451ED42A002",
INIT_36 => X"00000000000000000000B55EAAA100AA1D0F6F480B6A555A2A57A002A3D5FDB6",
INIT_37 => X"5EFAAAAB5E1AF3AABFF45592E88A0AFE80A8B0A0000000000000000000000000",
INIT_38 => X"65F520EBE9EF67D7BEA1FD5D556ABEF5D557FEBA55022A3F70C6B405F4D2AE97",
INIT_39 => X"C114728007521170821CE0FDE69411A8DED57CE1055555E5F58EFFC01FE2CACB",
INIT_3A => X"42341D5DEEBEF55080034E0A592A4AD0079C75D6070CC5CBB0280C029ABAA3EB",
INIT_3B => X"7F353AAF6C77F7F20D968BF57812A95E02A2AAB5EB0F280800EFAEE9F5D18F31",
INIT_3C => X"C91565455C141E41887D58AC448B69C30E02116220415A9540AA854140A0A204",
INIT_3D => X"DE6BE93172D7D625B556EEAB157ABEBE1B4D792A4AD1183454180DD3FDCAAAB7",
INIT_3E => X"F0000001FF0000001FF0000001FF0000001FF01EABC4B8014174FF7DA80F52FE",
INIT_3F => X"FF0000001FF0000001FF0000001FF0000001FF0000001FF0000001FF0000001F")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_2,               -- Port A enable input
WEA      => wbe_a_hi_1024_2(0),               -- Port A write enable input
DIA(0)   => data_write_a(0),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_2(0),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_2,               -- Port B enable input
WEB      => wbe_b_hi_1024_2(0),               -- Port B write enable input
DIB(0)   => data_write_b(0),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_2(0),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_1_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"212C001411984004084D000508C53810A03D1450E839B003342114428A000803",
INIT_01 => X"00000019400B100A8196000000CC004400400002000000000000028001340000",
INIT_02 => X"052137AE8031800C0044009000000000061800001CD4019802AD04CCCFC20004",
INIT_03 => X"04514108C60C21008C6042108400000201440020505100000043C30E10E9F000",
INIT_04 => X"02104001011DEFE088805681920000008000004001900800004002108C280008",
INIT_05 => X"040002340105000200000000080001900010000108040000000008411600401C",
INIT_06 => X"1034001042800808201000000001000820020000102000040000000000800180",
INIT_07 => X"64BF81A15EDFDE8031800C00843060C19E030022103600000450020800040004",
INIT_08 => X"00008004691687AA840008000090248CC84E000046000311555521F183060AC5",
INIT_09 => X"0820800D08100171000DB000154440C800400500000852020011200201012021",
INIT_0A => X"02000040001000880A2A04445004000102002041000001008208001440004140",
INIT_0B => X"4820018A1140440078050040511000102000A008183000010002404400000000",
INIT_0C => X"1000C80008000C030030880C2A030A00C28030A80C2A030A00C28018D4061401",
INIT_0D => X"10040802050080200284401C0022880F009E08008205C0020118088018000000",
INIT_0E => X"0F03C00280000000420860C60C0C0B92C0000000004000010042000040102008",
INIT_0F => X"001E078005000108400005E11C0610000000288058000003C0F000A000100000",
INIT_10 => X"F10E0380000000C202300000008D187038000000480800000781E00140002000",
INIT_11 => X"806302380C870010000004400100110800007861E0180000000C400680000001",
INIT_12 => X"023E00000000018000580C308000050000610C30800005000215006800000101",
INIT_13 => X"61E0000000018100B0001843812000014100B00016030C20000141002880026D",
INIT_14 => X"400A20009B404F80000000018400A20044096111C04000000304026000501580",
INIT_15 => X"0046820040082300218450C2800010094000482141E060190700100000002200",
INIT_16 => X"020080200802008020080200802008020080008008600500A82A1100A8000000",
INIT_17 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_18 => X"0080200802008020080200802008020080200802008020080200802008020080",
INIT_19 => X"81328A46BABEFC54A0810C7452B4428A14000000000000000000020080200802",
INIT_1A => X"AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA28A28A28A28A2A8218D2C0C924925",
INIT_1B => X"E974BA5D2E974BA5D2E974BA5D2E974BA5D2E975BADD6EB75BADD6EB75BAAAAA",
INIT_1C => X"FFFFFFFFFFFFFFFD8C6318C6318C6318C6318C63000002E974BA5D2E974BA5D2",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"70E1C3870E1C387FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"5555500000000000000000000000000000000000000000000070E1C3870E1C38",
INIT_28 => X"EBDF455D2EAABEFF7FFE8BFF5D0002155557FFFFFF007FC21EFA2FFD74AAAAD5",
INIT_29 => X"AA95400552AAAABAFFD1574105D7FD75FFAAAA800AAF7AA974BAFFFBE8B45F7A",
INIT_2A => X"0517DF555D2EAAA1055000015500557DF45AAD1400BAA2AE801550051555EFF7",
INIT_2B => X"FFD540155557FD5400F78028BFFFFFBEAB55F780020AAAA80020AA082EAAB550",
INIT_2C => X"AFF842ABEF5D517DF55552A974AAF7AE820AA0851574BAA2D1574AA5D7BFDEBA",
INIT_2D => X"EFAAD1575EF557FFFE10557FFFFFFFFD56AAAAFFFFD7555AAD168B45AAAEAAAB",
INIT_2E => X"0005D7FFDF4500043FE105D2E954BAF7AE80010082A97410557FEABFFAAFBE8B",
INIT_2F => X"51C7A2FBD5490BFD1C056A000000000000000000000000000000000000000000",
INIT_30 => X"974BAF7FFEFB45FFAABDF55492AA8BC2EBDFEAF7F1F840017D4975D2FEF147FC",
INIT_31 => X"080BEF495FC71D54124924385FAAA8AAAE3D145410F7F1D55D71C002DABAEBAA",
INIT_32 => X"002D082082AB8B6DBEDB7DF7F540E2AE85028B40155145F7AF6DBED5450AA1C2",
INIT_33 => X"78E021FF1471FDEAAFFD56F16D5571D2E28E38E0216FA2D1E8E80140F45082B4",
INIT_34 => X"A2DA3FB7DAAD4AAAAF487BC70BFA97F7AF6D417E92482BF84020BA495557E3FF",
INIT_35 => X"55554ADBD7A2FFC7BEFF6FFD7FC7002FD74951D71EDFFABFD16FAAAE92BD5545",
INIT_36 => X"00000000000000000000547AB8F550A8010E00492487482FFFE82A85EBAE2FFC",
INIT_37 => X"1EF005162BEF047FD5545AAFBF7400FBF9424F70000000000000000000000000",
INIT_38 => X"714F8338AAAA1D0AE974AAF7FFFDF55F7AABFF55082CA8B4DF6C1E8F5E540002",
INIT_39 => X"EABEF75550ACBB7582225FF5843404547184164AA5D2EBEEB0A2D555410D3555",
INIT_3A => X"FEAAEB083BC1000FF8409000512AEABFFDF79DCBF755962010BDCBBC21455D7F",
INIT_3B => X"801F8BA0C57740BDAA0688E5405D57D412F7D55F5E50C7F401BAAE8403CF5A3F",
INIT_3C => X"5D16BABAA3EBC3157ABD5FFE55F2AA9FEAFDF7F431A9F7FFE81FF013A8001AFF",
INIT_3D => X"FB863550229BCABEB7DA403FFFDA2FBF7FED2C7F955445079E280A00C56145EF",
INIT_3E => X"0000000000000000000000000000000000000596EBEF55080034E0A592A4AD00",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_2,               -- Port A enable input
WEA      => wbe_a_hi_1024_2(0),               -- Port A write enable input
DIA(0)   => data_write_a(1),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_2(1),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_2,               -- Port B enable input
WEB      => wbe_b_hi_1024_2(0),               -- Port B write enable input
DIB(0)   => data_write_b(1),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_2(1),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_2_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10E006600180111284380310006289800480032283E000A34301002001A0817",
INIT_01 => X"0005A00810790848048044A54E404350404000720885800802000906E4910200",
INIT_02 => X"407004208400408044C600C50AA055254010541A110222841200000002402544",
INIT_03 => X"0600011004182401004102408C28414043101000408118000145840440F5C415",
INIT_04 => X"5035855703A2900A000CD3088400F40688C9844409060850925E58A4081A0221",
INIT_05 => X"0200840D1021A15AC50494894850890540D1E12020C6E510818500440A280090",
INIT_06 => X"113044094002801020440090A8011A1224AB9380552102442884882A20004097",
INIT_07 => X"000100880004428400408044860000008C022402102100AA40004404B5075460",
INIT_08 => X"15C23440408C862A2A12382A8A5244145048C06085008010141521F000001240",
INIT_09 => X"400582B9033AA0E7AA4110B0506744810554542450694E710A836188C2C00222",
INIT_0A => X"443518360012C2210B020414109130A28038188096A06B8C120CA440A9C00802",
INIT_0B => X"1345E53300EC68005605002964AF222A5704004D080211121C80024200821780",
INIT_0C => X"181080C1110C882202211488452213C88472213C88472213488441109A442231",
INIT_0D => X"008204440210091341208041000810C00000300220201800A908000038AD0284",
INIT_0E => X"00040002804180300E88D28D206A40000554815500481440300000C44A081100",
INIT_0F => X"000008000500828700000000010000000002380000A00000010000A010050000",
INIT_10 => X"00010000000004CA000214000000020000000000684280000002000140200500",
INIT_11 => X"000000000020000000000442100002840000000800000000010C000026000000",
INIT_12 => X"00000000000805A4800000000000152300000000000015801272000100210020",
INIT_13 => X"000000000101C00000C000000000000940000120000000000009600004050000",
INIT_14 => X"0000130000000000000002018000106000000000000000002380000141000000",
INIT_15 => X"55000190000000000002000280000000011080C0000000000000000000002310",
INIT_16 => X"40902409064190641906419024090244902A9003004800415120D4A190804241",
INIT_17 => X"0900409004090641906419064190240902409024090641906419064190240902",
INIT_18 => X"9044090040900409004190441904419044090040900409004190441904419044",
INIT_19 => X"75960040138D70C030B51C50C7D100A2052F81F81F83F03F03F0419044190441",
INIT_1A => X"0410410410410410410410410410410410410410410410410248602081659659",
INIT_1B => X"5128944A25128944A25128944A25128944A25128944A25128944A25128941041",
INIT_1C => X"FFFFFFFFFFFFFFFE1084210842108421084210843FFF825128944A25128944A2",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"7FD5FF555815607FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"2AA000000000000000000000000000000000000000000000007FD5FF55581560",
INIT_28 => X"FC21EFA2FFD75EFAA8415410AA8415555087BFFF55A2AA800BAFFAE954000800",
INIT_29 => X"84155EFA2AEBDEAAA2FBEAABA5D7FE8B555551421455D0002145552EBFEBA007",
INIT_2A => X"2AEBDF555D2E954BAA2AA974BAFFFFE8B45552EBDF45FFAEAABFFF7FFE8B55F7",
INIT_2B => X"AAAAAAAAAFFD1574105D7FFFF555D2AAAAAA5D2E820BAA2FBEAB5555557DF55A",
INIT_2C => X"50055575EFFF84021555D043DEAA5D04021EF557FC21FFAA8428BFFAAAA954AA",
INIT_2D => X"10085568A00FF80175FFA2D17DFEFF7800215500557DF55AA80001FFAA800015",
INIT_2E => X"0005D00020AAAA80020AA082EAAB5500517DF555D042AA10A284154005D00154",
INIT_2F => X"00AAFFAA9543A080038A2A000000000000000000000000000000000000000000",
INIT_30 => X"0017D5D20B8EAA007FC51C7A2FBD55D2BE800042AFE8E1557D0075D2F45BEAA8",
INIT_31 => X"AA8BC7EBDFEAFEFFD00105FFBC20BDEAAA2FBF8AAA557BE8B6D5D5FFABEF4904",
INIT_32 => X"FFEFB6D555578F7DB6A0BDF7D480E174BFA02A974BAF7F5EFB455D2ABDF55492",
INIT_33 => X"ED1FDE90E3A497492B6AAADAAAE3D155E105571D55D71C002DABA5524820BAB6",
INIT_34 => X"BE8F401D7B6A0001470155C51D0092A071555D5E3AE821D00001FF0871C016DB",
INIT_35 => X"5BE8555400550A38428007FED000E3DA3DFD5E3DFFFBD5A38A021551C5F7AF6D",
INIT_36 => X"00000000000000000000410F45082B4002D082082AB8B6D1C5B7DF7FF78E075C",
INIT_37 => X"5EF005560B55F7AA800AAF7AA954AA00042AAA20000000000000000000000000",
INIT_38 => X"ABEF057D68F5F5A00021EF55042AAAA007FD5555AAFBD7545FBB8020A3F7AE97",
INIT_39 => X"7DF55D7AABFF5428ACA8F45A6C1E8F5EFF84165EFF7802BAB0A2FFEAABA557BE",
INIT_3A => X"CA8AA80800020AAF7FBFFFEF04552ABFFFF841FFE75CA882108202E974AAF7D5",
INIT_3B => X"00151FF0C57401E5F3D1E00A1A884174A8FFAEBFEB0A2D55541051555694F002",
INIT_3C => X"2AA801455D7FE8BFFF680800FFF7AAA155F595542455512A975455D3AA8A0055",
INIT_3D => X"5D79FCAF774AE005BE7895554005D2A8A0B882FFFFE10AAAAAB755A66B6AF56A",
INIT_3E => X"00000000000000000000000000000000000000C3BC1000FF8409000512AEABFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_2,               -- Port A enable input
WEA      => wbe_a_hi_1024_2(0),               -- Port A write enable input
DIA(0)   => data_write_a(2),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_2(2),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_2,               -- Port B enable input
WEB      => wbe_b_hi_1024_2(0),               -- Port B write enable input
DIB(0)   => data_write_b(2),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_2(2),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_3_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"210C00A20020000108430020001600B8156021104940741B3530400E02B92203",
INIT_01 => X"014C9BCA58B1296D24A402C992500B69404040028804A0080A000416A8D90A08",
INIT_02 => X"C12026A484318004404405C9C66E331352180D468B8203980300204442E02B34",
INIT_03 => X"04000748D60D24648D60524C88804D0215011020D15018148040C10A70E1D58C",
INIT_04 => X"18283333240FE41244187308C9104D70944852640901083801750EB0A418C220",
INIT_05 => X"0613142D01912CC2A1B4140528348900C612A104201C689044340ED413A07649",
INIT_06 => X"119000034019881822104C5E68035250A222829710A0A02C18C01A9920842413",
INIT_07 => X"402F00AB0016CA0431800444841020509D038B021230C1990001C644C8273200",
INIT_08 => X"16905000408482088290E8E64010248C4A5AA840C2000110001521F0810A92E7",
INIT_09 => X"0003CE6581BD016342A951AB146C4480530C3B2A8088D3542651670200C1826A",
INIT_0A => X"00735D36209A8A20020894004284B660821030C8990467401218004041020002",
INIT_0B => X"512445B740457154562F957CC08B00093700080D0A4851001D8302D20A0A1530",
INIT_0C => X"00508650008008021021A40861021840869021A408610218C0869810D6043095",
INIT_0D => X"1C8508438450801043A08090380A8834207007022209038080190000999C8F84",
INIT_0E => X"000400200000C0002A48A206204C4205F3304B33004C0041006240140A1C310A",
INIT_0F => X"0000080040000083800400000100000000008400018040000100080000510100",
INIT_10 => X"0001000000000800000244040000020000000100002A0080000200100000A702",
INIT_11 => X"000000000020000000200000080002C000800008000000000022000006808000",
INIT_12 => X"0000000000000A2281000000000040A3810000000000402001400000022002A0",
INIT_13 => X"000000000004200001C0400000000010200001C0400000000010000004490010",
INIT_14 => X"0001070004000000000000060000104C08000000000000001000000903008000",
INIT_15 => X"CC004050CA0C00020220200070040000010401C4000000000000000000100008",
INIT_16 => X"4310E4310A4210A4210A4210A4210A4210A8D0830A68010001B4DA881048061C",
INIT_17 => X"21084290A4210A4210A4210A4210A4210A4210A4210E4310E4310E4310E4310E",
INIT_18 => X"90A421084290A421084390E4310C4390E4310C4390E4310C4290A421084290A4",
INIT_19 => X"015303C0C78C706428A14C586291000A044001FFE000003FFC004290A4210842",
INIT_1A => X"2492492492492492492492492492492492410410410410412821600001249249",
INIT_1B => X"51A8D46A351A8D46A351A8D46A351A8D46A351A9D4EA753A9D4EA753A9D49249",
INIT_1C => X"FFFFFFFFFFFFFFFC00000000000000000000000038F56351A8D46A351A8D46A3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"55AB02055AB0207FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"420000000000000000000000000000000000000000000000007FFFAB57FFFAB5",
INIT_28 => X"A800BAFFAE9554508002AA00AA843DF55FFAA955EFA2D168B55557BEAA000055",
INIT_29 => X"002AB55AAAA955EF005568A00087BE8BFFA2D155410AA8415555087BFFF55A2A",
INIT_2A => X"AAABFF5508003FF555D0002145552ABFEBA007FC21EF007FD75FFAA841541008",
INIT_2B => X"082EBDEAAA2FBEAABA5D7FC0155005168B455D042AB45F7FFD741000042AA10A",
INIT_2C => X"FF7FBEAB55F7AABDEBA5D7FC2010A2D1575FFF7AA975555D2E80145F78415545",
INIT_2D => X"EF5555554AA087BC01FFFFAAAAB55552A954BAFFFFE8B55552EBDE00F7AEAABF",
INIT_2E => X"000082E820BAA2FBEAB5555557DF55A2AEBDF555D2E954BA002EAAABA002A821",
INIT_2F => X"FB7D5D7FEAA3808554203A000000000000000000000000000000000000000000",
INIT_30 => X"1557D1475FAF45BEAA800AAFFAA95578080038A2AA28E3AF55E3A0BA5D7AADB6",
INIT_31 => X"BD55D7BE80004AA1E8E2AB55B6A0925D7085F6AA10087FEABD7AAD57AEBAB68E",
INIT_32 => X"F5D0438140E2FA38B6AEBFF6D1D04AAFFA41040017D5D20B8EAA007FC51C7A2F",
INIT_33 => X"D0A901FFFF801557D1C20B8EAAA2FBE80AA557BE8B6D5D5FFABEF49002FB55FF",
INIT_34 => X"5D20BDE00EBAAA8BC7EBDFEAFEFAB8ABAE925D21C7010EADB525D7FFAE975C75",
INIT_35 => X"F002EADA921420871D74971D24820875C21D5EB8AA8FFF012A954BAFFF5EFB45",
INIT_36 => X"000000000000000000001C24820BAB6FFEFB6D555578F7DB6A0BDF7DEB8E125F",
INIT_37 => X"B55A28408145AAFFFFFFF5D7FEAABA0051400A20000000000000000000000000",
INIT_38 => X"AB55FAD568AA2AFAE975EF555168B55F7AA800BAF7AA955EF00042AAA2A2AEAA",
INIT_39 => X"2AAAA007FD55558A7BD7145FBB8020A35D2ABEF55F7800015F087FEAA00007FE",
INIT_3A => X"968F575D003FF55F7D5420BA5D2ABFEAAF7AE9DFF759A82AEF70800021EF5504",
INIT_3B => X"FFD5145FBAC9755F05040255FFD84175EF55002AAB0A2FFEAABA557BEA3EF057",
INIT_3C => X"82E974AAF7D57DF45552A3FF10AA8429F45A7D5EAF5FFBAEAAA10554155400AA",
INIT_3D => X"FF843FFE77C80825BC052ABFE10550415557085540000005156155FE90A8F5C0",
INIT_3E => X"00000000000000000000000000000000000005500020AAF7FBFFFEF04552ABFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_2,               -- Port A enable input
WEA      => wbe_a_hi_1024_2(0),               -- Port A write enable input
DIA(0)   => data_write_a(3),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_2(3),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_2,               -- Port B enable input
WEB      => wbe_b_hi_1024_2(0),               -- Port B write enable input
DIB(0)   => data_write_b(3),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_2(3),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_4_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"A108400020612C80284210081034849800A00030300004833522C82D04A16002",
INIT_01 => X"2043998A1839284D1CA0650E1E504368403008418984014902030806A0D10200",
INIT_02 => X"C120042200000000044441CE01E80F00A49043118680008002000000026208E4",
INIT_03 => X"040001020019200020011209CC0164C060000000690111040144800042F5C403",
INIT_04 => X"7029AF0F81A00010CCA47700CC513CAC0D0B8E02010740E19754080108988021",
INIT_05 => X"02139405007133C0712244CD20F20105D583000020E9892201D304D42A9835E1",
INIT_06 => X"9190440300078002014405D9EE814C0284A883B6D7038AE079059B7800048092",
INIT_07 => X"000100AA0004408000000004840400008D200102503000782000C00C8025C000",
INIT_08 => X"00728A00408403220811991E02120C044058080004000001101121F220000260",
INIT_09 => X"811001E1185B38AD23C3707AD46440818F3CF80EC423CA7D01D123C80200816A",
INIT_0A => X"45810810A01B40216361056D6150F41200280001900439001FD8A00041400000",
INIT_0B => X"11FC88076266E800D605402962A820211500024808010512C40106D222223B14",
INIT_0C => X"0408804116040B02C02C500B0C02C100B0C02C100B0402C300B0401618058611",
INIT_0D => X"040200050200501301208482200D00D0A0408402C4282200A84800009B878680",
INIT_0E => X"00000020000100024AC88300300060090F0D830F00025400300204D018000804",
INIT_0F => X"8000000040000206A2000800000000000000950002E010000000080000588040",
INIT_10 => X"0000000000000808000554000200000000000100006D0020000000100000BB00",
INIT_11 => X"0000400000000000002000001A0002504001000000000000002280000D800800",
INIT_12 => X"0800000000000E2C802000000000408D801000000000408012440000200110A0",
INIT_13 => X"000000000004680003A0040000000010280003800800000000102800000B0000",
INIT_14 => X"000005C0002000000000000620000158000010000000000010A0000B00000200",
INIT_15 => X"C30146200400104002602600400000000294004000000004000000000010001A",
INIT_16 => X"0080200000008020000000802000000080080000004090014134DA101288C6DB",
INIT_17 => X"0802000000000401806010040180601004018060100000802000000080200000",
INIT_18 => X"8060180601004010040080200802000000000000802008020000000000008020",
INIT_19 => X"C0A28A063807E0500014063450404882846FFE000003FFC00000010040100401",
INIT_1A => X"AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA28A28A28A28A2934C8D0CCD145144",
INIT_1B => X"68341A0D068341A0D068341A0D068341A0D068351A8D46A351A8D46A351AAAAA",
INIT_1C => X"FFFFFFFFFFFFFFFC0000000000000000000000001FE32068341A0D068341A0D0",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"408102040810207FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"800AA00000000000000000000000000000000000000000000040810204081020",
INIT_28 => X"168B55557BEAB4500554200000557FE10FFFBEAA10007FD7410FFAA97555082A",
INIT_29 => X"55574105D2A800AA00043FEBA5D7FEAA00007BE8AAAAA843DF55FFAA955EFA2D",
INIT_2A => X"57BC00AAA2FFEAAAAAA8415555087BFFF55A2AA800BAFFAE9555508002AA0000",
INIT_2B => X"A2AA955EF005568A00087BE8BFFA2D17DE1000517FE10AAAAA8AAA002E975455",
INIT_2C => X"FAA8417410A2D140000F7FBC2010A2D157400AAAE974AAAAAA974BA08002AB55",
INIT_2D => X"EFA2AABDEAA087BEAAAAA2FBD54BA080002145552ABFEAA007FC21EF007FD75F",
INIT_2E => X"00055042AB45F7FFD741000042AA10AAAABFF5508003FF55F7D568A00552EA8B",
INIT_2F => X"5400F7A49057D0824850B8000000000000000000000000000000000000000000",
INIT_30 => X"3AF55F7A0925D7AADB6FB7D5D7FEAB7808554203A145178E00FFFBE8A101475D",
INIT_31 => X"A9557D080038AAA145157428492E8008200043FE925571EFA380871C7028A28E",
INIT_32 => X"AEA8A9200249056D4175C5092AAF5FDA38BE8E1557D1475FAF45BEAA800AAFFA",
INIT_33 => X"AA4954281C0E2FB55B6A0925D7085F6AA10087FEABD7AAD57AEBA08517DE00AA",
INIT_34 => X"007FC51C7007BD55D7BE80004AAFEDB42028EBFBC2028BED152438AAA092492A",
INIT_35 => X"AF7DF6AA00412EAABFFAA803DEBA0875EDA80BEF1C743840040017D5520B8EAA",
INIT_36 => X"0000000000000000000041002FB55FFF5D0438140E2FA38B6AEBFF6DBE84AAEB",
INIT_37 => X"A00FFFFEAA105D5155410FF84021EF0800154B20000000000000000000000000",
INIT_38 => X"DEBA0851574B2AAAEAAB55F78400145AAFFFFFEF5D7FEABFF0051400A25D5568",
INIT_39 => X"68B55F7AA800BAF7AA955EF00042AAA25555410BA082E8201000043FE005D517",
INIT_3A => X"568AA200557DE00AAAAAAA000804001FF005575408AA557FEB2FFAE975EF5551",
INIT_3B => X"D1550AAAA8002010F2AC154B25F2ABFF55F7800015F087FEAA00007FEAB55FAD",
INIT_3C => X"800021EF55042AAAA007FD5555087BD6145FAAC000A2A6FBC00BAAAFBC00BAF7",
INIT_3D => X"F7AEBDFF779A82AA43F7FBE8A00082EA8BFFAA843FEBA08517DE00F3F9574B30",
INIT_3E => X"000000000000000000000000000000000000008003FF55F7D5420BA5D2ABFEAA",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_2,               -- Port A enable input
WEA      => wbe_a_hi_1024_2(0),               -- Port A write enable input
DIA(0)   => data_write_a(4),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_2(4),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_2,               -- Port B enable input
WEB      => wbe_b_hi_1024_2(0),               -- Port B write enable input
DIB(0)   => data_write_b(4),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_2(4),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_5_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50DF4A0791B3FCB694379283C81FD996A091832102004A336A20E03C040C002",
INIT_01 => X"805FBDC69830A84D5C6A60000C34C26841280A00084000C8C212892EEAD53235",
INIT_02 => X"3B2026B578918E640A4F01CF8011FF0002080000082CA9998276DF7772C7C80D",
INIT_03 => X"37134108420D700084205702A4008A1D9100002171C0E0051554D93A11F5D140",
INIT_04 => X"8A41A0FC03A56DA000425A819410E3816C086198A388B702A8CA1210844A0C4C",
INIT_05 => X"B1808A062E8BC835F5E84532D708238A282F00A9291224800A2861490343082C",
INIT_06 => X"903FB8483A90581859050424100940825C6184401CDC451B860A6507160C4100",
INIT_07 => X"D26F068BCC96CDF8918E640E96D1A3469D6300E2FFEA27F8E4D23248130E259C",
INIT_08 => X"0BFA82E568442B2A082C0A7E3014250D49DA37A2420619000002AFF48D1222E5",
INIT_09 => X"3F005001E40969289429360416DCD1C46083030604B1CA20C03DF83B0A2C60A5",
INIT_0A => X"14613C71005A10492B888120288F480D58858449026145B3830F449449062B4F",
INIT_0B => X"11AC04934AC648BFD727C031E64170A137D5AA5C3E4B0F8A3C58C34C002290E3",
INIT_0C => X"CA29C6CC50384B6AC6AC86AB31AACA6AB39AAC86AB39AACA6AB3055643559C31",
INIT_0D => X"C673E33CF28F38603855401985228A0614BD30A0A2819852011E5AC2B87F9182",
INIT_0E => X"FF87C002F87A803E460B2516510CA594FF0044FFA4B08BAC4BB2CD0F09CF84E3",
INIT_0F => X"0DFF0F8005F0F5100DFFF5E15D06101C55EB29F1E00BE53FE1F000BE1E802F94",
INIT_10 => X"F12F0380231F17D78FC029FFF58D9A70380230F2FE0017C37FC3E0017C3D005F",
INIT_11 => X"FC7F023C0CA700125C0F8F7E43F1F001BFFE7C69E01804E1E7CCF8FC003FF5F1",
INIT_12 => X"023E00017C1FC1A4BFD82C3081C5BD27BFE30C3081C5BD00C02365D645CEEF5B",
INIT_13 => X"61E0042787F181E9C1EFD8CB8120C5AF41E9C18FD60F0C20666F41E9F009FFFD",
INIT_14 => X"7A7C077FFF404F80005F07F187A7D14BFFC96111C048278DEB074F9930FF9D80",
INIT_15 => X"C064014B8B652E2B3120C81284641D3E8DBF7D636FE860190700132C1F0EFB80",
INIT_16 => X"38CE1384E3384E338CE138CE1384E33C4E3ECE32E128882551349A1CBAA44103",
INIT_17 => X"84E3384E3384E3384E338CE138CE1384E3384E338CE138CE1384E3384E338CE1",
INIT_18 => X"CE138CE138CE138CE1384E3384E3384E3384E338CE138CE138CE138CE1384E33",
INIT_19 => X"F5E5BB4E7F7B9DB7FF3A1B6DB7E8410A8C000000000000000000384E3384E338",
INIT_1A => X"BEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEF9F7CFDFDDCF3CF3D",
INIT_1B => X"BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEFBEF",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000001711C7BBDDEEF77BBDDEEF77",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"FDFFF00000000000000000000000000000000000000000000080000000000000",
INIT_28 => X"FD7410FFAA97410082A800AAAAAE955450055421FFFFFBC0010AAD5574BA557F",
INIT_29 => X"7FD74000055574BA5D7FD7555A2D5575EF55517FF5500557FE10FFFBEAA10007",
INIT_2A => X"0002AABA5D2ABFFFFAA843DF55FFAA955EFA2D168B55557BEAB5500554200000",
INIT_2B => X"5D2A800AA00043FEBA5D7FEAA00007BC00AAAAAEBDF45A28428B45FFD168BFF0",
INIT_2C => X"5080028A00A2FFFDE00F7D57FEBAFF80174BAAAD1555EF555555555005557410",
INIT_2D => X"BA5D2E821FFA2D5554BA557BD75FFAA8415555087BFFF55A2AA800BAFFAE9555",
INIT_2E => X"00000517FE10AAAAA8AAA002E97545557BC00AAA2FFEAAAA082A97545F7D5420",
INIT_2F => X"7010BEDF524AA5571FDFEF000000000000000000000000000000000000000000",
INIT_30 => X"78E00EBFBE8A101475D5400F7A49043D0824850B8A2AE9756D145B401FFFFFFC",
INIT_31 => X"FEAB7D0855420BA1471D74380851524BA5571D757DB6D5525EF555178F6D1451",
INIT_32 => X"8A28B6DEBDF6DBEF1C0A28AAA5524BFFFFA28E3AF55F7A0925D7AADB6FB7D5D7",
INIT_33 => X"5555057D145152428492E8008200043FE925571EFA380871C7028B6AEBDF45B6",
INIT_34 => X"BEAA800AAFFAA9557D080038AAAA2FBF8E10EBD578EAAFF8415482BED1555EF5",
INIT_35 => X"81C209256DFFDF420BA552A821FFB6DF574A85575C55EFBE8E1557D1475FAF45",
INIT_36 => X"0000000000000000000008517DE00AAAEA8A9200249056D4175C50920875FDA3",
INIT_37 => X"5FF5D7BC21EFF7FBD7400F7FBC00BA55557DFF70000000000000000000000000",
INIT_38 => X"01FF5D5568BE7555568A00AAFFEAA105D5155410FF84020AA0800154B2AAAA97",
INIT_39 => X"00145AAFFFFFEF5D7FEABFF0051400A25551554BA0051400BA5551575EFF7D14",
INIT_3A => X"1574B2FFAABFF45FFAAAABFFAAFFFDFFF552EA8AAA55043DFF7AAAEAAB55F784",
INIT_3B => X"8002410FFD5575EF5555421E75555400BA082E8201000043FE005D517DEBA085",
INIT_3C => X"FAE975EF555168B55F7AA800BAF7AA955EF00002AAA2A2FBE8A00A2D16AAAAFF",
INIT_3D => X"0055554088A557FEB25D00021FFFFFFC00BA552A821EFFFFFD74BA5D51575F7F",
INIT_3E => X"000000000000000000000000000000000000000557DE00AAAAAAA000804001FF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_2,               -- Port A enable input
WEA      => wbe_a_hi_1024_2(0),               -- Port A write enable input
DIA(0)   => data_write_a(5),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_2(5),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_2,               -- Port B enable input
WEB      => wbe_b_hi_1024_2(0),               -- Port B write enable input
DIB(0)   => data_write_b(5),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_2(5),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_6_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10800B0061A01002840002C03002818000402322520070B313301C4389B2082",
INIT_01 => X"250041CA3839684D18A160000C52426841000000090800090210080008110200",
INIT_02 => X"0020042080010000044654C0000C008010000000001020900200200002620814",
INIT_03 => X"060881021088200021080200E4000A0891000020610111500104C00000F14400",
INIT_04 => X"0880000100000002000052288144004281C050400100280000C8100000080001",
INIT_05 => X"928080840001100A08009000280201000850E022401400002028214043410820",
INIT_06 => X"10100518090012122100C808049310002040000410A0001400000200120840D2",
INIT_07 => X"000100800004400001000000860408108C22000A502010074120044800040001",
INIT_08 => X"50000040D0C4E2088003FD01C01004044058082004000000000121F020408244",
INIT_09 => X"00BF17E9001205A5204911F814444080400100020000D200DFD16400C2A40AA0",
INIT_0A => X"04611C17849000022862A1596C8B5DF04834948900000100220C244840000880",
INIT_0B => X"03AD0413424E4044D665C070C22602291504400D084915020448114080201000",
INIT_0C => X"5E08864011088B22D22C008B0022C408B1022C208B0822C608B1111600458010",
INIT_0D => X"4251A12CD28A300429688001000800000020280204001000A00804309A002182",
INIT_0E => X"0000000280402400420800000000006200FC10002442042429324294014E8CA7",
INIT_0F => X"A40000000500800840000800000000000002280018001480000000A010100052",
INIT_10 => X"00000000000004C2003000010240000000000000680800290000000140202000",
INIT_11 => X"2000C0000000000000000442000001080001000000000000010C000280001804",
INIT_12 => X"08000000000801C300A010000000156000902000000015101200002800000000",
INIT_13 => X"000000000101800038002408000000094000386028040000000940000ED40000",
INIT_14 => X"0003B000002000000000020180002A24005010000000000023000060C7000A40",
INIT_15 => X"3F0280090321000040A410C28108000160008094000810040000000000002300",
INIT_16 => X"284A5284A728CA5284A528CA728CA52C4A5A0A32A300940101349A0408240818",
INIT_17 => X"9CA1294A329CA5284A728CA7284A5284A728CA5284A528CA728CA5284A728CA7",
INIT_18 => X"CA3294A129CA3294A129CA1294A329CA1294A3294A129CA3294A129CA3294A32",
INIT_19 => X"F5F78BCE7F8FF0F4FA955F7CF7F40A80145D55555556AAAAAAAAA94A329CA129",
INIT_1A => X"8E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E39B6CEDECDDF7DF7D",
INIT_1B => X"F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE38E3",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000001A1A33F9FCFE7F3F9FCFE7F3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"555FF00000000000000000000000000000000000000000000080000000000000",
INIT_28 => X"BC0010AAD5574BA557FFDFFF087BFDF45F7AA974AAAAAA97555F784174BAF7D5",
INIT_29 => X"515555508043FE00F7AA97555A2FBD7410AA8428AAAAAAE955450055421FFFFF",
INIT_2A => X"7D1575EFFFAA9555500557FE10FFFBEAA10007FD7410FFAA97400082A800AA08",
INIT_2B => X"0055574BA5D7FD7555A2D5575EF55517FF55A2AA97400552AAAB45082E80155F",
INIT_2C => X"500554200000003DE10FFD5401FFF7AAA8A10082EAAB45A2FFC2000007FD7400",
INIT_2D => X"10AA803FE105D516AABAFF843FFFFAA843DF55FFAA955EFA2D168B55557BEAB5",
INIT_2E => X"000AAAEBDF45A28428B45FFD168BFF00002AABA5D2ABFFFF087BD5545007BFDE",
INIT_2F => X"256DEB84104BAFFD1525FF000000000000000000000000000000000000000000",
INIT_30 => X"9756D145B401FFFFFFC7010BEDF524AA5571FDFEF1C7BFFF55FFA095482B6A49",
INIT_31 => X"4904380824850381C5B5057D1C003DE28F7A49057DAAF5D2428A2842AAAAA2AE",
INIT_32 => X"2AAFB451C2A8017DE3DF525FFFFA49756D145178E00EBFBE8A101475D5400F7A",
INIT_33 => X"2F1C50381471D74380851524BA5571D757DB6D5525EF555178F6DAAA49542841",
INIT_34 => X"AADB6FB7D5D7FEAB7D0855420BA1C0E3FE00E3DB471EFE3AAAAA00082EA8B6DA",
INIT_35 => X"F1C7BD057D1C71FFE10A28038E1049516AAB8FF8428FEFA28E3AF55F7A0925D7",
INIT_36 => X"00000000000000000000B6AEBDF45B68A28B6DEBDF6DBEF1C0A28AAA5524BFFF",
INIT_37 => X"F55F78017400F780001FFAA84000AAFFD1401E70000000000000000000000000",
INIT_38 => X"20BAAA8428AA2AAAA975FF5D7BC21EFF7FBD7400F7FBC00BA55557DFF7557BFD",
INIT_39 => X"EAA105D5155410FF84020AA0800154B2557FC01EF55043FEAAFF80021EFA2D14",
INIT_3A => X"568BE7AA80174AA082ABDF555D2A821EFAAFBC01FFF780155F7555568A00AAFF",
INIT_3B => X"AEA8A10082EA8BEFAAD5554B25551554BA0051400BA5551575EFF7D1401FF5D5",
INIT_3C => X"AAEAAB55F78400145AAFFFFFEF5D7FEABFF0051400A25D2EBFE10AAFFD55EFA2",
INIT_3D => X"552EA8AAA55043DFF7557BC01EF55557DE00AA842AA0000516AABAFF8428BE7A",
INIT_3E => X"0000000000000000000000000000000000000FFAABFF45FFAAAABFFAAFFFDFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_2,               -- Port A enable input
WEA      => wbe_a_hi_1024_2(0),               -- Port A write enable input
DIA(0)   => data_write_a(6),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_2(6),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_2,               -- Port B enable input
WEB      => wbe_b_hi_1024_2(0),               -- Port B write enable input
DIB(0)   => data_write_b(6),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_2(6),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_7_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10844B00482258A2842112C02450418800002300500030B313300C418992002",
INIT_01 => X"000009CA3839684D1CA0E0000E51424840000000080000080200080008510204",
INIT_02 => X"0120042086010000044600C00008000004100000000260900200000002402004",
INIT_03 => X"8628A10000082400000002408400080011000000610008000208C00000E14400",
INIT_04 => X"0911800100A000000000524084000040000050001140200100C8100000080102",
INIT_05 => X"0300812401011000000000002000114008008060441000000020024093000000",
INIT_06 => X"9190431C0D4010100000880804010010800000041080081000000200010424B2",
INIT_07 => X"000100AA0004408601000004860000008C02000A103010006928040800062481",
INIT_08 => X"84000048D484C20888000A0002120484C048007004000000000021F000000244",
INIT_09 => X"00A06009881201A520491004106C48A04040002400A15A208001650004001020",
INIT_0A => X"C99E1060201002044809C1040140A001004808810000459033189C0A400118A0",
INIT_0B => X"102000024040484050050041648A0041140C500B08821054C000264120000400",
INIT_0C => X"0404A083260E0832132011880462011880462051881462051881D31018C40620",
INIT_0D => X"0001000080001000813094801A8F80F00A600B52602801A88848011118003700",
INIT_0E => X"000003C007C002808228010410082042C000C000000004001002000400040002",
INIT_0F => X"A4000007800F80C840000800009864038A1200081C0014800000F001F0200052",
INIT_10 => X"00002C0E00E0E4004038000102400002C0E00E0D20100029000001E003E04000",
INIT_11 => X"2000C04031100E0403D0700300080908000100000661801E1900040380001804",
INIT_12 => X"0840878083E8003780A01043203A101780902043203A10082410082880000000",
INIT_13 => X"0601E0187900181035E0240806483248181035E0280410C8198818100DDD0000",
INIT_14 => X"0403774000201021E020FA006040376C00501022131210722060806D47000A40",
INIT_15 => X"00928A0002000110888600C032128201519480D40009902430160403E0E00506",
INIT_16 => X"01000000020080601802000000000405000A0020020081014134928820480010",
INIT_17 => X"0802018040000000006018020080200804010000000000806018020080000004",
INIT_18 => X"0000000001806008020000001006008020080001004008020080201004000020",
INIT_19 => X"0000000000000000000000000000400A004618618618C30C30C3000020180600",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000000B0840000000000000000000",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"1555500000000000000000000000000000000000000000000080000000000000",
INIT_28 => X"A97555F784174BAF7D5555FFF780155EFAAAEA8ABAAAFBFDE0055556AA005D04",
INIT_29 => X"55555EFAAFFFDFEFAAAAAAB455D556AA00FFAE95555087BFDF45F7AA974AAAAA",
INIT_2A => X"02EAAAAA082EA8A00AAAE955450055421FFFFFBC0010AAD5574BA557FFDFFF55",
INIT_2B => X"08043FE00F7AA97555A2FBD7410AA8428AAA557BFDFFF55003DFFFF7FBEAA000",
INIT_2C => X"0082A800AAF7AE975FFA28000010552EBDE00007BEAAAAA2D140000085155555",
INIT_2D => X"45087FEAB455D516AB55557BD55FF00557FE10FFFBEAA10007FD7410FFAA9740",
INIT_2E => X"000A2AA97400552AAAB45082E80155F7D1575EFFFAA955555D51574AAAAFFD55",
INIT_2F => X"AE105D556AA10410E17555000000000000000000000000000000000000000000",
INIT_30 => X"FFF55FFA095482B6A49256DEB84104BAFFD1525FFFF8E175C7A2AAAAA82A2F1F",
INIT_31 => X"F524AA5571FDFEF415B575D7AAF1FFFD7AAAAAFB7D495F6AA10E3AE905551C7B",
INIT_32 => X"003AFEFEBFBEAA001C2EA8A821C2EAAA00A2AE9756D145B401FFFFFFC7010BED",
INIT_33 => X"EDB470101C5B5057D1C003DE28F7A49057DAAF5D2428A2842AAAA497BFAFFF49",
INIT_34 => X"1475D5400F7A490438082485038F7A4905C7A28A070384120BDE100075EAA82B",
INIT_35 => X"D495150492BEF1D2555087BE8B7D555F6AB57417BC05D7145178E00EBFBE8A10",
INIT_36 => X"00000000000000000000AAA495428412AAFB451C2A8017DE3DF525FFFFA49756",
INIT_37 => X"555A2AEA8A10AAD568A00555168A10002E9754D0000000000000000000000000",
INIT_38 => X"8A10AAAE8215D557BFDF55F78017400F780001FFAA84000AAFFD1401E7FFAA97",
INIT_39 => X"C21EFF7FBD7400F7FBC00BA55557DFF7007BD5555AAD57DF55AAAEBDFEF007BE",
INIT_3A => X"428AA2007FE8BFF080028BFFAAFFEAA105D2EAAA005D2AAAA18AAAA975FF5D7B",
INIT_3B => X"043DE0000516AA10F7FBD7408557FC01EF55043FEAAFF80021EFA2D1420BAAA8",
INIT_3C => X"55568A00AAFFEAA105D5155410FF84020AA0800154B2FF8402145A2AA954AA00",
INIT_3D => X"AAFBC01FFF780155F7005140000FFD140145007FE8BEF557BEAB55087FC215D5",
INIT_3E => X"0000000000000000000000000000000000000AA80174AA082ABDF555D2A821EF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_2,               -- Port A enable input
WEA      => wbe_a_hi_1024_2(0),               -- Port A write enable input
DIA(0)   => data_write_a(7),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_2(7),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_2,               -- Port B enable input
WEB      => wbe_b_hi_1024_2(0),               -- Port B write enable input
DIB(0)   => data_write_b(7),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_2(7),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_8_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00000648E2840112C00000418000002700500030B3132000400812082",
INIT_01 => X"100008480009004C04A100000252024840000000180800080200010040110204",
INIT_02 => X"0020042000490000004600804008000005100000000024900200000002400004",
INIT_03 => X"0A0C33400008082400000080A4004B0891000020610112000040C00000E5C000",
INIT_04 => X"18800001000000000000512080000040800150400824280110C8100000120200",
INIT_05 => X"908084A10100100200004080280008240810802206940000012C214451610800",
INIT_06 => X"81B000080860109021400008040000202048020414A0021400040200322824C1",
INIT_07 => X"000000080004408049000004860000008402001A50208000630C040800062483",
INIT_08 => X"440000428644212280800A00021004044048002124000000000021F000000244",
INIT_09 => X"00004009001001010008100414644410400102228000D20080114502006409A2",
INIT_0A => X"000051312000042200294429148A4801C80C8C81000045907118040340020832",
INIT_0B => X"4020000240404140004D0544C4AA0001150410090302500011C813428A000400",
INIT_0C => X"46501090008820240240409000240009000240009000240009000120204808A5",
INIT_0D => X"42D1A168D09A301468402480004780F00140080860280004085904309A002196",
INIT_0E => X"00783FC00044340242280000000000020000C0000442106419120004034685A3",
INIT_0F => X"8000F07F800088A80000081EA2F9EC0000064004081010001E0FF00011104040",
INIT_10 => X"0ED0FC7E00000422201080000202658FC7E0000021882020003C1FE000222080",
INIT_11 => X"018059C3F350FE0C00000002A0040500000103961FE780000110010090000800",
INIT_12 => X"FD41FF80000830200021C1CF600012200010D1CF600012121600100810000004",
INIT_13 => X"9E1FE000010A1802100004343ED8000898021000087073D80008980200800002",
INIT_14 => X"0080200000BEB07FE00002086008020000209AEE3F300000246020200000620B",
INIT_15 => X"0088881903210000440610C8000A808040000208901786E4F0FE0C0000000166",
INIT_16 => X"685A1685A769DA368DA368DA769DA36CDA121A11A141800011309284002C0810",
INIT_17 => X"95A5685A1685A5695A368DA368DA769DA368DA368DA7695A1685A1685A5695A1",
INIT_18 => X"5A1695A568DA368DA369DA768DA1685A1695A5685A168DA369DA768DA368DA16",
INIT_19 => X"A4028A0A543EBC57A10A1E75D64108080468618618630C30C30C69DA5685A168",
INIT_1A => X"9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7BF3CCD8DF5B2DB2C",
INIT_1B => X"F87D3E1F4F87D3E1F4F87D3E1F4F87D3E1F4F87C3E1F0F87C3E1F0F87C3E79E7",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000006A6D4F87D3E1F4F87D3E1F4",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"155FF00000000000000000000000000000000000000000000080000000000000",
INIT_28 => X"BFDE0055556AA005D0415555080000000087BEAA10F7803DE00FFAEBFFFF0800",
INIT_29 => X"2AA8AAA557FC0010F780154105D7FC2145005155555F780155EFAAAEA8ABAAAF",
INIT_2A => X"7FFFFF55AA80155FF087BFDF45F7AA974AAAAAA97555F784174BAF7D5555FF55",
INIT_2B => X"AAFFFDFEFAAAAAAB455D556AA00FFAE95555AAFFE8A00552EBFE00F7D17FF45F",
INIT_2C => X"A557FFDFFF5504000AAAAAAA8B55F7D140010552E821EFAAAABDF555555555EF",
INIT_2D => X"55AA8028A00A2D57FF45557BE8A00AAAE955450055421FFFFFBC0010AAD5574B",
INIT_2E => X"000557BFDFFF55003DFFFF7FBEAA00002EAAAAA082EA8A00002AA8A10F784021",
INIT_2F => X"FE10F7AEBAFFF080A175D7000000000000000000000000000000000000000000",
INIT_30 => X"175C7A2AAAAA82A2F1FAE105D556AA10410E17555080E000280071E8A00EB8E3",
INIT_31 => X"4104BAFFD1525FF492EA8AAA5571C2000FF8A17400557FC015514555757DFF8E",
INIT_32 => X"2ABDE10EBDF7AF6DE3FFF8F7DB68A105D71C7BFFF55FFA095482B6A49256DEB8",
INIT_33 => X"AA0BDF6D415B575D7AAF1FFFD7AAAAAFB7D495F6AA10E3AE90555A2FBE8A3849",
INIT_34 => X"FFFFC7010BEDF524AA5571FDFEF550E00082B6A0AFB55F7D1420104124821D7A",
INIT_35 => X"01C2EA8A00F7800017DA2842FA00B6D578F6D557FFDA00A2AE9756D145B401FF",
INIT_36 => X"00000000000000000000497BFAFFF49003AFEFEBFBEAA001C2EA8A821C2EAAA0",
INIT_37 => X"0BA08556AA00AAAABFE00F7AEAABEF082E955450000000000000000000000000",
INIT_38 => X"21555D51575EFFFAA97555A2AEA8A10AAD568A00555168A10002E9754D082E82",
INIT_39 => X"17400F780001FFAA84000AAFFD1401E7082EAAABA5D5140010F7AE974105D7BC",
INIT_3A => X"E8215DA2FFE8ABA082ABFE00AAFBEABFFAAFBEABFFF7AA80145557BFDF55F780",
INIT_3B => X"D540000000402145AA843FFFF007BD5555AAD57DF55AAAEBDFEF007BE8A10AAA",
INIT_3C => X"AAA975FF5D7BC21EFF7FBD7400F7FBC00BA55557DFF75D2E82010F7843DF45FF",
INIT_3D => X"5D2EAAA005D2AAAA185D2AAAA10F780021FFA2803DE10FFD16ABFF5D7BFDE10A",
INIT_3E => X"0000000000000000000000000000000000000007FE8BFF080028BFFAAFFEAA10",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_2,               -- Port A enable input
WEA      => wbe_a_hi_1024_2(1),               -- Port A write enable input
DIA(0)   => data_write_a(8),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_2(8),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_2,               -- Port B enable input
WEB      => wbe_b_hi_1024_2(1),               -- Port B write enable input
DIB(0)   => data_write_b(8),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_2(8),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_9_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00018248A2840112C00002C18000002300500030B3132000400812006",
INIT_01 => X"400008000000004C0020000000100248413C0A61590001D90213C10008110204",
INIT_02 => X"01A0042080010000054600C04008000004100000001020900200200002420804",
INIT_03 => X"024003400008012400000010E4004B0891000020610310000144C00000F5C000",
INIT_04 => X"1801800100E000000000510084000040010050020810200000C8900000320200",
INIT_05 => X"918004311104100000000000200008100800002000100000002C234415610820",
INIT_06 => X"81B00008080010100000980804000008800042041080001000100200322C2481",
INIT_07 => X"0000811800044080010000058600000086020002502080006000040800062C80",
INIT_08 => X"0000004001D4618008800A00061004044048002004000000000061F000000244",
INIT_09 => X"000040090802009420409004104444084001022400214A2080014400026401A2",
INIT_0A => X"04000071200000A003CA294140200800C80C8C8100004590111C040040120800",
INIT_0B => X"12210002404848502847040164880021150400080222000200C8034200000000",
INIT_0C => X"4610088010080421021040841021000841021000841021000841010800420820",
INIT_0D => X"42D0A16C529A321068500484000500D10042080040284000084900001A002196",
INIT_0E => X"00000002804000004228010410082002C000C0002400046419120410034285A1",
INIT_0F => X"A00000000500800800000800000000000002290008001080000000A010100042",
INIT_10 => X"00000000000004C2001000000240000000000000680800280000000140202000",
INIT_11 => X"0000C0000000000000000442020001000001000000000000010C800080000804",
INIT_12 => X"08000000000801A7802010000000152780102000000015000600000800000000",
INIT_13 => X"000000000101900011E0240000000009500011E0280000000009500004DD0000",
INIT_14 => X"000137400020000000000201C000136C00101000000000002340002947000240",
INIT_15 => X"0080881901210000000600C280028000419480D4000010040000000000002304",
INIT_16 => X"68DA368DA1685A1685A1685A1685A16C5A121A13A141950051309284A82C0010",
INIT_17 => X"85A1685A1685A1685A368DA368DA368DA368DA368DA368DA368DA368DA368DA3",
INIT_18 => X"5A1685A168DA368DA368DA368DA368DA368DA368DA3685A1685A1685A1685A16",
INIT_19 => X"0157344CCCF48DE68A895C38E2540A8010100000000000000000685A1685A168",
INIT_1A => X"14514514514514514514514514514514514D34D34D34D34D28E1004039248209",
INIT_1B => X"D268341A4D268341A0D069349A0D069349A0D068341A0D068341A0D068345145",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000014D490D069349A0D068341A4",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"EAABA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"03DE00FFAEBFFFF0800155FFAAFBE8B45002A974AAAA803DFFFAA843DF45FFFF",
INIT_29 => X"7BFDE00A2FBD7400F7FBFDFFFA2AEBDE00AAFBEAABA080000000087BEAA10F78",
INIT_2A => X"055401FFF7AEAAA10F780155EFAAAEA8ABAAAFBFDE0055556AA005D041555508",
INIT_2B => X"557FC0010F780154105D7FC2145005155555557BE8BEF007FFDEAAAAD1555EF0",
INIT_2C => X"AF7D5555FFF780154AA5D2AA8A10F7AA974AA082E80010A2AAAAA10552AA8AAA",
INIT_2D => X"BAF7D17FEBAA2AEBDF45002EAAABA087BFDF45F7AA974AAAAAA97555F784174B",
INIT_2E => X"000AAFFE8A00552EBFE00F7D17FF45F7FFFFF55AA80155FF080400145FFFBEAA",
INIT_2F => X"8FC7BE8A3DF7DF7F5E8A92000000000000000000000000000000000000000000",
INIT_30 => X"000280071E8A00EB8E3FE10F7AEBAFFF080A175D7BEF1E8B6D002090482B68E3",
INIT_31 => X"56AA10410E175550871FFE00A2FBD0400FFF5FDFC7B6A0BDE38B6F5E8A92080E",
INIT_32 => X"7BFAE82A2DB555C71C5B451D7FFAAA8A38FF8E175C7A2AAAAA82A2F1FAE105D5",
INIT_33 => X"2AEADA38492EA8AAA5571C2000FF8A17400557FC015514555757D5D71E8BEF14",
INIT_34 => X"B6A49256DEB84104BAFFD1525FFFF84174BA5D20AAA00E3AA904BA142A87010A",
INIT_35 => X"7000400155FFFBEDA82FFD57DEBAAAA0BFF7D0024ADA921C7BFFF55FFA095482",
INIT_36 => X"00000000000000000000A2FBE8A38492ABDE10EBDF7AF6DE3FFF8F7DB68A105D",
INIT_37 => X"BEF080402000F7AAA8B55FFAABDFEFF7D16AA000000000000000000000000000",
INIT_38 => X"FEAAFFD16AA00082E820BA08556AA00AAAABFE00F7AEAABEF082E95545F7D568",
INIT_39 => X"A8A10AAD568A00555168A10002E9754D00517DE00A2FFC2000F7D17FF55FF803",
INIT_3A => X"1575EF555568BEF5D7FE8A10AAFFD55555D7FD5555FFAAA8AAAFFAA97555A2AE",
INIT_3B => X"AE800AA552A97400A2AEBDEAA082EAAABA5D5140010F7AE974105D7BC21555D5",
INIT_3C => X"57BFDF55F78017400F780001FFAA84000AAFFD1401E7FF80174AA5D0028A00AA",
INIT_3D => X"AAFBEABFFF7AA80145080002145F7FBFFE00FFD17FEAAA2803DFEF08043FE005",
INIT_3E => X"0000000000000000000000000000000000000A2FFE8ABA082ABFE00AAFBEABFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_2,               -- Port A enable input
WEA      => wbe_a_hi_1024_2(1),               -- Port A write enable input
DIA(0)   => data_write_a(9),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_2(9),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_2,               -- Port B enable input
WEB      => wbe_b_hi_1024_2(1),               -- Port B write enable input
DIB(0)   => data_write_b(9),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_2(9),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_10_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00018248A2840112C00002C18000202300500030B3132000400992006",
INIT_01 => X"254008000000004C002000000010026840000000080000080200010008110204",
INIT_02 => X"0020042000010000004455800008000004100000000000900200000002400004",
INIT_03 => X"020001021089000021081000C400090011000000610001540104C00000F14400",
INIT_04 => X"0811800101A00002000050088554004200C840000000200080C8100000000001",
INIT_05 => X"030080001000100800009400200000000840E020201000000024024001200020",
INIT_06 => X"81B00008080012120004CC080492500280208004148000100000020020042493",
INIT_07 => X"0000000800044080010000048404081085020002502000006000040800062480",
INIT_08 => X"100202400084410808000A00021004044048000004000000000021F020408264",
INIT_09 => X"010040090002008420401004144440004040022484214A2080110108C2C00320",
INIT_0A => X"04004166A48A0001080000000000080080181881000045901118044040020800",
INIT_0B => X"1201000200484910000F0105602622291404020902005002018002400A022000",
INIT_0C => X"0440001011808020120004801120044800120004801120044800110002400884",
INIT_0D => X"008000440210100041308480800F82F00040180260A808008848000018002104",
INIT_0E => X"000000028040000002280104100820020000400020000440100204100A000100",
INIT_0F => X"040000000500800800000000000000000002280008000400000000A010100010",
INIT_10 => X"00000000000004C2001000010000000000000000680800010000000140202000",
INIT_11 => X"200000000000000000000442000001000000000000000000010C000080001000",
INIT_12 => X"00000000000801C0008000000000154000800000000015000410000800000000",
INIT_13 => X"0000000001019800180000080000000958001800000400000009580002800000",
INIT_14 => X"0000A0000000000000000201E0000A0000400000000000002360002080000800",
INIT_15 => X"0080881000000000000600C28102800060000000000800000000000000002306",
INIT_16 => X"401004010040100401004010040100441020D0030008840051309A90BA884010",
INIT_17 => X"0902409024090240900401004010040100401004010040100401004010040100",
INIT_18 => X"1004010040902409024090240902409024090240902409024090240902409024",
INIT_19 => X"F546890A940FE0D3971243555205428290100000000000000000401004010040",
INIT_1A => X"8A28A28A28A28A28A28A28A28A28A28A28A28A28A28A28A29554199854514514",
INIT_1B => X"2B95CAE532994CA6532995CAE572B94CA6532994CA6532994CA6532994CA28A2",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000002718E72B94CA6532994CA657",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"FDE1000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"03DFFFAA843DF45FFFFEAABA007FC2155F7D155545AA80001EFAAFBEAB45557F",
INIT_29 => X"042AB55FFD168B55AA8000010FFFBE8BFFF78402155AAFBE8B45002A974AAAA8",
INIT_2A => X"AD16AABA002ABDE10080000000087BEAA10F7803DE00FFAEBFFFF0800155FF00",
INIT_2B => X"A2FBD7400F7FBFDFFFA2AEBDE00AAFBEAABAA2FFD741055003DFEFF7AA801FFA",
INIT_2C => X"05D0415555007FD74105555555EFF7FBC0145F78028A00A2D142155087BFDE00",
INIT_2D => X"55AAD168ABA002A975FFF7AEBDEBAF780155EFAAAEA8ABAAAFBFDE0055556AA0",
INIT_2E => X"000557BE8BEF007FFDEAAAAD1555EF0055401FFF7AEAAA105D042ABFF5D556AB",
INIT_2F => X"71D7AAFBEFB455D71F8E00000000000000000000000000000000000000000000",
INIT_30 => X"E8B6D002090482B68E38FC7BE8A3DF7DF7F5E8A92007BC217DEBDB55555AA8E0",
INIT_31 => X"EBAFFF080A175D700042AB7DEBDB6DB55BE8E05000EBFFE8BC7E38E07145BEF1",
INIT_32 => X"0A3DFD7F7A4821D7A2D16FA82142EB8E00080E000280071E8A00EB8E3FE10F7A",
INIT_33 => X"ED1421450871FFE00A2FBD0400FFF5FDFC7B6A0BDE38B6F5E8A92B6FBD541049",
INIT_34 => X"A2F1FAE105D556AA10410E175550071D54104951555D7EBF5C5155E3842AA00B",
INIT_35 => X"8410E2ABD749516FB55BED16FA820820955EFE3AEBDEAAFF8E175C7A2AAAAA82",
INIT_36 => X"000000000000000000005D71E8BEF147BFAE82A2DB555C71C5B451D7FFAAA8A3",
INIT_37 => X"1EFA2FFD7545AAAE97555A2FBFDF455D556AA000000000000000000000000000",
INIT_38 => X"8B45AAAA95545F7D568BEF080402000F7AAA8B55FFAABDFEFF7D16AA00087FC0",
INIT_39 => X"6AA00AAAABFE00F7AEAABEF082E9554500042ABFFA2FFFFF45F7AE97400AAFFE",
INIT_3A => X"16AA00FFFBD5400082EBFF45F78400155A2D57FE00552EA8A00082E820BA0855",
INIT_3B => X"D557555A2802AA10FFD54214500517DE00A2FFC2000F7D17FF55FF803FEAAFFD",
INIT_3C => X"FAA97555A2AEA8A10AAD568A00555168A10002E9754D085155410085557555AA",
INIT_3D => X"5D7FD5555FFAAA8AAA002AAAB4508557DF55F7D17FE000804155FFAAAABDEAAF",
INIT_3E => X"0000000000000000000000000000000000000555568BEF5D7FE8A10AAFFD5555",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_2,               -- Port A enable input
WEA      => wbe_a_hi_1024_2(1),               -- Port A write enable input
DIA(0)   => data_write_a(10),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_2(10),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_2,               -- Port B enable input
WEB      => wbe_b_hi_1024_2(1),               -- Port B write enable input
DIB(0)   => data_write_b(10),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_2(10),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_11_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"A101C4B05A0034CA2840712C2D001419000002300500030B31B20084EC992002",
INIT_01 => X"90000986B83028491800E0000C26426040000000080000088200080802512224",
INIT_02 => X"1A2004205E010640024D00800008000004100000040EC090820018003241A00C",
INIT_03 => X"28639100000C5C00000045C08400C8001100000061806A001618C03001E54400",
INIT_04 => X"1A800001000009A0804059A190000040400040008058220008C8100000120D4E",
INIT_05 => X"02000E81080250010000002022000058080400000E1200000020004401000004",
INIT_06 => X"819435143F20101010001008040800B8100102041088011100022200000024B2",
INIT_07 => X"90640D280884453E01064002944180008402001295BA100022E4340800062D82",
INIT_08 => X"400000093204802200280A0012160585C1D808D004000000000323F40C102244",
INIT_09 => X"380040098010001100009204107C5950400000220080C200800900020C006827",
INIT_0A => X"80007100004016EA080801010000080D00200081000045B0511D289940103399",
INIT_0B => X"002000024040410A000D0104408810C115D9C008050042400100D04E88000002",
INIT_0C => X"00655010009264201200C7B421ED0C7B421ED0C7B431ED087B43176843DA1085",
INIT_0D => X"0401020080400A10012494881A4F80F209500BB2602881A488485C1318002000",
INIT_0E => X"6619A540124814800228010410082022C00040002020090020220C9600040802",
INIT_0F => X"ACCC334A802491600C587949B6D0141B4CC600D5761B1599865A500490B86A56",
INIT_10 => X"BAC845542056A61686EC81E3A6CB68AA2C622C9A251C352B330CB4A0092170D8",
INIT_11 => X"BCCAD0B5A81536080CC6B21A21B1FC09CB0F1076D4A200B2AD4068F4101639B5",
INIT_12 => X"4D2CC281E31AA0103AB8D5514066380804B268A2E060901204112566F10AC418",
INIT_13 => X"D551443C47281002540B2C9AAAA8662A1152B202AE3554403028115AA88201A1",
INIT_14 => X"548A20A0492A2724A0621620402A020141F172FB182A32AB6845AB6200251BC9",
INIT_15 => X"00C00A000200074044E6801832728080D00A380B753952C4877E0104DDE4D124",
INIT_16 => X"0080200802008020080200802008020480080022020081010124988800400010",
INIT_17 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_18 => X"0000000000802008020080200802008020080200802008020080200802008020",
INIT_19 => X"55062608804180C0B10A42104201400204000000000000000000000000000000",
INIT_1A => X"00000000000000000000000000000000000820820820820801C4149470000000",
INIT_1B => X"0000000000000000040200000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000007E0F0000000000000100800",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"000AA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0001EFAAFBEAB45557FFDE10082ABDF5508557DF45002ABDFFFF7803DE10AA80",
INIT_29 => X"AEBFF45FFAEBFEAA002A801FFF7FFE8A10A28000000007FC2155F7D155545AA8",
INIT_2A => X"2AABFE10082ABFFEFAAFBE8B45002A974AAAA803DFFFAA843DF45FFFFEAABAA2",
INIT_2B => X"FFD168B55AA8000010FFFBE8BFFF78402155AAD155555A28428BFF002ABDE00A",
INIT_2C => X"F0800155FF00557FF45557FC2010002A80010A2842AAAA007BFFF4500042AB55",
INIT_2D => X"FF5D00154BAF7FBE8BEFFFD540000080000000087BEAA10F7803DE00FFAEBFFF",
INIT_2E => X"000A2FFD741055003DFEFF7AA801FFAAD16AABA002ABDE10A2D168A10A284021",
INIT_2F => X"DFC7F78E3FE28B684070AA000000000000000000000000000000000000000000",
INIT_30 => X"C217DEBDB55555AA8E071D7AAFBEFB455D71F8E00002EBDF6D005B78F7D142AB",
INIT_31 => X"A3DF7DF7F5E8A92BEAEBFF7DEBA0BDEAA1C2A801C7E3FFEFA10B68407038007B",
INIT_32 => X"8A28BFF082ABAE10B6AAB8E280820B8FEFBEF1E8B6D002090482B68E38FC7BE8",
INIT_33 => X"07FF8F7D00042AB7DEBDB6DB55BE8E05000EBFFE8BC7E38E07145B6D15756DA2",
INIT_34 => X"EB8E3FE10F7AEBAFFF080A175D708517DF7D497BC5028142A87000A28A2AA920",
INIT_35 => X"0B6DB6AA28A280001FF5D0A10482FFFFEFBC7E3DF42028080E000280071E8A00",
INIT_36 => X"00000000000000000000B6FBD5410490A3DFD7F7A4821D7A2D16FA82142EB8E0",
INIT_37 => X"FEF007BE8BFF5D2ABDF55F7AABDEAAF784154BA0000000000000000000000000",
INIT_38 => X"DE00FF84154BA087FC01EFA2FFD7545AAAE97555A2FBFDF455D556AA00082EBF",
INIT_39 => X"02000F7AAA8B55FFAABDFEFF7D16AA00FFAEBFFEFAA803DEBA5D2E82155A2FBF",
INIT_3A => X"A95545F7D5555FFAAAAA8BFF002AAAA00FFAAA8AAA080028BFFF7D568BEF0804",
INIT_3B => X"2E95400A2AEA8A00007FEABFF00042ABFFA2FFFFF45F7AE97400AAFFE8B45AAA",
INIT_3C => X"82E820BA08556AA00AAAABFE00F7AEAABEF082E9554508557DFFF007BD54BA5D",
INIT_3D => X"A2D57FE00552EA8A00FFFFE8AAAAA80001FF5D2E82000F7FFFFF45AAFFC20BA0",
INIT_3E => X"0000000000000000000000000000000000000FFFBD5400082EBFF45F78400155",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_2,               -- Port A enable input
WEA      => wbe_a_hi_1024_2(1),               -- Port A write enable input
DIA(0)   => data_write_a(11),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_2(11),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_2,               -- Port B enable input
WEB      => wbe_b_hi_1024_2(1),               -- Port B write enable input
DIB(0)   => data_write_b(11),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_2(11),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_12_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50080B01BC002006940202C0DE041196A83183000000023322287E0FC000006",
INIT_01 => X"75400D849830C84C5823E0000C17424840000000080000088200002802153231",
INIT_02 => X"18A026B43ED180040147558040090000061800000C06ED9802768F4472C52005",
INIT_03 => X"2A67E34A528D0524A52850528400C8001100000171C02B550618C91A10E55440",
INIT_04 => X"1BC0000100056C8280825DE98154004300C840800850240080CA921084520A07",
INIT_05 => X"02000F832000500C0000941024000852084060202E100001002000448100000C",
INIT_06 => X"819A1D1C3FE01A1A40045408049A50BA4020C6041090001200006200000000F2",
INIT_07 => X"C26A0719CC96CC6ED18A64019695A854870300FA3968B20068FC06080106249F",
INIT_08 => X"D002024B3E040800008C0A002610240D494A06F3460409000000E3F0AD5282E5",
INIT_09 => X"27A06009200040000400120412445D78400001000410420080218029CC807A27",
INIT_0A => X"18000006848A026F000000000000080000F010C100204593F11A6CDF48003BF8",
INIT_0B => X"000000820040402B28050400400432C9349DF21A31A00ACC0000F04F80020001",
INIT_0C => X"00357804611AE45D05D0833430CD0833420CD0C33420CD0833430668619A1000",
INIT_0D => X"0000000000000A74812DF00E87E80A079F9F90FA0280E87E800C7FF3B8002000",
INIT_0E => X"3B6B0E404D26160682082002000401EA0000C40000800A006002818808000000",
INIT_0F => X"A476D61C809A4DA84272592D6246FC1B17B541F97E1B348EDA93900B2B286C56",
INIT_10 => X"30C669E622DBC325CFD881A962454CFBE5403AB99594362B1DB52720165650D9",
INIT_11 => X"F8D2D39A3745261E4A95A110A3F855000E4B1D32BAB504BB7490FCFF912A3834",
INIT_12 => X"B90E9B018C7530200AB8F8BF41F9A22006B37DC8E1F9A21A70116D4C5080651C",
INIT_13 => X"118780319CCA08AB1001ACDF34B8F1C688AB1002AE3F7B807B6289F368828C4C",
INIT_14 => X"2AF020233376A5ECC016B1A827CDA21160F051DE610A34C50427E6E220323E4A",
INIT_15 => X"0077020000000439FDC05C5806781FAB46095A0B5199B0AC55521524F1864022",
INIT_16 => X"000000000000000000000000000000000026C000002884000130921092804010",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"8020080200000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0051B946088881360A95090CB054420290100000000000000000008020080200",
INIT_1A => X"041041041041041041041041041041041049249249249249200100002D451451",
INIT_1B => X"92C964B2592C964B2592C964B2592C964B2592C86432190C86432190C8641041",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000003800F592C964B2592C964B25",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"7DE1000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"ABDFFFF7803DE10AA80000AAAA843FE0008557DFFF0800020105D557FEAA0055",
INIT_29 => X"D5420000051555FFA2AA8200000557DFFFF7AA80000082ABDF5508557DF45002",
INIT_2A => X"82AA8AAAAAFFC00BA007FC2155F7D155545AA80001EFAAFBEAB45557FFDE10AA",
INIT_2B => X"FFAEBFEAA002A801FFF7FFE8A10A28000000A2D155410F7FFFFEBA08003FE000",
INIT_2C => X"5FFFFEAABA000028A105D2ABFE10A2AABFE1055516ABEF5D517DEAAA2AEBFF45",
INIT_2D => X"55002A820AA08557DFFFF7AA82155AAFBE8B45002A974AAAA803DFFFAA843DF4",
INIT_2E => X"000AAD155555A28428BFF002ABDE00A2AABFE10082ABFFEF0855420000004175",
INIT_2F => X"5010495B7AE921C517DE10000000000000000000000000000000000000000000",
INIT_30 => X"BDF6D005B78F7D142ABDFC7F78E3FE28B684070AABE803AE38145B78FD700000",
INIT_31 => X"BEFB455D71F8E00BED547038145B505FFB6A487000005F7AFD7F7A482038002E",
INIT_32 => X"F1FDE821C003FE001C2EAAAAAB6F5C2082007BC217DEBDB55555AA8E071D7AAF",
INIT_33 => X"D517DEAABEAEBFF7DEBA0BDEAA1C2A801C7E3FFEFA10B68407038B6D550428FF",
INIT_34 => X"B68E38FC7BE8A3DF7DF7F5E8A9200002FA285D20BDE28A2A4B8E10555B68BEF5",
INIT_35 => X"F085F47038140010555142082082005F7DFD7F7A482155BEF1E8B6D002090482",
INIT_36 => X"00000000000000000000B6D15756DA28A28BFF082ABAE10B6AAB8E280820B8FE",
INIT_37 => X"ABA5D7FEAB45080015410007FEAA0055517DE000000000000000000000000000",
INIT_38 => X"AB45F780020BA082EBFFEF007BE8BFF5D2ABDF55F7AABDEAAF784154BAF7802A",
INIT_39 => X"D7545AAAE97555A2FBFDF455D556AA00F7D1554BA5D7BC01FFFF8015410007FE",
INIT_3A => X"4154BAF7D1400BAFFD57FE005D043FE10552EAAAAAFFD140000087FC01EFA2FF",
INIT_3B => X"8428A105D7FEABEF55557DEBAFFAEBFFEFAA803DEBA5D2E82155A2FBFDE00FF8",
INIT_3C => X"7D568BEF080402000F7AAA8B55FFAABDFEFF7D16AA0008003FEBA55003DEBAA2",
INIT_3D => X"FFAAA8AAA080028BFF087BD54AA550402145550000010087FFFF45F78402145F",
INIT_3E => X"0000000000000000000000000000000000000F7D5555FFAAAAA8BFF002AAAA00",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_2,               -- Port A enable input
WEA      => wbe_a_hi_1024_2(1),               -- Port A write enable input
DIA(0)   => data_write_a(12),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_2(12),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_2,               -- Port B enable input
WEB      => wbe_b_hi_1024_2(1),               -- Port B write enable input
DIB(0)   => data_write_b(12),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_2(12),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_13_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10154A0441836CA2840512822007C18000E02700500030B31B300040081A042",
INIT_01 => X"00000804A000C04800020000000002404001000008220008A200100802110204",
INIT_02 => X"02200430000104000A4700804008000004100000000420918204D3033240400D",
INIT_03 => X"AA4003400008592400000590C40009141100000C6180C0000000C00001E14000",
INIT_04 => X"0800000102400120088054019000004160004190BAA0270000C8100000600206",
INIT_05 => X"21000012040610050040000227003AA0082400E94C1200000824424005220020",
INIT_06 => X"81963B180C001010580000080400000058000004109C00138000020024142581",
INIT_07 => X"002C8008000441600106400A9600010494020002B8AAA000EF003408000E2580",
INIT_08 => X"000000E48194408000A00A001210040441C80320040210000002ABF004102244",
INIT_09 => X"2A004009640040100400940412D4C4004000022000104200802D983000480120",
INIT_0A => X"8000202020401480000000000000080C90090881000145B0111A14004015080D",
INIT_0B => X"00000002004040AA08050400404040C11444000805200A402090024000008002",
INIT_0C => X"8410000A00280020020040800020040800020000801020000800010020400000",
INIT_0D => X"84A14250A055100050100490000500D00040080040290000084E4000B800610C",
INIT_0E => X"DCD13042BEDA36820228000000000000C000400081A08BC812A2092B02850942",
INIT_0F => X"89B9A260857DB400431969CA985D480949D32804A40AB137341C10B7D6A02EC0",
INIT_10 => X"E6ACA678001CE7D0296C213A460CA4271CA2168AEC1017606E6838216FAD4055",
INIT_11 => X"84AD4961C281B20213073C5FC0058008632D30D522CE80239DCC01AB013A4D20",
INIT_12 => X"2E6B13804A4B01D83461299900F6BD583A519104A0EEBD1A141010B2A4C8E116",
INIT_13 => X"89E5E40913419151EE0E94641828F72B5151EE0D184B321037AF5158BB02D085",
INIT_14 => X"562EC0B42162D68EE0073AE1C562EC13D521921A4170300B2B458B56B01C2280",
INIT_15 => X"00888A120240034000E6DC8285028014B82372011FC1E4F5E0A00929684EAF84",
INIT_16 => X"50942509425094250942509425094254940A1421420082020120908800480030",
INIT_17 => X"0942509425094250942509425094250942509425094250942509425094250942",
INIT_18 => X"9425094250942509425094250942509425094250942509425094250942509425",
INIT_19 => X"F7EFBBEEFF3F7DF7FF3E9F7DF7E2450228000000000000000000509425094250",
INIT_1A => X"BAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBF7DFDFDDD555555",
INIT_1B => X"EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAEBAE",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000000000F7EBF5FAFD7EBF5FAFD7",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"2ABEF00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0020105D557FEAA00557DE10AAD5554BA087FFFF55557BD54AAF7FBC01FFA280",
INIT_29 => X"7BD75EF087FFFFEF557BEAB45552E80155AA802AB45AA843FE0008557DFFF080",
INIT_2A => X"FAE820AA5D5557555082ABDF5508557DF45002ABDFFFF7803DE10AA80000AA08",
INIT_2B => X"0051555FFA2AA8200000557DFFFF7AA80000AAD1420AA087BD7555FFD168AAAF",
INIT_2C => X"5557FFDE10AAAEA8BFFA2FBD7545FFD157555085140010F7AEAABFFAAD542000",
INIT_2D => X"BA557BE8A10A284154BAFFAAAAB45007FC2155F7D155545AA80001EFAAFBEAB4",
INIT_2E => X"000A2D155410F7FFFFEBA08003FE00082AA8AAAAAFFC00BA00002AAAAF7D5574",
INIT_2F => X"0492E3F1C71C7BE8A2ABD7000000000000000000000000000000000000000000",
INIT_30 => X"3AE38145B78FD7000005010495B7AE921C517DE10A2DB50482147FFAF554971D",
INIT_31 => X"E3FE28B684070AA1C71D25D7007FFAFD7497BE8B5555208217DBE8A2AB45BE80",
INIT_32 => X"7FD257DFFD568A82FFA4870BA555F5056D002EBDF6D005B78F7D142ABDFC7F78",
INIT_33 => X"FAAAFBFFBED547038145B505FFB6A487000005F7AFD7F7A482038AADF4709214",
INIT_34 => X"AA8E071D7AAFBEFB455D71F8E00A2A0ADBC7A2FFD257DE3DF52555085142000F",
INIT_35 => X"21C002AA92FFDF574824171EAA10B680124BAFFAAAFB45007BC217DEBDB55555",
INIT_36 => X"00000000000000000000B6D550428FFF1FDE821C003FE001C2EAAAAAB6F5C208",
INIT_37 => X"0105D7BE8B55085142010AAD157545F7AEA8B550000000000000000000000000",
INIT_38 => X"01EFF7AAA8B55F7802AABA5D7FEAB45080015410007FEAA0055517DE00A2FFC0",
INIT_39 => X"E8BFF5D2ABDF55F7AABDEAAF784154BA5D5140145007BE8B55087BEAB555D040",
INIT_3A => X"0020BAA2FFD54105D7FC21EFFFD16AA10FF80174AA557FC21EF082EBFFEF007B",
INIT_3B => X"FBC0155085540000FFAEBFFEFF7D1554BA5D7BC01FFFF8015410007FEAB45F78",
INIT_3C => X"87FC01EFA2FFD7545AAAE97555A2FBFDF455D556AA00A2803FF45AAFFC21EFAA",
INIT_3D => X"552EAAAAAFFD1400005D042AA00F7FBD5410085568A10FF80020AAFFAABFF550",
INIT_3E => X"0000000000000000000000000000000000000F7D1400BAFFD57FE005D043FE10",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_2,               -- Port A enable input
WEA      => wbe_a_hi_1024_2(1),               -- Port A write enable input
DIA(0)   => data_write_a(13),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_2(13),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_2,               -- Port B enable input
WEB      => wbe_b_hi_1024_2(1),               -- Port B write enable input
DIB(0)   => data_write_b(13),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_2(13),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_14_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10020A000180000284008280000281800000030000000033022000000580002",
INIT_01 => X"000008020000204D006800000030824840000000084000084200090008510200",
INIT_02 => X"0220043170010A600A4D008040080000041000000028009002000F333240800C",
INIT_03 => X"111813400008002400000000C400090011000000610200001104D83000F14000",
INIT_04 => X"0801800100A000000000540084000040000040000800200000C8100000000748",
INIT_05 => X"0100000000001000000000002000080008000000001000000024024001200020",
INIT_06 => X"819EB84028001010000000080400000000000004108000100000020020040081",
INIT_07 => X"92040608000440100102400A94810206844200021DA2A0002000340800062C80",
INIT_08 => X"000000000084400008800A001214040441481500040000000000A7F408002244",
INIT_09 => X"0A0040090002008420401004104444004000020400214A208001000002400120",
INIT_0A => X"0400002020000000000000000000080C8008088100004590111B480040120000",
INIT_0B => X"1000000200404800000504016000002114000008020000020080024000000000",
INIT_0C => X"0410000010000000000040001000000000000040000000000001000000000000",
INIT_0D => X"04810244825010004010000000000000000000000000000000080000B8002104",
INIT_0E => X"0002C38280001202020800000000001000004000000000401022000002040902",
INIT_0F => X"20000587050001404E8084341CBA3404800828805200008000E0E0A000080002",
INIT_10 => X"4D18178E012010C00224004091C3514072C000444A0400080001C1C140001000",
INIT_11 => X"51709A07424142084458476001003809D0104B01C5710044020C4006010500C5",
INIT_12 => X"C26EE3803180C18006519462A00005001460E4730000050A1011004001060049",
INIT_13 => X"01F9E00660318000000538318740000140000001B4600CE80001400000002B62",
INIT_14 => X"0000000AD89857B0E0684411800000003799EB764D000330C300000000E3554B",
INIT_15 => X"0000021002002C000024008284001A0902000422E3F5960080480A0216A07240",
INIT_16 => X"4090240902409024090240902409024090081021020080015134920800480010",
INIT_17 => X"0902409024090240902409024090240902409024090240902409024090240902",
INIT_18 => X"9024090240902409024090240902409024090240902409024090240902409024",
INIT_19 => X"F5579B4E5C8FF0F7BE9D5F7DF650400200000000000000000000409024090240",
INIT_1A => X"9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7BF7DDDDDFCF3CF3D",
INIT_1B => X"F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE79E7",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000003FFF03F9FCFE7F3F9FCFE7F3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"420BA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"BD54AAF7FBC01FFA2802ABEFA2FBE8B55A2AE80000F7D5555555D2AAAABAAAD1",
INIT_29 => X"AA801FFA28402000AAAE955455500155EF0804155EFAAD5554BA087FFFF55557",
INIT_2A => X"7AEA8B45080417400AA843FE0008557DFFF0800020105D557FEAA00557DE10A2",
INIT_2B => X"087FFFFEF557BEAB45552E80155AA802AB4500516AA00A2AE800BAFFFFC20BAF",
INIT_2C => X"0AA80000AA005568ABAA28402010A2843FEBAFFFBD7410A2D168BFF087BD75EF",
INIT_2D => X"005D7FFDF4555517DFEF00043FEAA082ABDF5508557DF45002ABDFFFF7803DE1",
INIT_2E => X"000AAD1420AA087BD7555FFD168AAAFFAE820AA5D5557555002E80155A280000",
INIT_2F => X"0555412AA8ABAAADB40092000000000000000000000000000000000000000000",
INIT_30 => X"50482147FFAF554971D0492E3F1C71C7BE8A2ABD7A2FFEDB55B6A080038E3DB5",
INIT_31 => X"B7AE921C517DE10A2AE851FFB68402038AAAA955554900105FF0800175D7A2DB",
INIT_32 => X"A0800BAE3F1C0092EBAAADB6D080A12410BE803AE38145B78FD7000005010495",
INIT_33 => X"2D568BC71C71D25D7007FFAFD7497BE8B5555208217DBE8A2AB451C556FA00A2",
INIT_34 => X"142ABDFC7F78E3FE28B684070AA00516DABAA28402038B6803DE82F7F5D5410A",
INIT_35 => X"D002A80155B680000105D7FF8F455D5F78FD7000E3FEAA002EBDF6D005B78F7D",
INIT_36 => X"00000000000000000000AADF47092147FD257DFFD568A82FFA4870BA555F5056",
INIT_37 => X"F55FF84000AAAAFBC0145002AA8AAAAAFFC20000000000000000000000000000",
INIT_38 => X"01EF080417555A2FFC00105D7BE8B55085142010AAD157545F7AEA8B55A2FBFF",
INIT_39 => X"EAB45080015410007FEAA0055517DE00A2AA955FFFF80020BAAAAA9754508000",
INIT_3A => X"AA8B555D557FE00A280020BAAAD140000A2AEBFFEF082A82010F7802AABA5D7F",
INIT_3B => X"803DE00FFD557400AAD56AB455D5140145007BE8B55087BEAB555D04001EFF7A",
INIT_3C => X"82EBFFEF007BE8BFF5D2ABDF55F7AABDEAAF784154BA08557FEAAA284000AAFF",
INIT_3D => X"FF80174AA557FC21EF082A80145F780020105D7BEAB45557BE8B45082EBFEBA0",
INIT_3E => X"0000000000000000000000000000000000000A2FFD54105D7FC21EFFFD16AA10",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_2,               -- Port A enable input
WEA      => wbe_a_hi_1024_2(1),               -- Port A write enable input
DIA(0)   => data_write_a(14),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_2(14),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_2,               -- Port B enable input
WEB      => wbe_b_hi_1024_2(1),               -- Port B write enable input
DIB(0)   => data_write_b(14),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_2(14),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_15_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000A000000000284000280000001800020030000000033022000000180002",
INIT_01 => X"8000080000000048000000000000026040000000080000080200000000110200",
INIT_02 => X"0020042004010E60004C0080000800000410000000020090020000300245E005",
INIT_03 => X"0000010000080400000000408400480111000000610008000000C00000E54400",
INIT_04 => X"980000010000000088C2550080000040000040000008A00028C8100000120000",
INIT_05 => X"020004012E025000000001322000000A28008000011000000220004D41000000",
INIT_06 => X"819588000800101000011008040000100001060418800510000A620000000092",
INIT_07 => X"0000000800044004010C20008440810284020002102220002000340800062480",
INIT_08 => X"0000000001140800002C0A001214050540C800400406180000002DF004000244",
INIT_09 => X"1E00400900000000000016041044400440000000000042008001000000000022",
INIT_0A => X"0000000000000220000000000000080C00000081000045901118000040000000",
INIT_0B => X"0000000200404000010500004000000114000009000000000000004200000000",
INIT_0C => X"0000000000000000000040001000040001000000000000000001000020000800",
INIT_0D => X"000000000000001001208000180800000000030200000180800C400030002000",
INIT_0E => X"0000000000002600020800000000001080004000000000000002000000000000",
INIT_0F => X"A400000000000000000008000000000000000000000014800000000000000052",
INIT_10 => X"0000000000000000000000010240000000000000000000290000000000000000",
INIT_11 => X"2001C05838120800000000000000000000010000000000000000000000001804",
INIT_12 => X"081004000000000000A010000000000000902000000000180010002020000000",
INIT_13 => X"6600000000000000000024080000000000000000280400000000000000000000",
INIT_14 => X"0000000000200801000000000000000000501001920000000000000000000A40",
INIT_15 => X"0000020000000000000000003000000000000000000A101C3614000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000080000120980000000010",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000400200000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"28BEF00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"5555555D2AAAABAAAD1420BAFF8000010082A954BA00003DFEF085155400F784",
INIT_29 => X"AE95555A2FBE8BEFA2843DE00AA8015400FF84001EFA2FBE8B55A2AE80000F7D",
INIT_2A => X"2FBEAB45F7D56AABAAAD5554BA087FFFF55557BD54AAF7FBC01FFA2802ABEFF7",
INIT_2B => X"A28402000AAAE955455500155EF0804155EFFFFBE8BFF0800174AA557BFDE10A",
INIT_2C => X"A00557DE10F7D1574AAA2D16AB55FFD568BEF087FE8A1055003FE00A2AA801FF",
INIT_2D => X"00AA802AA00AAAE800BA5D0015545AA843FE0008557DFFF0800020105D557FEA",
INIT_2E => X"00000516AA00A2AE800BAFFFFC20BAF7AEA8B45080417400FFFFC21450800154",
INIT_2F => X"8FD7005150438F78A2DBFF000000000000000000000000000000000000000000",
INIT_30 => X"EDB55B6A080038E3DB50555412AA8ABAAADB40092E38E070280024904AA1C043",
INIT_31 => X"1C71C7BE8A2ABD7E3AA9257DA2FFE8BC7BE8E38E10A28017400E38A051FFA2FF",
INIT_32 => X"00124AA557FFDE10A2FBEDB6DF7D16AABAA2DB50482147FFAF554971D0492E3F",
INIT_33 => X"10038E38A2AE851FFB68402038AAAA955554900105FF0800175D7E3FFEFBD700",
INIT_34 => X"000005010495B7AE921C517DE10FFDF50482A2DB6AB45FFD56DBD7087BEAA384",
INIT_35 => X"0FFF1C017D140410400BE8E28A10AAA085082550A1057DBE803AE38145B78FD7",
INIT_36 => X"000000000000000000001C556FA00A2A0800BAE3F1C0092EBAAADB6D080A1241",
INIT_37 => X"4AA0800020BA550028B550855400AAF7AEBDFEF0000000000000000000000000",
INIT_38 => X"7400AAAE975EFA2FBFFF55FF84000AAAAFBC0145002AA8AAAAAFFC2000AAAA97",
INIT_39 => X"E8B55085142010AAD157545F7AEA8B55AAAE821EFAAFBEAB55F7AAA8A00AA841",
INIT_3A => X"417555AAFFFDF450804020AA557BFFE10A2FFFFFEFF7D568ABAA2FFC00105D7B",
INIT_3B => X"D17DF45007FE8AAA08002AAAAA2AA955FFFF80020BAAAAA975450800001EF080",
INIT_3C => X"7802AABA5D7FEAB45080015410007FEAA0055517DE00FFFBC2000AAFBE8B55F7",
INIT_3D => X"A2AEBFFEF082A82010FFD5421EF5D0000010F7AAA8A10AA8017400552A801EFF",
INIT_3E => X"00000000000000000000000000000000000005D557FE00A280020BAAAD140000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_2,               -- Port A enable input
WEA      => wbe_a_hi_1024_2(1),               -- Port A write enable input
DIA(0)   => data_write_a(15),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_2(15),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_2,               -- Port B enable input
WEB      => wbe_b_hi_1024_2(1),               -- Port B write enable input
DIB(0)   => data_write_b(15),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_2(15),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_16_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"DA22C618B1000482B688B186588884862A400438255FC38381441205BA803003",
INIT_01 => X"7045A80028404C211203A952A90341080B173340412000E1005D628000820484",
INIT_02 => X"428406A4000850848330118D0AAC55001349B108818005460229044001C01784",
INIT_03 => X"092C4020000500020000500986812C405000001A48202050000A214AC0650115",
INIT_04 => X"4804A55440256F504025E003A054F46415A4E62B6FE3307943965A00001A1152",
INIT_05 => X"0000001C40A5B950ADB8EA097057ECE14C86D2B7F85AAD17F4B100000B88148C",
INIT_06 => X"415401DCDCF2C0A8030140BCB0820A200342A1C641C1E8782F508F2B00003584",
INIT_07 => X"002701881A3202080AE00480A2002840BE1480FA004342AA6F12000054004867",
INIT_08 => X"08C54828091002000002B32A8C19064E486A8001510000014140C1E2A14891E0",
INIT_09 => X"015452B103020814004088B64102680B6596594800400413CAC0208944800000",
INIT_0A => X"96AA000484094C000000000000012C9000A0000D0A80000BF8028E87C1B99270",
INIT_0B => X"014808A02004200E540480212000A448C0082024AE50064B44000000000002A2",
INIT_0C => X"0004000D5846256AAEA811150445411150445411150445411150422A088A8200",
INIT_0D => X"00000004010042A204A0C5817D00005034052E40000817D00440004004AD3240",
INIT_0E => X"632B2673FA4587978A2004102800809225545155121740000004900090000000",
INIT_0F => X"00C6564CE7F4EA4B940076D296D003030800462CBD320018CAAAACFE9164C800",
INIT_10 => X"28834ADB1440A114793A4A30A40839AA14910D08DCB2640031955559FD3AC990",
INIT_11 => X"594AB0B1A025371CA0E034E8443C097A800EB090D4AAC91208ED2FA0CE5E09B1",
INIT_12 => X"7B50446083001B94BB38C540EBE61284BB304880E3E4579EDC00992980D58033",
INIT_13 => X"5511121840E7A2CD952ECC12ABC3E6ACB3DFB12ECE315000F61FF1727A85FDBC",
INIT_14 => X"75DEB07F6F2E7084517F126F8395CB2BEFBAB8BA8AF698228CC5E2F08ECA5159",
INIT_15 => X"5580A840A8009F8B108C80A1021B080AFC0DF6422C6077F4A77F20D0C0E21084",
INIT_16 => X"0000000000000000000000000000000000044000102A0001148442A110810359",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"558D11544C690DA64C1C4F68A360400000000000000000000000000000000000",
INIT_1A => X"14D14D14D14D14D14D14D14D14D14D14D14514514514514529E5F87869E79E78",
INIT_1B => X"D1E8F47A3D1E8F47A7D3E9F4FA7D3E9F4FA7D3E9F47A7D1E9F47A7D1E9F4D14D",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000007D3E9F4FA7D3E8F47A3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"C00AA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"03DFEF085155400F78428BEF087FFFFEFF7D168B55AAD17FFFF552EBFE00007F",
INIT_29 => X"2E975EFF7D568BFFFF80175EF0004000BA552A821FFFF8000010082A954BA000",
INIT_2A => X"55540000082EAABFFA2FBE8B55A2AE80000F7D5555555D2AAAABAAAD1420BA5D",
INIT_2B => X"A2FBE8BEFA2843DE00AA8015400FF84001EF0000020AA5D00154005D043FF455",
INIT_2C => X"FA2802ABEF557BEABEF5D0415410087FD74BAAAAEBFFEF557FC00AAF7AE95555",
INIT_2D => X"FFFFAABFEAAFF84001FF002A821FFAAD5554BA087FFFF55557BD54AAF7FBC01F",
INIT_2E => X"000FFFBE8BFF0800174AA557BFDE10A2FBEAB45F7D56AABA082A97545F7D16AB",
INIT_2F => X"FFEF552AB8E38087FC2092000000000000000000000000000000000000000000",
INIT_30 => X"070280024904AA1C0438FD7005150438F78A2DBFF0871F8FC7E3D56AB6DBEDB7",
INIT_31 => X"AA8ABAAADB400924920925EFF7D16ABFFE38E175EF1400000BA412E871FFE38E",
INIT_32 => X"0A1240055003FF6D5551420101C2EAFBD7A2FFEDB55B6A080038E3DB50555412",
INIT_33 => X"57FC00BAE3AA9257DA2FFE8BC7BE8E38E10A28017400E38A051FF0804050BA41",
INIT_34 => X"4971D0492E3F1C71C7BE8A2ABD74975EDBC7550E12410087FD74AAB6AABFFC75",
INIT_35 => X"A08249756DF7D168BC7F7AABAEAAF780051C70824851D7A2DB50482147FFAF55",
INIT_36 => X"00000000000000000000E3FFEFBD70000124AA557FFDE10A2FBEDB6DF7D16AAB",
INIT_37 => X"B55A2D16ABEFFFFBFDFFF552AAAAAA007BC00000000000000000000000000000",
INIT_38 => X"20AA002A955EFAAAA974AA0800020BA550028B550855400AAF7AEBDFEF08516A",
INIT_39 => X"000AAAAFBC0145002AA8AAAAAFFC20000000021EFF7D568BFFA2AA955FF5D040",
INIT_3A => X"E975EF0800174BA002E820105D003DFEF5D51420005D2ABFF45A2FBFFF55FF84",
INIT_3B => X"7BD74AAF7AEBDF455D7BC20BAAAAE821EFAAFBEAB55F7AAA8A00AA8417400AAA",
INIT_3C => X"2FFC00105D7BE8B55085142010AAD157545F7AEA8B5500557DF45552A8200000",
INIT_3D => X"A2FFFFFEFF7D568ABA0804155FFF7D568B55FFAAAAABAFF8415545000015555A",
INIT_3E => X"0000000000000000000000000000000000000AAFFFDF450804020AA557BFFE10",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_2,               -- Port A enable input
WEA      => wbe_a_hi_1024_2(2),               -- Port A write enable input
DIA(0)   => data_write_a(16),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_2(16),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_2,               -- Port B enable input
WEB      => wbe_b_hi_1024_2(2),               -- Port B write enable input
DIB(0)   => data_write_b(16),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_2(16),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_17_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"5284CE4FB7BD2C8994A13392DBD02E14006B82AC7E800D44D3DD2FD5F9B961C0",
INIT_01 => X"2EACD01F7E03FC6793F2199B39FC233C11D93AE6F3BB92B32091DBC339B24542",
INIT_02 => X"E63CCCC00A82C08092A2AFAE667033DB50853379C10BFDC5C6F4044443C817C6",
INIT_03 => X"7FF183635AEF9E3635AEF9E18E237040404446965C0607EE6DB7854AC4DE060C",
INIT_04 => X"D78AC33FB604488B000892EF17BE6D84196482236FE100294152E294350FB697",
INIT_05 => X"081B5F9B409420D0CDB47A05403F6CE0C08A4AB7F840EDB6F48100DFC8081081",
INIT_06 => X"768465354781CBC30316367077B4BDB50646E8D87100A8201ED01C19C020F71A",
INIT_07 => X"4002A110C922480A82D0841147162C48EBB9537A0022DC67987042EE976ABEA7",
INIT_08 => X"DB931BFEF91C00002CC0E019C0C82A4E4820C15A2330E004401891181168C4D1",
INIT_09 => X"09F3A1BC11EFBC66DB65307071477FF1030C397C060B4254064302042F803A69",
INIT_0A => X"3F330802162F3B7EE3F3EC7C7DEF207000F00059D2ED56D7EED2ED3C9A867DC0",
INIT_0B => X"185C44B91BC1740B7605040BE0018CFC7429F326B9E822FFC00074D5A0AB033A",
INIT_0C => X"00367A28FC1B7F7FEFFCFBFF3EFFCFBFF3EFFCFBFF3EFFCFBFF3EFFE7DFF9E00",
INIT_0D => X"0000000008004BA78428C7AD7FC94B533F5B4FFBD2FAD7FCCA786D43FE67C218",
INIT_0E => X"BA494CEBFD4F2667ABB6F68B29760593F33FA0CF170F40006001B1A05C000000",
INIT_0F => X"7F749299D7FAEB237DFE5865B6D2BF23265CBACE542A6FEE92333AFF33E0A9BF",
INIT_10 => X"F6C24B6D18C3C9F8E2881F3F787D776B5DB94A09955054DFDD246675FE7AC153",
INIT_11 => X"BFB349E08FF9A27EDE9FA8AEFD9E7467BFCB195CFEB56A1A70D34D1706FFFA3E",
INIT_12 => X"6FE219CA80725B875EED723FF7FCB2875EDAAFEAF7FD929BFD55BBC71D79F639",
INIT_13 => X"546670D018E7A6E581D7B6AB75FDFCECA6E581D7BB5DDFC6FF0EB7D7E859FDB5",
INIT_14 => X"B978177F6D6AF5ECDB5FB76A5F5FA165B456E0FB308710C49FCFB741598B9C7E",
INIT_15 => X"CFDAAB00AC00A8BBFC8B501CF7A0FED9A540EA1952586CEB54D143ACFF9A3BA9",
INIT_16 => X"000000000000000000000000000000000026E100002F382DBD9ECFE117805F20",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"4372003009EDCC4052E917114F981800C0000000000000000000000000000000",
INIT_1A => X"BA69A69AEBA69AEBA69A69AEBA69AEBA69A69A69A69A69A68698686981D75D74",
INIT_1B => X"6A351A8D46A351A8D068341A0D068341A0D068341A0D46A341A0D46A341A69AE",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000000000046A351A8D46A351A8D4",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"7FEAA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"17FFFF552EBFE00007FC00AA087FFFFFFFFFFFFFEFF7FBEAB450804001EFAAD5",
INIT_29 => X"D168A000004020AA5D7BE8B450051401EF087FD74AA087FFFFEFF7D168B55AAD",
INIT_2A => X"D7FEAB55FF80175EFFF8000010082A954BA00003DFEF085155400F78428BEFAA",
INIT_2B => X"F7D568BFFFF80175EF0004000BA552A821FF5D00020BA552A82000552A821555",
INIT_2C => X"AAAD1420BAFFFFFDF45AAD17FFFFAAFBC01EF5D0015555557BFDEBA5D2E975EF",
INIT_2D => X"BA007FEABEF005555555A2D1554BAA2FBE8B55A2AE80000F7D5555555D2AAAAB",
INIT_2E => X"0000000020AA5D00154005D043FF45555540000082EAABFF00516AA10552E820",
INIT_2F => X"8B550000071EFB6DF7AE92000000000000000000000000000000000000000000",
INIT_30 => X"F8FC7E3D56AB6DBEDB7FFEF552AB8E38087FC2092147FFFFFFFFFBFDFC7EBF5E",
INIT_31 => X"150438F78A2DBFFBED16AA381C0A07082497FEFB6D1451471EF007BD04920871",
INIT_32 => X"2A850105D2A80155417BEFB6DEB8E175FFE38E070280024904AA1C0438FD7005",
INIT_33 => X"D7BFAEBA4920925EFF7D16ABFFE38E175EF1400000BA412E871FF550A0009249",
INIT_34 => X"E3DB50555412AA8ABAAADB40092FFF5FFF6DAADF7FFD7B6F1C71EF55001756D5",
INIT_35 => X"7145B6AA28492487082007FEDBD700515556DA2DF50492A2FFEDB55B6A080038",
INIT_36 => X"000000000000000000000804050BA410A1240055003FF6D5551420101C2EAFBD",
INIT_37 => X"FEFF7FBFFF55A2D16AB550000175EFFFFBEAA000000000000000000000000000",
INIT_38 => X"55EF087FC200008516AB55A2D16ABEFFFFBFDFFF552AAAAAA007BC0000557FFD",
INIT_39 => X"020BA550028B550855400AAF7AEBDFEFF7D568AAA5D2A97410007BFFFFF55515",
INIT_3A => X"A955EF5D2E80010002A954005D2A82155087FFFFEFAAAA975EFAAAA974AA0800",
INIT_3B => X"D1575FF5504175EF5D7FEAAAA0000021EFF7D568BFFA2AA955FF5D04020AA002",
INIT_3C => X"2FBFFF55FF84000AAAAFBC0145002AA8AAAAAFFC2000FFD57DFFFAAFFFDF55FF",
INIT_3D => X"5D51420005D2ABFF45557FE8AAA000415410007BFFF450051555EFA2FBC0000A",
INIT_3E => X"00000000000000000000000000000000000000800174BA002E820105D003DFEF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_2,               -- Port A enable input
WEA      => wbe_a_hi_1024_2(2),               -- Port A write enable input
DIA(0)   => data_write_a(17),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_2(17),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_2,               -- Port B enable input
WEB      => wbe_b_hi_1024_2(2),               -- Port B write enable input
DIB(0)   => data_write_b(17),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_2(17),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_18_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"69844019080000A21A611406840014122A641074155FC28A2024001001801003",
INIT_01 => X"7443D920034004180005E9E3C90360C0041C0181002001602025800008440084",
INIT_02 => X"E2DCCCE61D5C008103F2000781FC0FEDEAC2161B0B8FB0008620044443006010",
INIT_03 => X"884E300802006900802006995C896D605200000856E24A040000640052141103",
INIT_04 => X"480520FC026125AC0025C9122644E3E40EC8E2001001302281841A009038A86A",
INIT_05 => X"432000040089983070019400F01010004C8DB841405A80A100B586200FAC24AE",
INIT_06 => X"09044359DC7040000000002C109B0E0A00A1104641C0803804000707284600E1",
INIT_07 => X"400D10100400481D5EB08501620000007500CE801241021FE78E404860140060",
INIT_08 => X"00880C0106A0528020019307CC082A0A4A6A01ED725021400040D028000A9729",
INIT_09 => X"00117063038000282081402E4106400B6186128040600C10C1C0200950508110",
INIT_0A => X"C0C30C2E21580C874004008080003C32A10A19090C02010E1022944061688000",
INIT_0B => X"0180A8062026000DC425C0301311324AA2373088479105D044A1022000001835",
INIT_0C => X"0D89844703649000000200000000000000000000000000000000000000000010",
INIT_0D => X"0D8306C182701404C1973010802020404084001E00010802046092B5001FB365",
INIT_0E => X"528EB314068AB8B803DB00002900800400FC503F08180050942E4200020C1B06",
INIT_0F => X"40A51D66280D6032C5F96D3C51555D5D7D5AA87285820814A3CCC501C2A60820",
INIT_10 => X"8B35A3FEBF1FEDFD9C2B30E0468AAAD5D48F37E8FC1304102947998A03984C10",
INIT_11 => X"440FE1DD772D37A0A321BC6968F32658BF2D4F2A80BF8FE3F9FE3AC362080529",
INIT_12 => X"5487910D7E5A6D961A28456A1832E5161A100DD5182BC54020EA67A189C6ED36",
INIT_13 => X"AA444CAF91EDD1B725868403BE06323551B725868A100ABD119753B70964122B",
INIT_14 => X"EDC259048ACD868EE3803D65CEDC258A8F80D55E007C3F8EBB56F4C5362C978F",
INIT_15 => X"3F240014BE84370001B6922070440556B15F7FABBC0031BCF2257C41634B14D4",
INIT_16 => X"C1B06C1B06C1B06C1B06C1B06C1B06C1B0491069068000004060300A005A0118",
INIT_17 => X"1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06",
INIT_18 => X"B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C",
INIT_19 => X"B28BBECEB80EE173C2300F7DF16000000000000000000000000041B06C1B06C1",
INIT_1A => X"8A28A28AAAAAAA28A28A28AAAAAAA28A28A28A28A28A28A2910591505C104104",
INIT_1B => X"28944A25128944A25128944A25128944A25128944A2552A954AA5128944AAAA2",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000128944A25128944A251",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"9540000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"BEAB450804001EFAAD57FEAA087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974BA082E",
INIT_29 => X"7FFFFFFFFFBFDF45AAD568B55080028B55002E82000087FFFFFFFFFFFFFEFF7F",
INIT_2A => X"0043DE10AA843DE00087FFFFEFF7D168B55AAD17FFFF552EBFE00007FC00AA08",
INIT_2B => X"0004020AA5D7BE8B450051401EF087FD74AAAAFFFDF45A2D16AB55F7FFFFFFF0",
INIT_2C => X"0F78428BEFAA80000000804154BA55042ABEF5D7FD75FFAAD540145AAD168A00",
INIT_2D => X"00082E95555085168A10557FD7545FF8000010082A954BA00003DFEF08515540",
INIT_2E => X"0005D00020BA552A82000552A821555D7FEAB55FF80175EF5D00020105D2A974",
INIT_2F => X"DFFF5D2A954AA082A92428000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFBFDFC7EBF5E8B550000071EFB6DF7AE921C7FFFFFFFFFFFFFFFF7FBF",
INIT_31 => X"AB8E38087FC2092087FFDFC7E3F1FAF55A2DF6DB7D1C002AB7D002A82028147F",
INIT_32 => X"DF6DB7DE3F5FAFC708003DE28B68E38E280871F8FC7E3D56AB6DBEDB7FFEF552",
INIT_33 => X"ADF4516DBED16AA381C0A07082497FEFB6D1451471EF007BD0492B6F1F8F55AA",
INIT_34 => X"1C0438FD7005150438F78A2DBFFA28407038140410492550A2ABC7497BD25FFA",
INIT_35 => X"F5D0E05000492097428002E9557D1C516FA28417BD5545E38E070280024904AA",
INIT_36 => X"00000000000000000000550A00092492A850105D2A80155417BEFB6DEB8E175F",
INIT_37 => X"FFFFFFFFDFEFF7FBFFFEF552E974AA082A820AA0000000000000000000000000",
INIT_38 => X"ABEF002A800AA557FFDFEFF7FBFFF55A2D16AB550000175EFFFFBEAA00557FFF",
INIT_39 => X"6ABEFFFFBFDFFF552AAAAAA007BC0000087BFDF45AAD568B55AAFBFDFEF55042",
INIT_3A => X"FC2000FFD56AB45A2FFFDFFFAAD16AB4500043DEAAFFAEAAAAA08516AB55A2D1",
INIT_3B => X"2AA8B45087FC01EFA2FFD55EFF7D568AAA5D2A97410007BFFFFF5551555EF087",
INIT_3C => X"AAA974AA0800020BA550028B550855400AAF7AEBDFEFA280154BA55040000055",
INIT_3D => X"087FFFFEFAAAA975EF5D2E974000804154BA082A975EF5D517DEAA007BD5545A",
INIT_3E => X"00000000000000000000000000000000000005D2E80010002A954005D2A82155",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_2,               -- Port A enable input
WEA      => wbe_a_hi_1024_2(2),               -- Port A write enable input
DIA(0)   => data_write_a(18),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_2(18),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_2,               -- Port B enable input
WEB      => wbe_b_hi_1024_2(2),               -- Port B write enable input
DIB(0)   => data_write_b(18),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_2(18),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_19_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"042200000000000041088001001AA00000000000000000000000500802000003",
INIT_01 => X"040048000024000000000404000000000A22000800000800004A200000000001",
INIT_02 => X"200C8840085EB00480060000001C008002489E0F000405EA0004040404000000",
INIT_03 => X"24004000000000000000000900002C4050000000000069500208400002E14100",
INIT_04 => X"4800200C0000000044002000C80020E40000E200000130200188000000800100",
INIT_05 => X"000000000080181000000000701000004C8000000058800000B1000009880480",
INIT_06 => X"80500081081040000000002C100040400000004641C080380400070100000000",
INIT_07 => X"4020109801A4CE005C00048380142810010564C4100114012002402028044808",
INIT_08 => X"0070700000000000000083004C3902420062000020E0000100004082A140102B",
INIT_09 => X"001150200000000000000026400000016186100000000010C04002C000000000",
INIT_0A => X"007C00008082C0002000000000002C3000000004050001030102040000000000",
INIT_0B => X"0000000000000000000000000000010000800011000000000000000000000BC0",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"000000000000000000000000000000042000760000000000000000010004B200",
INIT_0E => X"0D74002280300F0002FB069040000060000C5003000800000000000000000000",
INIT_0F => X"C01AE8004500744C780687DBA828008080A5FC0D385598035D0008A00C015660",
INIT_10 => X"39D8140040201BF861F0E7D693E6170022408116DFE0AB3006BA0011401D02AC",
INIT_11 => X"5412E4997F5249FD005043B8680CC98F00D0F2DD0140100406FE053A98F6ECC7",
INIT_12 => X"7418663001858040E153888000010840E165D0000000285C246A181C03FE4662",
INIT_13 => X"8199830066F0020858385974000001260208583854E2200000660208D6B1423F",
INIT_14 => X"8235AC508FCE8811042040F008235AE04420C040CF00C031C80009B8F224978B",
INIT_15 => X"030004E00000C220010808C10D9A92A74CD7CF4A09051110AD5A3C9200B7F280",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000118",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"07208BBA3F0C7010C660C7441920000000000000000000000000000000000000",
INIT_1A => X"861869A61861861861869A61861861861861861861861861A8208C4C1534D34C",
INIT_1B => X"984C26130984C26130984C26130984C26130984D26930984C26130984C261861",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000984C26130984C26130",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"174BA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFDFEF5D2A974BA082E95400F7FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0004",
INIT_29 => X"FFFFFFFFFFFFFFFFF7FBFDFFF552E974BAA2FFFFE10087FFFFFFFFFFFFFFFFFF",
INIT_2A => X"004001EFAAAEA8ABA087FFFFFFFFFFFFFEFF7FBEAB450804001EFAAD57FEAAF7",
INIT_2B => X"FFFBFDF45AAD568B55080028B55002E82000F7FFFFFFFFFFFFDFEFA2D568B550",
INIT_2C => X"0007FC00AAF7FFFFFFFF7FBE8B55AAD16ABEF5D2ABFF55080402010087FFFFFF",
INIT_2D => X"55A2FFFDFEF5D2EBFE00AAFFFFEBA087FFFFEFF7D168B55AAD17FFFF552EBFE0",
INIT_2E => X"000AAFFFDF45A2D16AB55F7FFFFFFF00043DE10AA843DE00557FFDFEFA2D16AB",
INIT_2F => X"FFEF552A974AA0000104AA000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFF7FBFDFFF5D2A954AA082A92428E3FFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"0071EFB6DF7AE92EBFFFFFFFFFFFFDFEFF7F5FAFC7492A974AAB6F5F8E101C7F",
INIT_32 => X"F1F8FD7AAD16AB450000001FFBEA4A8AAA147FFFFFFFFFBFDFC7EBF5E8B55000",
INIT_33 => X"00000010087FFDFC7E3F1FAF55A2DF6DB7D1C002AB7D002A82028FFFFFFFEFF7",
INIT_34 => X"BEDB7FFEF552AB8E38087FC2092F7FBF8FC7E3F5EAB45B6DF6FBEF5D2AB8F7D0",
INIT_35 => X"84971F8FC7AAD56DB6DBEF5F8FD7412ABFE28B6F5F8E820871F8FC7E3D56AB6D",
INIT_36 => X"00000000000000000000B6F1F8F55AADF6DB7DE3F5FAFC708003DE28B68E38E2",
INIT_37 => X"FFFFFFFFFFFFFFFFFDFEF552E954AA0004000AA0000000000000000000000000",
INIT_38 => X"54AAF7D568A00557FFFFFFFFFFFDFEFF7FBFFFEF552E974AA082A820AAA2FFFF",
INIT_39 => X"FFF55A2D16AB550000175EFFFFBEAA00A2FFFFFFFF7FBFDFFFFFD568B55002A9",
INIT_3A => X"A800AAF7FBFDFEFF7D56AB45AAD56AB450004001EFFF842AAAA557FFDFEFF7FB",
INIT_3B => X"FFFFFFF552AA8BEF080402000087BFDF45AAD568B55AAFBFDFEF55042ABEF002",
INIT_3C => X"8516AB55A2D16ABEFFFFBFDFFF552AAAAAA007BC0000FFFBE8B55AAD168B55F7",
INIT_3D => X"00043DEAAFFAEAAAAA08556AB55A2D57FFFFF7D568B45002ABDEAAFFD16AA000",
INIT_3E => X"0000000000000000000000000000000000000FFD56AB45A2FFFDFFFAAD16AB45",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_2,               -- Port A enable input
WEA      => wbe_a_hi_1024_2(2),               -- Port A write enable input
DIA(0)   => data_write_a(19),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_2(19),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_2,               -- Port B enable input
WEB      => wbe_b_hi_1024_2(2),               -- Port B write enable input
DIB(0)   => data_write_b(19),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_2(19),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_20_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000003",
INIT_01 => X"F55FF80000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"E05022020800008400F655001FFCFF80018FA804400000000000004400000001",
INIT_03 => X"00000000000000000000000900002CC07000000000000000000000000000013F",
INIT_04 => X"68002FFE40900010000180000001FFEC0012EE0C001370F40780000000000000",
INIT_05 => X"0840000880FCBBF0100E204DF0F88311DD8005080679800000F3000029980580",
INIT_06 => X"001000030817C8E8840155FDF9001001050023F6C3C3D0F87FA19F7F011000E4",
INIT_07 => X"000000090492260800008000EE00000000000000002101FF2002C00000004018",
INIT_08 => X"2A040001071004000013FF7FCA302C0C0008214800002101554031F800000000",
INIT_09 => X"801F57F200000090000489FEC0000001EFBEF0040008023FDFC0000000004006",
INIT_0A => X"0000000008000000000000000000ADF000000200000008000008028300110230",
INIT_0B => X"0000000000000800080000000000000000000000000000000800800A40000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"000000040900005C848538000020000000800000080000020000800101FFB600",
INIT_0E => X"00800000003A010003000000000000600FFC53FF001800000002004080000000",
INIT_0F => X"0001000000007408040000004000000004E9000008020000200000000E800800",
INIT_10 => X"00200000000313100010002000008000000000129600040000400000001D0010",
INIT_11 => X"81C012060000000000218F7840000100800004000000000066C0000080080000",
INIT_12 => X"800000000017C000100000000001A800080000000001A8040000002840008185",
INIT_13 => X"0000000006F00000100200000000012600001004000000000066000000801040",
INIT_14 => X"0000200410100000000005F00000020080090A0000000085C800002000586000",
INIT_15 => X"FF00400000000000020020020001000040283024E4F2860400008000030ED080",
INIT_16 => X"00000000000000000000000000000004010201001003020200000000000127DB",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"A0700030038200010089120104D2040020000000000000000000000000000000",
INIT_1A => X"2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2C30C30C30C30C306982121A1E79E79",
INIT_1B => X"32190C86432190C86432190C86432190C86432190C86432190C86432190CB2CB",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000432190C86432190C864",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0201000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF552A974AA0004174BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA0804",
INIT_29 => X"7FFFFFFFFFFFFFFFFFFFFFFEF552E954AA000400000F7FFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E954BA007FC00BA087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974BA082E9540000",
INIT_2B => X"FFFFFFFFFF7FBFDFFF552E974BAA2FFFFE10FFFFFFFFFFFFFFFFFFFFFBFDFFF5",
INIT_2C => X"FAAD57FEAA007FFFFFFFFFFFFFEFF7FBFFF550800020BAAAD56AAAAF7FFFFFFF",
INIT_2D => X"EFF7D56AB450000021EFA2D57DE10087FFFFFFFFFFFFFEFF7FBEAB450804001E",
INIT_2E => X"000F7FFFFFFFFFFFFDFEFA2D568B550004001EFAAAEA8ABA5D7FFFFFFFFFFFDF",
INIT_2F => X"FFFF5D2E954AA080005000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFEF552A974AA0000104AAFFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"A954AA082A92428087FFFFFFFFFFFFFFFFFFBFDFEF5D2E974AA000A07000E3FF",
INIT_32 => X"FFFFFEFF7FBFFFFF552E974AA0071C50BA1C7FFFFFFFFFFFFFFFF7FBFDFFF5D2",
INIT_33 => X"EDF6FABAEBFFFFFFFFFFFFDFEFF7F5FAFC7492A974AAB6F5F8E10E3FFFFFFFFF",
INIT_34 => X"EBF5E8B550000071EFB6DF7AE921C7FFFFFFFFFBFDFEFE3F5F8F450004050AAB",
INIT_35 => X"A497FFFFFFF7FBF8FC7EBD168B450804021FFB6D57DE28147FFFFFFFFFBFDFC7",
INIT_36 => X"00000000000000000000FFFFFFFEFF7F1F8FD7AAD16AB450000001FFBEA4A8AA",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2A954AA0800174100000000000000000000000000",
INIT_38 => X"74AA002E95410A2FFFFFFFFFFFFFFFFFFFFFDFEF552E954AA0004000AAFFFFFF",
INIT_39 => X"FDFEFF7FBFFFEF552E974AA082A820AA087FFFFFFFFFFFFFEFF7FBFDFFF5D2A9",
INIT_3A => X"568A00AAFFFFFFFFFFBFDFEFFFFFFDFEF5D2E954AA0051554BA557FFFFFFFFFF",
INIT_3B => X"D16AB450804174AAFFFFFFEBAA2FFFFFFFF7FBFDFFFFFD568B55002A954AAF7D",
INIT_3C => X"57FFDFEFF7FBFFF55A2D16AB550000175EFFFFBEAA005D7FFFFEFF7FBFDFFFAA",
INIT_3D => X"0004001EFFF842AAAA087BFDFEFF7FFEAB45A2D568B550804001EFF7D57DEBA5",
INIT_3E => X"0000000000000000000000000000000000000F7FBFDFEFF7D56AB45AAD56AB45",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_2,               -- Port A enable input
WEA      => wbe_a_hi_1024_2(2),               -- Port A write enable input
DIA(0)   => data_write_a(20),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_2(20),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_2,               -- Port B enable input
WEB      => wbe_b_hi_1024_2(2),               -- Port B write enable input
DIB(0)   => data_write_b(20),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_2(20),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_21_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"4A302428B824900A128C090A5C1800261500213C005FE812D10420054085A202",
INIT_01 => X"001FFE3440B609703B0427F801A40B8115BC4F655300340288A40D30040E4DD8",
INIT_02 => X"E00424256888D8819801000F9FFFFFFFF149FF1FCA448046C60A0D2437C517F9",
INIT_03 => X"20030640003250640003250F06002CC1740002019824E001CD357832440001FF",
INIT_04 => X"EA2C3FFD400006E04401A8837001FFFC004AEF00080B70E08FB5789421007C5C",
INIT_05 => X"00011A0C40F9FFF80920954FF0F00809DF84A0202879800000F3000029980780",
INIT_06 => X"0805984B7A1FC0A0000101FFF0480080002281F7C3C381F87C03DFFF00009004",
INIT_07 => X"B424068086A205481A60A19000908204A855B000A08A61FF20C3D004D331D340",
INIT_08 => X"1BFA0001600802000023F7FFC08D234B40C2028253000040114200000D0226C0",
INIT_09 => X"EF1F5FF054096C6ADBA169FFC202B1C1FFBEF0440021083DFFCE22DC2880E24D",
INIT_0A => X"45FF0C004041D84862A28C54518DBFF00020004C0A6044901112A0908AA0A300",
INIT_0B => X"018C241102068006C620C03882019480E63180855A492712CC01C49C20201BFE",
INIT_0C => X"08A9464116544302C02D92236488D92236488D92236488D922366446C911B210",
INIT_0D => X"08800444021048034004001890000806002804A0822189000900D80621FFBE00",
INIT_0E => X"060580261013813A2CC396506102C4053FFD5BFF00A04A00200602CA52001100",
INIT_0F => X"080C0B004C202621A85C09411500135844C196D3606941018150098404C1A304",
INIT_10 => X"B02901013416181C96C2C9C600890A2028172192C460D1820302A0130809834A",
INIT_11 => X"9C5E803408250180AC268D185DB3F4350B811068C00049A0A4AA68F05C96A001",
INIT_12 => X"002C006560138F032B1804101244C883052208209040CC849063A747512B7678",
INIT_13 => X"41401E240665750440C9488280254530314080C2C601040420352148A00501B1",
INIT_14 => X"500811204D000700114204A70422016149916011008CAA8858850B00C32591C0",
INIT_15 => X"FFC06E60AC0496022300233104663040808E991765205000070121D41D18D098",
INIT_16 => X"40100401004010040100401004010040102090010008000001C0E010020007DF",
INIT_17 => X"0100401004010040100401004010040100401004010040100401004010040100",
INIT_18 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_19 => X"FFEF9FEEFF7FFDF7FF3E3DFDF7E0000000000000000000000000401004010040",
INIT_1A => X"BEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBFFDFDFFFCF3CF3F",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFEFF7FBFDFEFF7FBFDFEFBEF",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000FFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0001000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E954AA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0004",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA0004154BAFFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"52E974BA0804000AAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0004174BAFF",
INIT_2B => X"FFFFFFFFFFFFFFFFEF552E954AA000400000007FFFFFFFFFFFFFFFFFFFFFFEF5",
INIT_2C => X"A082E95400007FFFFFFFFFFFFFFFFFFFFDFEF5D2E974BA002E97400007FFFFFF",
INIT_2D => X"FFFFFBFDFEF5D2A954AA002E974BA087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFBFDFFF5D2E954BA007FC00BA5D7FFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA000002000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080005000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"A974AA0000104AAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974BA0000174AAFFFF",
INIT_32 => X"FFFFFFFFFFFFDFEF552E954BA080A000AAE3FFFFFFFFFFFFFFFFFFFFFFFEF552",
INIT_33 => X"02A95400087FFFFFFFFFFFFFFFFFFBFDFEF5D2E974AA000A07000007FFFFFFFF",
INIT_34 => X"F7FBFDFFF5D2A954AA082A924281C7FFFFFFFFFFFFFFFFFFBFDFEF5D2A974BA0",
INIT_35 => X"A557FFFFFFFFFFFFFFFF7FBFDFFF552E974BA0020924BA1C7FFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000E3FFFFFFFFFFFFFFEFF7FBFFFFF552E974AA0071C50B",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0000020000000000000000000000000000",
INIT_38 => X"74BA0000174BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954AA080017410FFFFFF",
INIT_39 => X"FFFFFFFFFFDFEF552E954AA0004000AAF7FFFFFFFFFFFFFFFFFFFFFFFEF552A9",
INIT_3A => X"E95410087FFFFFFFFFFFFFFFF7FBFDFEF5D2A954BA082E800AAA2FFFFFFFFFFF",
INIT_3B => X"FBFFFFF552E954BA002E97410087FFFFFFFFFFFFFEFF7FBFDFFF5D2A974AA002",
INIT_3C => X"57FFFFFFFFFFFDFEFF7FBFFFEF552E974AA082A820AA557FFFFFFFFFFFFFEFF7",
INIT_3D => X"5D2E954AA0051554BA5D7FFFFFFFFFBFDFEFF7FFFFFEF5D2A974BA0000020AA5",
INIT_3E => X"0000000000000000000000000000000000000AAFFFFFFFFFFBFDFEFFFFFFDFEF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_2,               -- Port A enable input
WEA      => wbe_a_hi_1024_2(2),               -- Port A write enable input
DIA(0)   => data_write_a(21),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_2(21),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_2,               -- Port B enable input
WEB      => wbe_b_hi_1024_2(2),               -- Port B write enable input
DIB(0)   => data_write_b(21),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_2(21),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_22_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"5290F4CDE914905A14A43D33F488243E17122300F55FEB189B343A1140548380",
INIT_01 => X"A54007B259F6A975386262000C344BA9573C6FF57B18A5FB0ABFCD3C2C5F4F0C",
INIT_02 => X"021DFF8C38B3C009D203551040030071869D0040180AA2DC53DB89BEA8204001",
INIT_03 => X"2603475A969D0475A969D0460EAA401005111011BD506954EDB40F5EF41434C0",
INIT_04 => X"922D9002100ED69E443D988B0D5400103E48003D0800011E803B06B5B9125A15",
INIT_05 => X"281B5A0C06000408F4DF9422010D8802022F2124A8022492580040440002021C",
INIT_06 => X"F780C4C052881ADA0E05440205DA50930FA182010004700083E220800440B588",
INIT_07 => X"049D028B93FB561833D8094A02F5EA92FD7247E10305C40040D136E6A023F7FC",
INIT_08 => X"00028241680A0E002A9400803A884B5B5206B7C2E53CA25144009007A64EBD64",
INIT_09 => X"41008810240240C6694008010392354010000560141801002028A83D2A08E06D",
INIT_0A => X"34000000848BCA6902A29C54539C020E11810098D4067EFF9FF284D483E2AB41",
INIT_0B => X"500001840000C80B410014088040F4A944B1AA313C0022AA0011C0DC00028001",
INIT_0C => X"80B14004D158C8CA24A1C2A870AA1C2A870AA1C2A870AA1C2A872550E1543800",
INIT_0D => X"80A14050A01509E050854498B5281A1C34E506A2C6898B52A154DAC6B6000850",
INIT_0E => X"0B03001A483A4146603050080410089180008800143D83888281A2034A850142",
INIT_0F => X"A4160600349075238473F1210006133835E92273612B3482C090068A0E84AC56",
INIT_10 => X"30060181BA1B13959DC08DA902458870201970B29602562B0581200D141D0959",
INIT_11 => X"E042021C040D0152C8058B3840F044708E7E1C20A0106EA166C13AFC14AA3804",
INIT_12 => X"080E004B0C17C1439A9838301DC1A8438EA32C009DC1A8255300650458A1D588",
INIT_13 => X"018010E186F110A908E3A8CB0026C9A610A908E6A60F0807626610E160589C4C",
INIT_14 => X"2A701667334005800B1605F043858125E0D04110408D2485CA034681E43A1E40",
INIT_15 => X"00646002304244A91102C93A2D608D2A258DF8034188200C050171A41108F084",
INIT_16 => X"110441104411044110441104411044110466C440446CA06951D4EA8010009804",
INIT_17 => X"0040100401004411044110441104411044110441104411044110441104411044",
INIT_18 => X"0401004010040100401004010040100401004010040100401004010040100401",
INIT_19 => X"F7DFBFDEFE8FF1F7DEBDDF7DF7D05122890000000003FFFFFFFF900401004010",
INIT_1A => X"9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7BFFDFD7DDDF7DF7D",
INIT_1B => X"F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE79E7",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000003F9FCFE7F3F9FCFE7F3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA000400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0800",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000002000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2A954BA000015400FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080402010FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2A954BA0004154BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A0004174BAFFFFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0800154AAFFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF552A974AA0000174BAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974A",
INIT_2E => X"000007FFFFFFFFFFFFFFFFFFFFFFEF552E974BA0804000AAA2FFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080400010000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E954AA080005000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000402010FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2A954BA000417410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"804154BAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974BA0000174AAFFFFFFFFFFF",
INIT_34 => X"FFFFFFFEF552A974AA0000104AAE3FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0",
INIT_35 => X"AA2FFFFFFFFFFFFFFFFFFFFFFFEF552E954BA000E124BAE3FFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000007FFFFFFFFFFFFFFFFFFFFDFEF552E954BA080A000A",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804000100000000000000000000000000",
INIT_38 => X"54AA000400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2A954AA080017410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"0174BAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A954BA000415400FFFFFFFFFFFFF",
INIT_3B => X"FFFDFEF552E974AA0804174AAF7FFFFFFFFFFFFFFFFFFFFFFFEF552A974BA000",
INIT_3C => X"2FFFFFFFFFFFFFFFFFFFFFDFEF552E954AA0004000AAA2FFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2A954BA082E800AAAAFFFFFFFFFFFFFFFFFFFBFDFEF5D2E954BA002A820BAA",
INIT_3E => X"0000000000000000000000000000000000000087FFFFFFFFFFFFFFFF7FBFDFEF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_2,               -- Port A enable input
WEA      => wbe_a_hi_1024_2(2),               -- Port A write enable input
DIA(0)   => data_write_a(22),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_2(22),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_2,               -- Port B enable input
WEB      => wbe_b_hi_1024_2(2),               -- Port B write enable input
DIB(0)   => data_write_b(22),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_2(22),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_23_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"EF20906D902424807BC8241BC81801B97D38AD3C0800103362A6741C80A12A02",
INIT_01 => X"001FFF8409F089003B4422000D80C80106804A7951C5B9D1C828043EA28838F9",
INIT_02 => X"E01CEE21649C82C40800000F9FFEFF8E72CA7F5FC2E22809925A0D3611C877F8",
INIT_03 => X"24000400402670400402670D48222DC1764446838624000080007460C40001BF",
INIT_04 => X"68403FFC020560E0443E21037C01FFFC0002EE00628BF0E02FAD781014085014",
INIT_05 => X"0112000202FBFFF00920017FF0F0628BFF8488890979800002F702002BB807A0",
INIT_06 => X"EF85788B681FC000000001FFF0010000000001F7CBC385F87C0BFFFF20040001",
INIT_07 => X"F6E200000000C1440E3AE408009120071070FA07A1CB23FFA403F0C4D23BF7C0",
INIT_08 => X"0BF87CA400804000003FF7FFD8880A034AC09662305AB10555421006891A1089",
INIT_09 => X"BE1F5FEA10092C0896A243FFC0008087FFBEF2000000001DFFC612C0C0400100",
INIT_0A => X"41FF0C2060501000600000000001BFFA800808189A657EF81DD0C00079CC8001",
INIT_0B => X"018C24110A860006C620C0312241C482B20400CC52492710CC80060020A81BFE",
INIT_0C => X"0C08866907048320C20C10030400C10030400C10030400C10030400608018210",
INIT_0D => X"040002000041500300100040000500C000801000C02400000952800001FFBF04",
INIT_0E => X"FC850015385380380CDB86106502C5043FFD5FFF00A04BC010A7724B10000800",
INIT_0F => X"89F90A002A70A710A51C01C05904014861433602A1CAF13F2110055614C72FC0",
INIT_10 => X"E02D02001C1E14981B43253EE50C8220180F1082E06397E07E42200AAC298E57",
INIT_11 => X"8421802400A90022B0070FAE18019214A380344920080B21A58B02AC60BACDF0",
INIT_12 => X"0A2A000C480B0704B54028101AC49C84BB4100009AC49C80857A82D20CE8CB22",
INIT_13 => X"01E00C8103416445C12ED0400027C5292445C12D500B0005A62D344CB241D095",
INIT_14 => X"132C907425604680038706A35132C94BDD011010404428886AC91B11311C8280",
INIT_15 => X"FF000470BE0692020328CA0028042054A92771C50FC070110001C1680809591D",
INIT_16 => X"00802008020080200802008020080200800800200200000000000008004807DF",
INIT_17 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_18 => X"8020080200802008020080200802008020080200802008020080200802008020",
INIT_19 => X"0000000000000000000000000000000000000000000000000000008020080200",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080002010FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974AA000400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000400010FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974AA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080000010FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E954AA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954A",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA000015400FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080002010FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974AA000400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000402010FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E954AA080005000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA080407000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA00041741",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080000010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000402010FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2A954AA080002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954AA080017410FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"552A954BA000415400F7FFFFFFFFFFFFFFFFFFFFFFFFF552A954BA080015410F",
INIT_3E => X"0000000000000000000000000000000000000F7FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_2,               -- Port A enable input
WEA      => wbe_a_hi_1024_2(2),               -- Port A write enable input
DIA(0)   => data_write_a(23),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_2(23),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_2,               -- Port B enable input
WEB      => wbe_b_hi_1024_2(2),               -- Port B write enable input
DIB(0)   => data_write_b(23),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_2(23),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_24_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100600007FFF000080108004000800020000840041000080808",
INIT_02 => X"FC5CA803400EB8209000000F9FFEFF8E7240FF1FC22409EA04018E50074017F0",
INIT_03 => X"11100400000000400000000D00002CC07400000090C080019001010A000001BF",
INIT_04 => X"68003FFC00040000000000008001FFFC0002EE00000370E007A100000000E468",
INIT_05 => X"0000000000F8BFF00920004DF0F00001DF8000000079800000F3000029980780",
INIT_06 => X"6E461803081FC000000001FFF0000000000001F7C3C380F87C019FFF00000000",
INIT_07 => X"600C2400013649609C8000980040814210254000A00B21FF2003F2A80D500000",
INIT_08 => X"0BF80000000000000003F7FFD88D2B4A02C0940062EC2804001610020408178B",
INIT_09 => X"8E1F5FE010092C0892A041FFC0000001FFBEF0000000001DFFC002C000000000",
INIT_0A => X"41FF0C0000000000600000000001BFFA0000005501AA00000CE2000009400000",
INIT_0B => X"018C0411020600048620C030020502000200000400490510CC00040020201BF4",
INIT_0C => X"0808064106040300C00C10030400C10030400C10030400C10030400608018210",
INIT_0D => X"0000000000004003000000000000001200580000000000000000000001FFBE00",
INIT_0E => X"0086C022005381380FDB96516140C6043FFD5BFF000041000000004110000000",
INIT_0F => X"80010D804400A7240C840C201D0210840043B4804012500021E0088014C04940",
INIT_10 => X"4109038041021C980200D06410C1924030008142E06024A00043C01100298092",
INIT_11 => X"587CC200002100C14428090A1D02348190814C09C010104025AA40041A0D8005",
INIT_12 => X"022E0030300B0E46177004208000D8C61D7004300000D884817B00011306B2D9",
INIT_13 => X"01E003060344710009875C018100013831000985DC000C20003C310006143B70",
INIT_14 => X"4001850EDC004780144806A64400186CBF8961104000C3807884000846EB9500",
INIT_15 => X"FF0006E08C063C0220002201490418082010A57263E0100008000290161E711C",
INIT_16 => X"00000000000000000000000000000000000000000000000000000000000007DF",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"F2D0AEEAF6E7CC1132CDB4441990000000000000000000000000000000000000",
INIT_1A => X"BEFBE79E79E79E79E79EFBEFBEFBEFBEFBEF9EF9EF9EF9EFA69861219575D75F",
INIT_1B => X"783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1EFBEF",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000783C1E0F0783C1E0F0",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0201000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A000400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA000400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000400000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402010000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"00002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080002010FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000400010FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA00040000",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020100000000000000000000000000",
INIT_38 => X"74BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"000010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA000002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974AA000402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000002010F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_2,               -- Port A enable input
WEA      => wbe_a_hi_1024_2(3),               -- Port A write enable input
DIA(0)   => data_write_a(24),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_2(24),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_2,               -- Port B enable input
WEB      => wbe_b_hi_1024_2(3),               -- Port B write enable input
DIB(0)   => data_write_b(24),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_2(24),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_25_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100200002000000080100004000000020000800041000080808",
INIT_02 => X"FC400086000000800000000F9FFEFF8E738FFF1FC204010000000111568DD7F8",
INIT_03 => X"00000400000000400000000D00002CC4740000008000000080000000000001BF",
INIT_04 => X"68003FFF64A564AC000000000001FFFE0082EF00010370E007A1000000004000",
INIT_05 => X"0A00040148F8BFF80920804DF0F00101DFC040000079C92484F30499299837C1",
INIT_06 => X"66041803081FC0E0801101FFFD000E41002299F7E3C380F87C019FFF81200096",
INIT_07 => X"000000080480AE00000080000000000000000000A00B21FF2003E00000000000",
INIT_08 => X"1BF80000400A02000003F7FFFA0008000200A0400008A0000014100200081000",
INIT_09 => X"8E1F5FFA53EFBCACB2E369FFE0010001FFBEF80C40630C7DFFEEBAF000800202",
INIT_0A => X"41FF0C0600000000600000000001BFFE00301000000000000CC020000140000C",
INIT_0B => X"01DCCC31222730A49620C030020100000200000400490D10EC00040220201BF4",
INIT_0C => X"0808064106240300C00C10030400C10030400C10030400C10030400608018210",
INIT_0D => X"0883044582114013412080000000000000000000000000000012800001FFBE00",
INIT_0E => X"00040020000180380FC386106140C6043FFD5BFF00A04B80608003CB120C1106",
INIT_0F => X"0000080040000200040400000100000000009480000240000100080000400900",
INIT_10 => X"0001000000000808000000240000020000000100006004800002001000008012",
INIT_11 => X"0001001808220000002004001900000080800008000000000022400000088000",
INIT_12 => X"0010000000000E00110000000000408009000000000040808063004000008200",
INIT_13 => X"6000000000046100000240000000001021000004400000000010210000001010",
INIT_14 => X"4000000404000800000000060400000088000001800000001084000000088000",
INIT_15 => X"FF800C608C041002000002000006100000002100000000180600000000100018",
INIT_16 => X"4110441104411044110441104411044510629041040D180400000010028047DF",
INIT_17 => X"1104411044110441104411044110441104411044110441104411044110441104",
INIT_18 => X"1044110441104411044110441104411044110441104411044110441104411044",
INIT_19 => X"FBA2894A196A8C5A2932EC15DA080800002FFFFFFFFFFFFFFFFFC11044110441",
INIT_1A => X"2492492492492492492410410410410410410492410492412000531215A69A6B",
INIT_1B => X"158AC562B158AC562B158AC562B158AC562B1588C46231188C46231188C49249",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000B158AC562B158AC562B",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080000010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000010FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08000000",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_2,               -- Port A enable input
WEA      => wbe_a_hi_1024_2(3),               -- Port A write enable input
DIA(0)   => data_write_a(25),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_2(25),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_2,               -- Port B enable input
WEB      => wbe_b_hi_1024_2(3),               -- Port B write enable input
DIB(0)   => data_write_b(25),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_2(25),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_26_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"E9264EAB20190CA3BA4997AA9002AE9C001006B0778015CFA17E0811039879C7",
INIT_01 => X"2FFFF9BB1F773C7F9BB07DFFFDD863FC5FFF3FEFFBBF9FFB22FFFBC7B9F30686",
INIT_02 => X"E06CCC62052E708180F6FFBFFFFCFFFFF9C7FF7FC24332E642090000074037F6",
INIT_03 => X"428003739CD9863739CD9869FE2B7DEAF300029E4E300DFE69A6E644E6FF473F",
INIT_04 => X"7C2FEFFFF5BA124F003DD31EAFFFFFEE9FF7EE6F4C0770FFD7DC7CA53997B2B1",
INIT_05 => X"DFFB5421C1F8BBFAFDBFFACDF0FFCC05DDDBFF3690F9EDB7F5F7AFF639BD7DE3",
INIT_06 => X"EFD044ABC817C3E3A74667FDFFB6FF5727CC3BFEF7C3FAF87FF59F7FFBFEF69F",
INIT_07 => X"00003002132462052E708180EF060C18E5BEFB051225CDFF7002C4EEDE77F6E0",
INIT_08 => X"3FFF7D5000EC75088ED3FF7FC8790E46426CE06CB1F8E041051831FA3068D77E",
INIT_09 => X"C05FD7FF9BEFBDCEFBEE59FEF44F6603EFBEFAFCC2E35E7FDFD147CCF3F583FA",
INIT_0A => X"67FF1C7FBFADEB31E35768E8ED6BFDF3EB3EBF9DDBCE7FDC1DF8A760F3EACC02",
INIT_0B => X"5BDDCC3B336F7C548667D47B7737AF3FD62601EDC25B3533DCEB07F262213FFC",
INIT_0C => X"5F9A06E19F4D93A0EA0F78C35E30D78C35E30D78C35E30D78C35E986BC61AE31",
INIT_0D => X"5FD7AFEFDFFAF59B6FF28FE1D80D73D840607307DCFE1D80EF69A004DFFFF7FF",
INIT_0E => X"0004001F8041897B2FFFC6D86D70CE04FFFFF3FF1F5F5475BD7F72E4D75EBFAF",
INIT_0F => X"F60008003F008237B0040A00010003E020023E0201F45EC0010007E01047D17B",
INIT_10 => X"00010001DC0004C81003DE050A700200001DC0006863E8BD8002000FC0208FA2",
INIT_11 => X"2200E400002801E1A00004C21C0206F60081800800007B00010F02007EC09A0E",
INIT_12 => X"0880007E000807C7C1A612001E0015C7C19C22001E0015C59DFE82011A311AA0",
INIT_13 => X"00001BC00101F60409F0670840070809760409F06984800780097604067D0010",
INIT_14 => X"81019F40042100001F800203D81019EC085614000085C80023D81009CF008A74",
INIT_15 => X"FF802FFDFFAFD082003B032FB987E04021D481D4000819060801E0D00001231D",
INIT_16 => X"EBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEFFBFBFBFBBFCFBB0FFDFEFFEF2DFFFFFB",
INIT_17 => X"BFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAF",
INIT_18 => X"FAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFE",
INIT_19 => X"475B15BCF491E166CC8553F86EDB5C88646FFFFFFFFFFFFFFFFFEBFAFEBFAFEB",
INIT_1A => X"861861861861861861861861861861861861869A69A61861AFBD54D5F871C71D",
INIT_1B => X"984C26130984C26130984C26130984C26130984C26130984C26130984C261861",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000984C26130984C26130",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040201",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_2,               -- Port A enable input
WEA      => wbe_a_hi_1024_2(3),               -- Port A write enable input
DIA(0)   => data_write_a(26),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_2(26),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_2,               -- Port B enable input
WEB      => wbe_b_hi_1024_2(3),               -- Port B write enable input
DIB(0)   => data_write_b(26),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_2(26),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_27_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"00080A40000A41248002029000050A088000008242A0004404480002000A1155",
INIT_01 => X"2FFFF1C11F781C129C107DFFFE0860941E81258CA2B71C2220EC1B86E1A00002",
INIT_02 => X"E1000000810000014400FF6FFFF0FFFFF8007F1FC21110005080200000221FF0",
INIT_03 => X"4080026318C18226318C1821302232EAE00002BE001115FE48620040840A863F",
INIT_04 => X"643D4FFC2530000F003D821C0BFFFF8E9EF79E6D440748FED70060842105B0B0",
INIT_05 => X"D6F39020D1F8A3FAFDBFBACDC8FDC405D1DB7F1490E5EDB7D5CBADB2385D79C3",
INIT_06 => X"6FE000A38007C3032646EFF1F0B6FF46A78C39F8E723F2E47FE59C7F9ADA2612",
INIT_07 => X"00002820000000810000014401060C180190310540118DFF1000C0849673F6C0",
INIT_08 => X"3FF779100062B12A8EC3F47FC80208808210880C00082050000110023068D030",
INIT_09 => X"005F07E09BFFBD07FBAC09F8E42922038F7DF8BEC2E39C5F1FD047CEF1B582D8",
INIT_0A => X"63FF5D5F9FADE911E81C09818109E1F16B16B71092CE7ED81CF403601228C402",
INIT_0B => X"1BFDCC39732F3554866AD57C37BEAF1C152201A4C05B7531D56B05B06A213FF8",
INIT_0C => X"5BCA06F18FC59380F00E34430D10C34430D10C34430D10C34430F0861A2186B5",
INIT_0D => X"5B56ADAB5FAAE58B2F628EA0C80FA3F04040510768EA0C80CC61A0044DFFC6EB",
INIT_0E => X"0004001D800188792CE79715710AE4047FFD23FF315D54358D593474955AB6AD",
INIT_0F => X"520008003B000297B0040200010003E020001F0201E44A400100076000579129",
INIT_10 => X"00010001DC00004A10035E0408300200001DC000086BC8948002000EC000AF22",
INIT_11 => X"02002400002801E1A00000C01E0202F60080800800007B00000782006EC0820A",
INIT_12 => X"0080007E000006A7C10602001E0001A7C10C02001E0001C18DE282010A311AA0",
INIT_13 => X"00001BC00000FE0401F04300400708007E0401F04180800780007E04047D0010",
INIT_14 => X"81011F40040100001F800002F81011EC080604000085C80001F810094F008034",
INIT_15 => X"FF800C6DDDAFD082001B03249887E04001D481D4000009020801E0D00001021F",
INIT_16 => X"AB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6BF1EBDABD8E270BF84A25C6ACB777E3",
INIT_17 => X"B6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6AD",
INIT_18 => X"6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADA",
INIT_19 => X"490E2168100481CA860402104A471688747FFFFFFFFFFFFFFFFFAB6ADAB6ADAB",
INIT_1A => X"000000000000000000000000000000000008200000000000200072F210000001",
INIT_1B => X"05028140A05028140A05028140A05028140A0500804020100804020100800000",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000A05028140A05028140A",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040201",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_2,               -- Port A enable input
WEA      => wbe_a_hi_1024_2(3),               -- Port A write enable input
DIA(0)   => data_write_a(27),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_2(27),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_2,               -- Port B enable input
WEB      => wbe_b_hi_1024_2(3),               -- Port B write enable input
DIB(0)   => data_write_b(27),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_2(27),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_28_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"02200AA400180030808802A900002A08001280A08A801044104A1000001818C3",
INIT_01 => X"0AA00011460214428114180000882214413D0A71592A01D92213D28005210202",
INIT_02 => X"0451110A012100884000AA30200000000C100040104112101100008888200000",
INIT_03 => X"448000318C52A20318C52A20148810200111100C211004AA00034204200A2200",
INIT_04 => X"04004001001A90110000121402AA0000003C00000500000040080421080D0080",
INIT_05 => X"4060000C8001000000002E000000050000001610300000010000802202040012",
INIT_06 => X"1000002080001111001222000425A1040026A008000000000000000009328280",
INIT_07 => X"2491008A00491201210088400122448908A20402000408001000040820000000",
INIT_08 => X"20058310402A160026500000028040101004200C840082115554000112244814",
INIT_09 => X"4140000800000060000720000102028000000490160801020002200011100010",
INIT_0A => X"020000081B34211082B694D4D294000020020381040000000200032040004400",
INIT_0B => X"4800210C19808400500010009110091500020B408810000100200020408B0000",
INIT_0C => X"01028000080118020023604858121604858121604858121604858090B0242C00",
INIT_0D => X"010000800920040804020A6058003108402043058C460580653020005A004039",
INIT_0E => X"00000002800008014004104104420A00C000200005000010040A0020CC000200",
INIT_0F => X"520000000500000010000200000000000000280000040A40000000A000001029",
INIT_10 => X"00000000000000C0000002000830000000000000480008148000000140000020",
INIT_11 => X"020024000000000000000440000000020000800000000000000C00000040020A",
INIT_12 => X"00800000000001804006020000000500400C0200000005400A90000000100000",
INIT_13 => X"0000000000018200001003004000000142000010018080000001420000200000",
INIT_14 => X"8000080000010000000000018800008000060400000000000310000008000034",
INIT_15 => X"000002040080000000110006B081400000400000000009020000000000002200",
INIT_16 => X"802008020080200802008020080200802101210810C39A66A90A85420413A820",
INIT_17 => X"0200802008020080200802008020080200802008020080200802008020080200",
INIT_18 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_19 => X"DE21102C110A00246972BD89A40A0C22E1000000000000000000002008020080",
INIT_1A => X"2082082082082082082082082082082082082082082082080D35050758C30C31",
INIT_1B => X"0582C160B0582C160B0582C160B0582C160B0580C06030180C06030180C08208",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000B0582C160B0582C160B",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_2,               -- Port A enable input
WEA      => wbe_a_hi_1024_2(3),               -- Port A write enable input
DIA(0)   => data_write_a(28),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_2(28),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_2,               -- Port B enable input
WEB      => wbe_b_hi_1024_2(3),               -- Port B write enable input
DIB(0)   => data_write_b(28),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_2(28),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_29_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"79964E4BA01DACAB9E659792D00AAE160002829C7FDFEFCEE97C2815039D70C3",
INIT_01 => X"0ABFF9AB0775343F9AB01DF80D5821FC0FFF3FEFD1AF9FF1207FFBC7B9720586",
INIT_02 => X"002CCC60050E700080F6AAA7BFFC007189C7FF2FC00330E602800000074037F6",
INIT_03 => X"468003210868A63210868A68DA017D207200021C4E200CAA6186A40042FF4300",
INIT_04 => X"7C2FE002F0900001003C5316A6ABFFE21F36E02F0D03701F47D41800109FB281",
INIT_05 => X"4979440580F9B808F49F6A4DF00F8D01DC4B97369078249370F482E62BA41462",
INIT_06 => X"B250442BC81001E1870223FC0BF7F11507C423FE33C078F803F19F00E936721D",
INIT_07 => X"00011080012460050E700080EF020408EC8CFA01122149FF700200665A35D260",
INIT_08 => X"2BFD055040A452000443FF00007906464068406C31F84000000831FA1028575A",
INIT_09 => X"805FD017102690AA694551FE30444681E0820AD40201423FC00122C493500172",
INIT_0A => X"0600002AFFBE2330815568A8AD6ABC02A02A0B0CCB463B4C0748A720B1EA4C00",
INIT_0B => X"0850400A11414C005005000B51158936D20601A98A10200308A002E240010BFC",
INIT_0C => X"05928020194918A22A2268C81A32068C81A32068C81A32068C81A99034640C00",
INIT_0D => X"058102C48970541944B20FA1580561D040406305587A158046282000DBFFF13D",
INIT_0E => X"000000028040890327DCD28928324400DFFFF0001F1F0050342D42A086040B02",
INIT_0F => X"F60000000500802010000A000000000000022A0000141EC0000000A01000507B",
INIT_10 => X"00000000000004C0000082010A700000000000006800283D80000001402000A0",
INIT_11 => X"2200E4000000000000000442040004020001800000000000010D000010401A0E",
INIT_12 => X"08800000000801C040A6120000001540409C2200000015441DAC800010100000",
INIT_13 => X"0000000001019600081027084000000956000810298480000009560002200000",
INIT_14 => X"800088000021000000000201D800088000561400000000002358000088000A74",
INIT_15 => X"00802594A282C0000033010FB181E00020400000000819060000000000002305",
INIT_16 => X"C0B02C0B02C0B02C0B02C0B02C0B02C4B12B312912831A27FCFE7FFB175B6FF8",
INIT_17 => X"0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02",
INIT_18 => X"B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C",
INIT_19 => X"BBCF9F96EE7FFDF7FE783FFDFFEA0C00602FFFFFFFFFFFFFFFFFC0B02C0B02C0",
INIT_1A => X"EFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEEBAEBAEBAEBAEBBFFDF9FBEFFFFFFE",
INIT_1B => X"BFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFBEFB",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000FBFDFEFF7FBFDFEFF7F",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_2,               -- Port A enable input
WEA      => wbe_a_hi_1024_2(3),               -- Port A write enable input
DIA(0)   => data_write_a(29),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_2(29),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_2,               -- Port B enable input
WEB      => wbe_b_hi_1024_2(3),               -- Port B write enable input
DIB(0)   => data_write_b(29),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_2(29),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_30_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"F7FFBFFEFF9FE1F7FFBFFFFDFFD0000000000000000000000000000000000000",
INIT_1A => X"9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7AFBD75F5FDF7DF7F",
INIT_1B => X"F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE79E7",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000003F9FCFE7F3F9FCFE7F3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_2,               -- Port A enable input
WEA      => wbe_a_hi_1024_2(3),               -- Port A write enable input
DIA(0)   => data_write_a(30),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_2(30),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_2,               -- Port B enable input
WEB      => wbe_b_hi_1024_2(3),               -- Port B write enable input
DIB(0)   => data_write_b(30),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_2(30),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_31_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"129000008004A00804A40000400800020000000C005FEA005800200400050100",
INIT_01 => X"255FF18019700810180065FFFC0040801E80258CA2951C2200EC0906A0804140",
INIT_02 => X"E0000000000000011000550FDFF0FFFFF0007F1FC200000044000000000817F0",
INIT_03 => X"0000024210A30024210A3001002220C06044469200040154482000408400043F",
INIT_04 => X"602D0FFC2420000E003D80080955FF8E1ECA8E2D400340FE870060842100B030",
INIT_05 => X"0213100040F8A3F8FDBF944DC0FDC001D1CB6904A061EDB6D4C30490281831C1",
INIT_06 => X"6FC000830007C202060445F1F0D25E4207A099F0E303F0E07FE19C7F80402412",
INIT_07 => X"0000200000000000000001100004081001103107000185FF0000C0849673F6C0",
INIT_08 => X"1BF27A00000000000883F47FC800080002008000000820440000100220489020",
INIT_09 => X"011F07E013EFBC06FBA009F8E00120038F3CF82C44630C5D1FC002CCE0808248",
INIT_0A => X"61FF0C06C48BC801600000000001A1F00110101092CE7ED81CF0004012288000",
INIT_0B => X"11DCCC31222730048620C4382204A608142002A440492530C401049020221BF8",
INIT_0C => X"0888066187448380E00C10030400C10030400C10030400C10030600608018210",
INIT_0D => X"080204010200418301208480800D02D00040100240A808008840800405FF8640",
INIT_0E => X"0004001D000180780CE386106100C4043FFD03FF101D40008001304018081004",
INIT_0F => X"000008003A000217A0040000010003E02000160201E040000100074000478100",
INIT_10 => X"00010001DC00000810035C0400000200001DC0000063C0800002000E80008F02",
INIT_11 => X"00000000002801E1A00000801C0202F40080000800007B00000302006E808000",
INIT_12 => X"0000007E00000607810000001E000087810000001E000081846282010A211AA0",
INIT_13 => X"00001BC00000740401E0400000070800340401E04000000780003404045D0010",
INIT_14 => X"01011740040000001F8000025010116C080000000085C80000C8100947008000",
INIT_15 => X"FF800C609C06D082000A03200806A040019481D4000000000801E0D00001001D",
INIT_16 => X"010040100401004010040100401004010060C040040C200950402090128057C3",
INIT_17 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_18 => X"0040100401004010040100401004010040100401004010040100401004010040",
INIT_19 => X"00000000000000000000000000001000802FFFFFFFFFFFFFFFFF810040100401",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_2,               -- Port A enable input
WEA      => wbe_a_hi_1024_2(3),               -- Port A write enable input
DIA(0)   => data_write_a(31),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_2(31),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_2,               -- Port B enable input
WEB      => wbe_b_hi_1024_2(3),               -- Port B write enable input
DIB(0)   => data_write_b(31),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_2(31),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_0_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"ED39BA795990D275FB4A6E96ACC4731DEA4598B0AFB54867F6EE4618C3749803",
INIT_01 => X"8AA0047D8607944AC7DA180001ECA2444042106208408208C20022E9173734B3",
INIT_02 => X"1A7DDD79F9A73E6CCA7DAAF00001000008478020113D98E382FEDF333027C80F",
INIT_03 => X"75D341110C58F31110C58F32A208921F8051500147A0E4AB3493FB3A01EBE240",
INIT_04 => X"86424001531009B100425A97B2AA0001E03501D0A39C8F0078420001106D0C4C",
INIT_05 => X"BCC8CA2EBF03400700402BB20F00239E20341699198600000B08694B16434804",
INIT_06 => X"103FB860B2800161F8432200012DA185F80F24081C3C0707800E600056881308",
INIT_07 => X"B24197ABCDA467F9A73E6CCAFDC3870EEEEC44E2BDFE220094D03022210C011C",
INIT_08 => X"240581B5695EAA80262C080032BF07C7C1FC3F8E94F65B11555EAFFC1C306758",
INIT_09 => X"7E40000BEC004170040DB60017FED1CC0001045002984202003DB931192D60A5",
INIT_0A => X"120071411A74315881A28C141118000C5A85A60444210123820B43B40804674D",
INIT_0B => X"0820008E514045BB514F0106D1D8599581D3A958BC104A89215AC14C48898403",
INIT_0C => X"C261C01C48B1584A0CA3E2687A9A1E2687A9A1E2687A9A1E26870CD061343885",
INIT_0D => X"D274E93A758FA8683AC54B287522E10A74AF4AA59C568752662F5AC218000002",
INIT_0E => X"FF83C002783A0904231C70470C7E0B92800224008AE09FAD4BD48D1FC5D3A4E9",
INIT_0F => X"5BFF078004F075885DFBF7E15C06101C55E921F1F80FAB7FE0F0009E0E903EAD",
INIT_10 => X"F12E0380231F13978FF023FAFDBD9870380230F2D6081F56FFC1E0013C1D207D",
INIT_11 => X"DE7F263C0C8700125C0F8F3C43F1F10BBF7EFC61E01804E1E6C8F8FE807F67FB",
INIT_12 => X"02BE00017C17C1007E5E2E3081C5AC007E6F0E3081C5AC44418D65FE45DEE55B",
INIT_13 => X"61E0042786F103E9F01F9BC3C120C5A703E9F01F978B8C20666703E9F8A0FFED",
INIT_14 => X"FA7E283FFB414F80005F05F10FA7E283F78F6511C048278DCA174FF038FF15B4",
INIT_15 => X"0066A20B61692F293185D8D724E15D3FCC6B7C236FE0691B0700132C1F0EF880",
INIT_16 => X"3A4E93A4E93A4E93A4E93A4E93A4E93A4F942F92E9628540AD2A91442525A000",
INIT_17 => X"A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E9",
INIT_18 => X"4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93",
INIT_19 => X"55F3898E09B56C74DAB15D1CF13501AA495000000000000000003A4E93A4E93A",
INIT_1A => X"082082082082082082082082082082082082082082082082082084E41DC71C71",
INIT_1B => X"E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F82082",
INIT_1C => X"FFFFFFFFFFFFFFF94A5294A5294A5294A5294A52800003E1F0F87C3E1F0F87C3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"3060C183060C187FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"BDEBA0000000000000000000000000000000000000000000003060C183060C18",
INIT_28 => X"168ABA002E82145085155545F7AA975EFFFAABDE00FFAEBDFFF5D2EAAAAAF7AE",
INIT_29 => X"7FFFE10005542145557FD5545FF8000155087FC0155F7D168B55007BFDF45085",
INIT_2A => X"7FFC0010080017555555568AAAFFFFD7545AA8028A00A2802AABAFF8028BEF5D",
INIT_2B => X"FF842AABAA2AE95545FFD168ABAF7AEAAAAAA2FFFDF4500043FE105D2E954BAF",
INIT_2C => X"5007FD7400550415410002E974BA5D5168A00A2D142155005142010FFAE820AA",
INIT_2D => X"FFF780000BA007FE8AAAFF803FFFF5D2A821550000000BA007FD55FF5D7FC014",
INIT_2E => X"000AAFBEAA00007BFDFFF082EBDF455D5142000082E82145FFD17DFEFFFD168B",
INIT_2F => X"DFD75D2AA8A80EA8E2FE3F000000000000000000000000000000000000000000",
INIT_30 => X"68B551475FAF6D1C556F0AA1C24AABEA495FC716F002A975FFE3AA95E00EBAEB",
INIT_31 => X"42A0070071C50BAFEF1FAE0016D56A16D557BC257D415E0216FA3F1E8FC0145B",
INIT_32 => X"8010E004924874825D7FEAA85487FD24AFE3D02DAAAE12BD5545A2803AA00005",
INIT_33 => X"120155EA568E870BAEB8A05A2AEA8B50F55A2F150005A3A438BD04AFAB8F550A",
INIT_34 => X"545E055FFBE81D0BE8EA8A3AA05A2A5504001C74BA42A1571E8028E3DB7816D0",
INIT_35 => X"A5C7E3DFFFE90B45B47ABA497A82FFAFD2A82485FD2415A105C21451ED42A002",
INIT_36 => X"00000000000000000000B55EAAA100AA1D0F6F480B6A555A2A57A002A3D5FDB6",
INIT_37 => X"5EFAAAAB5E1AF3AABFF45592E88A0AFE80A8B0A0000000000000000000000000",
INIT_38 => X"65F520EBE9EF67D7BEA1FD5D556ABEF5D557FEBA55022A3F70C6B405F4D2AE97",
INIT_39 => X"C114728007521170821CE0FDE69411A8DED57CE1055555E5F58EFFC01FE2CACB",
INIT_3A => X"42341D5DEEBEF55080034E0A592A4AD0079C75D6070CC5CBB0280C029ABAA3EB",
INIT_3B => X"7F353AAF6C77F7F20D968BF57812A95E02A2AAB5EB0F280800EFAEE9F5D18F31",
INIT_3C => X"C91565455C141E41887D58AC448B69C30E02116220415A9540AA854140A0A204",
INIT_3D => X"DE6BE93172D7D625B556EEAB157ABEBE1B4D792A4AD1183454180DD3FDCAAAB7",
INIT_3E => X"F0000001FF0000001FF0000001FF0000001FF01EABC4B8014174FF7DA80F52FE",
INIT_3F => X"FF0000001FF0000001FF0000001FF0000001FF0000001FF0000001FF0000001F")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_3,               -- Port A enable input
WEA      => wbe_a_lo_1024_3(0),               -- Port A write enable input
DIA(0)   => data_write_a(0),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_3(0),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_3,               -- Port B enable input
WEB      => wbe_b_lo_1024_3(0),               -- Port B write enable input
DIB(0)   => data_write_b(0),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_3(0),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_1_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"212C001411984004084D000508C53810A03D1450E839B003342114428A000803",
INIT_01 => X"00000019400B100A8196000000CC004400400002000000000000028001340000",
INIT_02 => X"052137AE8031800C0044009000000000061800001CD4019802AD04CCCFC20004",
INIT_03 => X"04514108C60C21008C6042108400000201440020505100000043C30E10E9F000",
INIT_04 => X"02104001011DEFE088805681920000008000004001900800004002108C280008",
INIT_05 => X"040002340105000200000000080001900010000108040000000008411600401C",
INIT_06 => X"1034001042800808201000000001000820020000102000040000000000800180",
INIT_07 => X"64BF81A15EDFDE8031800C00843060C19E030022103600000450020800040004",
INIT_08 => X"00008004691687AA840008000090248CC84E000046000311555521F183060AC5",
INIT_09 => X"0820800D08100171000DB000154440C800400500000852020011200201012021",
INIT_0A => X"02000040001000880A2A04445004000102002041000001008208001440004140",
INIT_0B => X"4820018A1140440078050040511000102000A008183000010002404400000000",
INIT_0C => X"1000C80008000C030030880C2A030A00C28030A80C2A030A00C28018D4061401",
INIT_0D => X"10040802050080200284401C0022880F009E08008205C0020118088018000000",
INIT_0E => X"0F03C00280000000420860C60C0C0B92C0000000004000010042000040102008",
INIT_0F => X"001E078005000108400005E11C0610000000288058000003C0F000A000100000",
INIT_10 => X"F10E0380000000C202300000008D187038000000480800000781E00140002000",
INIT_11 => X"806302380C870010000004400100110800007861E0180000000C400680000001",
INIT_12 => X"023E00000000018000580C308000050000610C30800005000215006800000101",
INIT_13 => X"61E0000000018100B0001843812000014100B00016030C20000141002880026D",
INIT_14 => X"400A20009B404F80000000018400A20044096111C04000000304026000501580",
INIT_15 => X"0046820040082300218450C2800010094000482141E060190700100000002200",
INIT_16 => X"020080200802008020080200802008020080008008600500A82A1100A8000000",
INIT_17 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_18 => X"0080200802008020080200802008020080200802008020080200802008020080",
INIT_19 => X"81328A46BABEFC54A0810C7452B4428A14000000000000000000020080200802",
INIT_1A => X"AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA28A28A28A28A2A8218D2C0C924925",
INIT_1B => X"E974BA5D2E974BA5D2E974BA5D2E974BA5D2E975BADD6EB75BADD6EB75BAAAAA",
INIT_1C => X"FFFFFFFFFFFFFFFD8C6318C6318C6318C6318C63000002E974BA5D2E974BA5D2",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"70E1C3870E1C387FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"5555500000000000000000000000000000000000000000000070E1C3870E1C38",
INIT_28 => X"EBDF455D2EAABEFF7FFE8BFF5D0002155557FFFFFF007FC21EFA2FFD74AAAAD5",
INIT_29 => X"AA95400552AAAABAFFD1574105D7FD75FFAAAA800AAF7AA974BAFFFBE8B45F7A",
INIT_2A => X"0517DF555D2EAAA1055000015500557DF45AAD1400BAA2AE801550051555EFF7",
INIT_2B => X"FFD540155557FD5400F78028BFFFFFBEAB55F780020AAAA80020AA082EAAB550",
INIT_2C => X"AFF842ABEF5D517DF55552A974AAF7AE820AA0851574BAA2D1574AA5D7BFDEBA",
INIT_2D => X"EFAAD1575EF557FFFE10557FFFFFFFFD56AAAAFFFFD7555AAD168B45AAAEAAAB",
INIT_2E => X"0005D7FFDF4500043FE105D2E954BAF7AE80010082A97410557FEABFFAAFBE8B",
INIT_2F => X"51C7A2FBD5490BFD1C056A000000000000000000000000000000000000000000",
INIT_30 => X"974BAF7FFEFB45FFAABDF55492AA8BC2EBDFEAF7F1F840017D4975D2FEF147FC",
INIT_31 => X"080BEF495FC71D54124924385FAAA8AAAE3D145410F7F1D55D71C002DABAEBAA",
INIT_32 => X"002D082082AB8B6DBEDB7DF7F540E2AE85028B40155145F7AF6DBED5450AA1C2",
INIT_33 => X"78E021FF1471FDEAAFFD56F16D5571D2E28E38E0216FA2D1E8E80140F45082B4",
INIT_34 => X"A2DA3FB7DAAD4AAAAF487BC70BFA97F7AF6D417E92482BF84020BA495557E3FF",
INIT_35 => X"55554ADBD7A2FFC7BEFF6FFD7FC7002FD74951D71EDFFABFD16FAAAE92BD5545",
INIT_36 => X"00000000000000000000547AB8F550A8010E00492487482FFFE82A85EBAE2FFC",
INIT_37 => X"1EF005162BEF047FD5545AAFBF7400FBF9424F70000000000000000000000000",
INIT_38 => X"714F8338AAAA1D0AE974AAF7FFFDF55F7AABFF55082CA8B4DF6C1E8F5E540002",
INIT_39 => X"EABEF75550ACBB7582225FF5843404547184164AA5D2EBEEB0A2D555410D3555",
INIT_3A => X"FEAAEB083BC1000FF8409000512AEABFFDF79DCBF755962010BDCBBC21455D7F",
INIT_3B => X"801F8BA0C57740BDAA0688E5405D57D412F7D55F5E50C7F401BAAE8403CF5A3F",
INIT_3C => X"5D16BABAA3EBC3157ABD5FFE55F2AA9FEAFDF7F431A9F7FFE81FF013A8001AFF",
INIT_3D => X"FB863550229BCABEB7DA403FFFDA2FBF7FED2C7F955445079E280A00C56145EF",
INIT_3E => X"0000000000000000000000000000000000000596EBEF55080034E0A592A4AD00",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_3,               -- Port A enable input
WEA      => wbe_a_lo_1024_3(0),               -- Port A write enable input
DIA(0)   => data_write_a(1),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_3(1),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_3,               -- Port B enable input
WEB      => wbe_b_lo_1024_3(0),               -- Port B write enable input
DIB(0)   => data_write_b(1),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_3(1),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_2_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10E006600180111284380310006289800480032283E000A34301002001A0817",
INIT_01 => X"0005A00810790848048044A54E404350404000720885800802000906E4910200",
INIT_02 => X"407004208400408044C600C50AA055254010541A110222841200000002402544",
INIT_03 => X"0600011004182401004102408C28414043101000408118000145840440F5C415",
INIT_04 => X"5035855703A2900A000CD3088400F40688C9844409060850925E58A4081A0221",
INIT_05 => X"0200840D1021A15AC50494894850890540D1E12020C6E510818500440A280090",
INIT_06 => X"113044094002801020440090A8011A1224AB9380552102442884882A20004097",
INIT_07 => X"000100880004428400408044860000008C022402102100AA40004404B5075460",
INIT_08 => X"15C23440408C862A2A12382A8A5244145048C06085008010141521F000001240",
INIT_09 => X"400582B9033AA0E7AA4110B0506744810554542450694E710A836188C2C00222",
INIT_0A => X"443518360012C2210B020414109130A28038188096A06B8C120CA440A9C00802",
INIT_0B => X"1345E53300EC68005605002964AF222A5704004D080211121C80024200821780",
INIT_0C => X"181080C1110C882202211488452213C88472213C88472213488441109A442231",
INIT_0D => X"008204440210091341208041000810C00000300220201800A908000038AD0284",
INIT_0E => X"00040002804180300E88D28D206A40000554815500481440300000C44A081100",
INIT_0F => X"000008000500828700000000010000000002380000A00000010000A010050000",
INIT_10 => X"00010000000004CA000214000000020000000000684280000002000140200500",
INIT_11 => X"000000000020000000000442100002840000000800000000010C000026000000",
INIT_12 => X"00000000000805A4800000000000152300000000000015801272000100210020",
INIT_13 => X"000000000101C00000C000000000000940000120000000000009600004050000",
INIT_14 => X"0000130000000000000002018000106000000000000000002380000141000000",
INIT_15 => X"55000190000000000002000280000000011080C0000000000000000000002310",
INIT_16 => X"40902409064190641906419024090244902A9003004800415120D4A190804241",
INIT_17 => X"0900409004090641906419064190240902409024090641906419064190240902",
INIT_18 => X"9044090040900409004190441904419044090040900409004190441904419044",
INIT_19 => X"75960040138D70C030B51C50C7D100A2052F81F81F83F03F03F0419044190441",
INIT_1A => X"0410410410410410410410410410410410410410410410410248602081659659",
INIT_1B => X"5128944A25128944A25128944A25128944A25128944A25128944A25128941041",
INIT_1C => X"FFFFFFFFFFFFFFFE1084210842108421084210843FFF825128944A25128944A2",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"7FD5FF555815607FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"2AA000000000000000000000000000000000000000000000007FD5FF55581560",
INIT_28 => X"FC21EFA2FFD75EFAA8415410AA8415555087BFFF55A2AA800BAFFAE954000800",
INIT_29 => X"84155EFA2AEBDEAAA2FBEAABA5D7FE8B555551421455D0002145552EBFEBA007",
INIT_2A => X"2AEBDF555D2E954BAA2AA974BAFFFFE8B45552EBDF45FFAEAABFFF7FFE8B55F7",
INIT_2B => X"AAAAAAAAAFFD1574105D7FFFF555D2AAAAAA5D2E820BAA2FBEAB5555557DF55A",
INIT_2C => X"50055575EFFF84021555D043DEAA5D04021EF557FC21FFAA8428BFFAAAA954AA",
INIT_2D => X"10085568A00FF80175FFA2D17DFEFF7800215500557DF55AA80001FFAA800015",
INIT_2E => X"0005D00020AAAA80020AA082EAAB5500517DF555D042AA10A284154005D00154",
INIT_2F => X"00AAFFAA9543A080038A2A000000000000000000000000000000000000000000",
INIT_30 => X"0017D5D20B8EAA007FC51C7A2FBD55D2BE800042AFE8E1557D0075D2F45BEAA8",
INIT_31 => X"AA8BC7EBDFEAFEFFD00105FFBC20BDEAAA2FBF8AAA557BE8B6D5D5FFABEF4904",
INIT_32 => X"FFEFB6D555578F7DB6A0BDF7D480E174BFA02A974BAF7F5EFB455D2ABDF55492",
INIT_33 => X"ED1FDE90E3A497492B6AAADAAAE3D155E105571D55D71C002DABA5524820BAB6",
INIT_34 => X"BE8F401D7B6A0001470155C51D0092A071555D5E3AE821D00001FF0871C016DB",
INIT_35 => X"5BE8555400550A38428007FED000E3DA3DFD5E3DFFFBD5A38A021551C5F7AF6D",
INIT_36 => X"00000000000000000000410F45082B4002D082082AB8B6D1C5B7DF7FF78E075C",
INIT_37 => X"5EF005560B55F7AA800AAF7AA954AA00042AAA20000000000000000000000000",
INIT_38 => X"ABEF057D68F5F5A00021EF55042AAAA007FD5555AAFBD7545FBB8020A3F7AE97",
INIT_39 => X"7DF55D7AABFF5428ACA8F45A6C1E8F5EFF84165EFF7802BAB0A2FFEAABA557BE",
INIT_3A => X"CA8AA80800020AAF7FBFFFEF04552ABFFFF841FFE75CA882108202E974AAF7D5",
INIT_3B => X"00151FF0C57401E5F3D1E00A1A884174A8FFAEBFEB0A2D55541051555694F002",
INIT_3C => X"2AA801455D7FE8BFFF680800FFF7AAA155F595542455512A975455D3AA8A0055",
INIT_3D => X"5D79FCAF774AE005BE7895554005D2A8A0B882FFFFE10AAAAAB755A66B6AF56A",
INIT_3E => X"00000000000000000000000000000000000000C3BC1000FF8409000512AEABFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_3,               -- Port A enable input
WEA      => wbe_a_lo_1024_3(0),               -- Port A write enable input
DIA(0)   => data_write_a(2),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_3(2),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_3,               -- Port B enable input
WEB      => wbe_b_lo_1024_3(0),               -- Port B write enable input
DIB(0)   => data_write_b(2),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_3(2),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_3_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"210C00A20020000108430020001600B8156021104940741B3530400E02B92203",
INIT_01 => X"014C9BCA58B1296D24A402C992500B69404040028804A0080A000416A8D90A08",
INIT_02 => X"C12026A484318004404405C9C66E331352180D468B8203980300204442E02B34",
INIT_03 => X"04000748D60D24648D60524C88804D0215011020D15018148040C10A70E1D58C",
INIT_04 => X"18283333240FE41244187308C9104D70944852640901083801750EB0A418C220",
INIT_05 => X"0613142D01912CC2A1B4140528348900C612A104201C689044340ED413A07649",
INIT_06 => X"119000034019881822104C5E68035250A222829710A0A02C18C01A9920842413",
INIT_07 => X"402F00AB0016CA0431800444841020509D038B021230C1990001C644C8273200",
INIT_08 => X"16905000408482088290E8E64010248C4A5AA840C2000110001521F0810A92E7",
INIT_09 => X"0003CE6581BD016342A951AB146C4480530C3B2A8088D3542651670200C1826A",
INIT_0A => X"00735D36209A8A20020894004284B660821030C8990467401218004041020002",
INIT_0B => X"512445B740457154562F957CC08B00093700080D0A4851001D8302D20A0A1530",
INIT_0C => X"00508650008008021021A40861021840869021A408610218C0869810D6043095",
INIT_0D => X"1C8508438450801043A08090380A8834207007022209038080190000999C8F84",
INIT_0E => X"000400200000C0002A48A206204C4205F3304B33004C0041006240140A1C310A",
INIT_0F => X"0000080040000083800400000100000000008400018040000100080000510100",
INIT_10 => X"0001000000000800000244040000020000000100002A0080000200100000A702",
INIT_11 => X"000000000020000000200000080002C000800008000000000022000006808000",
INIT_12 => X"0000000000000A2281000000000040A3810000000000402001400000022002A0",
INIT_13 => X"000000000004200001C0400000000010200001C0400000000010000004490010",
INIT_14 => X"0001070004000000000000060000104C08000000000000001000000903008000",
INIT_15 => X"CC004050CA0C00020220200070040000010401C4000000000000000000100008",
INIT_16 => X"4310E4310A4210A4210A4210A4210A4210A8D0830A68010001B4DA881048061C",
INIT_17 => X"21084290A4210A4210A4210A4210A4210A4210A4210E4310E4310E4310E4310E",
INIT_18 => X"90A421084290A421084390E4310C4390E4310C4390E4310C4290A421084290A4",
INIT_19 => X"015303C0C78C706428A14C586291000A044001FFE000003FFC004290A4210842",
INIT_1A => X"2492492492492492492492492492492492410410410410412821600001249249",
INIT_1B => X"51A8D46A351A8D46A351A8D46A351A8D46A351A9D4EA753A9D4EA753A9D49249",
INIT_1C => X"FFFFFFFFFFFFFFFC00000000000000000000000038F56351A8D46A351A8D46A3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"55AB02055AB0207FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"420000000000000000000000000000000000000000000000007FFFAB57FFFAB5",
INIT_28 => X"A800BAFFAE9554508002AA00AA843DF55FFAA955EFA2D168B55557BEAA000055",
INIT_29 => X"002AB55AAAA955EF005568A00087BE8BFFA2D155410AA8415555087BFFF55A2A",
INIT_2A => X"AAABFF5508003FF555D0002145552ABFEBA007FC21EF007FD75FFAA841541008",
INIT_2B => X"082EBDEAAA2FBEAABA5D7FC0155005168B455D042AB45F7FFD741000042AA10A",
INIT_2C => X"FF7FBEAB55F7AABDEBA5D7FC2010A2D1575FFF7AA975555D2E80145F78415545",
INIT_2D => X"EF5555554AA087BC01FFFFAAAAB55552A954BAFFFFE8B55552EBDE00F7AEAABF",
INIT_2E => X"000082E820BAA2FBEAB5555557DF55A2AEBDF555D2E954BA002EAAABA002A821",
INIT_2F => X"FB7D5D7FEAA3808554203A000000000000000000000000000000000000000000",
INIT_30 => X"1557D1475FAF45BEAA800AAFFAA95578080038A2AA28E3AF55E3A0BA5D7AADB6",
INIT_31 => X"BD55D7BE80004AA1E8E2AB55B6A0925D7085F6AA10087FEABD7AAD57AEBAB68E",
INIT_32 => X"F5D0438140E2FA38B6AEBFF6D1D04AAFFA41040017D5D20B8EAA007FC51C7A2F",
INIT_33 => X"D0A901FFFF801557D1C20B8EAAA2FBE80AA557BE8B6D5D5FFABEF49002FB55FF",
INIT_34 => X"5D20BDE00EBAAA8BC7EBDFEAFEFAB8ABAE925D21C7010EADB525D7FFAE975C75",
INIT_35 => X"F002EADA921420871D74971D24820875C21D5EB8AA8FFF012A954BAFFF5EFB45",
INIT_36 => X"000000000000000000001C24820BAB6FFEFB6D555578F7DB6A0BDF7DEB8E125F",
INIT_37 => X"B55A28408145AAFFFFFFF5D7FEAABA0051400A20000000000000000000000000",
INIT_38 => X"AB55FAD568AA2AFAE975EF555168B55F7AA800BAF7AA955EF00042AAA2A2AEAA",
INIT_39 => X"2AAAA007FD55558A7BD7145FBB8020A35D2ABEF55F7800015F087FEAA00007FE",
INIT_3A => X"968F575D003FF55F7D5420BA5D2ABFEAAF7AE9DFF759A82AEF70800021EF5504",
INIT_3B => X"FFD5145FBAC9755F05040255FFD84175EF55002AAB0A2FFEAABA557BEA3EF057",
INIT_3C => X"82E974AAF7D57DF45552A3FF10AA8429F45A7D5EAF5FFBAEAAA10554155400AA",
INIT_3D => X"FF843FFE77C80825BC052ABFE10550415557085540000005156155FE90A8F5C0",
INIT_3E => X"00000000000000000000000000000000000005500020AAF7FBFFFEF04552ABFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_3,               -- Port A enable input
WEA      => wbe_a_lo_1024_3(0),               -- Port A write enable input
DIA(0)   => data_write_a(3),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_3(3),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_3,               -- Port B enable input
WEB      => wbe_b_lo_1024_3(0),               -- Port B write enable input
DIB(0)   => data_write_b(3),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_3(3),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_4_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A108400020612C80284210081034849800A00030300004833522C82D04A16002",
INIT_01 => X"2043998A1839284D1CA0650E1E504368403008418984014902030806A0D10200",
INIT_02 => X"C120042200000000044441CE01E80F00A49043118680008002000000026208E4",
INIT_03 => X"040001020019200020011209CC0164C060000000690111040144800042F5C403",
INIT_04 => X"7029AF0F81A00010CCA47700CC513CAC0D0B8E02010740E19754080108988021",
INIT_05 => X"02139405007133C0712244CD20F20105D583000020E9892201D304D42A9835E1",
INIT_06 => X"9190440300078002014405D9EE814C0284A883B6D7038AE079059B7800048092",
INIT_07 => X"000100AA0004408000000004840400008D200102503000782000C00C8025C000",
INIT_08 => X"00728A00408403220811991E02120C044058080004000001101121F220000260",
INIT_09 => X"811001E1185B38AD23C3707AD46440818F3CF80EC423CA7D01D123C80200816A",
INIT_0A => X"45810810A01B40216361056D6150F41200280001900439001FD8A00041400000",
INIT_0B => X"11FC88076266E800D605402962A820211500024808010512C40106D222223B14",
INIT_0C => X"0408804116040B02C02C500B0C02C100B0C02C100B0402C300B0401618058611",
INIT_0D => X"040200050200501301208482200D00D0A0408402C4282200A84800009B878680",
INIT_0E => X"00000020000100024AC88300300060090F0D830F00025400300204D018000804",
INIT_0F => X"8000000040000206A2000800000000000000950002E010000000080000588040",
INIT_10 => X"0000000000000808000554000200000000000100006D0020000000100000BB00",
INIT_11 => X"0000400000000000002000001A0002504001000000000000002280000D800800",
INIT_12 => X"0800000000000E2C802000000000408D801000000000408012440000200110A0",
INIT_13 => X"000000000004680003A0040000000010280003800800000000102800000B0000",
INIT_14 => X"000005C0002000000000000620000158000010000000000010A0000B00000200",
INIT_15 => X"C30146200400104002602600400000000294004000000004000000000010001A",
INIT_16 => X"0080200000008020000000802000000080080000004090014134DA101288C6DB",
INIT_17 => X"0802000000000401806010040180601004018060100000802000000080200000",
INIT_18 => X"8060180601004010040080200802000000000000802008020000000000008020",
INIT_19 => X"C0A28A063807E0500014063450404882846FFE000003FFC00000010040100401",
INIT_1A => X"AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA28A28A28A28A2934C8D0CCD145144",
INIT_1B => X"68341A0D068341A0D068341A0D068341A0D068351A8D46A351A8D46A351AAAAA",
INIT_1C => X"FFFFFFFFFFFFFFFC0000000000000000000000001FE32068341A0D068341A0D0",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"408102040810207FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"800AA00000000000000000000000000000000000000000000040810204081020",
INIT_28 => X"168B55557BEAB4500554200000557FE10FFFBEAA10007FD7410FFAA97555082A",
INIT_29 => X"55574105D2A800AA00043FEBA5D7FEAA00007BE8AAAAA843DF55FFAA955EFA2D",
INIT_2A => X"57BC00AAA2FFEAAAAAA8415555087BFFF55A2AA800BAFFAE9555508002AA0000",
INIT_2B => X"A2AA955EF005568A00087BE8BFFA2D17DE1000517FE10AAAAA8AAA002E975455",
INIT_2C => X"FAA8417410A2D140000F7FBC2010A2D157400AAAE974AAAAAA974BA08002AB55",
INIT_2D => X"EFA2AABDEAA087BEAAAAA2FBD54BA080002145552ABFEAA007FC21EF007FD75F",
INIT_2E => X"00055042AB45F7FFD741000042AA10AAAABFF5508003FF55F7D568A00552EA8B",
INIT_2F => X"5400F7A49057D0824850B8000000000000000000000000000000000000000000",
INIT_30 => X"3AF55F7A0925D7AADB6FB7D5D7FEAB7808554203A145178E00FFFBE8A101475D",
INIT_31 => X"A9557D080038AAA145157428492E8008200043FE925571EFA380871C7028A28E",
INIT_32 => X"AEA8A9200249056D4175C5092AAF5FDA38BE8E1557D1475FAF45BEAA800AAFFA",
INIT_33 => X"AA4954281C0E2FB55B6A0925D7085F6AA10087FEABD7AAD57AEBA08517DE00AA",
INIT_34 => X"007FC51C7007BD55D7BE80004AAFEDB42028EBFBC2028BED152438AAA092492A",
INIT_35 => X"AF7DF6AA00412EAABFFAA803DEBA0875EDA80BEF1C743840040017D5520B8EAA",
INIT_36 => X"0000000000000000000041002FB55FFF5D0438140E2FA38B6AEBFF6DBE84AAEB",
INIT_37 => X"A00FFFFEAA105D5155410FF84021EF0800154B20000000000000000000000000",
INIT_38 => X"DEBA0851574B2AAAEAAB55F78400145AAFFFFFEF5D7FEABFF0051400A25D5568",
INIT_39 => X"68B55F7AA800BAF7AA955EF00042AAA25555410BA082E8201000043FE005D517",
INIT_3A => X"568AA200557DE00AAAAAAA000804001FF005575408AA557FEB2FFAE975EF5551",
INIT_3B => X"D1550AAAA8002010F2AC154B25F2ABFF55F7800015F087FEAA00007FEAB55FAD",
INIT_3C => X"800021EF55042AAAA007FD5555087BD6145FAAC000A2A6FBC00BAAAFBC00BAF7",
INIT_3D => X"F7AEBDFF779A82AA43F7FBE8A00082EA8BFFAA843FEBA08517DE00F3F9574B30",
INIT_3E => X"000000000000000000000000000000000000008003FF55F7D5420BA5D2ABFEAA",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_3,               -- Port A enable input
WEA      => wbe_a_lo_1024_3(0),               -- Port A write enable input
DIA(0)   => data_write_a(4),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_3(4),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_3,               -- Port B enable input
WEB      => wbe_b_lo_1024_3(0),               -- Port B write enable input
DIB(0)   => data_write_b(4),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_3(4),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_5_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50DF4A0791B3FCB694379283C81FD996A091832102004A336A20E03C040C002",
INIT_01 => X"805FBDC69830A84D5C6A60000C34C26841280A00084000C8C212892EEAD53235",
INIT_02 => X"3B2026B578918E640A4F01CF8011FF0002080000082CA9998276DF7772C7C80D",
INIT_03 => X"37134108420D700084205702A4008A1D9100002171C0E0051554D93A11F5D140",
INIT_04 => X"8A41A0FC03A56DA000425A819410E3816C086198A388B702A8CA1210844A0C4C",
INIT_05 => X"B1808A062E8BC835F5E84532D708238A282F00A9291224800A2861490343082C",
INIT_06 => X"903FB8483A90581859050424100940825C6184401CDC451B860A6507160C4100",
INIT_07 => X"D26F068BCC96CDF8918E640E96D1A3469D6300E2FFEA27F8E4D23248130E259C",
INIT_08 => X"0BFA82E568442B2A082C0A7E3014250D49DA37A2420619000002AFF48D1222E5",
INIT_09 => X"3F005001E40969289429360416DCD1C46083030604B1CA20C03DF83B0A2C60A5",
INIT_0A => X"14613C71005A10492B888120288F480D58858449026145B3830F449449062B4F",
INIT_0B => X"11AC04934AC648BFD727C031E64170A137D5AA5C3E4B0F8A3C58C34C002290E3",
INIT_0C => X"CA29C6CC50384B6AC6AC86AB31AACA6AB39AAC86AB39AACA6AB3055643559C31",
INIT_0D => X"C673E33CF28F38603855401985228A0614BD30A0A2819852011E5AC2B87F9182",
INIT_0E => X"FF87C002F87A803E460B2516510CA594FF0044FFA4B08BAC4BB2CD0F09CF84E3",
INIT_0F => X"0DFF0F8005F0F5100DFFF5E15D06101C55EB29F1E00BE53FE1F000BE1E802F94",
INIT_10 => X"F12F0380231F17D78FC029FFF58D9A70380230F2FE0017C37FC3E0017C3D005F",
INIT_11 => X"FC7F023C0CA700125C0F8F7E43F1F001BFFE7C69E01804E1E7CCF8FC003FF5F1",
INIT_12 => X"023E00017C1FC1A4BFD82C3081C5BD27BFE30C3081C5BD00C02365D645CEEF5B",
INIT_13 => X"61E0042787F181E9C1EFD8CB8120C5AF41E9C18FD60F0C20666F41E9F009FFFD",
INIT_14 => X"7A7C077FFF404F80005F07F187A7D14BFFC96111C048278DEB074F9930FF9D80",
INIT_15 => X"C064014B8B652E2B3120C81284641D3E8DBF7D636FE860190700132C1F0EFB80",
INIT_16 => X"38CE1384E3384E338CE138CE1384E33C4E3ECE32E128882551349A1CBAA44103",
INIT_17 => X"84E3384E3384E3384E338CE138CE1384E3384E338CE138CE1384E3384E338CE1",
INIT_18 => X"CE138CE138CE138CE1384E3384E3384E3384E338CE138CE138CE138CE1384E33",
INIT_19 => X"F5E5BB4E7F7B9DB7FF3A1B6DB7E8410A8C000000000000000000384E3384E338",
INIT_1A => X"BEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEF9F7CFDFDDCF3CF3D",
INIT_1B => X"BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEFBEF",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000001711C7BBDDEEF77BBDDEEF77",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"FDFFF00000000000000000000000000000000000000000000080000000000000",
INIT_28 => X"FD7410FFAA97410082A800AAAAAE955450055421FFFFFBC0010AAD5574BA557F",
INIT_29 => X"7FD74000055574BA5D7FD7555A2D5575EF55517FF5500557FE10FFFBEAA10007",
INIT_2A => X"0002AABA5D2ABFFFFAA843DF55FFAA955EFA2D168B55557BEAB5500554200000",
INIT_2B => X"5D2A800AA00043FEBA5D7FEAA00007BC00AAAAAEBDF45A28428B45FFD168BFF0",
INIT_2C => X"5080028A00A2FFFDE00F7D57FEBAFF80174BAAAD1555EF555555555005557410",
INIT_2D => X"BA5D2E821FFA2D5554BA557BD75FFAA8415555087BFFF55A2AA800BAFFAE9555",
INIT_2E => X"00000517FE10AAAAA8AAA002E97545557BC00AAA2FFEAAAA082A97545F7D5420",
INIT_2F => X"7010BEDF524AA5571FDFEF000000000000000000000000000000000000000000",
INIT_30 => X"78E00EBFBE8A101475D5400F7A49043D0824850B8A2AE9756D145B401FFFFFFC",
INIT_31 => X"FEAB7D0855420BA1471D74380851524BA5571D757DB6D5525EF555178F6D1451",
INIT_32 => X"8A28B6DEBDF6DBEF1C0A28AAA5524BFFFFA28E3AF55F7A0925D7AADB6FB7D5D7",
INIT_33 => X"5555057D145152428492E8008200043FE925571EFA380871C7028B6AEBDF45B6",
INIT_34 => X"BEAA800AAFFAA9557D080038AAAA2FBF8E10EBD578EAAFF8415482BED1555EF5",
INIT_35 => X"81C209256DFFDF420BA552A821FFB6DF574A85575C55EFBE8E1557D1475FAF45",
INIT_36 => X"0000000000000000000008517DE00AAAEA8A9200249056D4175C50920875FDA3",
INIT_37 => X"5FF5D7BC21EFF7FBD7400F7FBC00BA55557DFF70000000000000000000000000",
INIT_38 => X"01FF5D5568BE7555568A00AAFFEAA105D5155410FF84020AA0800154B2AAAA97",
INIT_39 => X"00145AAFFFFFEF5D7FEABFF0051400A25551554BA0051400BA5551575EFF7D14",
INIT_3A => X"1574B2FFAABFF45FFAAAABFFAAFFFDFFF552EA8AAA55043DFF7AAAEAAB55F784",
INIT_3B => X"8002410FFD5575EF5555421E75555400BA082E8201000043FE005D517DEBA085",
INIT_3C => X"FAE975EF555168B55F7AA800BAF7AA955EF00002AAA2A2FBE8A00A2D16AAAAFF",
INIT_3D => X"0055554088A557FEB25D00021FFFFFFC00BA552A821EFFFFFD74BA5D51575F7F",
INIT_3E => X"000000000000000000000000000000000000000557DE00AAAAAAA000804001FF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_3,               -- Port A enable input
WEA      => wbe_a_lo_1024_3(0),               -- Port A write enable input
DIA(0)   => data_write_a(5),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_3(5),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_3,               -- Port B enable input
WEB      => wbe_b_lo_1024_3(0),               -- Port B write enable input
DIB(0)   => data_write_b(5),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_3(5),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_6_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10800B0061A01002840002C03002818000402322520070B313301C4389B2082",
INIT_01 => X"250041CA3839684D18A160000C52426841000000090800090210080008110200",
INIT_02 => X"0020042080010000044654C0000C008010000000001020900200200002620814",
INIT_03 => X"060881021088200021080200E4000A0891000020610111500104C00000F14400",
INIT_04 => X"0880000100000002000052288144004281C050400100280000C8100000080001",
INIT_05 => X"928080840001100A08009000280201000850E022401400002028214043410820",
INIT_06 => X"10100518090012122100C808049310002040000410A0001400000200120840D2",
INIT_07 => X"000100800004400001000000860408108C22000A502010074120044800040001",
INIT_08 => X"50000040D0C4E2088003FD01C01004044058082004000000000121F020408244",
INIT_09 => X"00BF17E9001205A5204911F814444080400100020000D200DFD16400C2A40AA0",
INIT_0A => X"04611C17849000022862A1596C8B5DF04834948900000100220C244840000880",
INIT_0B => X"03AD0413424E4044D665C070C22602291504400D084915020448114080201000",
INIT_0C => X"5E08864011088B22D22C008B0022C408B1022C208B0822C608B1111600458010",
INIT_0D => X"4251A12CD28A300429688001000800000020280204001000A00804309A002182",
INIT_0E => X"0000000280402400420800000000006200FC10002442042429324294014E8CA7",
INIT_0F => X"A40000000500800840000800000000000002280018001480000000A010100052",
INIT_10 => X"00000000000004C2003000010240000000000000680800290000000140202000",
INIT_11 => X"2000C0000000000000000442000001080001000000000000010C000280001804",
INIT_12 => X"08000000000801C300A010000000156000902000000015101200002800000000",
INIT_13 => X"000000000101800038002408000000094000386028040000000940000ED40000",
INIT_14 => X"0003B000002000000000020180002A24005010000000000023000060C7000A40",
INIT_15 => X"3F0280090321000040A410C28108000160008094000810040000000000002300",
INIT_16 => X"284A5284A728CA5284A528CA728CA52C4A5A0A32A300940101349A0408240818",
INIT_17 => X"9CA1294A329CA5284A728CA7284A5284A728CA5284A528CA728CA5284A728CA7",
INIT_18 => X"CA3294A129CA3294A129CA1294A329CA1294A3294A129CA3294A129CA3294A32",
INIT_19 => X"F5F78BCE7F8FF0F4FA955F7CF7F40A80145D55555556AAAAAAAAA94A329CA129",
INIT_1A => X"8E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E39B6CEDECDDF7DF7D",
INIT_1B => X"F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE38E3",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000001A1A33F9FCFE7F3F9FCFE7F3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"555FF00000000000000000000000000000000000000000000080000000000000",
INIT_28 => X"BC0010AAD5574BA557FFDFFF087BFDF45F7AA974AAAAAA97555F784174BAF7D5",
INIT_29 => X"515555508043FE00F7AA97555A2FBD7410AA8428AAAAAAE955450055421FFFFF",
INIT_2A => X"7D1575EFFFAA9555500557FE10FFFBEAA10007FD7410FFAA97400082A800AA08",
INIT_2B => X"0055574BA5D7FD7555A2D5575EF55517FF55A2AA97400552AAAB45082E80155F",
INIT_2C => X"500554200000003DE10FFD5401FFF7AAA8A10082EAAB45A2FFC2000007FD7400",
INIT_2D => X"10AA803FE105D516AABAFF843FFFFAA843DF55FFAA955EFA2D168B55557BEAB5",
INIT_2E => X"000AAAEBDF45A28428B45FFD168BFF00002AABA5D2ABFFFF087BD5545007BFDE",
INIT_2F => X"256DEB84104BAFFD1525FF000000000000000000000000000000000000000000",
INIT_30 => X"9756D145B401FFFFFFC7010BEDF524AA5571FDFEF1C7BFFF55FFA095482B6A49",
INIT_31 => X"4904380824850381C5B5057D1C003DE28F7A49057DAAF5D2428A2842AAAAA2AE",
INIT_32 => X"2AAFB451C2A8017DE3DF525FFFFA49756D145178E00EBFBE8A101475D5400F7A",
INIT_33 => X"2F1C50381471D74380851524BA5571D757DB6D5525EF555178F6DAAA49542841",
INIT_34 => X"AADB6FB7D5D7FEAB7D0855420BA1C0E3FE00E3DB471EFE3AAAAA00082EA8B6DA",
INIT_35 => X"F1C7BD057D1C71FFE10A28038E1049516AAB8FF8428FEFA28E3AF55F7A0925D7",
INIT_36 => X"00000000000000000000B6AEBDF45B68A28B6DEBDF6DBEF1C0A28AAA5524BFFF",
INIT_37 => X"F55F78017400F780001FFAA84000AAFFD1401E70000000000000000000000000",
INIT_38 => X"20BAAA8428AA2AAAA975FF5D7BC21EFF7FBD7400F7FBC00BA55557DFF7557BFD",
INIT_39 => X"EAA105D5155410FF84020AA0800154B2557FC01EF55043FEAAFF80021EFA2D14",
INIT_3A => X"568BE7AA80174AA082ABDF555D2A821EFAAFBC01FFF780155F7555568A00AAFF",
INIT_3B => X"AEA8A10082EA8BEFAAD5554B25551554BA0051400BA5551575EFF7D1401FF5D5",
INIT_3C => X"AAEAAB55F78400145AAFFFFFEF5D7FEABFF0051400A25D2EBFE10AAFFD55EFA2",
INIT_3D => X"552EA8AAA55043DFF7557BC01EF55557DE00AA842AA0000516AABAFF8428BE7A",
INIT_3E => X"0000000000000000000000000000000000000FFAABFF45FFAAAABFFAAFFFDFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_3,               -- Port A enable input
WEA      => wbe_a_lo_1024_3(0),               -- Port A write enable input
DIA(0)   => data_write_a(6),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_3(6),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_3,               -- Port B enable input
WEB      => wbe_b_lo_1024_3(0),               -- Port B write enable input
DIB(0)   => data_write_b(6),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_3(6),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_7_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10844B00482258A2842112C02450418800002300500030B313300C418992002",
INIT_01 => X"000009CA3839684D1CA0E0000E51424840000000080000080200080008510204",
INIT_02 => X"0120042086010000044600C00008000004100000000260900200000002402004",
INIT_03 => X"8628A10000082400000002408400080011000000610008000208C00000E14400",
INIT_04 => X"0911800100A000000000524084000040000050001140200100C8100000080102",
INIT_05 => X"0300812401011000000000002000114008008060441000000020024093000000",
INIT_06 => X"9190431C0D4010100000880804010010800000041080081000000200010424B2",
INIT_07 => X"000100AA0004408601000004860000008C02000A103010006928040800062481",
INIT_08 => X"84000048D484C20888000A0002120484C048007004000000000021F000000244",
INIT_09 => X"00A06009881201A520491004106C48A04040002400A15A208001650004001020",
INIT_0A => X"C99E1060201002044809C1040140A001004808810000459033189C0A400118A0",
INIT_0B => X"102000024040484050050041648A0041140C500B08821054C000264120000400",
INIT_0C => X"0404A083260E0832132011880462011880462051881462051881D31018C40620",
INIT_0D => X"0001000080001000813094801A8F80F00A600B52602801A88848011118003700",
INIT_0E => X"000003C007C002808228010410082042C000C000000004001002000400040002",
INIT_0F => X"A4000007800F80C840000800009864038A1200081C0014800000F001F0200052",
INIT_10 => X"00002C0E00E0E4004038000102400002C0E00E0D20100029000001E003E04000",
INIT_11 => X"2000C04031100E0403D0700300080908000100000661801E1900040380001804",
INIT_12 => X"0840878083E8003780A01043203A101780902043203A10082410082880000000",
INIT_13 => X"0601E0187900181035E0240806483248181035E0280410C8198818100DDD0000",
INIT_14 => X"0403774000201021E020FA006040376C00501022131210722060806D47000A40",
INIT_15 => X"00928A0002000110888600C032128201519480D40009902430160403E0E00506",
INIT_16 => X"01000000020080601802000000000405000A0020020081014134928820480010",
INIT_17 => X"0802018040000000006018020080200804010000000000806018020080000004",
INIT_18 => X"0000000001806008020000001006008020080001004008020080201004000020",
INIT_19 => X"0000000000000000000000000000400A004618618618C30C30C3000020180600",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000000B0840000000000000000000",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"1555500000000000000000000000000000000000000000000080000000000000",
INIT_28 => X"A97555F784174BAF7D5555FFF780155EFAAAEA8ABAAAFBFDE0055556AA005D04",
INIT_29 => X"55555EFAAFFFDFEFAAAAAAB455D556AA00FFAE95555087BFDF45F7AA974AAAAA",
INIT_2A => X"02EAAAAA082EA8A00AAAE955450055421FFFFFBC0010AAD5574BA557FFDFFF55",
INIT_2B => X"08043FE00F7AA97555A2FBD7410AA8428AAA557BFDFFF55003DFFFF7FBEAA000",
INIT_2C => X"0082A800AAF7AE975FFA28000010552EBDE00007BEAAAAA2D140000085155555",
INIT_2D => X"45087FEAB455D516AB55557BD55FF00557FE10FFFBEAA10007FD7410FFAA9740",
INIT_2E => X"000A2AA97400552AAAB45082E80155F7D1575EFFFAA955555D51574AAAAFFD55",
INIT_2F => X"AE105D556AA10410E17555000000000000000000000000000000000000000000",
INIT_30 => X"FFF55FFA095482B6A49256DEB84104BAFFD1525FFFF8E175C7A2AAAAA82A2F1F",
INIT_31 => X"F524AA5571FDFEF415B575D7AAF1FFFD7AAAAAFB7D495F6AA10E3AE905551C7B",
INIT_32 => X"003AFEFEBFBEAA001C2EA8A821C2EAAA00A2AE9756D145B401FFFFFFC7010BED",
INIT_33 => X"EDB470101C5B5057D1C003DE28F7A49057DAAF5D2428A2842AAAA497BFAFFF49",
INIT_34 => X"1475D5400F7A490438082485038F7A4905C7A28A070384120BDE100075EAA82B",
INIT_35 => X"D495150492BEF1D2555087BE8B7D555F6AB57417BC05D7145178E00EBFBE8A10",
INIT_36 => X"00000000000000000000AAA495428412AAFB451C2A8017DE3DF525FFFFA49756",
INIT_37 => X"555A2AEA8A10AAD568A00555168A10002E9754D0000000000000000000000000",
INIT_38 => X"8A10AAAE8215D557BFDF55F78017400F780001FFAA84000AAFFD1401E7FFAA97",
INIT_39 => X"C21EFF7FBD7400F7FBC00BA55557DFF7007BD5555AAD57DF55AAAEBDFEF007BE",
INIT_3A => X"428AA2007FE8BFF080028BFFAAFFEAA105D2EAAA005D2AAAA18AAAA975FF5D7B",
INIT_3B => X"043DE0000516AA10F7FBD7408557FC01EF55043FEAAFF80021EFA2D1420BAAA8",
INIT_3C => X"55568A00AAFFEAA105D5155410FF84020AA0800154B2FF8402145A2AA954AA00",
INIT_3D => X"AAFBC01FFF780155F7005140000FFD140145007FE8BEF557BEAB55087FC215D5",
INIT_3E => X"0000000000000000000000000000000000000AA80174AA082ABDF555D2A821EF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_3,               -- Port A enable input
WEA      => wbe_a_lo_1024_3(0),               -- Port A write enable input
DIA(0)   => data_write_a(7),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_3(7),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_3,               -- Port B enable input
WEB      => wbe_b_lo_1024_3(0),               -- Port B write enable input
DIB(0)   => data_write_b(7),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_3(7),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_8_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00000648E2840112C00000418000002700500030B3132000400812082",
INIT_01 => X"100008480009004C04A100000252024840000000180800080200010040110204",
INIT_02 => X"0020042000490000004600804008000005100000000024900200000002400004",
INIT_03 => X"0A0C33400008082400000080A4004B0891000020610112000040C00000E5C000",
INIT_04 => X"18800001000000000000512080000040800150400824280110C8100000120200",
INIT_05 => X"908084A10100100200004080280008240810802206940000012C214451610800",
INIT_06 => X"81B000080860109021400008040000202048020414A0021400040200322824C1",
INIT_07 => X"000000080004408049000004860000008402001A50208000630C040800062483",
INIT_08 => X"440000428644212280800A00021004044048002124000000000021F000000244",
INIT_09 => X"00004009001001010008100414644410400102228000D20080114502006409A2",
INIT_0A => X"000051312000042200294429148A4801C80C8C81000045907118040340020832",
INIT_0B => X"4020000240404140004D0544C4AA0001150410090302500011C813428A000400",
INIT_0C => X"46501090008820240240409000240009000240009000240009000120204808A5",
INIT_0D => X"42D1A168D09A301468402480004780F00140080860280004085904309A002196",
INIT_0E => X"00783FC00044340242280000000000020000C0000442106419120004034685A3",
INIT_0F => X"8000F07F800088A80000081EA2F9EC0000064004081010001E0FF00011104040",
INIT_10 => X"0ED0FC7E00000422201080000202658FC7E0000021882020003C1FE000222080",
INIT_11 => X"018059C3F350FE0C00000002A0040500000103961FE780000110010090000800",
INIT_12 => X"FD41FF80000830200021C1CF600012200010D1CF600012121600100810000004",
INIT_13 => X"9E1FE000010A1802100004343ED8000898021000087073D80008980200800002",
INIT_14 => X"0080200000BEB07FE00002086008020000209AEE3F300000246020200000620B",
INIT_15 => X"0088881903210000440610C8000A808040000208901786E4F0FE0C0000000166",
INIT_16 => X"685A1685A769DA368DA368DA769DA36CDA121A11A141800011309284002C0810",
INIT_17 => X"95A5685A1685A5695A368DA368DA769DA368DA368DA7695A1685A1685A5695A1",
INIT_18 => X"5A1695A568DA368DA369DA768DA1685A1695A5685A168DA369DA768DA368DA16",
INIT_19 => X"A4028A0A543EBC57A10A1E75D64108080468618618630C30C30C69DA5685A168",
INIT_1A => X"9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7BF3CCD8DF5B2DB2C",
INIT_1B => X"F87D3E1F4F87D3E1F4F87D3E1F4F87D3E1F4F87C3E1F0F87C3E1F0F87C3E79E7",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000006A6D4F87D3E1F4F87D3E1F4",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"155FF00000000000000000000000000000000000000000000080000000000000",
INIT_28 => X"BFDE0055556AA005D0415555080000000087BEAA10F7803DE00FFAEBFFFF0800",
INIT_29 => X"2AA8AAA557FC0010F780154105D7FC2145005155555F780155EFAAAEA8ABAAAF",
INIT_2A => X"7FFFFF55AA80155FF087BFDF45F7AA974AAAAAA97555F784174BAF7D5555FF55",
INIT_2B => X"AAFFFDFEFAAAAAAB455D556AA00FFAE95555AAFFE8A00552EBFE00F7D17FF45F",
INIT_2C => X"A557FFDFFF5504000AAAAAAA8B55F7D140010552E821EFAAAABDF555555555EF",
INIT_2D => X"55AA8028A00A2D57FF45557BE8A00AAAE955450055421FFFFFBC0010AAD5574B",
INIT_2E => X"000557BFDFFF55003DFFFF7FBEAA00002EAAAAA082EA8A00002AA8A10F784021",
INIT_2F => X"FE10F7AEBAFFF080A175D7000000000000000000000000000000000000000000",
INIT_30 => X"175C7A2AAAAA82A2F1FAE105D556AA10410E17555080E000280071E8A00EB8E3",
INIT_31 => X"4104BAFFD1525FF492EA8AAA5571C2000FF8A17400557FC015514555757DFF8E",
INIT_32 => X"2ABDE10EBDF7AF6DE3FFF8F7DB68A105D71C7BFFF55FFA095482B6A49256DEB8",
INIT_33 => X"AA0BDF6D415B575D7AAF1FFFD7AAAAAFB7D495F6AA10E3AE90555A2FBE8A3849",
INIT_34 => X"FFFFC7010BEDF524AA5571FDFEF550E00082B6A0AFB55F7D1420104124821D7A",
INIT_35 => X"01C2EA8A00F7800017DA2842FA00B6D578F6D557FFDA00A2AE9756D145B401FF",
INIT_36 => X"00000000000000000000497BFAFFF49003AFEFEBFBEAA001C2EA8A821C2EAAA0",
INIT_37 => X"0BA08556AA00AAAABFE00F7AEAABEF082E955450000000000000000000000000",
INIT_38 => X"21555D51575EFFFAA97555A2AEA8A10AAD568A00555168A10002E9754D082E82",
INIT_39 => X"17400F780001FFAA84000AAFFD1401E7082EAAABA5D5140010F7AE974105D7BC",
INIT_3A => X"E8215DA2FFE8ABA082ABFE00AAFBEABFFAAFBEABFFF7AA80145557BFDF55F780",
INIT_3B => X"D540000000402145AA843FFFF007BD5555AAD57DF55AAAEBDFEF007BE8A10AAA",
INIT_3C => X"AAA975FF5D7BC21EFF7FBD7400F7FBC00BA55557DFF75D2E82010F7843DF45FF",
INIT_3D => X"5D2EAAA005D2AAAA185D2AAAA10F780021FFA2803DE10FFD16ABFF5D7BFDE10A",
INIT_3E => X"0000000000000000000000000000000000000007FE8BFF080028BFFAAFFEAA10",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_3,               -- Port A enable input
WEA      => wbe_a_lo_1024_3(1),               -- Port A write enable input
DIA(0)   => data_write_a(8),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_3(8),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_3,               -- Port B enable input
WEB      => wbe_b_lo_1024_3(1),               -- Port B write enable input
DIB(0)   => data_write_b(8),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_3(8),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_9_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00018248A2840112C00002C18000002300500030B3132000400812006",
INIT_01 => X"400008000000004C0020000000100248413C0A61590001D90213C10008110204",
INIT_02 => X"01A0042080010000054600C04008000004100000001020900200200002420804",
INIT_03 => X"024003400008012400000010E4004B0891000020610310000144C00000F5C000",
INIT_04 => X"1801800100E000000000510084000040010050020810200000C8900000320200",
INIT_05 => X"918004311104100000000000200008100800002000100000002C234415610820",
INIT_06 => X"81B00008080010100000980804000008800042041080001000100200322C2481",
INIT_07 => X"0000811800044080010000058600000086020002502080006000040800062C80",
INIT_08 => X"0000004001D4618008800A00061004044048002004000000000061F000000244",
INIT_09 => X"000040090802009420409004104444084001022400214A2080014400026401A2",
INIT_0A => X"04000071200000A003CA294140200800C80C8C8100004590111C040040120800",
INIT_0B => X"12210002404848502847040164880021150400080222000200C8034200000000",
INIT_0C => X"4610088010080421021040841021000841021000841021000841010800420820",
INIT_0D => X"42D0A16C529A321068500484000500D10042080040284000084900001A002196",
INIT_0E => X"00000002804000004228010410082002C000C0002400046419120410034285A1",
INIT_0F => X"A00000000500800800000800000000000002290008001080000000A010100042",
INIT_10 => X"00000000000004C2001000000240000000000000680800280000000140202000",
INIT_11 => X"0000C0000000000000000442020001000001000000000000010C800080000804",
INIT_12 => X"08000000000801A7802010000000152780102000000015000600000800000000",
INIT_13 => X"000000000101900011E0240000000009500011E0280000000009500004DD0000",
INIT_14 => X"000137400020000000000201C000136C00101000000000002340002947000240",
INIT_15 => X"0080881901210000000600C280028000419480D4000010040000000000002304",
INIT_16 => X"68DA368DA1685A1685A1685A1685A16C5A121A13A141950051309284A82C0010",
INIT_17 => X"85A1685A1685A1685A368DA368DA368DA368DA368DA368DA368DA368DA368DA3",
INIT_18 => X"5A1685A168DA368DA368DA368DA368DA368DA368DA3685A1685A1685A1685A16",
INIT_19 => X"0157344CCCF48DE68A895C38E2540A8010100000000000000000685A1685A168",
INIT_1A => X"14514514514514514514514514514514514D34D34D34D34D28E1004039248209",
INIT_1B => X"D268341A4D268341A0D069349A0D069349A0D068341A0D068341A0D068345145",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000014D490D069349A0D068341A4",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"EAABA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"03DE00FFAEBFFFF0800155FFAAFBE8B45002A974AAAA803DFFFAA843DF45FFFF",
INIT_29 => X"7BFDE00A2FBD7400F7FBFDFFFA2AEBDE00AAFBEAABA080000000087BEAA10F78",
INIT_2A => X"055401FFF7AEAAA10F780155EFAAAEA8ABAAAFBFDE0055556AA005D041555508",
INIT_2B => X"557FC0010F780154105D7FC2145005155555557BE8BEF007FFDEAAAAD1555EF0",
INIT_2C => X"AF7D5555FFF780154AA5D2AA8A10F7AA974AA082E80010A2AAAAA10552AA8AAA",
INIT_2D => X"BAF7D17FEBAA2AEBDF45002EAAABA087BFDF45F7AA974AAAAAA97555F784174B",
INIT_2E => X"000AAFFE8A00552EBFE00F7D17FF45F7FFFFF55AA80155FF080400145FFFBEAA",
INIT_2F => X"8FC7BE8A3DF7DF7F5E8A92000000000000000000000000000000000000000000",
INIT_30 => X"000280071E8A00EB8E3FE10F7AEBAFFF080A175D7BEF1E8B6D002090482B68E3",
INIT_31 => X"56AA10410E175550871FFE00A2FBD0400FFF5FDFC7B6A0BDE38B6F5E8A92080E",
INIT_32 => X"7BFAE82A2DB555C71C5B451D7FFAAA8A38FF8E175C7A2AAAAA82A2F1FAE105D5",
INIT_33 => X"2AEADA38492EA8AAA5571C2000FF8A17400557FC015514555757D5D71E8BEF14",
INIT_34 => X"B6A49256DEB84104BAFFD1525FFFF84174BA5D20AAA00E3AA904BA142A87010A",
INIT_35 => X"7000400155FFFBEDA82FFD57DEBAAAA0BFF7D0024ADA921C7BFFF55FFA095482",
INIT_36 => X"00000000000000000000A2FBE8A38492ABDE10EBDF7AF6DE3FFF8F7DB68A105D",
INIT_37 => X"BEF080402000F7AAA8B55FFAABDFEFF7D16AA000000000000000000000000000",
INIT_38 => X"FEAAFFD16AA00082E820BA08556AA00AAAABFE00F7AEAABEF082E95545F7D568",
INIT_39 => X"A8A10AAD568A00555168A10002E9754D00517DE00A2FFC2000F7D17FF55FF803",
INIT_3A => X"1575EF555568BEF5D7FE8A10AAFFD55555D7FD5555FFAAA8AAAFFAA97555A2AE",
INIT_3B => X"AE800AA552A97400A2AEBDEAA082EAAABA5D5140010F7AE974105D7BC21555D5",
INIT_3C => X"57BFDF55F78017400F780001FFAA84000AAFFD1401E7FF80174AA5D0028A00AA",
INIT_3D => X"AAFBEABFFF7AA80145080002145F7FBFFE00FFD17FEAAA2803DFEF08043FE005",
INIT_3E => X"0000000000000000000000000000000000000A2FFE8ABA082ABFE00AAFBEABFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_3,               -- Port A enable input
WEA      => wbe_a_lo_1024_3(1),               -- Port A write enable input
DIA(0)   => data_write_a(9),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_3(9),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_3,               -- Port B enable input
WEB      => wbe_b_lo_1024_3(1),               -- Port B write enable input
DIB(0)   => data_write_b(9),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_3(9),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_10_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00018248A2840112C00002C18000202300500030B3132000400992006",
INIT_01 => X"254008000000004C002000000010026840000000080000080200010008110204",
INIT_02 => X"0020042000010000004455800008000004100000000000900200000002400004",
INIT_03 => X"020001021089000021081000C400090011000000610001540104C00000F14400",
INIT_04 => X"0811800101A00002000050088554004200C840000000200080C8100000000001",
INIT_05 => X"030080001000100800009400200000000840E020201000000024024001200020",
INIT_06 => X"81B00008080012120004CC080492500280208004148000100000020020042493",
INIT_07 => X"0000000800044080010000048404081085020002502000006000040800062480",
INIT_08 => X"100202400084410808000A00021004044048000004000000000021F020408264",
INIT_09 => X"010040090002008420401004144440004040022484214A2080110108C2C00320",
INIT_0A => X"04004166A48A0001080000000000080080181881000045901118044040020800",
INIT_0B => X"1201000200484910000F0105602622291404020902005002018002400A022000",
INIT_0C => X"0440001011808020120004801120044800120004801120044800110002400884",
INIT_0D => X"008000440210100041308480800F82F00040180260A808008848000018002104",
INIT_0E => X"000000028040000002280104100820020000400020000440100204100A000100",
INIT_0F => X"040000000500800800000000000000000002280008000400000000A010100010",
INIT_10 => X"00000000000004C2001000010000000000000000680800010000000140202000",
INIT_11 => X"200000000000000000000442000001000000000000000000010C000080001000",
INIT_12 => X"00000000000801C0008000000000154000800000000015000410000800000000",
INIT_13 => X"0000000001019800180000080000000958001800000400000009580002800000",
INIT_14 => X"0000A0000000000000000201E0000A0000400000000000002360002080000800",
INIT_15 => X"0080881000000000000600C28102800060000000000800000000000000002306",
INIT_16 => X"401004010040100401004010040100441020D0030008840051309A90BA884010",
INIT_17 => X"0902409024090240900401004010040100401004010040100401004010040100",
INIT_18 => X"1004010040902409024090240902409024090240902409024090240902409024",
INIT_19 => X"F546890A940FE0D3971243555205428290100000000000000000401004010040",
INIT_1A => X"8A28A28A28A28A28A28A28A28A28A28A28A28A28A28A28A29554199854514514",
INIT_1B => X"2B95CAE532994CA6532995CAE572B94CA6532994CA6532994CA6532994CA28A2",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000002718E72B94CA6532994CA657",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"FDE1000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"03DFFFAA843DF45FFFFEAABA007FC2155F7D155545AA80001EFAAFBEAB45557F",
INIT_29 => X"042AB55FFD168B55AA8000010FFFBE8BFFF78402155AAFBE8B45002A974AAAA8",
INIT_2A => X"AD16AABA002ABDE10080000000087BEAA10F7803DE00FFAEBFFFF0800155FF00",
INIT_2B => X"A2FBD7400F7FBFDFFFA2AEBDE00AAFBEAABAA2FFD741055003DFEFF7AA801FFA",
INIT_2C => X"05D0415555007FD74105555555EFF7FBC0145F78028A00A2D142155087BFDE00",
INIT_2D => X"55AAD168ABA002A975FFF7AEBDEBAF780155EFAAAEA8ABAAAFBFDE0055556AA0",
INIT_2E => X"000557BE8BEF007FFDEAAAAD1555EF0055401FFF7AEAAA105D042ABFF5D556AB",
INIT_2F => X"71D7AAFBEFB455D71F8E00000000000000000000000000000000000000000000",
INIT_30 => X"E8B6D002090482B68E38FC7BE8A3DF7DF7F5E8A92007BC217DEBDB55555AA8E0",
INIT_31 => X"EBAFFF080A175D700042AB7DEBDB6DB55BE8E05000EBFFE8BC7E38E07145BEF1",
INIT_32 => X"0A3DFD7F7A4821D7A2D16FA82142EB8E00080E000280071E8A00EB8E3FE10F7A",
INIT_33 => X"ED1421450871FFE00A2FBD0400FFF5FDFC7B6A0BDE38B6F5E8A92B6FBD541049",
INIT_34 => X"A2F1FAE105D556AA10410E175550071D54104951555D7EBF5C5155E3842AA00B",
INIT_35 => X"8410E2ABD749516FB55BED16FA820820955EFE3AEBDEAAFF8E175C7A2AAAAA82",
INIT_36 => X"000000000000000000005D71E8BEF147BFAE82A2DB555C71C5B451D7FFAAA8A3",
INIT_37 => X"1EFA2FFD7545AAAE97555A2FBFDF455D556AA000000000000000000000000000",
INIT_38 => X"8B45AAAA95545F7D568BEF080402000F7AAA8B55FFAABDFEFF7D16AA00087FC0",
INIT_39 => X"6AA00AAAABFE00F7AEAABEF082E9554500042ABFFA2FFFFF45F7AE97400AAFFE",
INIT_3A => X"16AA00FFFBD5400082EBFF45F78400155A2D57FE00552EA8A00082E820BA0855",
INIT_3B => X"D557555A2802AA10FFD54214500517DE00A2FFC2000F7D17FF55FF803FEAAFFD",
INIT_3C => X"FAA97555A2AEA8A10AAD568A00555168A10002E9754D085155410085557555AA",
INIT_3D => X"5D7FD5555FFAAA8AAA002AAAB4508557DF55F7D17FE000804155FFAAAABDEAAF",
INIT_3E => X"0000000000000000000000000000000000000555568BEF5D7FE8A10AAFFD5555",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_3,               -- Port A enable input
WEA      => wbe_a_lo_1024_3(1),               -- Port A write enable input
DIA(0)   => data_write_a(10),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_3(10),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_3,               -- Port B enable input
WEB      => wbe_b_lo_1024_3(1),               -- Port B write enable input
DIB(0)   => data_write_b(10),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_3(10),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_11_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A101C4B05A0034CA2840712C2D001419000002300500030B31B20084EC992002",
INIT_01 => X"90000986B83028491800E0000C26426040000000080000088200080802512224",
INIT_02 => X"1A2004205E010640024D00800008000004100000040EC090820018003241A00C",
INIT_03 => X"28639100000C5C00000045C08400C8001100000061806A001618C03001E54400",
INIT_04 => X"1A800001000009A0804059A190000040400040008058220008C8100000120D4E",
INIT_05 => X"02000E81080250010000002022000058080400000E1200000020004401000004",
INIT_06 => X"819435143F20101010001008040800B8100102041088011100022200000024B2",
INIT_07 => X"90640D280884453E01064002944180008402001295BA100022E4340800062D82",
INIT_08 => X"400000093204802200280A0012160585C1D808D004000000000323F40C102244",
INIT_09 => X"380040098010001100009204107C5950400000220080C200800900020C006827",
INIT_0A => X"80007100004016EA080801010000080D00200081000045B0511D289940103399",
INIT_0B => X"002000024040410A000D0104408810C115D9C008050042400100D04E88000002",
INIT_0C => X"00655010009264201200C7B421ED0C7B421ED0C7B431ED087B43176843DA1085",
INIT_0D => X"0401020080400A10012494881A4F80F209500BB2602881A488485C1318002000",
INIT_0E => X"6619A540124814800228010410082022C00040002020090020220C9600040802",
INIT_0F => X"ACCC334A802491600C587949B6D0141B4CC600D5761B1599865A500490B86A56",
INIT_10 => X"BAC845542056A61686EC81E3A6CB68AA2C622C9A251C352B330CB4A0092170D8",
INIT_11 => X"BCCAD0B5A81536080CC6B21A21B1FC09CB0F1076D4A200B2AD4068F4101639B5",
INIT_12 => X"4D2CC281E31AA0103AB8D5514066380804B268A2E060901204112566F10AC418",
INIT_13 => X"D551443C47281002540B2C9AAAA8662A1152B202AE3554403028115AA88201A1",
INIT_14 => X"548A20A0492A2724A0621620402A020141F172FB182A32AB6845AB6200251BC9",
INIT_15 => X"00C00A000200074044E6801832728080D00A380B753952C4877E0104DDE4D124",
INIT_16 => X"0080200802008020080200802008020480080022020081010124988800400010",
INIT_17 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_18 => X"0000000000802008020080200802008020080200802008020080200802008020",
INIT_19 => X"55062608804180C0B10A42104201400204000000000000000000000000000000",
INIT_1A => X"00000000000000000000000000000000000820820820820801C4149470000000",
INIT_1B => X"0000000000000000040200000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000007E0F0000000000000100800",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"000AA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0001EFAAFBEAB45557FFDE10082ABDF5508557DF45002ABDFFFF7803DE10AA80",
INIT_29 => X"AEBFF45FFAEBFEAA002A801FFF7FFE8A10A28000000007FC2155F7D155545AA8",
INIT_2A => X"2AABFE10082ABFFEFAAFBE8B45002A974AAAA803DFFFAA843DF45FFFFEAABAA2",
INIT_2B => X"FFD168B55AA8000010FFFBE8BFFF78402155AAD155555A28428BFF002ABDE00A",
INIT_2C => X"F0800155FF00557FF45557FC2010002A80010A2842AAAA007BFFF4500042AB55",
INIT_2D => X"FF5D00154BAF7FBE8BEFFFD540000080000000087BEAA10F7803DE00FFAEBFFF",
INIT_2E => X"000A2FFD741055003DFEFF7AA801FFAAD16AABA002ABDE10A2D168A10A284021",
INIT_2F => X"DFC7F78E3FE28B684070AA000000000000000000000000000000000000000000",
INIT_30 => X"C217DEBDB55555AA8E071D7AAFBEFB455D71F8E00002EBDF6D005B78F7D142AB",
INIT_31 => X"A3DF7DF7F5E8A92BEAEBFF7DEBA0BDEAA1C2A801C7E3FFEFA10B68407038007B",
INIT_32 => X"8A28BFF082ABAE10B6AAB8E280820B8FEFBEF1E8B6D002090482B68E38FC7BE8",
INIT_33 => X"07FF8F7D00042AB7DEBDB6DB55BE8E05000EBFFE8BC7E38E07145B6D15756DA2",
INIT_34 => X"EB8E3FE10F7AEBAFFF080A175D708517DF7D497BC5028142A87000A28A2AA920",
INIT_35 => X"0B6DB6AA28A280001FF5D0A10482FFFFEFBC7E3DF42028080E000280071E8A00",
INIT_36 => X"00000000000000000000B6FBD5410490A3DFD7F7A4821D7A2D16FA82142EB8E0",
INIT_37 => X"FEF007BE8BFF5D2ABDF55F7AABDEAAF784154BA0000000000000000000000000",
INIT_38 => X"DE00FF84154BA087FC01EFA2FFD7545AAAE97555A2FBFDF455D556AA00082EBF",
INIT_39 => X"02000F7AAA8B55FFAABDFEFF7D16AA00FFAEBFFEFAA803DEBA5D2E82155A2FBF",
INIT_3A => X"A95545F7D5555FFAAAAA8BFF002AAAA00FFAAA8AAA080028BFFF7D568BEF0804",
INIT_3B => X"2E95400A2AEA8A00007FEABFF00042ABFFA2FFFFF45F7AE97400AAFFE8B45AAA",
INIT_3C => X"82E820BA08556AA00AAAABFE00F7AEAABEF082E9554508557DFFF007BD54BA5D",
INIT_3D => X"A2D57FE00552EA8A00FFFFE8AAAAA80001FF5D2E82000F7FFFFF45AAFFC20BA0",
INIT_3E => X"0000000000000000000000000000000000000FFFBD5400082EBFF45F78400155",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_3,               -- Port A enable input
WEA      => wbe_a_lo_1024_3(1),               -- Port A write enable input
DIA(0)   => data_write_a(11),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_3(11),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_3,               -- Port B enable input
WEB      => wbe_b_lo_1024_3(1),               -- Port B write enable input
DIB(0)   => data_write_b(11),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_3(11),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_12_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50080B01BC002006940202C0DE041196A83183000000023322287E0FC000006",
INIT_01 => X"75400D849830C84C5823E0000C17424840000000080000088200002802153231",
INIT_02 => X"18A026B43ED180040147558040090000061800000C06ED9802768F4472C52005",
INIT_03 => X"2A67E34A528D0524A52850528400C8001100000171C02B550618C91A10E55440",
INIT_04 => X"1BC0000100056C8280825DE98154004300C840800850240080CA921084520A07",
INIT_05 => X"02000F832000500C0000941024000852084060202E100001002000448100000C",
INIT_06 => X"819A1D1C3FE01A1A40045408049A50BA4020C6041090001200006200000000F2",
INIT_07 => X"C26A0719CC96CC6ED18A64019695A854870300FA3968B20068FC06080106249F",
INIT_08 => X"D002024B3E040800008C0A002610240D494A06F3460409000000E3F0AD5282E5",
INIT_09 => X"27A06009200040000400120412445D78400001000410420080218029CC807A27",
INIT_0A => X"18000006848A026F000000000000080000F010C100204593F11A6CDF48003BF8",
INIT_0B => X"000000820040402B28050400400432C9349DF21A31A00ACC0000F04F80020001",
INIT_0C => X"00357804611AE45D05D0833430CD0833420CD0C33420CD0833430668619A1000",
INIT_0D => X"0000000000000A74812DF00E87E80A079F9F90FA0280E87E800C7FF3B8002000",
INIT_0E => X"3B6B0E404D26160682082002000401EA0000C40000800A006002818808000000",
INIT_0F => X"A476D61C809A4DA84272592D6246FC1B17B541F97E1B348EDA93900B2B286C56",
INIT_10 => X"30C669E622DBC325CFD881A962454CFBE5403AB99594362B1DB52720165650D9",
INIT_11 => X"F8D2D39A3745261E4A95A110A3F855000E4B1D32BAB504BB7490FCFF912A3834",
INIT_12 => X"B90E9B018C7530200AB8F8BF41F9A22006B37DC8E1F9A21A70116D4C5080651C",
INIT_13 => X"118780319CCA08AB1001ACDF34B8F1C688AB1002AE3F7B807B6289F368828C4C",
INIT_14 => X"2AF020233376A5ECC016B1A827CDA21160F051DE610A34C50427E6E220323E4A",
INIT_15 => X"0077020000000439FDC05C5806781FAB46095A0B5199B0AC55521524F1864022",
INIT_16 => X"000000000000000000000000000000000026C000002884000130921092804010",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"8020080200000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0051B946088881360A95090CB054420290100000000000000000008020080200",
INIT_1A => X"041041041041041041041041041041041049249249249249200100002D451451",
INIT_1B => X"92C964B2592C964B2592C964B2592C964B2592C86432190C86432190C8641041",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000003800F592C964B2592C964B25",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"7DE1000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"ABDFFFF7803DE10AA80000AAAA843FE0008557DFFF0800020105D557FEAA0055",
INIT_29 => X"D5420000051555FFA2AA8200000557DFFFF7AA80000082ABDF5508557DF45002",
INIT_2A => X"82AA8AAAAAFFC00BA007FC2155F7D155545AA80001EFAAFBEAB45557FFDE10AA",
INIT_2B => X"FFAEBFEAA002A801FFF7FFE8A10A28000000A2D155410F7FFFFEBA08003FE000",
INIT_2C => X"5FFFFEAABA000028A105D2ABFE10A2AABFE1055516ABEF5D517DEAAA2AEBFF45",
INIT_2D => X"55002A820AA08557DFFFF7AA82155AAFBE8B45002A974AAAA803DFFFAA843DF4",
INIT_2E => X"000AAD155555A28428BFF002ABDE00A2AABFE10082ABFFEF0855420000004175",
INIT_2F => X"5010495B7AE921C517DE10000000000000000000000000000000000000000000",
INIT_30 => X"BDF6D005B78F7D142ABDFC7F78E3FE28B684070AABE803AE38145B78FD700000",
INIT_31 => X"BEFB455D71F8E00BED547038145B505FFB6A487000005F7AFD7F7A482038002E",
INIT_32 => X"F1FDE821C003FE001C2EAAAAAB6F5C2082007BC217DEBDB55555AA8E071D7AAF",
INIT_33 => X"D517DEAABEAEBFF7DEBA0BDEAA1C2A801C7E3FFEFA10B68407038B6D550428FF",
INIT_34 => X"B68E38FC7BE8A3DF7DF7F5E8A9200002FA285D20BDE28A2A4B8E10555B68BEF5",
INIT_35 => X"F085F47038140010555142082082005F7DFD7F7A482155BEF1E8B6D002090482",
INIT_36 => X"00000000000000000000B6D15756DA28A28BFF082ABAE10B6AAB8E280820B8FE",
INIT_37 => X"ABA5D7FEAB45080015410007FEAA0055517DE000000000000000000000000000",
INIT_38 => X"AB45F780020BA082EBFFEF007BE8BFF5D2ABDF55F7AABDEAAF784154BAF7802A",
INIT_39 => X"D7545AAAE97555A2FBFDF455D556AA00F7D1554BA5D7BC01FFFF8015410007FE",
INIT_3A => X"4154BAF7D1400BAFFD57FE005D043FE10552EAAAAAFFD140000087FC01EFA2FF",
INIT_3B => X"8428A105D7FEABEF55557DEBAFFAEBFFEFAA803DEBA5D2E82155A2FBFDE00FF8",
INIT_3C => X"7D568BEF080402000F7AAA8B55FFAABDFEFF7D16AA0008003FEBA55003DEBAA2",
INIT_3D => X"FFAAA8AAA080028BFF087BD54AA550402145550000010087FFFF45F78402145F",
INIT_3E => X"0000000000000000000000000000000000000F7D5555FFAAAAA8BFF002AAAA00",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_3,               -- Port A enable input
WEA      => wbe_a_lo_1024_3(1),               -- Port A write enable input
DIA(0)   => data_write_a(12),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_3(12),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_3,               -- Port B enable input
WEB      => wbe_b_lo_1024_3(1),               -- Port B write enable input
DIB(0)   => data_write_b(12),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_3(12),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_13_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10154A0441836CA2840512822007C18000E02700500030B31B300040081A042",
INIT_01 => X"00000804A000C04800020000000002404001000008220008A200100802110204",
INIT_02 => X"02200430000104000A4700804008000004100000000420918204D3033240400D",
INIT_03 => X"AA4003400008592400000590C40009141100000C6180C0000000C00001E14000",
INIT_04 => X"0800000102400120088054019000004160004190BAA0270000C8100000600206",
INIT_05 => X"21000012040610050040000227003AA0082400E94C1200000824424005220020",
INIT_06 => X"81963B180C001010580000080400000058000004109C00138000020024142581",
INIT_07 => X"002C8008000441600106400A9600010494020002B8AAA000EF003408000E2580",
INIT_08 => X"000000E48194408000A00A001210040441C80320040210000002ABF004102244",
INIT_09 => X"2A004009640040100400940412D4C4004000022000104200802D983000480120",
INIT_0A => X"8000202020401480000000000000080C90090881000145B0111A14004015080D",
INIT_0B => X"00000002004040AA08050400404040C11444000805200A402090024000008002",
INIT_0C => X"8410000A00280020020040800020040800020000801020000800010020400000",
INIT_0D => X"84A14250A055100050100490000500D00040080040290000084E4000B800610C",
INIT_0E => X"DCD13042BEDA36820228000000000000C000400081A08BC812A2092B02850942",
INIT_0F => X"89B9A260857DB400431969CA985D480949D32804A40AB137341C10B7D6A02EC0",
INIT_10 => X"E6ACA678001CE7D0296C213A460CA4271CA2168AEC1017606E6838216FAD4055",
INIT_11 => X"84AD4961C281B20213073C5FC0058008632D30D522CE80239DCC01AB013A4D20",
INIT_12 => X"2E6B13804A4B01D83461299900F6BD583A519104A0EEBD1A141010B2A4C8E116",
INIT_13 => X"89E5E40913419151EE0E94641828F72B5151EE0D184B321037AF5158BB02D085",
INIT_14 => X"562EC0B42162D68EE0073AE1C562EC13D521921A4170300B2B458B56B01C2280",
INIT_15 => X"00888A120240034000E6DC8285028014B82372011FC1E4F5E0A00929684EAF84",
INIT_16 => X"50942509425094250942509425094254940A1421420082020120908800480030",
INIT_17 => X"0942509425094250942509425094250942509425094250942509425094250942",
INIT_18 => X"9425094250942509425094250942509425094250942509425094250942509425",
INIT_19 => X"F7EFBBEEFF3F7DF7FF3E9F7DF7E2450228000000000000000000509425094250",
INIT_1A => X"BAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBF7DFDFDDD555555",
INIT_1B => X"EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAEBAE",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000000000F7EBF5FAFD7EBF5FAFD7",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"2ABEF00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0020105D557FEAA00557DE10AAD5554BA087FFFF55557BD54AAF7FBC01FFA280",
INIT_29 => X"7BD75EF087FFFFEF557BEAB45552E80155AA802AB45AA843FE0008557DFFF080",
INIT_2A => X"FAE820AA5D5557555082ABDF5508557DF45002ABDFFFF7803DE10AA80000AA08",
INIT_2B => X"0051555FFA2AA8200000557DFFFF7AA80000AAD1420AA087BD7555FFD168AAAF",
INIT_2C => X"5557FFDE10AAAEA8BFFA2FBD7545FFD157555085140010F7AEAABFFAAD542000",
INIT_2D => X"BA557BE8A10A284154BAFFAAAAB45007FC2155F7D155545AA80001EFAAFBEAB4",
INIT_2E => X"000A2D155410F7FFFFEBA08003FE00082AA8AAAAAFFC00BA00002AAAAF7D5574",
INIT_2F => X"0492E3F1C71C7BE8A2ABD7000000000000000000000000000000000000000000",
INIT_30 => X"3AE38145B78FD7000005010495B7AE921C517DE10A2DB50482147FFAF554971D",
INIT_31 => X"E3FE28B684070AA1C71D25D7007FFAFD7497BE8B5555208217DBE8A2AB45BE80",
INIT_32 => X"7FD257DFFD568A82FFA4870BA555F5056D002EBDF6D005B78F7D142ABDFC7F78",
INIT_33 => X"FAAAFBFFBED547038145B505FFB6A487000005F7AFD7F7A482038AADF4709214",
INIT_34 => X"AA8E071D7AAFBEFB455D71F8E00A2A0ADBC7A2FFD257DE3DF52555085142000F",
INIT_35 => X"21C002AA92FFDF574824171EAA10B680124BAFFAAAFB45007BC217DEBDB55555",
INIT_36 => X"00000000000000000000B6D550428FFF1FDE821C003FE001C2EAAAAAB6F5C208",
INIT_37 => X"0105D7BE8B55085142010AAD157545F7AEA8B550000000000000000000000000",
INIT_38 => X"01EFF7AAA8B55F7802AABA5D7FEAB45080015410007FEAA0055517DE00A2FFC0",
INIT_39 => X"E8BFF5D2ABDF55F7AABDEAAF784154BA5D5140145007BE8B55087BEAB555D040",
INIT_3A => X"0020BAA2FFD54105D7FC21EFFFD16AA10FF80174AA557FC21EF082EBFFEF007B",
INIT_3B => X"FBC0155085540000FFAEBFFEFF7D1554BA5D7BC01FFFF8015410007FEAB45F78",
INIT_3C => X"87FC01EFA2FFD7545AAAE97555A2FBFDF455D556AA00A2803FF45AAFFC21EFAA",
INIT_3D => X"552EAAAAAFFD1400005D042AA00F7FBD5410085568A10FF80020AAFFAABFF550",
INIT_3E => X"0000000000000000000000000000000000000F7D1400BAFFD57FE005D043FE10",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_3,               -- Port A enable input
WEA      => wbe_a_lo_1024_3(1),               -- Port A write enable input
DIA(0)   => data_write_a(13),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_3(13),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_3,               -- Port B enable input
WEB      => wbe_b_lo_1024_3(1),               -- Port B write enable input
DIB(0)   => data_write_b(13),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_3(13),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_14_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10020A000180000284008280000281800000030000000033022000000580002",
INIT_01 => X"000008020000204D006800000030824840000000084000084200090008510200",
INIT_02 => X"0220043170010A600A4D008040080000041000000028009002000F333240800C",
INIT_03 => X"111813400008002400000000C400090011000000610200001104D83000F14000",
INIT_04 => X"0801800100A000000000540084000040000040000800200000C8100000000748",
INIT_05 => X"0100000000001000000000002000080008000000001000000024024001200020",
INIT_06 => X"819EB84028001010000000080400000000000004108000100000020020040081",
INIT_07 => X"92040608000440100102400A94810206844200021DA2A0002000340800062C80",
INIT_08 => X"000000000084400008800A001214040441481500040000000000A7F408002244",
INIT_09 => X"0A0040090002008420401004104444004000020400214A208001000002400120",
INIT_0A => X"0400002020000000000000000000080C8008088100004590111B480040120000",
INIT_0B => X"1000000200404800000504016000002114000008020000020080024000000000",
INIT_0C => X"0410000010000000000040001000000000000040000000000001000000000000",
INIT_0D => X"04810244825010004010000000000000000000000000000000080000B8002104",
INIT_0E => X"0002C38280001202020800000000001000004000000000401022000002040902",
INIT_0F => X"20000587050001404E8084341CBA3404800828805200008000E0E0A000080002",
INIT_10 => X"4D18178E012010C00224004091C3514072C000444A0400080001C1C140001000",
INIT_11 => X"51709A07424142084458476001003809D0104B01C5710044020C4006010500C5",
INIT_12 => X"C26EE3803180C18006519462A00005001460E4730000050A1011004001060049",
INIT_13 => X"01F9E00660318000000538318740000140000001B4600CE80001400000002B62",
INIT_14 => X"0000000AD89857B0E0684411800000003799EB764D000330C300000000E3554B",
INIT_15 => X"0000021002002C000024008284001A0902000422E3F5960080480A0216A07240",
INIT_16 => X"4090240902409024090240902409024090081021020080015134920800480010",
INIT_17 => X"0902409024090240902409024090240902409024090240902409024090240902",
INIT_18 => X"9024090240902409024090240902409024090240902409024090240902409024",
INIT_19 => X"F5579B4E5C8FF0F7BE9D5F7DF650400200000000000000000000409024090240",
INIT_1A => X"9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7BF7DDDDDFCF3CF3D",
INIT_1B => X"F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE79E7",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000003FFF03F9FCFE7F3F9FCFE7F3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"420BA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"BD54AAF7FBC01FFA2802ABEFA2FBE8B55A2AE80000F7D5555555D2AAAABAAAD1",
INIT_29 => X"AA801FFA28402000AAAE955455500155EF0804155EFAAD5554BA087FFFF55557",
INIT_2A => X"7AEA8B45080417400AA843FE0008557DFFF0800020105D557FEAA00557DE10A2",
INIT_2B => X"087FFFFEF557BEAB45552E80155AA802AB4500516AA00A2AE800BAFFFFC20BAF",
INIT_2C => X"0AA80000AA005568ABAA28402010A2843FEBAFFFBD7410A2D168BFF087BD75EF",
INIT_2D => X"005D7FFDF4555517DFEF00043FEAA082ABDF5508557DF45002ABDFFFF7803DE1",
INIT_2E => X"000AAD1420AA087BD7555FFD168AAAFFAE820AA5D5557555002E80155A280000",
INIT_2F => X"0555412AA8ABAAADB40092000000000000000000000000000000000000000000",
INIT_30 => X"50482147FFAF554971D0492E3F1C71C7BE8A2ABD7A2FFEDB55B6A080038E3DB5",
INIT_31 => X"B7AE921C517DE10A2AE851FFB68402038AAAA955554900105FF0800175D7A2DB",
INIT_32 => X"A0800BAE3F1C0092EBAAADB6D080A12410BE803AE38145B78FD7000005010495",
INIT_33 => X"2D568BC71C71D25D7007FFAFD7497BE8B5555208217DBE8A2AB451C556FA00A2",
INIT_34 => X"142ABDFC7F78E3FE28B684070AA00516DABAA28402038B6803DE82F7F5D5410A",
INIT_35 => X"D002A80155B680000105D7FF8F455D5F78FD7000E3FEAA002EBDF6D005B78F7D",
INIT_36 => X"00000000000000000000AADF47092147FD257DFFD568A82FFA4870BA555F5056",
INIT_37 => X"F55FF84000AAAAFBC0145002AA8AAAAAFFC20000000000000000000000000000",
INIT_38 => X"01EF080417555A2FFC00105D7BE8B55085142010AAD157545F7AEA8B55A2FBFF",
INIT_39 => X"EAB45080015410007FEAA0055517DE00A2AA955FFFF80020BAAAAA9754508000",
INIT_3A => X"AA8B555D557FE00A280020BAAAD140000A2AEBFFEF082A82010F7802AABA5D7F",
INIT_3B => X"803DE00FFD557400AAD56AB455D5140145007BE8B55087BEAB555D04001EFF7A",
INIT_3C => X"82EBFFEF007BE8BFF5D2ABDF55F7AABDEAAF784154BA08557FEAAA284000AAFF",
INIT_3D => X"FF80174AA557FC21EF082A80145F780020105D7BEAB45557BE8B45082EBFEBA0",
INIT_3E => X"0000000000000000000000000000000000000A2FFD54105D7FC21EFFFD16AA10",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_3,               -- Port A enable input
WEA      => wbe_a_lo_1024_3(1),               -- Port A write enable input
DIA(0)   => data_write_a(14),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_3(14),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_3,               -- Port B enable input
WEB      => wbe_b_lo_1024_3(1),               -- Port B write enable input
DIB(0)   => data_write_b(14),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_3(14),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_15_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000A000000000284000280000001800020030000000033022000000180002",
INIT_01 => X"8000080000000048000000000000026040000000080000080200000000110200",
INIT_02 => X"0020042004010E60004C0080000800000410000000020090020000300245E005",
INIT_03 => X"0000010000080400000000408400480111000000610008000000C00000E54400",
INIT_04 => X"980000010000000088C2550080000040000040000008A00028C8100000120000",
INIT_05 => X"020004012E025000000001322000000A28008000011000000220004D41000000",
INIT_06 => X"819588000800101000011008040000100001060418800510000A620000000092",
INIT_07 => X"0000000800044004010C20008440810284020002102220002000340800062480",
INIT_08 => X"0000000001140800002C0A001214050540C800400406180000002DF004000244",
INIT_09 => X"1E00400900000000000016041044400440000000000042008001000000000022",
INIT_0A => X"0000000000000220000000000000080C00000081000045901118000040000000",
INIT_0B => X"0000000200404000010500004000000114000009000000000000004200000000",
INIT_0C => X"0000000000000000000040001000040001000000000000000001000020000800",
INIT_0D => X"000000000000001001208000180800000000030200000180800C400030002000",
INIT_0E => X"0000000000002600020800000000001080004000000000000002000000000000",
INIT_0F => X"A400000000000000000008000000000000000000000014800000000000000052",
INIT_10 => X"0000000000000000000000010240000000000000000000290000000000000000",
INIT_11 => X"2001C05838120800000000000000000000010000000000000000000000001804",
INIT_12 => X"081004000000000000A010000000000000902000000000180010002020000000",
INIT_13 => X"6600000000000000000024080000000000000000280400000000000000000000",
INIT_14 => X"0000000000200801000000000000000000501001920000000000000000000A40",
INIT_15 => X"0000020000000000000000003000000000000000000A101C3614000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000080000120980000000010",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000400200000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"28BEF00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"5555555D2AAAABAAAD1420BAFF8000010082A954BA00003DFEF085155400F784",
INIT_29 => X"AE95555A2FBE8BEFA2843DE00AA8015400FF84001EFA2FBE8B55A2AE80000F7D",
INIT_2A => X"2FBEAB45F7D56AABAAAD5554BA087FFFF55557BD54AAF7FBC01FFA2802ABEFF7",
INIT_2B => X"A28402000AAAE955455500155EF0804155EFFFFBE8BFF0800174AA557BFDE10A",
INIT_2C => X"A00557DE10F7D1574AAA2D16AB55FFD568BEF087FE8A1055003FE00A2AA801FF",
INIT_2D => X"00AA802AA00AAAE800BA5D0015545AA843FE0008557DFFF0800020105D557FEA",
INIT_2E => X"00000516AA00A2AE800BAFFFFC20BAF7AEA8B45080417400FFFFC21450800154",
INIT_2F => X"8FD7005150438F78A2DBFF000000000000000000000000000000000000000000",
INIT_30 => X"EDB55B6A080038E3DB50555412AA8ABAAADB40092E38E070280024904AA1C043",
INIT_31 => X"1C71C7BE8A2ABD7E3AA9257DA2FFE8BC7BE8E38E10A28017400E38A051FFA2FF",
INIT_32 => X"00124AA557FFDE10A2FBEDB6DF7D16AABAA2DB50482147FFAF554971D0492E3F",
INIT_33 => X"10038E38A2AE851FFB68402038AAAA955554900105FF0800175D7E3FFEFBD700",
INIT_34 => X"000005010495B7AE921C517DE10FFDF50482A2DB6AB45FFD56DBD7087BEAA384",
INIT_35 => X"0FFF1C017D140410400BE8E28A10AAA085082550A1057DBE803AE38145B78FD7",
INIT_36 => X"000000000000000000001C556FA00A2A0800BAE3F1C0092EBAAADB6D080A1241",
INIT_37 => X"4AA0800020BA550028B550855400AAF7AEBDFEF0000000000000000000000000",
INIT_38 => X"7400AAAE975EFA2FBFFF55FF84000AAAAFBC0145002AA8AAAAAFFC2000AAAA97",
INIT_39 => X"E8B55085142010AAD157545F7AEA8B55AAAE821EFAAFBEAB55F7AAA8A00AA841",
INIT_3A => X"417555AAFFFDF450804020AA557BFFE10A2FFFFFEFF7D568ABAA2FFC00105D7B",
INIT_3B => X"D17DF45007FE8AAA08002AAAAA2AA955FFFF80020BAAAAA975450800001EF080",
INIT_3C => X"7802AABA5D7FEAB45080015410007FEAA0055517DE00FFFBC2000AAFBE8B55F7",
INIT_3D => X"A2AEBFFEF082A82010FFD5421EF5D0000010F7AAA8A10AA8017400552A801EFF",
INIT_3E => X"00000000000000000000000000000000000005D557FE00A280020BAAAD140000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_3,               -- Port A enable input
WEA      => wbe_a_lo_1024_3(1),               -- Port A write enable input
DIA(0)   => data_write_a(15),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_3(15),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_3,               -- Port B enable input
WEB      => wbe_b_lo_1024_3(1),               -- Port B write enable input
DIB(0)   => data_write_b(15),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_3(15),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_16_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"DA22C618B1000482B688B186588884862A400438255FC38381441205BA803003",
INIT_01 => X"7045A80028404C211203A952A90341080B173340412000E1005D628000820484",
INIT_02 => X"428406A4000850848330118D0AAC55001349B108818005460229044001C01784",
INIT_03 => X"092C4020000500020000500986812C405000001A48202050000A214AC0650115",
INIT_04 => X"4804A55440256F504025E003A054F46415A4E62B6FE3307943965A00001A1152",
INIT_05 => X"0000001C40A5B950ADB8EA097057ECE14C86D2B7F85AAD17F4B100000B88148C",
INIT_06 => X"415401DCDCF2C0A8030140BCB0820A200342A1C641C1E8782F508F2B00003584",
INIT_07 => X"002701881A3202080AE00480A2002840BE1480FA004342AA6F12000054004867",
INIT_08 => X"08C54828091002000002B32A8C19064E486A8001510000014140C1E2A14891E0",
INIT_09 => X"015452B103020814004088B64102680B6596594800400413CAC0208944800000",
INIT_0A => X"96AA000484094C000000000000012C9000A0000D0A80000BF8028E87C1B99270",
INIT_0B => X"014808A02004200E540480212000A448C0082024AE50064B44000000000002A2",
INIT_0C => X"0004000D5846256AAEA811150445411150445411150445411150422A088A8200",
INIT_0D => X"00000004010042A204A0C5817D00005034052E40000817D00440004004AD3240",
INIT_0E => X"632B2673FA4587978A2004102800809225545155121740000004900090000000",
INIT_0F => X"00C6564CE7F4EA4B940076D296D003030800462CBD320018CAAAACFE9164C800",
INIT_10 => X"28834ADB1440A114793A4A30A40839AA14910D08DCB2640031955559FD3AC990",
INIT_11 => X"594AB0B1A025371CA0E034E8443C097A800EB090D4AAC91208ED2FA0CE5E09B1",
INIT_12 => X"7B50446083001B94BB38C540EBE61284BB304880E3E4579EDC00992980D58033",
INIT_13 => X"5511121840E7A2CD952ECC12ABC3E6ACB3DFB12ECE315000F61FF1727A85FDBC",
INIT_14 => X"75DEB07F6F2E7084517F126F8395CB2BEFBAB8BA8AF698228CC5E2F08ECA5159",
INIT_15 => X"5580A840A8009F8B108C80A1021B080AFC0DF6422C6077F4A77F20D0C0E21084",
INIT_16 => X"0000000000000000000000000000000000044000102A0001148442A110810359",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"558D11544C690DA64C1C4F68A360400000000000000000000000000000000000",
INIT_1A => X"14D14D14D14D14D14D14D14D14D14D14D14514514514514529E5F87869E79E78",
INIT_1B => X"D1E8F47A3D1E8F47A7D3E9F4FA7D3E9F4FA7D3E9F47A7D1E9F47A7D1E9F4D14D",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000007D3E9F4FA7D3E8F47A3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"C00AA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"03DFEF085155400F78428BEF087FFFFEFF7D168B55AAD17FFFF552EBFE00007F",
INIT_29 => X"2E975EFF7D568BFFFF80175EF0004000BA552A821FFFF8000010082A954BA000",
INIT_2A => X"55540000082EAABFFA2FBE8B55A2AE80000F7D5555555D2AAAABAAAD1420BA5D",
INIT_2B => X"A2FBE8BEFA2843DE00AA8015400FF84001EF0000020AA5D00154005D043FF455",
INIT_2C => X"FA2802ABEF557BEABEF5D0415410087FD74BAAAAEBFFEF557FC00AAF7AE95555",
INIT_2D => X"FFFFAABFEAAFF84001FF002A821FFAAD5554BA087FFFF55557BD54AAF7FBC01F",
INIT_2E => X"000FFFBE8BFF0800174AA557BFDE10A2FBEAB45F7D56AABA082A97545F7D16AB",
INIT_2F => X"FFEF552AB8E38087FC2092000000000000000000000000000000000000000000",
INIT_30 => X"070280024904AA1C0438FD7005150438F78A2DBFF0871F8FC7E3D56AB6DBEDB7",
INIT_31 => X"AA8ABAAADB400924920925EFF7D16ABFFE38E175EF1400000BA412E871FFE38E",
INIT_32 => X"0A1240055003FF6D5551420101C2EAFBD7A2FFEDB55B6A080038E3DB50555412",
INIT_33 => X"57FC00BAE3AA9257DA2FFE8BC7BE8E38E10A28017400E38A051FF0804050BA41",
INIT_34 => X"4971D0492E3F1C71C7BE8A2ABD74975EDBC7550E12410087FD74AAB6AABFFC75",
INIT_35 => X"A08249756DF7D168BC7F7AABAEAAF780051C70824851D7A2DB50482147FFAF55",
INIT_36 => X"00000000000000000000E3FFEFBD70000124AA557FFDE10A2FBEDB6DF7D16AAB",
INIT_37 => X"B55A2D16ABEFFFFBFDFFF552AAAAAA007BC00000000000000000000000000000",
INIT_38 => X"20AA002A955EFAAAA974AA0800020BA550028B550855400AAF7AEBDFEF08516A",
INIT_39 => X"000AAAAFBC0145002AA8AAAAAFFC20000000021EFF7D568BFFA2AA955FF5D040",
INIT_3A => X"E975EF0800174BA002E820105D003DFEF5D51420005D2ABFF45A2FBFFF55FF84",
INIT_3B => X"7BD74AAF7AEBDF455D7BC20BAAAAE821EFAAFBEAB55F7AAA8A00AA8417400AAA",
INIT_3C => X"2FFC00105D7BE8B55085142010AAD157545F7AEA8B5500557DF45552A8200000",
INIT_3D => X"A2FFFFFEFF7D568ABA0804155FFF7D568B55FFAAAAABAFF8415545000015555A",
INIT_3E => X"0000000000000000000000000000000000000AAFFFDF450804020AA557BFFE10",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_3,               -- Port A enable input
WEA      => wbe_a_lo_1024_3(2),               -- Port A write enable input
DIA(0)   => data_write_a(16),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_3(16),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_3,               -- Port B enable input
WEB      => wbe_b_lo_1024_3(2),               -- Port B write enable input
DIB(0)   => data_write_b(16),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_3(16),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_17_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"5284CE4FB7BD2C8994A13392DBD02E14006B82AC7E800D44D3DD2FD5F9B961C0",
INIT_01 => X"2EACD01F7E03FC6793F2199B39FC233C11D93AE6F3BB92B32091DBC339B24542",
INIT_02 => X"E63CCCC00A82C08092A2AFAE667033DB50853379C10BFDC5C6F4044443C817C6",
INIT_03 => X"7FF183635AEF9E3635AEF9E18E237040404446965C0607EE6DB7854AC4DE060C",
INIT_04 => X"D78AC33FB604488B000892EF17BE6D84196482236FE100294152E294350FB697",
INIT_05 => X"081B5F9B409420D0CDB47A05403F6CE0C08A4AB7F840EDB6F48100DFC8081081",
INIT_06 => X"768465354781CBC30316367077B4BDB50646E8D87100A8201ED01C19C020F71A",
INIT_07 => X"4002A110C922480A82D0841147162C48EBB9537A0022DC67987042EE976ABEA7",
INIT_08 => X"DB931BFEF91C00002CC0E019C0C82A4E4820C15A2330E004401891181168C4D1",
INIT_09 => X"09F3A1BC11EFBC66DB65307071477FF1030C397C060B4254064302042F803A69",
INIT_0A => X"3F330802162F3B7EE3F3EC7C7DEF207000F00059D2ED56D7EED2ED3C9A867DC0",
INIT_0B => X"185C44B91BC1740B7605040BE0018CFC7429F326B9E822FFC00074D5A0AB033A",
INIT_0C => X"00367A28FC1B7F7FEFFCFBFF3EFFCFBFF3EFFCFBFF3EFFCFBFF3EFFE7DFF9E00",
INIT_0D => X"0000000008004BA78428C7AD7FC94B533F5B4FFBD2FAD7FCCA786D43FE67C218",
INIT_0E => X"BA494CEBFD4F2667ABB6F68B29760593F33FA0CF170F40006001B1A05C000000",
INIT_0F => X"7F749299D7FAEB237DFE5865B6D2BF23265CBACE542A6FEE92333AFF33E0A9BF",
INIT_10 => X"F6C24B6D18C3C9F8E2881F3F787D776B5DB94A09955054DFDD246675FE7AC153",
INIT_11 => X"BFB349E08FF9A27EDE9FA8AEFD9E7467BFCB195CFEB56A1A70D34D1706FFFA3E",
INIT_12 => X"6FE219CA80725B875EED723FF7FCB2875EDAAFEAF7FD929BFD55BBC71D79F639",
INIT_13 => X"546670D018E7A6E581D7B6AB75FDFCECA6E581D7BB5DDFC6FF0EB7D7E859FDB5",
INIT_14 => X"B978177F6D6AF5ECDB5FB76A5F5FA165B456E0FB308710C49FCFB741598B9C7E",
INIT_15 => X"CFDAAB00AC00A8BBFC8B501CF7A0FED9A540EA1952586CEB54D143ACFF9A3BA9",
INIT_16 => X"000000000000000000000000000000000026E100002F382DBD9ECFE117805F20",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"4372003009EDCC4052E917114F981800C0000000000000000000000000000000",
INIT_1A => X"BA69A69AEBA69AEBA69A69AEBA69AEBA69A69A69A69A69A68698686981D75D74",
INIT_1B => X"6A351A8D46A351A8D068341A0D068341A0D068341A0D46A341A0D46A341A69AE",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000000000046A351A8D46A351A8D4",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"7FEAA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"17FFFF552EBFE00007FC00AA087FFFFFFFFFFFFFEFF7FBEAB450804001EFAAD5",
INIT_29 => X"D168A000004020AA5D7BE8B450051401EF087FD74AA087FFFFEFF7D168B55AAD",
INIT_2A => X"D7FEAB55FF80175EFFF8000010082A954BA00003DFEF085155400F78428BEFAA",
INIT_2B => X"F7D568BFFFF80175EF0004000BA552A821FF5D00020BA552A82000552A821555",
INIT_2C => X"AAAD1420BAFFFFFDF45AAD17FFFFAAFBC01EF5D0015555557BFDEBA5D2E975EF",
INIT_2D => X"BA007FEABEF005555555A2D1554BAA2FBE8B55A2AE80000F7D5555555D2AAAAB",
INIT_2E => X"0000000020AA5D00154005D043FF45555540000082EAABFF00516AA10552E820",
INIT_2F => X"8B550000071EFB6DF7AE92000000000000000000000000000000000000000000",
INIT_30 => X"F8FC7E3D56AB6DBEDB7FFEF552AB8E38087FC2092147FFFFFFFFFBFDFC7EBF5E",
INIT_31 => X"150438F78A2DBFFBED16AA381C0A07082497FEFB6D1451471EF007BD04920871",
INIT_32 => X"2A850105D2A80155417BEFB6DEB8E175FFE38E070280024904AA1C0438FD7005",
INIT_33 => X"D7BFAEBA4920925EFF7D16ABFFE38E175EF1400000BA412E871FF550A0009249",
INIT_34 => X"E3DB50555412AA8ABAAADB40092FFF5FFF6DAADF7FFD7B6F1C71EF55001756D5",
INIT_35 => X"7145B6AA28492487082007FEDBD700515556DA2DF50492A2FFEDB55B6A080038",
INIT_36 => X"000000000000000000000804050BA410A1240055003FF6D5551420101C2EAFBD",
INIT_37 => X"FEFF7FBFFF55A2D16AB550000175EFFFFBEAA000000000000000000000000000",
INIT_38 => X"55EF087FC200008516AB55A2D16ABEFFFFBFDFFF552AAAAAA007BC0000557FFD",
INIT_39 => X"020BA550028B550855400AAF7AEBDFEFF7D568AAA5D2A97410007BFFFFF55515",
INIT_3A => X"A955EF5D2E80010002A954005D2A82155087FFFFEFAAAA975EFAAAA974AA0800",
INIT_3B => X"D1575FF5504175EF5D7FEAAAA0000021EFF7D568BFFA2AA955FF5D04020AA002",
INIT_3C => X"2FBFFF55FF84000AAAAFBC0145002AA8AAAAAFFC2000FFD57DFFFAAFFFDF55FF",
INIT_3D => X"5D51420005D2ABFF45557FE8AAA000415410007BFFF450051555EFA2FBC0000A",
INIT_3E => X"00000000000000000000000000000000000000800174BA002E820105D003DFEF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_3,               -- Port A enable input
WEA      => wbe_a_lo_1024_3(2),               -- Port A write enable input
DIA(0)   => data_write_a(17),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_3(17),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_3,               -- Port B enable input
WEB      => wbe_b_lo_1024_3(2),               -- Port B write enable input
DIB(0)   => data_write_b(17),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_3(17),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_18_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"69844019080000A21A611406840014122A641074155FC28A2024001001801003",
INIT_01 => X"7443D920034004180005E9E3C90360C0041C0181002001602025800008440084",
INIT_02 => X"E2DCCCE61D5C008103F2000781FC0FEDEAC2161B0B8FB0008620044443006010",
INIT_03 => X"884E300802006900802006995C896D605200000856E24A040000640052141103",
INIT_04 => X"480520FC026125AC0025C9122644E3E40EC8E2001001302281841A009038A86A",
INIT_05 => X"432000040089983070019400F01010004C8DB841405A80A100B586200FAC24AE",
INIT_06 => X"09044359DC7040000000002C109B0E0A00A1104641C0803804000707284600E1",
INIT_07 => X"400D10100400481D5EB08501620000007500CE801241021FE78E404860140060",
INIT_08 => X"00880C0106A0528020019307CC082A0A4A6A01ED725021400040D028000A9729",
INIT_09 => X"00117063038000282081402E4106400B6186128040600C10C1C0200950508110",
INIT_0A => X"C0C30C2E21580C874004008080003C32A10A19090C02010E1022944061688000",
INIT_0B => X"0180A8062026000DC425C0301311324AA2373088479105D044A1022000001835",
INIT_0C => X"0D89844703649000000200000000000000000000000000000000000000000010",
INIT_0D => X"0D8306C182701404C1973010802020404084001E00010802046092B5001FB365",
INIT_0E => X"528EB314068AB8B803DB00002900800400FC503F08180050942E4200020C1B06",
INIT_0F => X"40A51D66280D6032C5F96D3C51555D5D7D5AA87285820814A3CCC501C2A60820",
INIT_10 => X"8B35A3FEBF1FEDFD9C2B30E0468AAAD5D48F37E8FC1304102947998A03984C10",
INIT_11 => X"440FE1DD772D37A0A321BC6968F32658BF2D4F2A80BF8FE3F9FE3AC362080529",
INIT_12 => X"5487910D7E5A6D961A28456A1832E5161A100DD5182BC54020EA67A189C6ED36",
INIT_13 => X"AA444CAF91EDD1B725868403BE06323551B725868A100ABD119753B70964122B",
INIT_14 => X"EDC259048ACD868EE3803D65CEDC258A8F80D55E007C3F8EBB56F4C5362C978F",
INIT_15 => X"3F240014BE84370001B6922070440556B15F7FABBC0031BCF2257C41634B14D4",
INIT_16 => X"C1B06C1B06C1B06C1B06C1B06C1B06C1B0491069068000004060300A005A0118",
INIT_17 => X"1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06",
INIT_18 => X"B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C",
INIT_19 => X"B28BBECEB80EE173C2300F7DF16000000000000000000000000041B06C1B06C1",
INIT_1A => X"8A28A28AAAAAAA28A28A28AAAAAAA28A28A28A28A28A28A2910591505C104104",
INIT_1B => X"28944A25128944A25128944A25128944A25128944A2552A954AA5128944AAAA2",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000128944A25128944A251",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"9540000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"BEAB450804001EFAAD57FEAA087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974BA082E",
INIT_29 => X"7FFFFFFFFFBFDF45AAD568B55080028B55002E82000087FFFFFFFFFFFFFEFF7F",
INIT_2A => X"0043DE10AA843DE00087FFFFEFF7D168B55AAD17FFFF552EBFE00007FC00AA08",
INIT_2B => X"0004020AA5D7BE8B450051401EF087FD74AAAAFFFDF45A2D16AB55F7FFFFFFF0",
INIT_2C => X"0F78428BEFAA80000000804154BA55042ABEF5D7FD75FFAAD540145AAD168A00",
INIT_2D => X"00082E95555085168A10557FD7545FF8000010082A954BA00003DFEF08515540",
INIT_2E => X"0005D00020BA552A82000552A821555D7FEAB55FF80175EF5D00020105D2A974",
INIT_2F => X"DFFF5D2A954AA082A92428000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFBFDFC7EBF5E8B550000071EFB6DF7AE921C7FFFFFFFFFFFFFFFF7FBF",
INIT_31 => X"AB8E38087FC2092087FFDFC7E3F1FAF55A2DF6DB7D1C002AB7D002A82028147F",
INIT_32 => X"DF6DB7DE3F5FAFC708003DE28B68E38E280871F8FC7E3D56AB6DBEDB7FFEF552",
INIT_33 => X"ADF4516DBED16AA381C0A07082497FEFB6D1451471EF007BD0492B6F1F8F55AA",
INIT_34 => X"1C0438FD7005150438F78A2DBFFA28407038140410492550A2ABC7497BD25FFA",
INIT_35 => X"F5D0E05000492097428002E9557D1C516FA28417BD5545E38E070280024904AA",
INIT_36 => X"00000000000000000000550A00092492A850105D2A80155417BEFB6DEB8E175F",
INIT_37 => X"FFFFFFFFDFEFF7FBFFFEF552E974AA082A820AA0000000000000000000000000",
INIT_38 => X"ABEF002A800AA557FFDFEFF7FBFFF55A2D16AB550000175EFFFFBEAA00557FFF",
INIT_39 => X"6ABEFFFFBFDFFF552AAAAAA007BC0000087BFDF45AAD568B55AAFBFDFEF55042",
INIT_3A => X"FC2000FFD56AB45A2FFFDFFFAAD16AB4500043DEAAFFAEAAAAA08516AB55A2D1",
INIT_3B => X"2AA8B45087FC01EFA2FFD55EFF7D568AAA5D2A97410007BFFFFF5551555EF087",
INIT_3C => X"AAA974AA0800020BA550028B550855400AAF7AEBDFEFA280154BA55040000055",
INIT_3D => X"087FFFFEFAAAA975EF5D2E974000804154BA082A975EF5D517DEAA007BD5545A",
INIT_3E => X"00000000000000000000000000000000000005D2E80010002A954005D2A82155",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_3,               -- Port A enable input
WEA      => wbe_a_lo_1024_3(2),               -- Port A write enable input
DIA(0)   => data_write_a(18),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_3(18),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_3,               -- Port B enable input
WEB      => wbe_b_lo_1024_3(2),               -- Port B write enable input
DIB(0)   => data_write_b(18),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_3(18),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_19_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"042200000000000041088001001AA00000000000000000000000500802000003",
INIT_01 => X"040048000024000000000404000000000A22000800000800004A200000000001",
INIT_02 => X"200C8840085EB00480060000001C008002489E0F000405EA0004040404000000",
INIT_03 => X"24004000000000000000000900002C4050000000000069500208400002E14100",
INIT_04 => X"4800200C0000000044002000C80020E40000E200000130200188000000800100",
INIT_05 => X"000000000080181000000000701000004C8000000058800000B1000009880480",
INIT_06 => X"80500081081040000000002C100040400000004641C080380400070100000000",
INIT_07 => X"4020109801A4CE005C00048380142810010564C4100114012002402028044808",
INIT_08 => X"0070700000000000000083004C3902420062000020E0000100004082A140102B",
INIT_09 => X"001150200000000000000026400000016186100000000010C04002C000000000",
INIT_0A => X"007C00008082C0002000000000002C3000000004050001030102040000000000",
INIT_0B => X"0000000000000000000000000000010000800011000000000000000000000BC0",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"000000000000000000000000000000042000760000000000000000010004B200",
INIT_0E => X"0D74002280300F0002FB069040000060000C5003000800000000000000000000",
INIT_0F => X"C01AE8004500744C780687DBA828008080A5FC0D385598035D0008A00C015660",
INIT_10 => X"39D8140040201BF861F0E7D693E6170022408116DFE0AB3006BA0011401D02AC",
INIT_11 => X"5412E4997F5249FD005043B8680CC98F00D0F2DD0140100406FE053A98F6ECC7",
INIT_12 => X"7418663001858040E153888000010840E165D0000000285C246A181C03FE4662",
INIT_13 => X"8199830066F0020858385974000001260208583854E2200000660208D6B1423F",
INIT_14 => X"8235AC508FCE8811042040F008235AE04420C040CF00C031C80009B8F224978B",
INIT_15 => X"030004E00000C220010808C10D9A92A74CD7CF4A09051110AD5A3C9200B7F280",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000118",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"07208BBA3F0C7010C660C7441920000000000000000000000000000000000000",
INIT_1A => X"861869A61861861861869A61861861861861861861861861A8208C4C1534D34C",
INIT_1B => X"984C26130984C26130984C26130984C26130984D26930984C26130984C261861",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000984C26130984C26130",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"174BA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFDFEF5D2A974BA082E95400F7FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0004",
INIT_29 => X"FFFFFFFFFFFFFFFFF7FBFDFFF552E974BAA2FFFFE10087FFFFFFFFFFFFFFFFFF",
INIT_2A => X"004001EFAAAEA8ABA087FFFFFFFFFFFFFEFF7FBEAB450804001EFAAD57FEAAF7",
INIT_2B => X"FFFBFDF45AAD568B55080028B55002E82000F7FFFFFFFFFFFFDFEFA2D568B550",
INIT_2C => X"0007FC00AAF7FFFFFFFF7FBE8B55AAD16ABEF5D2ABFF55080402010087FFFFFF",
INIT_2D => X"55A2FFFDFEF5D2EBFE00AAFFFFEBA087FFFFEFF7D168B55AAD17FFFF552EBFE0",
INIT_2E => X"000AAFFFDF45A2D16AB55F7FFFFFFF00043DE10AA843DE00557FFDFEFA2D16AB",
INIT_2F => X"FFEF552A974AA0000104AA000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFF7FBFDFFF5D2A954AA082A92428E3FFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"0071EFB6DF7AE92EBFFFFFFFFFFFFDFEFF7F5FAFC7492A974AAB6F5F8E101C7F",
INIT_32 => X"F1F8FD7AAD16AB450000001FFBEA4A8AAA147FFFFFFFFFBFDFC7EBF5E8B55000",
INIT_33 => X"00000010087FFDFC7E3F1FAF55A2DF6DB7D1C002AB7D002A82028FFFFFFFEFF7",
INIT_34 => X"BEDB7FFEF552AB8E38087FC2092F7FBF8FC7E3F5EAB45B6DF6FBEF5D2AB8F7D0",
INIT_35 => X"84971F8FC7AAD56DB6DBEF5F8FD7412ABFE28B6F5F8E820871F8FC7E3D56AB6D",
INIT_36 => X"00000000000000000000B6F1F8F55AADF6DB7DE3F5FAFC708003DE28B68E38E2",
INIT_37 => X"FFFFFFFFFFFFFFFFFDFEF552E954AA0004000AA0000000000000000000000000",
INIT_38 => X"54AAF7D568A00557FFFFFFFFFFFDFEFF7FBFFFEF552E974AA082A820AAA2FFFF",
INIT_39 => X"FFF55A2D16AB550000175EFFFFBEAA00A2FFFFFFFF7FBFDFFFFFD568B55002A9",
INIT_3A => X"A800AAF7FBFDFEFF7D56AB45AAD56AB450004001EFFF842AAAA557FFDFEFF7FB",
INIT_3B => X"FFFFFFF552AA8BEF080402000087BFDF45AAD568B55AAFBFDFEF55042ABEF002",
INIT_3C => X"8516AB55A2D16ABEFFFFBFDFFF552AAAAAA007BC0000FFFBE8B55AAD168B55F7",
INIT_3D => X"00043DEAAFFAEAAAAA08556AB55A2D57FFFFF7D568B45002ABDEAAFFD16AA000",
INIT_3E => X"0000000000000000000000000000000000000FFD56AB45A2FFFDFFFAAD16AB45",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_3,               -- Port A enable input
WEA      => wbe_a_lo_1024_3(2),               -- Port A write enable input
DIA(0)   => data_write_a(19),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_3(19),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_3,               -- Port B enable input
WEB      => wbe_b_lo_1024_3(2),               -- Port B write enable input
DIB(0)   => data_write_b(19),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_3(19),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_20_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000003",
INIT_01 => X"F55FF80000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"E05022020800008400F655001FFCFF80018FA804400000000000004400000001",
INIT_03 => X"00000000000000000000000900002CC07000000000000000000000000000013F",
INIT_04 => X"68002FFE40900010000180000001FFEC0012EE0C001370F40780000000000000",
INIT_05 => X"0840000880FCBBF0100E204DF0F88311DD8005080679800000F3000029980580",
INIT_06 => X"001000030817C8E8840155FDF9001001050023F6C3C3D0F87FA19F7F011000E4",
INIT_07 => X"000000090492260800008000EE00000000000000002101FF2002C00000004018",
INIT_08 => X"2A040001071004000013FF7FCA302C0C0008214800002101554031F800000000",
INIT_09 => X"801F57F200000090000489FEC0000001EFBEF0040008023FDFC0000000004006",
INIT_0A => X"0000000008000000000000000000ADF000000200000008000008028300110230",
INIT_0B => X"0000000000000800080000000000000000000000000000000800800A40000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"000000040900005C848538000020000000800000080000020000800101FFB600",
INIT_0E => X"00800000003A010003000000000000600FFC53FF001800000002004080000000",
INIT_0F => X"0001000000007408040000004000000004E9000008020000200000000E800800",
INIT_10 => X"00200000000313100010002000008000000000129600040000400000001D0010",
INIT_11 => X"81C012060000000000218F7840000100800004000000000066C0000080080000",
INIT_12 => X"800000000017C000100000000001A800080000000001A8040000002840008185",
INIT_13 => X"0000000006F00000100200000000012600001004000000000066000000801040",
INIT_14 => X"0000200410100000000005F00000020080090A0000000085C800002000586000",
INIT_15 => X"FF00400000000000020020020001000040283024E4F2860400008000030ED080",
INIT_16 => X"00000000000000000000000000000004010201001003020200000000000127DB",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"A0700030038200010089120104D2040020000000000000000000000000000000",
INIT_1A => X"2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2C30C30C30C30C306982121A1E79E79",
INIT_1B => X"32190C86432190C86432190C86432190C86432190C86432190C86432190CB2CB",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000432190C86432190C864",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0201000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF552A974AA0004174BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA0804",
INIT_29 => X"7FFFFFFFFFFFFFFFFFFFFFFEF552E954AA000400000F7FFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E954BA007FC00BA087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974BA082E9540000",
INIT_2B => X"FFFFFFFFFF7FBFDFFF552E974BAA2FFFFE10FFFFFFFFFFFFFFFFFFFFFBFDFFF5",
INIT_2C => X"FAAD57FEAA007FFFFFFFFFFFFFEFF7FBFFF550800020BAAAD56AAAAF7FFFFFFF",
INIT_2D => X"EFF7D56AB450000021EFA2D57DE10087FFFFFFFFFFFFFEFF7FBEAB450804001E",
INIT_2E => X"000F7FFFFFFFFFFFFDFEFA2D568B550004001EFAAAEA8ABA5D7FFFFFFFFFFFDF",
INIT_2F => X"FFFF5D2E954AA080005000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFEF552A974AA0000104AAFFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"A954AA082A92428087FFFFFFFFFFFFFFFFFFBFDFEF5D2E974AA000A07000E3FF",
INIT_32 => X"FFFFFEFF7FBFFFFF552E974AA0071C50BA1C7FFFFFFFFFFFFFFFF7FBFDFFF5D2",
INIT_33 => X"EDF6FABAEBFFFFFFFFFFFFDFEFF7F5FAFC7492A974AAB6F5F8E10E3FFFFFFFFF",
INIT_34 => X"EBF5E8B550000071EFB6DF7AE921C7FFFFFFFFFBFDFEFE3F5F8F450004050AAB",
INIT_35 => X"A497FFFFFFF7FBF8FC7EBD168B450804021FFB6D57DE28147FFFFFFFFFBFDFC7",
INIT_36 => X"00000000000000000000FFFFFFFEFF7F1F8FD7AAD16AB450000001FFBEA4A8AA",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2A954AA0800174100000000000000000000000000",
INIT_38 => X"74AA002E95410A2FFFFFFFFFFFFFFFFFFFFFDFEF552E954AA0004000AAFFFFFF",
INIT_39 => X"FDFEFF7FBFFFEF552E974AA082A820AA087FFFFFFFFFFFFFEFF7FBFDFFF5D2A9",
INIT_3A => X"568A00AAFFFFFFFFFFBFDFEFFFFFFDFEF5D2E954AA0051554BA557FFFFFFFFFF",
INIT_3B => X"D16AB450804174AAFFFFFFEBAA2FFFFFFFF7FBFDFFFFFD568B55002A954AAF7D",
INIT_3C => X"57FFDFEFF7FBFFF55A2D16AB550000175EFFFFBEAA005D7FFFFEFF7FBFDFFFAA",
INIT_3D => X"0004001EFFF842AAAA087BFDFEFF7FFEAB45A2D568B550804001EFF7D57DEBA5",
INIT_3E => X"0000000000000000000000000000000000000F7FBFDFEFF7D56AB45AAD56AB45",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_3,               -- Port A enable input
WEA      => wbe_a_lo_1024_3(2),               -- Port A write enable input
DIA(0)   => data_write_a(20),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_3(20),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_3,               -- Port B enable input
WEB      => wbe_b_lo_1024_3(2),               -- Port B write enable input
DIB(0)   => data_write_b(20),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_3(20),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_21_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"4A302428B824900A128C090A5C1800261500213C005FE812D10420054085A202",
INIT_01 => X"001FFE3440B609703B0427F801A40B8115BC4F655300340288A40D30040E4DD8",
INIT_02 => X"E00424256888D8819801000F9FFFFFFFF149FF1FCA448046C60A0D2437C517F9",
INIT_03 => X"20030640003250640003250F06002CC1740002019824E001CD357832440001FF",
INIT_04 => X"EA2C3FFD400006E04401A8837001FFFC004AEF00080B70E08FB5789421007C5C",
INIT_05 => X"00011A0C40F9FFF80920954FF0F00809DF84A0202879800000F3000029980780",
INIT_06 => X"0805984B7A1FC0A0000101FFF0480080002281F7C3C381F87C03DFFF00009004",
INIT_07 => X"B424068086A205481A60A19000908204A855B000A08A61FF20C3D004D331D340",
INIT_08 => X"1BFA0001600802000023F7FFC08D234B40C2028253000040114200000D0226C0",
INIT_09 => X"EF1F5FF054096C6ADBA169FFC202B1C1FFBEF0440021083DFFCE22DC2880E24D",
INIT_0A => X"45FF0C004041D84862A28C54518DBFF00020004C0A6044901112A0908AA0A300",
INIT_0B => X"018C241102068006C620C03882019480E63180855A492712CC01C49C20201BFE",
INIT_0C => X"08A9464116544302C02D92236488D92236488D92236488D922366446C911B210",
INIT_0D => X"08800444021048034004001890000806002804A0822189000900D80621FFBE00",
INIT_0E => X"060580261013813A2CC396506102C4053FFD5BFF00A04A00200602CA52001100",
INIT_0F => X"080C0B004C202621A85C09411500135844C196D3606941018150098404C1A304",
INIT_10 => X"B02901013416181C96C2C9C600890A2028172192C460D1820302A0130809834A",
INIT_11 => X"9C5E803408250180AC268D185DB3F4350B811068C00049A0A4AA68F05C96A001",
INIT_12 => X"002C006560138F032B1804101244C883052208209040CC849063A747512B7678",
INIT_13 => X"41401E240665750440C9488280254530314080C2C601040420352148A00501B1",
INIT_14 => X"500811204D000700114204A70422016149916011008CAA8858850B00C32591C0",
INIT_15 => X"FFC06E60AC0496022300233104663040808E991765205000070121D41D18D098",
INIT_16 => X"40100401004010040100401004010040102090010008000001C0E010020007DF",
INIT_17 => X"0100401004010040100401004010040100401004010040100401004010040100",
INIT_18 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_19 => X"FFEF9FEEFF7FFDF7FF3E3DFDF7E0000000000000000000000000401004010040",
INIT_1A => X"BEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBFFDFDFFFCF3CF3F",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFEFF7FBFDFEFF7FBFDFEFBEF",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000FFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0001000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E954AA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0004",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA0004154BAFFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"52E974BA0804000AAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0004174BAFF",
INIT_2B => X"FFFFFFFFFFFFFFFFEF552E954AA000400000007FFFFFFFFFFFFFFFFFFFFFFEF5",
INIT_2C => X"A082E95400007FFFFFFFFFFFFFFFFFFFFDFEF5D2E974BA002E97400007FFFFFF",
INIT_2D => X"FFFFFBFDFEF5D2A954AA002E974BA087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFBFDFFF5D2E954BA007FC00BA5D7FFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA000002000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080005000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"A974AA0000104AAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974BA0000174AAFFFF",
INIT_32 => X"FFFFFFFFFFFFDFEF552E954BA080A000AAE3FFFFFFFFFFFFFFFFFFFFFFFEF552",
INIT_33 => X"02A95400087FFFFFFFFFFFFFFFFFFBFDFEF5D2E974AA000A07000007FFFFFFFF",
INIT_34 => X"F7FBFDFFF5D2A954AA082A924281C7FFFFFFFFFFFFFFFFFFBFDFEF5D2A974BA0",
INIT_35 => X"A557FFFFFFFFFFFFFFFF7FBFDFFF552E974BA0020924BA1C7FFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000E3FFFFFFFFFFFFFFEFF7FBFFFFF552E974AA0071C50B",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0000020000000000000000000000000000",
INIT_38 => X"74BA0000174BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954AA080017410FFFFFF",
INIT_39 => X"FFFFFFFFFFDFEF552E954AA0004000AAF7FFFFFFFFFFFFFFFFFFFFFFFEF552A9",
INIT_3A => X"E95410087FFFFFFFFFFFFFFFF7FBFDFEF5D2A954BA082E800AAA2FFFFFFFFFFF",
INIT_3B => X"FBFFFFF552E954BA002E97410087FFFFFFFFFFFFFEFF7FBFDFFF5D2A974AA002",
INIT_3C => X"57FFFFFFFFFFFDFEFF7FBFFFEF552E974AA082A820AA557FFFFFFFFFFFFFEFF7",
INIT_3D => X"5D2E954AA0051554BA5D7FFFFFFFFFBFDFEFF7FFFFFEF5D2A974BA0000020AA5",
INIT_3E => X"0000000000000000000000000000000000000AAFFFFFFFFFFBFDFEFFFFFFDFEF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_3,               -- Port A enable input
WEA      => wbe_a_lo_1024_3(2),               -- Port A write enable input
DIA(0)   => data_write_a(21),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_3(21),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_3,               -- Port B enable input
WEB      => wbe_b_lo_1024_3(2),               -- Port B write enable input
DIB(0)   => data_write_b(21),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_3(21),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_22_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"5290F4CDE914905A14A43D33F488243E17122300F55FEB189B343A1140548380",
INIT_01 => X"A54007B259F6A975386262000C344BA9573C6FF57B18A5FB0ABFCD3C2C5F4F0C",
INIT_02 => X"021DFF8C38B3C009D203551040030071869D0040180AA2DC53DB89BEA8204001",
INIT_03 => X"2603475A969D0475A969D0460EAA401005111011BD506954EDB40F5EF41434C0",
INIT_04 => X"922D9002100ED69E443D988B0D5400103E48003D0800011E803B06B5B9125A15",
INIT_05 => X"281B5A0C06000408F4DF9422010D8802022F2124A8022492580040440002021C",
INIT_06 => X"F780C4C052881ADA0E05440205DA50930FA182010004700083E220800440B588",
INIT_07 => X"049D028B93FB561833D8094A02F5EA92FD7247E10305C40040D136E6A023F7FC",
INIT_08 => X"00028241680A0E002A9400803A884B5B5206B7C2E53CA25144009007A64EBD64",
INIT_09 => X"41008810240240C6694008010392354010000560141801002028A83D2A08E06D",
INIT_0A => X"34000000848BCA6902A29C54539C020E11810098D4067EFF9FF284D483E2AB41",
INIT_0B => X"500001840000C80B410014088040F4A944B1AA313C0022AA0011C0DC00028001",
INIT_0C => X"80B14004D158C8CA24A1C2A870AA1C2A870AA1C2A870AA1C2A872550E1543800",
INIT_0D => X"80A14050A01509E050854498B5281A1C34E506A2C6898B52A154DAC6B6000850",
INIT_0E => X"0B03001A483A4146603050080410089180008800143D83888281A2034A850142",
INIT_0F => X"A4160600349075238473F1210006133835E92273612B3482C090068A0E84AC56",
INIT_10 => X"30060181BA1B13959DC08DA902458870201970B29602562B0581200D141D0959",
INIT_11 => X"E042021C040D0152C8058B3840F044708E7E1C20A0106EA166C13AFC14AA3804",
INIT_12 => X"080E004B0C17C1439A9838301DC1A8438EA32C009DC1A8255300650458A1D588",
INIT_13 => X"018010E186F110A908E3A8CB0026C9A610A908E6A60F0807626610E160589C4C",
INIT_14 => X"2A701667334005800B1605F043858125E0D04110408D2485CA034681E43A1E40",
INIT_15 => X"00646002304244A91102C93A2D608D2A258DF8034188200C050171A41108F084",
INIT_16 => X"110441104411044110441104411044110466C440446CA06951D4EA8010009804",
INIT_17 => X"0040100401004411044110441104411044110441104411044110441104411044",
INIT_18 => X"0401004010040100401004010040100401004010040100401004010040100401",
INIT_19 => X"F7DFBFDEFE8FF1F7DEBDDF7DF7D05122890000000003FFFFFFFF900401004010",
INIT_1A => X"9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7BFFDFD7DDDF7DF7D",
INIT_1B => X"F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE79E7",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000003F9FCFE7F3F9FCFE7F3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA000400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0800",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000002000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2A954BA000015400FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080402010FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2A954BA0004154BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A0004174BAFFFFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0800154AAFFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF552A974AA0000174BAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974A",
INIT_2E => X"000007FFFFFFFFFFFFFFFFFFFFFFEF552E974BA0804000AAA2FFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080400010000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E954AA080005000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000402010FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2A954BA000417410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"804154BAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974BA0000174AAFFFFFFFFFFF",
INIT_34 => X"FFFFFFFEF552A974AA0000104AAE3FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0",
INIT_35 => X"AA2FFFFFFFFFFFFFFFFFFFFFFFEF552E954BA000E124BAE3FFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000007FFFFFFFFFFFFFFFFFFFFDFEF552E954BA080A000A",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804000100000000000000000000000000",
INIT_38 => X"54AA000400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2A954AA080017410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"0174BAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A954BA000415400FFFFFFFFFFFFF",
INIT_3B => X"FFFDFEF552E974AA0804174AAF7FFFFFFFFFFFFFFFFFFFFFFFEF552A974BA000",
INIT_3C => X"2FFFFFFFFFFFFFFFFFFFFFDFEF552E954AA0004000AAA2FFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2A954BA082E800AAAAFFFFFFFFFFFFFFFFFFFBFDFEF5D2E954BA002A820BAA",
INIT_3E => X"0000000000000000000000000000000000000087FFFFFFFFFFFFFFFF7FBFDFEF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_3,               -- Port A enable input
WEA      => wbe_a_lo_1024_3(2),               -- Port A write enable input
DIA(0)   => data_write_a(22),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_3(22),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_3,               -- Port B enable input
WEB      => wbe_b_lo_1024_3(2),               -- Port B write enable input
DIB(0)   => data_write_b(22),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_3(22),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_23_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"EF20906D902424807BC8241BC81801B97D38AD3C0800103362A6741C80A12A02",
INIT_01 => X"001FFF8409F089003B4422000D80C80106804A7951C5B9D1C828043EA28838F9",
INIT_02 => X"E01CEE21649C82C40800000F9FFEFF8E72CA7F5FC2E22809925A0D3611C877F8",
INIT_03 => X"24000400402670400402670D48222DC1764446838624000080007460C40001BF",
INIT_04 => X"68403FFC020560E0443E21037C01FFFC0002EE00628BF0E02FAD781014085014",
INIT_05 => X"0112000202FBFFF00920017FF0F0628BFF8488890979800002F702002BB807A0",
INIT_06 => X"EF85788B681FC000000001FFF0010000000001F7CBC385F87C0BFFFF20040001",
INIT_07 => X"F6E200000000C1440E3AE408009120071070FA07A1CB23FFA403F0C4D23BF7C0",
INIT_08 => X"0BF87CA400804000003FF7FFD8880A034AC09662305AB10555421006891A1089",
INIT_09 => X"BE1F5FEA10092C0896A243FFC0008087FFBEF2000000001DFFC612C0C0400100",
INIT_0A => X"41FF0C2060501000600000000001BFFA800808189A657EF81DD0C00079CC8001",
INIT_0B => X"018C24110A860006C620C0312241C482B20400CC52492710CC80060020A81BFE",
INIT_0C => X"0C08866907048320C20C10030400C10030400C10030400C10030400608018210",
INIT_0D => X"040002000041500300100040000500C000801000C02400000952800001FFBF04",
INIT_0E => X"FC850015385380380CDB86106502C5043FFD5FFF00A04BC010A7724B10000800",
INIT_0F => X"89F90A002A70A710A51C01C05904014861433602A1CAF13F2110055614C72FC0",
INIT_10 => X"E02D02001C1E14981B43253EE50C8220180F1082E06397E07E42200AAC298E57",
INIT_11 => X"8421802400A90022B0070FAE18019214A380344920080B21A58B02AC60BACDF0",
INIT_12 => X"0A2A000C480B0704B54028101AC49C84BB4100009AC49C80857A82D20CE8CB22",
INIT_13 => X"01E00C8103416445C12ED0400027C5292445C12D500B0005A62D344CB241D095",
INIT_14 => X"132C907425604680038706A35132C94BDD011010404428886AC91B11311C8280",
INIT_15 => X"FF000470BE0692020328CA0028042054A92771C50FC070110001C1680809591D",
INIT_16 => X"00802008020080200802008020080200800800200200000000000008004807DF",
INIT_17 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_18 => X"8020080200802008020080200802008020080200802008020080200802008020",
INIT_19 => X"0000000000000000000000000000000000000000000000000000008020080200",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080002010FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974AA000400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000400010FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974AA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080000010FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E954AA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954A",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA000015400FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080002010FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974AA000400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000402010FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E954AA080005000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA080407000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA00041741",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080000010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000402010FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2A954AA080002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954AA080017410FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"552A954BA000415400F7FFFFFFFFFFFFFFFFFFFFFFFFF552A954BA080015410F",
INIT_3E => X"0000000000000000000000000000000000000F7FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_3,               -- Port A enable input
WEA      => wbe_a_lo_1024_3(2),               -- Port A write enable input
DIA(0)   => data_write_a(23),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_3(23),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_3,               -- Port B enable input
WEB      => wbe_b_lo_1024_3(2),               -- Port B write enable input
DIB(0)   => data_write_b(23),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_3(23),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_24_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100600007FFF000080108004000800020000840041000080808",
INIT_02 => X"FC5CA803400EB8209000000F9FFEFF8E7240FF1FC22409EA04018E50074017F0",
INIT_03 => X"11100400000000400000000D00002CC07400000090C080019001010A000001BF",
INIT_04 => X"68003FFC00040000000000008001FFFC0002EE00000370E007A100000000E468",
INIT_05 => X"0000000000F8BFF00920004DF0F00001DF8000000079800000F3000029980780",
INIT_06 => X"6E461803081FC000000001FFF0000000000001F7C3C380F87C019FFF00000000",
INIT_07 => X"600C2400013649609C8000980040814210254000A00B21FF2003F2A80D500000",
INIT_08 => X"0BF80000000000000003F7FFD88D2B4A02C0940062EC2804001610020408178B",
INIT_09 => X"8E1F5FE010092C0892A041FFC0000001FFBEF0000000001DFFC002C000000000",
INIT_0A => X"41FF0C0000000000600000000001BFFA0000005501AA00000CE2000009400000",
INIT_0B => X"018C0411020600048620C030020502000200000400490510CC00040020201BF4",
INIT_0C => X"0808064106040300C00C10030400C10030400C10030400C10030400608018210",
INIT_0D => X"0000000000004003000000000000001200580000000000000000000001FFBE00",
INIT_0E => X"0086C022005381380FDB96516140C6043FFD5BFF000041000000004110000000",
INIT_0F => X"80010D804400A7240C840C201D0210840043B4804012500021E0088014C04940",
INIT_10 => X"4109038041021C980200D06410C1924030008142E06024A00043C01100298092",
INIT_11 => X"587CC200002100C14428090A1D02348190814C09C010104025AA40041A0D8005",
INIT_12 => X"022E0030300B0E46177004208000D8C61D7004300000D884817B00011306B2D9",
INIT_13 => X"01E003060344710009875C018100013831000985DC000C20003C310006143B70",
INIT_14 => X"4001850EDC004780144806A64400186CBF8961104000C3807884000846EB9500",
INIT_15 => X"FF0006E08C063C0220002201490418082010A57263E0100008000290161E711C",
INIT_16 => X"00000000000000000000000000000000000000000000000000000000000007DF",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"F2D0AEEAF6E7CC1132CDB4441990000000000000000000000000000000000000",
INIT_1A => X"BEFBE79E79E79E79E79EFBEFBEFBEFBEFBEF9EF9EF9EF9EFA69861219575D75F",
INIT_1B => X"783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1EFBEF",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000783C1E0F0783C1E0F0",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0201000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A000400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA000400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000400000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402010000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"00002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080002010FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000400010FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA00040000",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020100000000000000000000000000",
INIT_38 => X"74BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"000010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA000002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974AA000402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000002010F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_3,               -- Port A enable input
WEA      => wbe_a_lo_1024_3(3),               -- Port A write enable input
DIA(0)   => data_write_a(24),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_3(24),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_3,               -- Port B enable input
WEB      => wbe_b_lo_1024_3(3),               -- Port B write enable input
DIB(0)   => data_write_b(24),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_3(24),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_25_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100200002000000080100004000000020000800041000080808",
INIT_02 => X"FC400086000000800000000F9FFEFF8E738FFF1FC204010000000111568DD7F8",
INIT_03 => X"00000400000000400000000D00002CC4740000008000000080000000000001BF",
INIT_04 => X"68003FFF64A564AC000000000001FFFE0082EF00010370E007A1000000004000",
INIT_05 => X"0A00040148F8BFF80920804DF0F00101DFC040000079C92484F30499299837C1",
INIT_06 => X"66041803081FC0E0801101FFFD000E41002299F7E3C380F87C019FFF81200096",
INIT_07 => X"000000080480AE00000080000000000000000000A00B21FF2003E00000000000",
INIT_08 => X"1BF80000400A02000003F7FFFA0008000200A0400008A0000014100200081000",
INIT_09 => X"8E1F5FFA53EFBCACB2E369FFE0010001FFBEF80C40630C7DFFEEBAF000800202",
INIT_0A => X"41FF0C0600000000600000000001BFFE00301000000000000CC020000140000C",
INIT_0B => X"01DCCC31222730A49620C030020100000200000400490D10EC00040220201BF4",
INIT_0C => X"0808064106240300C00C10030400C10030400C10030400C10030400608018210",
INIT_0D => X"0883044582114013412080000000000000000000000000000012800001FFBE00",
INIT_0E => X"00040020000180380FC386106140C6043FFD5BFF00A04B80608003CB120C1106",
INIT_0F => X"0000080040000200040400000100000000009480000240000100080000400900",
INIT_10 => X"0001000000000808000000240000020000000100006004800002001000008012",
INIT_11 => X"0001001808220000002004001900000080800008000000000022400000088000",
INIT_12 => X"0010000000000E00110000000000408009000000000040808063004000008200",
INIT_13 => X"6000000000046100000240000000001021000004400000000010210000001010",
INIT_14 => X"4000000404000800000000060400000088000001800000001084000000088000",
INIT_15 => X"FF800C608C041002000002000006100000002100000000180600000000100018",
INIT_16 => X"4110441104411044110441104411044510629041040D180400000010028047DF",
INIT_17 => X"1104411044110441104411044110441104411044110441104411044110441104",
INIT_18 => X"1044110441104411044110441104411044110441104411044110441104411044",
INIT_19 => X"FBA2894A196A8C5A2932EC15DA080800002FFFFFFFFFFFFFFFFFC11044110441",
INIT_1A => X"2492492492492492492410410410410410410492410492412000531215A69A6B",
INIT_1B => X"158AC562B158AC562B158AC562B158AC562B1588C46231188C46231188C49249",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000B158AC562B158AC562B",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080000010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000010FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08000000",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_3,               -- Port A enable input
WEA      => wbe_a_lo_1024_3(3),               -- Port A write enable input
DIA(0)   => data_write_a(25),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_3(25),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_3,               -- Port B enable input
WEB      => wbe_b_lo_1024_3(3),               -- Port B write enable input
DIB(0)   => data_write_b(25),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_3(25),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_26_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"E9264EAB20190CA3BA4997AA9002AE9C001006B0778015CFA17E0811039879C7",
INIT_01 => X"2FFFF9BB1F773C7F9BB07DFFFDD863FC5FFF3FEFFBBF9FFB22FFFBC7B9F30686",
INIT_02 => X"E06CCC62052E708180F6FFBFFFFCFFFFF9C7FF7FC24332E642090000074037F6",
INIT_03 => X"428003739CD9863739CD9869FE2B7DEAF300029E4E300DFE69A6E644E6FF473F",
INIT_04 => X"7C2FEFFFF5BA124F003DD31EAFFFFFEE9FF7EE6F4C0770FFD7DC7CA53997B2B1",
INIT_05 => X"DFFB5421C1F8BBFAFDBFFACDF0FFCC05DDDBFF3690F9EDB7F5F7AFF639BD7DE3",
INIT_06 => X"EFD044ABC817C3E3A74667FDFFB6FF5727CC3BFEF7C3FAF87FF59F7FFBFEF69F",
INIT_07 => X"00003002132462052E708180EF060C18E5BEFB051225CDFF7002C4EEDE77F6E0",
INIT_08 => X"3FFF7D5000EC75088ED3FF7FC8790E46426CE06CB1F8E041051831FA3068D77E",
INIT_09 => X"C05FD7FF9BEFBDCEFBEE59FEF44F6603EFBEFAFCC2E35E7FDFD147CCF3F583FA",
INIT_0A => X"67FF1C7FBFADEB31E35768E8ED6BFDF3EB3EBF9DDBCE7FDC1DF8A760F3EACC02",
INIT_0B => X"5BDDCC3B336F7C548667D47B7737AF3FD62601EDC25B3533DCEB07F262213FFC",
INIT_0C => X"5F9A06E19F4D93A0EA0F78C35E30D78C35E30D78C35E30D78C35E986BC61AE31",
INIT_0D => X"5FD7AFEFDFFAF59B6FF28FE1D80D73D840607307DCFE1D80EF69A004DFFFF7FF",
INIT_0E => X"0004001F8041897B2FFFC6D86D70CE04FFFFF3FF1F5F5475BD7F72E4D75EBFAF",
INIT_0F => X"F60008003F008237B0040A00010003E020023E0201F45EC0010007E01047D17B",
INIT_10 => X"00010001DC0004C81003DE050A700200001DC0006863E8BD8002000FC0208FA2",
INIT_11 => X"2200E400002801E1A00004C21C0206F60081800800007B00010F02007EC09A0E",
INIT_12 => X"0880007E000807C7C1A612001E0015C7C19C22001E0015C59DFE82011A311AA0",
INIT_13 => X"00001BC00101F60409F0670840070809760409F06984800780097604067D0010",
INIT_14 => X"81019F40042100001F800203D81019EC085614000085C80023D81009CF008A74",
INIT_15 => X"FF802FFDFFAFD082003B032FB987E04021D481D4000819060801E0D00001231D",
INIT_16 => X"EBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEFFBFBFBFBBFCFBB0FFDFEFFEF2DFFFFFB",
INIT_17 => X"BFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAF",
INIT_18 => X"FAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFE",
INIT_19 => X"475B15BCF491E166CC8553F86EDB5C88646FFFFFFFFFFFFFFFFFEBFAFEBFAFEB",
INIT_1A => X"861861861861861861861861861861861861869A69A61861AFBD54D5F871C71D",
INIT_1B => X"984C26130984C26130984C26130984C26130984C26130984C26130984C261861",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000984C26130984C26130",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040201",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_3,               -- Port A enable input
WEA      => wbe_a_lo_1024_3(3),               -- Port A write enable input
DIA(0)   => data_write_a(26),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_3(26),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_3,               -- Port B enable input
WEB      => wbe_b_lo_1024_3(3),               -- Port B write enable input
DIB(0)   => data_write_b(26),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_3(26),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_27_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"00080A40000A41248002029000050A088000008242A0004404480002000A1155",
INIT_01 => X"2FFFF1C11F781C129C107DFFFE0860941E81258CA2B71C2220EC1B86E1A00002",
INIT_02 => X"E1000000810000014400FF6FFFF0FFFFF8007F1FC21110005080200000221FF0",
INIT_03 => X"4080026318C18226318C1821302232EAE00002BE001115FE48620040840A863F",
INIT_04 => X"643D4FFC2530000F003D821C0BFFFF8E9EF79E6D440748FED70060842105B0B0",
INIT_05 => X"D6F39020D1F8A3FAFDBFBACDC8FDC405D1DB7F1490E5EDB7D5CBADB2385D79C3",
INIT_06 => X"6FE000A38007C3032646EFF1F0B6FF46A78C39F8E723F2E47FE59C7F9ADA2612",
INIT_07 => X"00002820000000810000014401060C180190310540118DFF1000C0849673F6C0",
INIT_08 => X"3FF779100062B12A8EC3F47FC80208808210880C00082050000110023068D030",
INIT_09 => X"005F07E09BFFBD07FBAC09F8E42922038F7DF8BEC2E39C5F1FD047CEF1B582D8",
INIT_0A => X"63FF5D5F9FADE911E81C09818109E1F16B16B71092CE7ED81CF403601228C402",
INIT_0B => X"1BFDCC39732F3554866AD57C37BEAF1C152201A4C05B7531D56B05B06A213FF8",
INIT_0C => X"5BCA06F18FC59380F00E34430D10C34430D10C34430D10C34430F0861A2186B5",
INIT_0D => X"5B56ADAB5FAAE58B2F628EA0C80FA3F04040510768EA0C80CC61A0044DFFC6EB",
INIT_0E => X"0004001D800188792CE79715710AE4047FFD23FF315D54358D593474955AB6AD",
INIT_0F => X"520008003B000297B0040200010003E020001F0201E44A400100076000579129",
INIT_10 => X"00010001DC00004A10035E0408300200001DC000086BC8948002000EC000AF22",
INIT_11 => X"02002400002801E1A00000C01E0202F60080800800007B00000782006EC0820A",
INIT_12 => X"0080007E000006A7C10602001E0001A7C10C02001E0001C18DE282010A311AA0",
INIT_13 => X"00001BC00000FE0401F04300400708007E0401F04180800780007E04047D0010",
INIT_14 => X"81011F40040100001F800002F81011EC080604000085C80001F810094F008034",
INIT_15 => X"FF800C6DDDAFD082001B03249887E04001D481D4000009020801E0D00001021F",
INIT_16 => X"AB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6BF1EBDABD8E270BF84A25C6ACB777E3",
INIT_17 => X"B6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6AD",
INIT_18 => X"6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADA",
INIT_19 => X"490E2168100481CA860402104A471688747FFFFFFFFFFFFFFFFFAB6ADAB6ADAB",
INIT_1A => X"000000000000000000000000000000000008200000000000200072F210000001",
INIT_1B => X"05028140A05028140A05028140A05028140A0500804020100804020100800000",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000A05028140A05028140A",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040201",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_3,               -- Port A enable input
WEA      => wbe_a_lo_1024_3(3),               -- Port A write enable input
DIA(0)   => data_write_a(27),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_3(27),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_3,               -- Port B enable input
WEB      => wbe_b_lo_1024_3(3),               -- Port B write enable input
DIB(0)   => data_write_b(27),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_3(27),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_28_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"02200AA400180030808802A900002A08001280A08A801044104A1000001818C3",
INIT_01 => X"0AA00011460214428114180000882214413D0A71592A01D92213D28005210202",
INIT_02 => X"0451110A012100884000AA30200000000C100040104112101100008888200000",
INIT_03 => X"448000318C52A20318C52A20148810200111100C211004AA00034204200A2200",
INIT_04 => X"04004001001A90110000121402AA0000003C00000500000040080421080D0080",
INIT_05 => X"4060000C8001000000002E000000050000001610300000010000802202040012",
INIT_06 => X"1000002080001111001222000425A1040026A008000000000000000009328280",
INIT_07 => X"2491008A00491201210088400122448908A20402000408001000040820000000",
INIT_08 => X"20058310402A160026500000028040101004200C840082115554000112244814",
INIT_09 => X"4140000800000060000720000102028000000490160801020002200011100010",
INIT_0A => X"020000081B34211082B694D4D294000020020381040000000200032040004400",
INIT_0B => X"4800210C19808400500010009110091500020B408810000100200020408B0000",
INIT_0C => X"01028000080118020023604858121604858121604858121604858090B0242C00",
INIT_0D => X"010000800920040804020A6058003108402043058C460580653020005A004039",
INIT_0E => X"00000002800008014004104104420A00C000200005000010040A0020CC000200",
INIT_0F => X"520000000500000010000200000000000000280000040A40000000A000001029",
INIT_10 => X"00000000000000C0000002000830000000000000480008148000000140000020",
INIT_11 => X"020024000000000000000440000000020000800000000000000C00000040020A",
INIT_12 => X"00800000000001804006020000000500400C0200000005400A90000000100000",
INIT_13 => X"0000000000018200001003004000000142000010018080000001420000200000",
INIT_14 => X"8000080000010000000000018800008000060400000000000310000008000034",
INIT_15 => X"000002040080000000110006B081400000400000000009020000000000002200",
INIT_16 => X"802008020080200802008020080200802101210810C39A66A90A85420413A820",
INIT_17 => X"0200802008020080200802008020080200802008020080200802008020080200",
INIT_18 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_19 => X"DE21102C110A00246972BD89A40A0C22E1000000000000000000002008020080",
INIT_1A => X"2082082082082082082082082082082082082082082082080D35050758C30C31",
INIT_1B => X"0582C160B0582C160B0582C160B0582C160B0580C06030180C06030180C08208",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000B0582C160B0582C160B",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_3,               -- Port A enable input
WEA      => wbe_a_lo_1024_3(3),               -- Port A write enable input
DIA(0)   => data_write_a(28),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_3(28),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_3,               -- Port B enable input
WEB      => wbe_b_lo_1024_3(3),               -- Port B write enable input
DIB(0)   => data_write_b(28),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_3(28),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_29_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"79964E4BA01DACAB9E659792D00AAE160002829C7FDFEFCEE97C2815039D70C3",
INIT_01 => X"0ABFF9AB0775343F9AB01DF80D5821FC0FFF3FEFD1AF9FF1207FFBC7B9720586",
INIT_02 => X"002CCC60050E700080F6AAA7BFFC007189C7FF2FC00330E602800000074037F6",
INIT_03 => X"468003210868A63210868A68DA017D207200021C4E200CAA6186A40042FF4300",
INIT_04 => X"7C2FE002F0900001003C5316A6ABFFE21F36E02F0D03701F47D41800109FB281",
INIT_05 => X"4979440580F9B808F49F6A4DF00F8D01DC4B97369078249370F482E62BA41462",
INIT_06 => X"B250442BC81001E1870223FC0BF7F11507C423FE33C078F803F19F00E936721D",
INIT_07 => X"00011080012460050E700080EF020408EC8CFA01122149FF700200665A35D260",
INIT_08 => X"2BFD055040A452000443FF00007906464068406C31F84000000831FA1028575A",
INIT_09 => X"805FD017102690AA694551FE30444681E0820AD40201423FC00122C493500172",
INIT_0A => X"0600002AFFBE2330815568A8AD6ABC02A02A0B0CCB463B4C0748A720B1EA4C00",
INIT_0B => X"0850400A11414C005005000B51158936D20601A98A10200308A002E240010BFC",
INIT_0C => X"05928020194918A22A2268C81A32068C81A32068C81A32068C81A99034640C00",
INIT_0D => X"058102C48970541944B20FA1580561D040406305587A158046282000DBFFF13D",
INIT_0E => X"000000028040890327DCD28928324400DFFFF0001F1F0050342D42A086040B02",
INIT_0F => X"F60000000500802010000A000000000000022A0000141EC0000000A01000507B",
INIT_10 => X"00000000000004C0000082010A700000000000006800283D80000001402000A0",
INIT_11 => X"2200E4000000000000000442040004020001800000000000010D000010401A0E",
INIT_12 => X"08800000000801C040A6120000001540409C2200000015441DAC800010100000",
INIT_13 => X"0000000001019600081027084000000956000810298480000009560002200000",
INIT_14 => X"800088000021000000000201D800088000561400000000002358000088000A74",
INIT_15 => X"00802594A282C0000033010FB181E00020400000000819060000000000002305",
INIT_16 => X"C0B02C0B02C0B02C0B02C0B02C0B02C4B12B312912831A27FCFE7FFB175B6FF8",
INIT_17 => X"0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02",
INIT_18 => X"B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C",
INIT_19 => X"BBCF9F96EE7FFDF7FE783FFDFFEA0C00602FFFFFFFFFFFFFFFFFC0B02C0B02C0",
INIT_1A => X"EFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEEBAEBAEBAEBAEBBFFDF9FBEFFFFFFE",
INIT_1B => X"BFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFBEFB",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000FBFDFEFF7FBFDFEFF7F",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_3,               -- Port A enable input
WEA      => wbe_a_lo_1024_3(3),               -- Port A write enable input
DIA(0)   => data_write_a(29),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_3(29),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_3,               -- Port B enable input
WEB      => wbe_b_lo_1024_3(3),               -- Port B write enable input
DIB(0)   => data_write_b(29),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_3(29),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_30_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"F7FFBFFEFF9FE1F7FFBFFFFDFFD0000000000000000000000000000000000000",
INIT_1A => X"9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7AFBD75F5FDF7DF7F",
INIT_1B => X"F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE79E7",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000003F9FCFE7F3F9FCFE7F3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_3,               -- Port A enable input
WEA      => wbe_a_lo_1024_3(3),               -- Port A write enable input
DIA(0)   => data_write_a(30),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_3(30),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_3,               -- Port B enable input
WEB      => wbe_b_lo_1024_3(3),               -- Port B write enable input
DIB(0)   => data_write_b(30),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_3(30),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_31_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"129000008004A00804A40000400800020000000C005FEA005800200400050100",
INIT_01 => X"255FF18019700810180065FFFC0040801E80258CA2951C2200EC0906A0804140",
INIT_02 => X"E0000000000000011000550FDFF0FFFFF0007F1FC200000044000000000817F0",
INIT_03 => X"0000024210A30024210A3001002220C06044469200040154482000408400043F",
INIT_04 => X"602D0FFC2420000E003D80080955FF8E1ECA8E2D400340FE870060842100B030",
INIT_05 => X"0213100040F8A3F8FDBF944DC0FDC001D1CB6904A061EDB6D4C30490281831C1",
INIT_06 => X"6FC000830007C202060445F1F0D25E4207A099F0E303F0E07FE19C7F80402412",
INIT_07 => X"0000200000000000000001100004081001103107000185FF0000C0849673F6C0",
INIT_08 => X"1BF27A00000000000883F47FC800080002008000000820440000100220489020",
INIT_09 => X"011F07E013EFBC06FBA009F8E00120038F3CF82C44630C5D1FC002CCE0808248",
INIT_0A => X"61FF0C06C48BC801600000000001A1F00110101092CE7ED81CF0004012288000",
INIT_0B => X"11DCCC31222730048620C4382204A608142002A440492530C401049020221BF8",
INIT_0C => X"0888066187448380E00C10030400C10030400C10030400C10030600608018210",
INIT_0D => X"080204010200418301208480800D02D00040100240A808008840800405FF8640",
INIT_0E => X"0004001D000180780CE386106100C4043FFD03FF101D40008001304018081004",
INIT_0F => X"000008003A000217A0040000010003E02000160201E040000100074000478100",
INIT_10 => X"00010001DC00000810035C0400000200001DC0000063C0800002000E80008F02",
INIT_11 => X"00000000002801E1A00000801C0202F40080000800007B00000302006E808000",
INIT_12 => X"0000007E00000607810000001E000087810000001E000081846282010A211AA0",
INIT_13 => X"00001BC00000740401E0400000070800340401E04000000780003404045D0010",
INIT_14 => X"01011740040000001F8000025010116C080000000085C80000C8100947008000",
INIT_15 => X"FF800C609C06D082000A03200806A040019481D4000000000801E0D00001001D",
INIT_16 => X"010040100401004010040100401004010060C040040C200950402090128057C3",
INIT_17 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_18 => X"0040100401004010040100401004010040100401004010040100401004010040",
INIT_19 => X"00000000000000000000000000001000802FFFFFFFFFFFFFFFFF810040100401",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_3,               -- Port A enable input
WEA      => wbe_a_lo_1024_3(3),               -- Port A write enable input
DIA(0)   => data_write_a(31),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_3(31),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_3,               -- Port B enable input
WEB      => wbe_b_lo_1024_3(3),               -- Port B write enable input
DIB(0)   => data_write_b(31),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_3(31),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_0_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"ED39BA795990D275FB4A6E96ACC4731DEA4598B0AFB54867F6EE4618C3749803",
INIT_01 => X"8AA0047D8607944AC7DA180001ECA2444042106208408208C20022E9173734B3",
INIT_02 => X"1A7DDD79F9A73E6CCA7DAAF00001000008478020113D98E382FEDF333027C80F",
INIT_03 => X"75D341110C58F31110C58F32A208921F8051500147A0E4AB3493FB3A01EBE240",
INIT_04 => X"86424001531009B100425A97B2AA0001E03501D0A39C8F0078420001106D0C4C",
INIT_05 => X"BCC8CA2EBF03400700402BB20F00239E20341699198600000B08694B16434804",
INIT_06 => X"103FB860B2800161F8432200012DA185F80F24081C3C0707800E600056881308",
INIT_07 => X"B24197ABCDA467F9A73E6CCAFDC3870EEEEC44E2BDFE220094D03022210C011C",
INIT_08 => X"240581B5695EAA80262C080032BF07C7C1FC3F8E94F65B11555EAFFC1C306758",
INIT_09 => X"7E40000BEC004170040DB60017FED1CC0001045002984202003DB931192D60A5",
INIT_0A => X"120071411A74315881A28C141118000C5A85A60444210123820B43B40804674D",
INIT_0B => X"0820008E514045BB514F0106D1D8599581D3A958BC104A89215AC14C48898403",
INIT_0C => X"C261C01C48B1584A0CA3E2687A9A1E2687A9A1E2687A9A1E26870CD061343885",
INIT_0D => X"D274E93A758FA8683AC54B287522E10A74AF4AA59C568752662F5AC218000002",
INIT_0E => X"FF83C002783A0904231C70470C7E0B92800224008AE09FAD4BD48D1FC5D3A4E9",
INIT_0F => X"5BFF078004F075885DFBF7E15C06101C55E921F1F80FAB7FE0F0009E0E903EAD",
INIT_10 => X"F12E0380231F13978FF023FAFDBD9870380230F2D6081F56FFC1E0013C1D207D",
INIT_11 => X"DE7F263C0C8700125C0F8F3C43F1F10BBF7EFC61E01804E1E6C8F8FE807F67FB",
INIT_12 => X"02BE00017C17C1007E5E2E3081C5AC007E6F0E3081C5AC44418D65FE45DEE55B",
INIT_13 => X"61E0042786F103E9F01F9BC3C120C5A703E9F01F978B8C20666703E9F8A0FFED",
INIT_14 => X"FA7E283FFB414F80005F05F10FA7E283F78F6511C048278DCA174FF038FF15B4",
INIT_15 => X"0066A20B61692F293185D8D724E15D3FCC6B7C236FE0691B0700132C1F0EF880",
INIT_16 => X"3A4E93A4E93A4E93A4E93A4E93A4E93A4F942F92E9628540AD2A91442525A000",
INIT_17 => X"A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E9",
INIT_18 => X"4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93",
INIT_19 => X"55F3898E09B56C74DAB15D1CF13501AA495000000000000000003A4E93A4E93A",
INIT_1A => X"082082082082082082082082082082082082082082082082082084E41DC71C71",
INIT_1B => X"E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F82082",
INIT_1C => X"FFFFFFFFFFFFFFF94A5294A5294A5294A5294A52800003E1F0F87C3E1F0F87C3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"3060C183060C187FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"BDEBA0000000000000000000000000000000000000000000003060C183060C18",
INIT_28 => X"168ABA002E82145085155545F7AA975EFFFAABDE00FFAEBDFFF5D2EAAAAAF7AE",
INIT_29 => X"7FFFE10005542145557FD5545FF8000155087FC0155F7D168B55007BFDF45085",
INIT_2A => X"7FFC0010080017555555568AAAFFFFD7545AA8028A00A2802AABAFF8028BEF5D",
INIT_2B => X"FF842AABAA2AE95545FFD168ABAF7AEAAAAAA2FFFDF4500043FE105D2E954BAF",
INIT_2C => X"5007FD7400550415410002E974BA5D5168A00A2D142155005142010FFAE820AA",
INIT_2D => X"FFF780000BA007FE8AAAFF803FFFF5D2A821550000000BA007FD55FF5D7FC014",
INIT_2E => X"000AAFBEAA00007BFDFFF082EBDF455D5142000082E82145FFD17DFEFFFD168B",
INIT_2F => X"DFD75D2AA8A80EA8E2FE3F000000000000000000000000000000000000000000",
INIT_30 => X"68B551475FAF6D1C556F0AA1C24AABEA495FC716F002A975FFE3AA95E00EBAEB",
INIT_31 => X"42A0070071C50BAFEF1FAE0016D56A16D557BC257D415E0216FA3F1E8FC0145B",
INIT_32 => X"8010E004924874825D7FEAA85487FD24AFE3D02DAAAE12BD5545A2803AA00005",
INIT_33 => X"120155EA568E870BAEB8A05A2AEA8B50F55A2F150005A3A438BD04AFAB8F550A",
INIT_34 => X"545E055FFBE81D0BE8EA8A3AA05A2A5504001C74BA42A1571E8028E3DB7816D0",
INIT_35 => X"A5C7E3DFFFE90B45B47ABA497A82FFAFD2A82485FD2415A105C21451ED42A002",
INIT_36 => X"00000000000000000000B55EAAA100AA1D0F6F480B6A555A2A57A002A3D5FDB6",
INIT_37 => X"5EFAAAAB5E1AF3AABFF45592E88A0AFE80A8B0A0000000000000000000000000",
INIT_38 => X"65F520EBE9EF67D7BEA1FD5D556ABEF5D557FEBA55022A3F70C6B405F4D2AE97",
INIT_39 => X"C114728007521170821CE0FDE69411A8DED57CE1055555E5F58EFFC01FE2CACB",
INIT_3A => X"42341D5DEEBEF55080034E0A592A4AD0079C75D6070CC5CBB0280C029ABAA3EB",
INIT_3B => X"7F353AAF6C77F7F20D968BF57812A95E02A2AAB5EB0F280800EFAEE9F5D18F31",
INIT_3C => X"C91565455C141E41887D58AC448B69C30E02116220415A9540AA854140A0A204",
INIT_3D => X"DE6BE93172D7D625B556EEAB157ABEBE1B4D792A4AD1183454180DD3FDCAAAB7",
INIT_3E => X"F0000001FF0000001FF0000001FF0000001FF01EABC4B8014174FF7DA80F52FE",
INIT_3F => X"FF0000001FF0000001FF0000001FF0000001FF0000001FF0000001FF0000001F")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_3,               -- Port A enable input
WEA      => wbe_a_hi_1024_3(0),               -- Port A write enable input
DIA(0)   => data_write_a(0),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_3(0),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_3,               -- Port B enable input
WEB      => wbe_b_hi_1024_3(0),               -- Port B write enable input
DIB(0)   => data_write_b(0),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_3(0),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_1_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"212C001411984004084D000508C53810A03D1450E839B003342114428A000803",
INIT_01 => X"00000019400B100A8196000000CC004400400002000000000000028001340000",
INIT_02 => X"052137AE8031800C0044009000000000061800001CD4019802AD04CCCFC20004",
INIT_03 => X"04514108C60C21008C6042108400000201440020505100000043C30E10E9F000",
INIT_04 => X"02104001011DEFE088805681920000008000004001900800004002108C280008",
INIT_05 => X"040002340105000200000000080001900010000108040000000008411600401C",
INIT_06 => X"1034001042800808201000000001000820020000102000040000000000800180",
INIT_07 => X"64BF81A15EDFDE8031800C00843060C19E030022103600000450020800040004",
INIT_08 => X"00008004691687AA840008000090248CC84E000046000311555521F183060AC5",
INIT_09 => X"0820800D08100171000DB000154440C800400500000852020011200201012021",
INIT_0A => X"02000040001000880A2A04445004000102002041000001008208001440004140",
INIT_0B => X"4820018A1140440078050040511000102000A008183000010002404400000000",
INIT_0C => X"1000C80008000C030030880C2A030A00C28030A80C2A030A00C28018D4061401",
INIT_0D => X"10040802050080200284401C0022880F009E08008205C0020118088018000000",
INIT_0E => X"0F03C00280000000420860C60C0C0B92C0000000004000010042000040102008",
INIT_0F => X"001E078005000108400005E11C0610000000288058000003C0F000A000100000",
INIT_10 => X"F10E0380000000C202300000008D187038000000480800000781E00140002000",
INIT_11 => X"806302380C870010000004400100110800007861E0180000000C400680000001",
INIT_12 => X"023E00000000018000580C308000050000610C30800005000215006800000101",
INIT_13 => X"61E0000000018100B0001843812000014100B00016030C20000141002880026D",
INIT_14 => X"400A20009B404F80000000018400A20044096111C04000000304026000501580",
INIT_15 => X"0046820040082300218450C2800010094000482141E060190700100000002200",
INIT_16 => X"020080200802008020080200802008020080008008600500A82A1100A8000000",
INIT_17 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_18 => X"0080200802008020080200802008020080200802008020080200802008020080",
INIT_19 => X"81328A46BABEFC54A0810C7452B4428A14000000000000000000020080200802",
INIT_1A => X"AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA28A28A28A28A2A8218D2C0C924925",
INIT_1B => X"E974BA5D2E974BA5D2E974BA5D2E974BA5D2E975BADD6EB75BADD6EB75BAAAAA",
INIT_1C => X"FFFFFFFFFFFFFFFD8C6318C6318C6318C6318C63000002E974BA5D2E974BA5D2",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"70E1C3870E1C387FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"5555500000000000000000000000000000000000000000000070E1C3870E1C38",
INIT_28 => X"EBDF455D2EAABEFF7FFE8BFF5D0002155557FFFFFF007FC21EFA2FFD74AAAAD5",
INIT_29 => X"AA95400552AAAABAFFD1574105D7FD75FFAAAA800AAF7AA974BAFFFBE8B45F7A",
INIT_2A => X"0517DF555D2EAAA1055000015500557DF45AAD1400BAA2AE801550051555EFF7",
INIT_2B => X"FFD540155557FD5400F78028BFFFFFBEAB55F780020AAAA80020AA082EAAB550",
INIT_2C => X"AFF842ABEF5D517DF55552A974AAF7AE820AA0851574BAA2D1574AA5D7BFDEBA",
INIT_2D => X"EFAAD1575EF557FFFE10557FFFFFFFFD56AAAAFFFFD7555AAD168B45AAAEAAAB",
INIT_2E => X"0005D7FFDF4500043FE105D2E954BAF7AE80010082A97410557FEABFFAAFBE8B",
INIT_2F => X"51C7A2FBD5490BFD1C056A000000000000000000000000000000000000000000",
INIT_30 => X"974BAF7FFEFB45FFAABDF55492AA8BC2EBDFEAF7F1F840017D4975D2FEF147FC",
INIT_31 => X"080BEF495FC71D54124924385FAAA8AAAE3D145410F7F1D55D71C002DABAEBAA",
INIT_32 => X"002D082082AB8B6DBEDB7DF7F540E2AE85028B40155145F7AF6DBED5450AA1C2",
INIT_33 => X"78E021FF1471FDEAAFFD56F16D5571D2E28E38E0216FA2D1E8E80140F45082B4",
INIT_34 => X"A2DA3FB7DAAD4AAAAF487BC70BFA97F7AF6D417E92482BF84020BA495557E3FF",
INIT_35 => X"55554ADBD7A2FFC7BEFF6FFD7FC7002FD74951D71EDFFABFD16FAAAE92BD5545",
INIT_36 => X"00000000000000000000547AB8F550A8010E00492487482FFFE82A85EBAE2FFC",
INIT_37 => X"1EF005162BEF047FD5545AAFBF7400FBF9424F70000000000000000000000000",
INIT_38 => X"714F8338AAAA1D0AE974AAF7FFFDF55F7AABFF55082CA8B4DF6C1E8F5E540002",
INIT_39 => X"EABEF75550ACBB7582225FF5843404547184164AA5D2EBEEB0A2D555410D3555",
INIT_3A => X"FEAAEB083BC1000FF8409000512AEABFFDF79DCBF755962010BDCBBC21455D7F",
INIT_3B => X"801F8BA0C57740BDAA0688E5405D57D412F7D55F5E50C7F401BAAE8403CF5A3F",
INIT_3C => X"5D16BABAA3EBC3157ABD5FFE55F2AA9FEAFDF7F431A9F7FFE81FF013A8001AFF",
INIT_3D => X"FB863550229BCABEB7DA403FFFDA2FBF7FED2C7F955445079E280A00C56145EF",
INIT_3E => X"0000000000000000000000000000000000000596EBEF55080034E0A592A4AD00",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_3,               -- Port A enable input
WEA      => wbe_a_hi_1024_3(0),               -- Port A write enable input
DIA(0)   => data_write_a(1),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_3(1),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_3,               -- Port B enable input
WEB      => wbe_b_hi_1024_3(0),               -- Port B write enable input
DIB(0)   => data_write_b(1),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_3(1),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_2_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10E006600180111284380310006289800480032283E000A34301002001A0817",
INIT_01 => X"0005A00810790848048044A54E404350404000720885800802000906E4910200",
INIT_02 => X"407004208400408044C600C50AA055254010541A110222841200000002402544",
INIT_03 => X"0600011004182401004102408C28414043101000408118000145840440F5C415",
INIT_04 => X"5035855703A2900A000CD3088400F40688C9844409060850925E58A4081A0221",
INIT_05 => X"0200840D1021A15AC50494894850890540D1E12020C6E510818500440A280090",
INIT_06 => X"113044094002801020440090A8011A1224AB9380552102442884882A20004097",
INIT_07 => X"000100880004428400408044860000008C022402102100AA40004404B5075460",
INIT_08 => X"15C23440408C862A2A12382A8A5244145048C06085008010141521F000001240",
INIT_09 => X"400582B9033AA0E7AA4110B0506744810554542450694E710A836188C2C00222",
INIT_0A => X"443518360012C2210B020414109130A28038188096A06B8C120CA440A9C00802",
INIT_0B => X"1345E53300EC68005605002964AF222A5704004D080211121C80024200821780",
INIT_0C => X"181080C1110C882202211488452213C88472213C88472213488441109A442231",
INIT_0D => X"008204440210091341208041000810C00000300220201800A908000038AD0284",
INIT_0E => X"00040002804180300E88D28D206A40000554815500481440300000C44A081100",
INIT_0F => X"000008000500828700000000010000000002380000A00000010000A010050000",
INIT_10 => X"00010000000004CA000214000000020000000000684280000002000140200500",
INIT_11 => X"000000000020000000000442100002840000000800000000010C000026000000",
INIT_12 => X"00000000000805A4800000000000152300000000000015801272000100210020",
INIT_13 => X"000000000101C00000C000000000000940000120000000000009600004050000",
INIT_14 => X"0000130000000000000002018000106000000000000000002380000141000000",
INIT_15 => X"55000190000000000002000280000000011080C0000000000000000000002310",
INIT_16 => X"40902409064190641906419024090244902A9003004800415120D4A190804241",
INIT_17 => X"0900409004090641906419064190240902409024090641906419064190240902",
INIT_18 => X"9044090040900409004190441904419044090040900409004190441904419044",
INIT_19 => X"75960040138D70C030B51C50C7D100A2052F81F81F83F03F03F0419044190441",
INIT_1A => X"0410410410410410410410410410410410410410410410410248602081659659",
INIT_1B => X"5128944A25128944A25128944A25128944A25128944A25128944A25128941041",
INIT_1C => X"FFFFFFFFFFFFFFFE1084210842108421084210843FFF825128944A25128944A2",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"7FD5FF555815607FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"2AA000000000000000000000000000000000000000000000007FD5FF55581560",
INIT_28 => X"FC21EFA2FFD75EFAA8415410AA8415555087BFFF55A2AA800BAFFAE954000800",
INIT_29 => X"84155EFA2AEBDEAAA2FBEAABA5D7FE8B555551421455D0002145552EBFEBA007",
INIT_2A => X"2AEBDF555D2E954BAA2AA974BAFFFFE8B45552EBDF45FFAEAABFFF7FFE8B55F7",
INIT_2B => X"AAAAAAAAAFFD1574105D7FFFF555D2AAAAAA5D2E820BAA2FBEAB5555557DF55A",
INIT_2C => X"50055575EFFF84021555D043DEAA5D04021EF557FC21FFAA8428BFFAAAA954AA",
INIT_2D => X"10085568A00FF80175FFA2D17DFEFF7800215500557DF55AA80001FFAA800015",
INIT_2E => X"0005D00020AAAA80020AA082EAAB5500517DF555D042AA10A284154005D00154",
INIT_2F => X"00AAFFAA9543A080038A2A000000000000000000000000000000000000000000",
INIT_30 => X"0017D5D20B8EAA007FC51C7A2FBD55D2BE800042AFE8E1557D0075D2F45BEAA8",
INIT_31 => X"AA8BC7EBDFEAFEFFD00105FFBC20BDEAAA2FBF8AAA557BE8B6D5D5FFABEF4904",
INIT_32 => X"FFEFB6D555578F7DB6A0BDF7D480E174BFA02A974BAF7F5EFB455D2ABDF55492",
INIT_33 => X"ED1FDE90E3A497492B6AAADAAAE3D155E105571D55D71C002DABA5524820BAB6",
INIT_34 => X"BE8F401D7B6A0001470155C51D0092A071555D5E3AE821D00001FF0871C016DB",
INIT_35 => X"5BE8555400550A38428007FED000E3DA3DFD5E3DFFFBD5A38A021551C5F7AF6D",
INIT_36 => X"00000000000000000000410F45082B4002D082082AB8B6D1C5B7DF7FF78E075C",
INIT_37 => X"5EF005560B55F7AA800AAF7AA954AA00042AAA20000000000000000000000000",
INIT_38 => X"ABEF057D68F5F5A00021EF55042AAAA007FD5555AAFBD7545FBB8020A3F7AE97",
INIT_39 => X"7DF55D7AABFF5428ACA8F45A6C1E8F5EFF84165EFF7802BAB0A2FFEAABA557BE",
INIT_3A => X"CA8AA80800020AAF7FBFFFEF04552ABFFFF841FFE75CA882108202E974AAF7D5",
INIT_3B => X"00151FF0C57401E5F3D1E00A1A884174A8FFAEBFEB0A2D55541051555694F002",
INIT_3C => X"2AA801455D7FE8BFFF680800FFF7AAA155F595542455512A975455D3AA8A0055",
INIT_3D => X"5D79FCAF774AE005BE7895554005D2A8A0B882FFFFE10AAAAAB755A66B6AF56A",
INIT_3E => X"00000000000000000000000000000000000000C3BC1000FF8409000512AEABFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_3,               -- Port A enable input
WEA      => wbe_a_hi_1024_3(0),               -- Port A write enable input
DIA(0)   => data_write_a(2),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_3(2),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_3,               -- Port B enable input
WEB      => wbe_b_hi_1024_3(0),               -- Port B write enable input
DIB(0)   => data_write_b(2),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_3(2),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_3_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"210C00A20020000108430020001600B8156021104940741B3530400E02B92203",
INIT_01 => X"014C9BCA58B1296D24A402C992500B69404040028804A0080A000416A8D90A08",
INIT_02 => X"C12026A484318004404405C9C66E331352180D468B8203980300204442E02B34",
INIT_03 => X"04000748D60D24648D60524C88804D0215011020D15018148040C10A70E1D58C",
INIT_04 => X"18283333240FE41244187308C9104D70944852640901083801750EB0A418C220",
INIT_05 => X"0613142D01912CC2A1B4140528348900C612A104201C689044340ED413A07649",
INIT_06 => X"119000034019881822104C5E68035250A222829710A0A02C18C01A9920842413",
INIT_07 => X"402F00AB0016CA0431800444841020509D038B021230C1990001C644C8273200",
INIT_08 => X"16905000408482088290E8E64010248C4A5AA840C2000110001521F0810A92E7",
INIT_09 => X"0003CE6581BD016342A951AB146C4480530C3B2A8088D3542651670200C1826A",
INIT_0A => X"00735D36209A8A20020894004284B660821030C8990467401218004041020002",
INIT_0B => X"512445B740457154562F957CC08B00093700080D0A4851001D8302D20A0A1530",
INIT_0C => X"00508650008008021021A40861021840869021A408610218C0869810D6043095",
INIT_0D => X"1C8508438450801043A08090380A8834207007022209038080190000999C8F84",
INIT_0E => X"000400200000C0002A48A206204C4205F3304B33004C0041006240140A1C310A",
INIT_0F => X"0000080040000083800400000100000000008400018040000100080000510100",
INIT_10 => X"0001000000000800000244040000020000000100002A0080000200100000A702",
INIT_11 => X"000000000020000000200000080002C000800008000000000022000006808000",
INIT_12 => X"0000000000000A2281000000000040A3810000000000402001400000022002A0",
INIT_13 => X"000000000004200001C0400000000010200001C0400000000010000004490010",
INIT_14 => X"0001070004000000000000060000104C08000000000000001000000903008000",
INIT_15 => X"CC004050CA0C00020220200070040000010401C4000000000000000000100008",
INIT_16 => X"4310E4310A4210A4210A4210A4210A4210A8D0830A68010001B4DA881048061C",
INIT_17 => X"21084290A4210A4210A4210A4210A4210A4210A4210E4310E4310E4310E4310E",
INIT_18 => X"90A421084290A421084390E4310C4390E4310C4390E4310C4290A421084290A4",
INIT_19 => X"015303C0C78C706428A14C586291000A044001FFE000003FFC004290A4210842",
INIT_1A => X"2492492492492492492492492492492492410410410410412821600001249249",
INIT_1B => X"51A8D46A351A8D46A351A8D46A351A8D46A351A9D4EA753A9D4EA753A9D49249",
INIT_1C => X"FFFFFFFFFFFFFFFC00000000000000000000000038F56351A8D46A351A8D46A3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"55AB02055AB0207FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"420000000000000000000000000000000000000000000000007FFFAB57FFFAB5",
INIT_28 => X"A800BAFFAE9554508002AA00AA843DF55FFAA955EFA2D168B55557BEAA000055",
INIT_29 => X"002AB55AAAA955EF005568A00087BE8BFFA2D155410AA8415555087BFFF55A2A",
INIT_2A => X"AAABFF5508003FF555D0002145552ABFEBA007FC21EF007FD75FFAA841541008",
INIT_2B => X"082EBDEAAA2FBEAABA5D7FC0155005168B455D042AB45F7FFD741000042AA10A",
INIT_2C => X"FF7FBEAB55F7AABDEBA5D7FC2010A2D1575FFF7AA975555D2E80145F78415545",
INIT_2D => X"EF5555554AA087BC01FFFFAAAAB55552A954BAFFFFE8B55552EBDE00F7AEAABF",
INIT_2E => X"000082E820BAA2FBEAB5555557DF55A2AEBDF555D2E954BA002EAAABA002A821",
INIT_2F => X"FB7D5D7FEAA3808554203A000000000000000000000000000000000000000000",
INIT_30 => X"1557D1475FAF45BEAA800AAFFAA95578080038A2AA28E3AF55E3A0BA5D7AADB6",
INIT_31 => X"BD55D7BE80004AA1E8E2AB55B6A0925D7085F6AA10087FEABD7AAD57AEBAB68E",
INIT_32 => X"F5D0438140E2FA38B6AEBFF6D1D04AAFFA41040017D5D20B8EAA007FC51C7A2F",
INIT_33 => X"D0A901FFFF801557D1C20B8EAAA2FBE80AA557BE8B6D5D5FFABEF49002FB55FF",
INIT_34 => X"5D20BDE00EBAAA8BC7EBDFEAFEFAB8ABAE925D21C7010EADB525D7FFAE975C75",
INIT_35 => X"F002EADA921420871D74971D24820875C21D5EB8AA8FFF012A954BAFFF5EFB45",
INIT_36 => X"000000000000000000001C24820BAB6FFEFB6D555578F7DB6A0BDF7DEB8E125F",
INIT_37 => X"B55A28408145AAFFFFFFF5D7FEAABA0051400A20000000000000000000000000",
INIT_38 => X"AB55FAD568AA2AFAE975EF555168B55F7AA800BAF7AA955EF00042AAA2A2AEAA",
INIT_39 => X"2AAAA007FD55558A7BD7145FBB8020A35D2ABEF55F7800015F087FEAA00007FE",
INIT_3A => X"968F575D003FF55F7D5420BA5D2ABFEAAF7AE9DFF759A82AEF70800021EF5504",
INIT_3B => X"FFD5145FBAC9755F05040255FFD84175EF55002AAB0A2FFEAABA557BEA3EF057",
INIT_3C => X"82E974AAF7D57DF45552A3FF10AA8429F45A7D5EAF5FFBAEAAA10554155400AA",
INIT_3D => X"FF843FFE77C80825BC052ABFE10550415557085540000005156155FE90A8F5C0",
INIT_3E => X"00000000000000000000000000000000000005500020AAF7FBFFFEF04552ABFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_3,               -- Port A enable input
WEA      => wbe_a_hi_1024_3(0),               -- Port A write enable input
DIA(0)   => data_write_a(3),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_3(3),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_3,               -- Port B enable input
WEB      => wbe_b_hi_1024_3(0),               -- Port B write enable input
DIB(0)   => data_write_b(3),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_3(3),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_4_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A108400020612C80284210081034849800A00030300004833522C82D04A16002",
INIT_01 => X"2043998A1839284D1CA0650E1E504368403008418984014902030806A0D10200",
INIT_02 => X"C120042200000000044441CE01E80F00A49043118680008002000000026208E4",
INIT_03 => X"040001020019200020011209CC0164C060000000690111040144800042F5C403",
INIT_04 => X"7029AF0F81A00010CCA47700CC513CAC0D0B8E02010740E19754080108988021",
INIT_05 => X"02139405007133C0712244CD20F20105D583000020E9892201D304D42A9835E1",
INIT_06 => X"9190440300078002014405D9EE814C0284A883B6D7038AE079059B7800048092",
INIT_07 => X"000100AA0004408000000004840400008D200102503000782000C00C8025C000",
INIT_08 => X"00728A00408403220811991E02120C044058080004000001101121F220000260",
INIT_09 => X"811001E1185B38AD23C3707AD46440818F3CF80EC423CA7D01D123C80200816A",
INIT_0A => X"45810810A01B40216361056D6150F41200280001900439001FD8A00041400000",
INIT_0B => X"11FC88076266E800D605402962A820211500024808010512C40106D222223B14",
INIT_0C => X"0408804116040B02C02C500B0C02C100B0C02C100B0402C300B0401618058611",
INIT_0D => X"040200050200501301208482200D00D0A0408402C4282200A84800009B878680",
INIT_0E => X"00000020000100024AC88300300060090F0D830F00025400300204D018000804",
INIT_0F => X"8000000040000206A2000800000000000000950002E010000000080000588040",
INIT_10 => X"0000000000000808000554000200000000000100006D0020000000100000BB00",
INIT_11 => X"0000400000000000002000001A0002504001000000000000002280000D800800",
INIT_12 => X"0800000000000E2C802000000000408D801000000000408012440000200110A0",
INIT_13 => X"000000000004680003A0040000000010280003800800000000102800000B0000",
INIT_14 => X"000005C0002000000000000620000158000010000000000010A0000B00000200",
INIT_15 => X"C30146200400104002602600400000000294004000000004000000000010001A",
INIT_16 => X"0080200000008020000000802000000080080000004090014134DA101288C6DB",
INIT_17 => X"0802000000000401806010040180601004018060100000802000000080200000",
INIT_18 => X"8060180601004010040080200802000000000000802008020000000000008020",
INIT_19 => X"C0A28A063807E0500014063450404882846FFE000003FFC00000010040100401",
INIT_1A => X"AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA28A28A28A28A2934C8D0CCD145144",
INIT_1B => X"68341A0D068341A0D068341A0D068341A0D068351A8D46A351A8D46A351AAAAA",
INIT_1C => X"FFFFFFFFFFFFFFFC0000000000000000000000001FE32068341A0D068341A0D0",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"408102040810207FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"800AA00000000000000000000000000000000000000000000040810204081020",
INIT_28 => X"168B55557BEAB4500554200000557FE10FFFBEAA10007FD7410FFAA97555082A",
INIT_29 => X"55574105D2A800AA00043FEBA5D7FEAA00007BE8AAAAA843DF55FFAA955EFA2D",
INIT_2A => X"57BC00AAA2FFEAAAAAA8415555087BFFF55A2AA800BAFFAE9555508002AA0000",
INIT_2B => X"A2AA955EF005568A00087BE8BFFA2D17DE1000517FE10AAAAA8AAA002E975455",
INIT_2C => X"FAA8417410A2D140000F7FBC2010A2D157400AAAE974AAAAAA974BA08002AB55",
INIT_2D => X"EFA2AABDEAA087BEAAAAA2FBD54BA080002145552ABFEAA007FC21EF007FD75F",
INIT_2E => X"00055042AB45F7FFD741000042AA10AAAABFF5508003FF55F7D568A00552EA8B",
INIT_2F => X"5400F7A49057D0824850B8000000000000000000000000000000000000000000",
INIT_30 => X"3AF55F7A0925D7AADB6FB7D5D7FEAB7808554203A145178E00FFFBE8A101475D",
INIT_31 => X"A9557D080038AAA145157428492E8008200043FE925571EFA380871C7028A28E",
INIT_32 => X"AEA8A9200249056D4175C5092AAF5FDA38BE8E1557D1475FAF45BEAA800AAFFA",
INIT_33 => X"AA4954281C0E2FB55B6A0925D7085F6AA10087FEABD7AAD57AEBA08517DE00AA",
INIT_34 => X"007FC51C7007BD55D7BE80004AAFEDB42028EBFBC2028BED152438AAA092492A",
INIT_35 => X"AF7DF6AA00412EAABFFAA803DEBA0875EDA80BEF1C743840040017D5520B8EAA",
INIT_36 => X"0000000000000000000041002FB55FFF5D0438140E2FA38B6AEBFF6DBE84AAEB",
INIT_37 => X"A00FFFFEAA105D5155410FF84021EF0800154B20000000000000000000000000",
INIT_38 => X"DEBA0851574B2AAAEAAB55F78400145AAFFFFFEF5D7FEABFF0051400A25D5568",
INIT_39 => X"68B55F7AA800BAF7AA955EF00042AAA25555410BA082E8201000043FE005D517",
INIT_3A => X"568AA200557DE00AAAAAAA000804001FF005575408AA557FEB2FFAE975EF5551",
INIT_3B => X"D1550AAAA8002010F2AC154B25F2ABFF55F7800015F087FEAA00007FEAB55FAD",
INIT_3C => X"800021EF55042AAAA007FD5555087BD6145FAAC000A2A6FBC00BAAAFBC00BAF7",
INIT_3D => X"F7AEBDFF779A82AA43F7FBE8A00082EA8BFFAA843FEBA08517DE00F3F9574B30",
INIT_3E => X"000000000000000000000000000000000000008003FF55F7D5420BA5D2ABFEAA",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_3,               -- Port A enable input
WEA      => wbe_a_hi_1024_3(0),               -- Port A write enable input
DIA(0)   => data_write_a(4),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_3(4),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_3,               -- Port B enable input
WEB      => wbe_b_hi_1024_3(0),               -- Port B write enable input
DIB(0)   => data_write_b(4),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_3(4),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_5_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50DF4A0791B3FCB694379283C81FD996A091832102004A336A20E03C040C002",
INIT_01 => X"805FBDC69830A84D5C6A60000C34C26841280A00084000C8C212892EEAD53235",
INIT_02 => X"3B2026B578918E640A4F01CF8011FF0002080000082CA9998276DF7772C7C80D",
INIT_03 => X"37134108420D700084205702A4008A1D9100002171C0E0051554D93A11F5D140",
INIT_04 => X"8A41A0FC03A56DA000425A819410E3816C086198A388B702A8CA1210844A0C4C",
INIT_05 => X"B1808A062E8BC835F5E84532D708238A282F00A9291224800A2861490343082C",
INIT_06 => X"903FB8483A90581859050424100940825C6184401CDC451B860A6507160C4100",
INIT_07 => X"D26F068BCC96CDF8918E640E96D1A3469D6300E2FFEA27F8E4D23248130E259C",
INIT_08 => X"0BFA82E568442B2A082C0A7E3014250D49DA37A2420619000002AFF48D1222E5",
INIT_09 => X"3F005001E40969289429360416DCD1C46083030604B1CA20C03DF83B0A2C60A5",
INIT_0A => X"14613C71005A10492B888120288F480D58858449026145B3830F449449062B4F",
INIT_0B => X"11AC04934AC648BFD727C031E64170A137D5AA5C3E4B0F8A3C58C34C002290E3",
INIT_0C => X"CA29C6CC50384B6AC6AC86AB31AACA6AB39AAC86AB39AACA6AB3055643559C31",
INIT_0D => X"C673E33CF28F38603855401985228A0614BD30A0A2819852011E5AC2B87F9182",
INIT_0E => X"FF87C002F87A803E460B2516510CA594FF0044FFA4B08BAC4BB2CD0F09CF84E3",
INIT_0F => X"0DFF0F8005F0F5100DFFF5E15D06101C55EB29F1E00BE53FE1F000BE1E802F94",
INIT_10 => X"F12F0380231F17D78FC029FFF58D9A70380230F2FE0017C37FC3E0017C3D005F",
INIT_11 => X"FC7F023C0CA700125C0F8F7E43F1F001BFFE7C69E01804E1E7CCF8FC003FF5F1",
INIT_12 => X"023E00017C1FC1A4BFD82C3081C5BD27BFE30C3081C5BD00C02365D645CEEF5B",
INIT_13 => X"61E0042787F181E9C1EFD8CB8120C5AF41E9C18FD60F0C20666F41E9F009FFFD",
INIT_14 => X"7A7C077FFF404F80005F07F187A7D14BFFC96111C048278DEB074F9930FF9D80",
INIT_15 => X"C064014B8B652E2B3120C81284641D3E8DBF7D636FE860190700132C1F0EFB80",
INIT_16 => X"38CE1384E3384E338CE138CE1384E33C4E3ECE32E128882551349A1CBAA44103",
INIT_17 => X"84E3384E3384E3384E338CE138CE1384E3384E338CE138CE1384E3384E338CE1",
INIT_18 => X"CE138CE138CE138CE1384E3384E3384E3384E338CE138CE138CE138CE1384E33",
INIT_19 => X"F5E5BB4E7F7B9DB7FF3A1B6DB7E8410A8C000000000000000000384E3384E338",
INIT_1A => X"BEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEF9F7CFDFDDCF3CF3D",
INIT_1B => X"BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEFBEF",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000001711C7BBDDEEF77BBDDEEF77",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"FDFFF00000000000000000000000000000000000000000000080000000000000",
INIT_28 => X"FD7410FFAA97410082A800AAAAAE955450055421FFFFFBC0010AAD5574BA557F",
INIT_29 => X"7FD74000055574BA5D7FD7555A2D5575EF55517FF5500557FE10FFFBEAA10007",
INIT_2A => X"0002AABA5D2ABFFFFAA843DF55FFAA955EFA2D168B55557BEAB5500554200000",
INIT_2B => X"5D2A800AA00043FEBA5D7FEAA00007BC00AAAAAEBDF45A28428B45FFD168BFF0",
INIT_2C => X"5080028A00A2FFFDE00F7D57FEBAFF80174BAAAD1555EF555555555005557410",
INIT_2D => X"BA5D2E821FFA2D5554BA557BD75FFAA8415555087BFFF55A2AA800BAFFAE9555",
INIT_2E => X"00000517FE10AAAAA8AAA002E97545557BC00AAA2FFEAAAA082A97545F7D5420",
INIT_2F => X"7010BEDF524AA5571FDFEF000000000000000000000000000000000000000000",
INIT_30 => X"78E00EBFBE8A101475D5400F7A49043D0824850B8A2AE9756D145B401FFFFFFC",
INIT_31 => X"FEAB7D0855420BA1471D74380851524BA5571D757DB6D5525EF555178F6D1451",
INIT_32 => X"8A28B6DEBDF6DBEF1C0A28AAA5524BFFFFA28E3AF55F7A0925D7AADB6FB7D5D7",
INIT_33 => X"5555057D145152428492E8008200043FE925571EFA380871C7028B6AEBDF45B6",
INIT_34 => X"BEAA800AAFFAA9557D080038AAAA2FBF8E10EBD578EAAFF8415482BED1555EF5",
INIT_35 => X"81C209256DFFDF420BA552A821FFB6DF574A85575C55EFBE8E1557D1475FAF45",
INIT_36 => X"0000000000000000000008517DE00AAAEA8A9200249056D4175C50920875FDA3",
INIT_37 => X"5FF5D7BC21EFF7FBD7400F7FBC00BA55557DFF70000000000000000000000000",
INIT_38 => X"01FF5D5568BE7555568A00AAFFEAA105D5155410FF84020AA0800154B2AAAA97",
INIT_39 => X"00145AAFFFFFEF5D7FEABFF0051400A25551554BA0051400BA5551575EFF7D14",
INIT_3A => X"1574B2FFAABFF45FFAAAABFFAAFFFDFFF552EA8AAA55043DFF7AAAEAAB55F784",
INIT_3B => X"8002410FFD5575EF5555421E75555400BA082E8201000043FE005D517DEBA085",
INIT_3C => X"FAE975EF555168B55F7AA800BAF7AA955EF00002AAA2A2FBE8A00A2D16AAAAFF",
INIT_3D => X"0055554088A557FEB25D00021FFFFFFC00BA552A821EFFFFFD74BA5D51575F7F",
INIT_3E => X"000000000000000000000000000000000000000557DE00AAAAAAA000804001FF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_3,               -- Port A enable input
WEA      => wbe_a_hi_1024_3(0),               -- Port A write enable input
DIA(0)   => data_write_a(5),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_3(5),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_3,               -- Port B enable input
WEB      => wbe_b_hi_1024_3(0),               -- Port B write enable input
DIB(0)   => data_write_b(5),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_3(5),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_6_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10800B0061A01002840002C03002818000402322520070B313301C4389B2082",
INIT_01 => X"250041CA3839684D18A160000C52426841000000090800090210080008110200",
INIT_02 => X"0020042080010000044654C0000C008010000000001020900200200002620814",
INIT_03 => X"060881021088200021080200E4000A0891000020610111500104C00000F14400",
INIT_04 => X"0880000100000002000052288144004281C050400100280000C8100000080001",
INIT_05 => X"928080840001100A08009000280201000850E022401400002028214043410820",
INIT_06 => X"10100518090012122100C808049310002040000410A0001400000200120840D2",
INIT_07 => X"000100800004400001000000860408108C22000A502010074120044800040001",
INIT_08 => X"50000040D0C4E2088003FD01C01004044058082004000000000121F020408244",
INIT_09 => X"00BF17E9001205A5204911F814444080400100020000D200DFD16400C2A40AA0",
INIT_0A => X"04611C17849000022862A1596C8B5DF04834948900000100220C244840000880",
INIT_0B => X"03AD0413424E4044D665C070C22602291504400D084915020448114080201000",
INIT_0C => X"5E08864011088B22D22C008B0022C408B1022C208B0822C608B1111600458010",
INIT_0D => X"4251A12CD28A300429688001000800000020280204001000A00804309A002182",
INIT_0E => X"0000000280402400420800000000006200FC10002442042429324294014E8CA7",
INIT_0F => X"A40000000500800840000800000000000002280018001480000000A010100052",
INIT_10 => X"00000000000004C2003000010240000000000000680800290000000140202000",
INIT_11 => X"2000C0000000000000000442000001080001000000000000010C000280001804",
INIT_12 => X"08000000000801C300A010000000156000902000000015101200002800000000",
INIT_13 => X"000000000101800038002408000000094000386028040000000940000ED40000",
INIT_14 => X"0003B000002000000000020180002A24005010000000000023000060C7000A40",
INIT_15 => X"3F0280090321000040A410C28108000160008094000810040000000000002300",
INIT_16 => X"284A5284A728CA5284A528CA728CA52C4A5A0A32A300940101349A0408240818",
INIT_17 => X"9CA1294A329CA5284A728CA7284A5284A728CA5284A528CA728CA5284A728CA7",
INIT_18 => X"CA3294A129CA3294A129CA1294A329CA1294A3294A129CA3294A129CA3294A32",
INIT_19 => X"F5F78BCE7F8FF0F4FA955F7CF7F40A80145D55555556AAAAAAAAA94A329CA129",
INIT_1A => X"8E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E39B6CEDECDDF7DF7D",
INIT_1B => X"F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE38E3",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000001A1A33F9FCFE7F3F9FCFE7F3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"555FF00000000000000000000000000000000000000000000080000000000000",
INIT_28 => X"BC0010AAD5574BA557FFDFFF087BFDF45F7AA974AAAAAA97555F784174BAF7D5",
INIT_29 => X"515555508043FE00F7AA97555A2FBD7410AA8428AAAAAAE955450055421FFFFF",
INIT_2A => X"7D1575EFFFAA9555500557FE10FFFBEAA10007FD7410FFAA97400082A800AA08",
INIT_2B => X"0055574BA5D7FD7555A2D5575EF55517FF55A2AA97400552AAAB45082E80155F",
INIT_2C => X"500554200000003DE10FFD5401FFF7AAA8A10082EAAB45A2FFC2000007FD7400",
INIT_2D => X"10AA803FE105D516AABAFF843FFFFAA843DF55FFAA955EFA2D168B55557BEAB5",
INIT_2E => X"000AAAEBDF45A28428B45FFD168BFF00002AABA5D2ABFFFF087BD5545007BFDE",
INIT_2F => X"256DEB84104BAFFD1525FF000000000000000000000000000000000000000000",
INIT_30 => X"9756D145B401FFFFFFC7010BEDF524AA5571FDFEF1C7BFFF55FFA095482B6A49",
INIT_31 => X"4904380824850381C5B5057D1C003DE28F7A49057DAAF5D2428A2842AAAAA2AE",
INIT_32 => X"2AAFB451C2A8017DE3DF525FFFFA49756D145178E00EBFBE8A101475D5400F7A",
INIT_33 => X"2F1C50381471D74380851524BA5571D757DB6D5525EF555178F6DAAA49542841",
INIT_34 => X"AADB6FB7D5D7FEAB7D0855420BA1C0E3FE00E3DB471EFE3AAAAA00082EA8B6DA",
INIT_35 => X"F1C7BD057D1C71FFE10A28038E1049516AAB8FF8428FEFA28E3AF55F7A0925D7",
INIT_36 => X"00000000000000000000B6AEBDF45B68A28B6DEBDF6DBEF1C0A28AAA5524BFFF",
INIT_37 => X"F55F78017400F780001FFAA84000AAFFD1401E70000000000000000000000000",
INIT_38 => X"20BAAA8428AA2AAAA975FF5D7BC21EFF7FBD7400F7FBC00BA55557DFF7557BFD",
INIT_39 => X"EAA105D5155410FF84020AA0800154B2557FC01EF55043FEAAFF80021EFA2D14",
INIT_3A => X"568BE7AA80174AA082ABDF555D2A821EFAAFBC01FFF780155F7555568A00AAFF",
INIT_3B => X"AEA8A10082EA8BEFAAD5554B25551554BA0051400BA5551575EFF7D1401FF5D5",
INIT_3C => X"AAEAAB55F78400145AAFFFFFEF5D7FEABFF0051400A25D2EBFE10AAFFD55EFA2",
INIT_3D => X"552EA8AAA55043DFF7557BC01EF55557DE00AA842AA0000516AABAFF8428BE7A",
INIT_3E => X"0000000000000000000000000000000000000FFAABFF45FFAAAABFFAAFFFDFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_3,               -- Port A enable input
WEA      => wbe_a_hi_1024_3(0),               -- Port A write enable input
DIA(0)   => data_write_a(6),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_3(6),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_3,               -- Port B enable input
WEB      => wbe_b_hi_1024_3(0),               -- Port B write enable input
DIB(0)   => data_write_b(6),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_3(6),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_7_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10844B00482258A2842112C02450418800002300500030B313300C418992002",
INIT_01 => X"000009CA3839684D1CA0E0000E51424840000000080000080200080008510204",
INIT_02 => X"0120042086010000044600C00008000004100000000260900200000002402004",
INIT_03 => X"8628A10000082400000002408400080011000000610008000208C00000E14400",
INIT_04 => X"0911800100A000000000524084000040000050001140200100C8100000080102",
INIT_05 => X"0300812401011000000000002000114008008060441000000020024093000000",
INIT_06 => X"9190431C0D4010100000880804010010800000041080081000000200010424B2",
INIT_07 => X"000100AA0004408601000004860000008C02000A103010006928040800062481",
INIT_08 => X"84000048D484C20888000A0002120484C048007004000000000021F000000244",
INIT_09 => X"00A06009881201A520491004106C48A04040002400A15A208001650004001020",
INIT_0A => X"C99E1060201002044809C1040140A001004808810000459033189C0A400118A0",
INIT_0B => X"102000024040484050050041648A0041140C500B08821054C000264120000400",
INIT_0C => X"0404A083260E0832132011880462011880462051881462051881D31018C40620",
INIT_0D => X"0001000080001000813094801A8F80F00A600B52602801A88848011118003700",
INIT_0E => X"000003C007C002808228010410082042C000C000000004001002000400040002",
INIT_0F => X"A4000007800F80C840000800009864038A1200081C0014800000F001F0200052",
INIT_10 => X"00002C0E00E0E4004038000102400002C0E00E0D20100029000001E003E04000",
INIT_11 => X"2000C04031100E0403D0700300080908000100000661801E1900040380001804",
INIT_12 => X"0840878083E8003780A01043203A101780902043203A10082410082880000000",
INIT_13 => X"0601E0187900181035E0240806483248181035E0280410C8198818100DDD0000",
INIT_14 => X"0403774000201021E020FA006040376C00501022131210722060806D47000A40",
INIT_15 => X"00928A0002000110888600C032128201519480D40009902430160403E0E00506",
INIT_16 => X"01000000020080601802000000000405000A0020020081014134928820480010",
INIT_17 => X"0802018040000000006018020080200804010000000000806018020080000004",
INIT_18 => X"0000000001806008020000001006008020080001004008020080201004000020",
INIT_19 => X"0000000000000000000000000000400A004618618618C30C30C3000020180600",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000000B0840000000000000000000",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"1555500000000000000000000000000000000000000000000080000000000000",
INIT_28 => X"A97555F784174BAF7D5555FFF780155EFAAAEA8ABAAAFBFDE0055556AA005D04",
INIT_29 => X"55555EFAAFFFDFEFAAAAAAB455D556AA00FFAE95555087BFDF45F7AA974AAAAA",
INIT_2A => X"02EAAAAA082EA8A00AAAE955450055421FFFFFBC0010AAD5574BA557FFDFFF55",
INIT_2B => X"08043FE00F7AA97555A2FBD7410AA8428AAA557BFDFFF55003DFFFF7FBEAA000",
INIT_2C => X"0082A800AAF7AE975FFA28000010552EBDE00007BEAAAAA2D140000085155555",
INIT_2D => X"45087FEAB455D516AB55557BD55FF00557FE10FFFBEAA10007FD7410FFAA9740",
INIT_2E => X"000A2AA97400552AAAB45082E80155F7D1575EFFFAA955555D51574AAAAFFD55",
INIT_2F => X"AE105D556AA10410E17555000000000000000000000000000000000000000000",
INIT_30 => X"FFF55FFA095482B6A49256DEB84104BAFFD1525FFFF8E175C7A2AAAAA82A2F1F",
INIT_31 => X"F524AA5571FDFEF415B575D7AAF1FFFD7AAAAAFB7D495F6AA10E3AE905551C7B",
INIT_32 => X"003AFEFEBFBEAA001C2EA8A821C2EAAA00A2AE9756D145B401FFFFFFC7010BED",
INIT_33 => X"EDB470101C5B5057D1C003DE28F7A49057DAAF5D2428A2842AAAA497BFAFFF49",
INIT_34 => X"1475D5400F7A490438082485038F7A4905C7A28A070384120BDE100075EAA82B",
INIT_35 => X"D495150492BEF1D2555087BE8B7D555F6AB57417BC05D7145178E00EBFBE8A10",
INIT_36 => X"00000000000000000000AAA495428412AAFB451C2A8017DE3DF525FFFFA49756",
INIT_37 => X"555A2AEA8A10AAD568A00555168A10002E9754D0000000000000000000000000",
INIT_38 => X"8A10AAAE8215D557BFDF55F78017400F780001FFAA84000AAFFD1401E7FFAA97",
INIT_39 => X"C21EFF7FBD7400F7FBC00BA55557DFF7007BD5555AAD57DF55AAAEBDFEF007BE",
INIT_3A => X"428AA2007FE8BFF080028BFFAAFFEAA105D2EAAA005D2AAAA18AAAA975FF5D7B",
INIT_3B => X"043DE0000516AA10F7FBD7408557FC01EF55043FEAAFF80021EFA2D1420BAAA8",
INIT_3C => X"55568A00AAFFEAA105D5155410FF84020AA0800154B2FF8402145A2AA954AA00",
INIT_3D => X"AAFBC01FFF780155F7005140000FFD140145007FE8BEF557BEAB55087FC215D5",
INIT_3E => X"0000000000000000000000000000000000000AA80174AA082ABDF555D2A821EF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_3,               -- Port A enable input
WEA      => wbe_a_hi_1024_3(0),               -- Port A write enable input
DIA(0)   => data_write_a(7),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_3(7),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_3,               -- Port B enable input
WEB      => wbe_b_hi_1024_3(0),               -- Port B write enable input
DIB(0)   => data_write_b(7),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_3(7),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_8_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00000648E2840112C00000418000002700500030B3132000400812082",
INIT_01 => X"100008480009004C04A100000252024840000000180800080200010040110204",
INIT_02 => X"0020042000490000004600804008000005100000000024900200000002400004",
INIT_03 => X"0A0C33400008082400000080A4004B0891000020610112000040C00000E5C000",
INIT_04 => X"18800001000000000000512080000040800150400824280110C8100000120200",
INIT_05 => X"908084A10100100200004080280008240810802206940000012C214451610800",
INIT_06 => X"81B000080860109021400008040000202048020414A0021400040200322824C1",
INIT_07 => X"000000080004408049000004860000008402001A50208000630C040800062483",
INIT_08 => X"440000428644212280800A00021004044048002124000000000021F000000244",
INIT_09 => X"00004009001001010008100414644410400102228000D20080114502006409A2",
INIT_0A => X"000051312000042200294429148A4801C80C8C81000045907118040340020832",
INIT_0B => X"4020000240404140004D0544C4AA0001150410090302500011C813428A000400",
INIT_0C => X"46501090008820240240409000240009000240009000240009000120204808A5",
INIT_0D => X"42D1A168D09A301468402480004780F00140080860280004085904309A002196",
INIT_0E => X"00783FC00044340242280000000000020000C0000442106419120004034685A3",
INIT_0F => X"8000F07F800088A80000081EA2F9EC0000064004081010001E0FF00011104040",
INIT_10 => X"0ED0FC7E00000422201080000202658FC7E0000021882020003C1FE000222080",
INIT_11 => X"018059C3F350FE0C00000002A0040500000103961FE780000110010090000800",
INIT_12 => X"FD41FF80000830200021C1CF600012200010D1CF600012121600100810000004",
INIT_13 => X"9E1FE000010A1802100004343ED8000898021000087073D80008980200800002",
INIT_14 => X"0080200000BEB07FE00002086008020000209AEE3F300000246020200000620B",
INIT_15 => X"0088881903210000440610C8000A808040000208901786E4F0FE0C0000000166",
INIT_16 => X"685A1685A769DA368DA368DA769DA36CDA121A11A141800011309284002C0810",
INIT_17 => X"95A5685A1685A5695A368DA368DA769DA368DA368DA7695A1685A1685A5695A1",
INIT_18 => X"5A1695A568DA368DA369DA768DA1685A1695A5685A168DA369DA768DA368DA16",
INIT_19 => X"A4028A0A543EBC57A10A1E75D64108080468618618630C30C30C69DA5685A168",
INIT_1A => X"9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7BF3CCD8DF5B2DB2C",
INIT_1B => X"F87D3E1F4F87D3E1F4F87D3E1F4F87D3E1F4F87C3E1F0F87C3E1F0F87C3E79E7",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000006A6D4F87D3E1F4F87D3E1F4",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"155FF00000000000000000000000000000000000000000000080000000000000",
INIT_28 => X"BFDE0055556AA005D0415555080000000087BEAA10F7803DE00FFAEBFFFF0800",
INIT_29 => X"2AA8AAA557FC0010F780154105D7FC2145005155555F780155EFAAAEA8ABAAAF",
INIT_2A => X"7FFFFF55AA80155FF087BFDF45F7AA974AAAAAA97555F784174BAF7D5555FF55",
INIT_2B => X"AAFFFDFEFAAAAAAB455D556AA00FFAE95555AAFFE8A00552EBFE00F7D17FF45F",
INIT_2C => X"A557FFDFFF5504000AAAAAAA8B55F7D140010552E821EFAAAABDF555555555EF",
INIT_2D => X"55AA8028A00A2D57FF45557BE8A00AAAE955450055421FFFFFBC0010AAD5574B",
INIT_2E => X"000557BFDFFF55003DFFFF7FBEAA00002EAAAAA082EA8A00002AA8A10F784021",
INIT_2F => X"FE10F7AEBAFFF080A175D7000000000000000000000000000000000000000000",
INIT_30 => X"175C7A2AAAAA82A2F1FAE105D556AA10410E17555080E000280071E8A00EB8E3",
INIT_31 => X"4104BAFFD1525FF492EA8AAA5571C2000FF8A17400557FC015514555757DFF8E",
INIT_32 => X"2ABDE10EBDF7AF6DE3FFF8F7DB68A105D71C7BFFF55FFA095482B6A49256DEB8",
INIT_33 => X"AA0BDF6D415B575D7AAF1FFFD7AAAAAFB7D495F6AA10E3AE90555A2FBE8A3849",
INIT_34 => X"FFFFC7010BEDF524AA5571FDFEF550E00082B6A0AFB55F7D1420104124821D7A",
INIT_35 => X"01C2EA8A00F7800017DA2842FA00B6D578F6D557FFDA00A2AE9756D145B401FF",
INIT_36 => X"00000000000000000000497BFAFFF49003AFEFEBFBEAA001C2EA8A821C2EAAA0",
INIT_37 => X"0BA08556AA00AAAABFE00F7AEAABEF082E955450000000000000000000000000",
INIT_38 => X"21555D51575EFFFAA97555A2AEA8A10AAD568A00555168A10002E9754D082E82",
INIT_39 => X"17400F780001FFAA84000AAFFD1401E7082EAAABA5D5140010F7AE974105D7BC",
INIT_3A => X"E8215DA2FFE8ABA082ABFE00AAFBEABFFAAFBEABFFF7AA80145557BFDF55F780",
INIT_3B => X"D540000000402145AA843FFFF007BD5555AAD57DF55AAAEBDFEF007BE8A10AAA",
INIT_3C => X"AAA975FF5D7BC21EFF7FBD7400F7FBC00BA55557DFF75D2E82010F7843DF45FF",
INIT_3D => X"5D2EAAA005D2AAAA185D2AAAA10F780021FFA2803DE10FFD16ABFF5D7BFDE10A",
INIT_3E => X"0000000000000000000000000000000000000007FE8BFF080028BFFAAFFEAA10",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_3,               -- Port A enable input
WEA      => wbe_a_hi_1024_3(1),               -- Port A write enable input
DIA(0)   => data_write_a(8),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_3(8),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_3,               -- Port B enable input
WEB      => wbe_b_hi_1024_3(1),               -- Port B write enable input
DIB(0)   => data_write_b(8),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_3(8),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_9_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00018248A2840112C00002C18000002300500030B3132000400812006",
INIT_01 => X"400008000000004C0020000000100248413C0A61590001D90213C10008110204",
INIT_02 => X"01A0042080010000054600C04008000004100000001020900200200002420804",
INIT_03 => X"024003400008012400000010E4004B0891000020610310000144C00000F5C000",
INIT_04 => X"1801800100E000000000510084000040010050020810200000C8900000320200",
INIT_05 => X"918004311104100000000000200008100800002000100000002C234415610820",
INIT_06 => X"81B00008080010100000980804000008800042041080001000100200322C2481",
INIT_07 => X"0000811800044080010000058600000086020002502080006000040800062C80",
INIT_08 => X"0000004001D4618008800A00061004044048002004000000000061F000000244",
INIT_09 => X"000040090802009420409004104444084001022400214A2080014400026401A2",
INIT_0A => X"04000071200000A003CA294140200800C80C8C8100004590111C040040120800",
INIT_0B => X"12210002404848502847040164880021150400080222000200C8034200000000",
INIT_0C => X"4610088010080421021040841021000841021000841021000841010800420820",
INIT_0D => X"42D0A16C529A321068500484000500D10042080040284000084900001A002196",
INIT_0E => X"00000002804000004228010410082002C000C0002400046419120410034285A1",
INIT_0F => X"A00000000500800800000800000000000002290008001080000000A010100042",
INIT_10 => X"00000000000004C2001000000240000000000000680800280000000140202000",
INIT_11 => X"0000C0000000000000000442020001000001000000000000010C800080000804",
INIT_12 => X"08000000000801A7802010000000152780102000000015000600000800000000",
INIT_13 => X"000000000101900011E0240000000009500011E0280000000009500004DD0000",
INIT_14 => X"000137400020000000000201C000136C00101000000000002340002947000240",
INIT_15 => X"0080881901210000000600C280028000419480D4000010040000000000002304",
INIT_16 => X"68DA368DA1685A1685A1685A1685A16C5A121A13A141950051309284A82C0010",
INIT_17 => X"85A1685A1685A1685A368DA368DA368DA368DA368DA368DA368DA368DA368DA3",
INIT_18 => X"5A1685A168DA368DA368DA368DA368DA368DA368DA3685A1685A1685A1685A16",
INIT_19 => X"0157344CCCF48DE68A895C38E2540A8010100000000000000000685A1685A168",
INIT_1A => X"14514514514514514514514514514514514D34D34D34D34D28E1004039248209",
INIT_1B => X"D268341A4D268341A0D069349A0D069349A0D068341A0D068341A0D068345145",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000014D490D069349A0D068341A4",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"EAABA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"03DE00FFAEBFFFF0800155FFAAFBE8B45002A974AAAA803DFFFAA843DF45FFFF",
INIT_29 => X"7BFDE00A2FBD7400F7FBFDFFFA2AEBDE00AAFBEAABA080000000087BEAA10F78",
INIT_2A => X"055401FFF7AEAAA10F780155EFAAAEA8ABAAAFBFDE0055556AA005D041555508",
INIT_2B => X"557FC0010F780154105D7FC2145005155555557BE8BEF007FFDEAAAAD1555EF0",
INIT_2C => X"AF7D5555FFF780154AA5D2AA8A10F7AA974AA082E80010A2AAAAA10552AA8AAA",
INIT_2D => X"BAF7D17FEBAA2AEBDF45002EAAABA087BFDF45F7AA974AAAAAA97555F784174B",
INIT_2E => X"000AAFFE8A00552EBFE00F7D17FF45F7FFFFF55AA80155FF080400145FFFBEAA",
INIT_2F => X"8FC7BE8A3DF7DF7F5E8A92000000000000000000000000000000000000000000",
INIT_30 => X"000280071E8A00EB8E3FE10F7AEBAFFF080A175D7BEF1E8B6D002090482B68E3",
INIT_31 => X"56AA10410E175550871FFE00A2FBD0400FFF5FDFC7B6A0BDE38B6F5E8A92080E",
INIT_32 => X"7BFAE82A2DB555C71C5B451D7FFAAA8A38FF8E175C7A2AAAAA82A2F1FAE105D5",
INIT_33 => X"2AEADA38492EA8AAA5571C2000FF8A17400557FC015514555757D5D71E8BEF14",
INIT_34 => X"B6A49256DEB84104BAFFD1525FFFF84174BA5D20AAA00E3AA904BA142A87010A",
INIT_35 => X"7000400155FFFBEDA82FFD57DEBAAAA0BFF7D0024ADA921C7BFFF55FFA095482",
INIT_36 => X"00000000000000000000A2FBE8A38492ABDE10EBDF7AF6DE3FFF8F7DB68A105D",
INIT_37 => X"BEF080402000F7AAA8B55FFAABDFEFF7D16AA000000000000000000000000000",
INIT_38 => X"FEAAFFD16AA00082E820BA08556AA00AAAABFE00F7AEAABEF082E95545F7D568",
INIT_39 => X"A8A10AAD568A00555168A10002E9754D00517DE00A2FFC2000F7D17FF55FF803",
INIT_3A => X"1575EF555568BEF5D7FE8A10AAFFD55555D7FD5555FFAAA8AAAFFAA97555A2AE",
INIT_3B => X"AE800AA552A97400A2AEBDEAA082EAAABA5D5140010F7AE974105D7BC21555D5",
INIT_3C => X"57BFDF55F78017400F780001FFAA84000AAFFD1401E7FF80174AA5D0028A00AA",
INIT_3D => X"AAFBEABFFF7AA80145080002145F7FBFFE00FFD17FEAAA2803DFEF08043FE005",
INIT_3E => X"0000000000000000000000000000000000000A2FFE8ABA082ABFE00AAFBEABFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_3,               -- Port A enable input
WEA      => wbe_a_hi_1024_3(1),               -- Port A write enable input
DIA(0)   => data_write_a(9),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_3(9),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_3,               -- Port B enable input
WEB      => wbe_b_hi_1024_3(1),               -- Port B write enable input
DIB(0)   => data_write_b(9),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_3(9),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_10_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00018248A2840112C00002C18000202300500030B3132000400992006",
INIT_01 => X"254008000000004C002000000010026840000000080000080200010008110204",
INIT_02 => X"0020042000010000004455800008000004100000000000900200000002400004",
INIT_03 => X"020001021089000021081000C400090011000000610001540104C00000F14400",
INIT_04 => X"0811800101A00002000050088554004200C840000000200080C8100000000001",
INIT_05 => X"030080001000100800009400200000000840E020201000000024024001200020",
INIT_06 => X"81B00008080012120004CC080492500280208004148000100000020020042493",
INIT_07 => X"0000000800044080010000048404081085020002502000006000040800062480",
INIT_08 => X"100202400084410808000A00021004044048000004000000000021F020408264",
INIT_09 => X"010040090002008420401004144440004040022484214A2080110108C2C00320",
INIT_0A => X"04004166A48A0001080000000000080080181881000045901118044040020800",
INIT_0B => X"1201000200484910000F0105602622291404020902005002018002400A022000",
INIT_0C => X"0440001011808020120004801120044800120004801120044800110002400884",
INIT_0D => X"008000440210100041308480800F82F00040180260A808008848000018002104",
INIT_0E => X"000000028040000002280104100820020000400020000440100204100A000100",
INIT_0F => X"040000000500800800000000000000000002280008000400000000A010100010",
INIT_10 => X"00000000000004C2001000010000000000000000680800010000000140202000",
INIT_11 => X"200000000000000000000442000001000000000000000000010C000080001000",
INIT_12 => X"00000000000801C0008000000000154000800000000015000410000800000000",
INIT_13 => X"0000000001019800180000080000000958001800000400000009580002800000",
INIT_14 => X"0000A0000000000000000201E0000A0000400000000000002360002080000800",
INIT_15 => X"0080881000000000000600C28102800060000000000800000000000000002306",
INIT_16 => X"401004010040100401004010040100441020D0030008840051309A90BA884010",
INIT_17 => X"0902409024090240900401004010040100401004010040100401004010040100",
INIT_18 => X"1004010040902409024090240902409024090240902409024090240902409024",
INIT_19 => X"F546890A940FE0D3971243555205428290100000000000000000401004010040",
INIT_1A => X"8A28A28A28A28A28A28A28A28A28A28A28A28A28A28A28A29554199854514514",
INIT_1B => X"2B95CAE532994CA6532995CAE572B94CA6532994CA6532994CA6532994CA28A2",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000002718E72B94CA6532994CA657",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"FDE1000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"03DFFFAA843DF45FFFFEAABA007FC2155F7D155545AA80001EFAAFBEAB45557F",
INIT_29 => X"042AB55FFD168B55AA8000010FFFBE8BFFF78402155AAFBE8B45002A974AAAA8",
INIT_2A => X"AD16AABA002ABDE10080000000087BEAA10F7803DE00FFAEBFFFF0800155FF00",
INIT_2B => X"A2FBD7400F7FBFDFFFA2AEBDE00AAFBEAABAA2FFD741055003DFEFF7AA801FFA",
INIT_2C => X"05D0415555007FD74105555555EFF7FBC0145F78028A00A2D142155087BFDE00",
INIT_2D => X"55AAD168ABA002A975FFF7AEBDEBAF780155EFAAAEA8ABAAAFBFDE0055556AA0",
INIT_2E => X"000557BE8BEF007FFDEAAAAD1555EF0055401FFF7AEAAA105D042ABFF5D556AB",
INIT_2F => X"71D7AAFBEFB455D71F8E00000000000000000000000000000000000000000000",
INIT_30 => X"E8B6D002090482B68E38FC7BE8A3DF7DF7F5E8A92007BC217DEBDB55555AA8E0",
INIT_31 => X"EBAFFF080A175D700042AB7DEBDB6DB55BE8E05000EBFFE8BC7E38E07145BEF1",
INIT_32 => X"0A3DFD7F7A4821D7A2D16FA82142EB8E00080E000280071E8A00EB8E3FE10F7A",
INIT_33 => X"ED1421450871FFE00A2FBD0400FFF5FDFC7B6A0BDE38B6F5E8A92B6FBD541049",
INIT_34 => X"A2F1FAE105D556AA10410E175550071D54104951555D7EBF5C5155E3842AA00B",
INIT_35 => X"8410E2ABD749516FB55BED16FA820820955EFE3AEBDEAAFF8E175C7A2AAAAA82",
INIT_36 => X"000000000000000000005D71E8BEF147BFAE82A2DB555C71C5B451D7FFAAA8A3",
INIT_37 => X"1EFA2FFD7545AAAE97555A2FBFDF455D556AA000000000000000000000000000",
INIT_38 => X"8B45AAAA95545F7D568BEF080402000F7AAA8B55FFAABDFEFF7D16AA00087FC0",
INIT_39 => X"6AA00AAAABFE00F7AEAABEF082E9554500042ABFFA2FFFFF45F7AE97400AAFFE",
INIT_3A => X"16AA00FFFBD5400082EBFF45F78400155A2D57FE00552EA8A00082E820BA0855",
INIT_3B => X"D557555A2802AA10FFD54214500517DE00A2FFC2000F7D17FF55FF803FEAAFFD",
INIT_3C => X"FAA97555A2AEA8A10AAD568A00555168A10002E9754D085155410085557555AA",
INIT_3D => X"5D7FD5555FFAAA8AAA002AAAB4508557DF55F7D17FE000804155FFAAAABDEAAF",
INIT_3E => X"0000000000000000000000000000000000000555568BEF5D7FE8A10AAFFD5555",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_3,               -- Port A enable input
WEA      => wbe_a_hi_1024_3(1),               -- Port A write enable input
DIA(0)   => data_write_a(10),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_3(10),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_3,               -- Port B enable input
WEB      => wbe_b_hi_1024_3(1),               -- Port B write enable input
DIB(0)   => data_write_b(10),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_3(10),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_11_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A101C4B05A0034CA2840712C2D001419000002300500030B31B20084EC992002",
INIT_01 => X"90000986B83028491800E0000C26426040000000080000088200080802512224",
INIT_02 => X"1A2004205E010640024D00800008000004100000040EC090820018003241A00C",
INIT_03 => X"28639100000C5C00000045C08400C8001100000061806A001618C03001E54400",
INIT_04 => X"1A800001000009A0804059A190000040400040008058220008C8100000120D4E",
INIT_05 => X"02000E81080250010000002022000058080400000E1200000020004401000004",
INIT_06 => X"819435143F20101010001008040800B8100102041088011100022200000024B2",
INIT_07 => X"90640D280884453E01064002944180008402001295BA100022E4340800062D82",
INIT_08 => X"400000093204802200280A0012160585C1D808D004000000000323F40C102244",
INIT_09 => X"380040098010001100009204107C5950400000220080C200800900020C006827",
INIT_0A => X"80007100004016EA080801010000080D00200081000045B0511D289940103399",
INIT_0B => X"002000024040410A000D0104408810C115D9C008050042400100D04E88000002",
INIT_0C => X"00655010009264201200C7B421ED0C7B421ED0C7B431ED087B43176843DA1085",
INIT_0D => X"0401020080400A10012494881A4F80F209500BB2602881A488485C1318002000",
INIT_0E => X"6619A540124814800228010410082022C00040002020090020220C9600040802",
INIT_0F => X"ACCC334A802491600C587949B6D0141B4CC600D5761B1599865A500490B86A56",
INIT_10 => X"BAC845542056A61686EC81E3A6CB68AA2C622C9A251C352B330CB4A0092170D8",
INIT_11 => X"BCCAD0B5A81536080CC6B21A21B1FC09CB0F1076D4A200B2AD4068F4101639B5",
INIT_12 => X"4D2CC281E31AA0103AB8D5514066380804B268A2E060901204112566F10AC418",
INIT_13 => X"D551443C47281002540B2C9AAAA8662A1152B202AE3554403028115AA88201A1",
INIT_14 => X"548A20A0492A2724A0621620402A020141F172FB182A32AB6845AB6200251BC9",
INIT_15 => X"00C00A000200074044E6801832728080D00A380B753952C4877E0104DDE4D124",
INIT_16 => X"0080200802008020080200802008020480080022020081010124988800400010",
INIT_17 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_18 => X"0000000000802008020080200802008020080200802008020080200802008020",
INIT_19 => X"55062608804180C0B10A42104201400204000000000000000000000000000000",
INIT_1A => X"00000000000000000000000000000000000820820820820801C4149470000000",
INIT_1B => X"0000000000000000040200000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000007E0F0000000000000100800",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"000AA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0001EFAAFBEAB45557FFDE10082ABDF5508557DF45002ABDFFFF7803DE10AA80",
INIT_29 => X"AEBFF45FFAEBFEAA002A801FFF7FFE8A10A28000000007FC2155F7D155545AA8",
INIT_2A => X"2AABFE10082ABFFEFAAFBE8B45002A974AAAA803DFFFAA843DF45FFFFEAABAA2",
INIT_2B => X"FFD168B55AA8000010FFFBE8BFFF78402155AAD155555A28428BFF002ABDE00A",
INIT_2C => X"F0800155FF00557FF45557FC2010002A80010A2842AAAA007BFFF4500042AB55",
INIT_2D => X"FF5D00154BAF7FBE8BEFFFD540000080000000087BEAA10F7803DE00FFAEBFFF",
INIT_2E => X"000A2FFD741055003DFEFF7AA801FFAAD16AABA002ABDE10A2D168A10A284021",
INIT_2F => X"DFC7F78E3FE28B684070AA000000000000000000000000000000000000000000",
INIT_30 => X"C217DEBDB55555AA8E071D7AAFBEFB455D71F8E00002EBDF6D005B78F7D142AB",
INIT_31 => X"A3DF7DF7F5E8A92BEAEBFF7DEBA0BDEAA1C2A801C7E3FFEFA10B68407038007B",
INIT_32 => X"8A28BFF082ABAE10B6AAB8E280820B8FEFBEF1E8B6D002090482B68E38FC7BE8",
INIT_33 => X"07FF8F7D00042AB7DEBDB6DB55BE8E05000EBFFE8BC7E38E07145B6D15756DA2",
INIT_34 => X"EB8E3FE10F7AEBAFFF080A175D708517DF7D497BC5028142A87000A28A2AA920",
INIT_35 => X"0B6DB6AA28A280001FF5D0A10482FFFFEFBC7E3DF42028080E000280071E8A00",
INIT_36 => X"00000000000000000000B6FBD5410490A3DFD7F7A4821D7A2D16FA82142EB8E0",
INIT_37 => X"FEF007BE8BFF5D2ABDF55F7AABDEAAF784154BA0000000000000000000000000",
INIT_38 => X"DE00FF84154BA087FC01EFA2FFD7545AAAE97555A2FBFDF455D556AA00082EBF",
INIT_39 => X"02000F7AAA8B55FFAABDFEFF7D16AA00FFAEBFFEFAA803DEBA5D2E82155A2FBF",
INIT_3A => X"A95545F7D5555FFAAAAA8BFF002AAAA00FFAAA8AAA080028BFFF7D568BEF0804",
INIT_3B => X"2E95400A2AEA8A00007FEABFF00042ABFFA2FFFFF45F7AE97400AAFFE8B45AAA",
INIT_3C => X"82E820BA08556AA00AAAABFE00F7AEAABEF082E9554508557DFFF007BD54BA5D",
INIT_3D => X"A2D57FE00552EA8A00FFFFE8AAAAA80001FF5D2E82000F7FFFFF45AAFFC20BA0",
INIT_3E => X"0000000000000000000000000000000000000FFFBD5400082EBFF45F78400155",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_3,               -- Port A enable input
WEA      => wbe_a_hi_1024_3(1),               -- Port A write enable input
DIA(0)   => data_write_a(11),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_3(11),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_3,               -- Port B enable input
WEB      => wbe_b_hi_1024_3(1),               -- Port B write enable input
DIB(0)   => data_write_b(11),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_3(11),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_12_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50080B01BC002006940202C0DE041196A83183000000023322287E0FC000006",
INIT_01 => X"75400D849830C84C5823E0000C17424840000000080000088200002802153231",
INIT_02 => X"18A026B43ED180040147558040090000061800000C06ED9802768F4472C52005",
INIT_03 => X"2A67E34A528D0524A52850528400C8001100000171C02B550618C91A10E55440",
INIT_04 => X"1BC0000100056C8280825DE98154004300C840800850240080CA921084520A07",
INIT_05 => X"02000F832000500C0000941024000852084060202E100001002000448100000C",
INIT_06 => X"819A1D1C3FE01A1A40045408049A50BA4020C6041090001200006200000000F2",
INIT_07 => X"C26A0719CC96CC6ED18A64019695A854870300FA3968B20068FC06080106249F",
INIT_08 => X"D002024B3E040800008C0A002610240D494A06F3460409000000E3F0AD5282E5",
INIT_09 => X"27A06009200040000400120412445D78400001000410420080218029CC807A27",
INIT_0A => X"18000006848A026F000000000000080000F010C100204593F11A6CDF48003BF8",
INIT_0B => X"000000820040402B28050400400432C9349DF21A31A00ACC0000F04F80020001",
INIT_0C => X"00357804611AE45D05D0833430CD0833420CD0C33420CD0833430668619A1000",
INIT_0D => X"0000000000000A74812DF00E87E80A079F9F90FA0280E87E800C7FF3B8002000",
INIT_0E => X"3B6B0E404D26160682082002000401EA0000C40000800A006002818808000000",
INIT_0F => X"A476D61C809A4DA84272592D6246FC1B17B541F97E1B348EDA93900B2B286C56",
INIT_10 => X"30C669E622DBC325CFD881A962454CFBE5403AB99594362B1DB52720165650D9",
INIT_11 => X"F8D2D39A3745261E4A95A110A3F855000E4B1D32BAB504BB7490FCFF912A3834",
INIT_12 => X"B90E9B018C7530200AB8F8BF41F9A22006B37DC8E1F9A21A70116D4C5080651C",
INIT_13 => X"118780319CCA08AB1001ACDF34B8F1C688AB1002AE3F7B807B6289F368828C4C",
INIT_14 => X"2AF020233376A5ECC016B1A827CDA21160F051DE610A34C50427E6E220323E4A",
INIT_15 => X"0077020000000439FDC05C5806781FAB46095A0B5199B0AC55521524F1864022",
INIT_16 => X"000000000000000000000000000000000026C000002884000130921092804010",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"8020080200000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0051B946088881360A95090CB054420290100000000000000000008020080200",
INIT_1A => X"041041041041041041041041041041041049249249249249200100002D451451",
INIT_1B => X"92C964B2592C964B2592C964B2592C964B2592C86432190C86432190C8641041",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000003800F592C964B2592C964B25",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"7DE1000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"ABDFFFF7803DE10AA80000AAAA843FE0008557DFFF0800020105D557FEAA0055",
INIT_29 => X"D5420000051555FFA2AA8200000557DFFFF7AA80000082ABDF5508557DF45002",
INIT_2A => X"82AA8AAAAAFFC00BA007FC2155F7D155545AA80001EFAAFBEAB45557FFDE10AA",
INIT_2B => X"FFAEBFEAA002A801FFF7FFE8A10A28000000A2D155410F7FFFFEBA08003FE000",
INIT_2C => X"5FFFFEAABA000028A105D2ABFE10A2AABFE1055516ABEF5D517DEAAA2AEBFF45",
INIT_2D => X"55002A820AA08557DFFFF7AA82155AAFBE8B45002A974AAAA803DFFFAA843DF4",
INIT_2E => X"000AAD155555A28428BFF002ABDE00A2AABFE10082ABFFEF0855420000004175",
INIT_2F => X"5010495B7AE921C517DE10000000000000000000000000000000000000000000",
INIT_30 => X"BDF6D005B78F7D142ABDFC7F78E3FE28B684070AABE803AE38145B78FD700000",
INIT_31 => X"BEFB455D71F8E00BED547038145B505FFB6A487000005F7AFD7F7A482038002E",
INIT_32 => X"F1FDE821C003FE001C2EAAAAAB6F5C2082007BC217DEBDB55555AA8E071D7AAF",
INIT_33 => X"D517DEAABEAEBFF7DEBA0BDEAA1C2A801C7E3FFEFA10B68407038B6D550428FF",
INIT_34 => X"B68E38FC7BE8A3DF7DF7F5E8A9200002FA285D20BDE28A2A4B8E10555B68BEF5",
INIT_35 => X"F085F47038140010555142082082005F7DFD7F7A482155BEF1E8B6D002090482",
INIT_36 => X"00000000000000000000B6D15756DA28A28BFF082ABAE10B6AAB8E280820B8FE",
INIT_37 => X"ABA5D7FEAB45080015410007FEAA0055517DE000000000000000000000000000",
INIT_38 => X"AB45F780020BA082EBFFEF007BE8BFF5D2ABDF55F7AABDEAAF784154BAF7802A",
INIT_39 => X"D7545AAAE97555A2FBFDF455D556AA00F7D1554BA5D7BC01FFFF8015410007FE",
INIT_3A => X"4154BAF7D1400BAFFD57FE005D043FE10552EAAAAAFFD140000087FC01EFA2FF",
INIT_3B => X"8428A105D7FEABEF55557DEBAFFAEBFFEFAA803DEBA5D2E82155A2FBFDE00FF8",
INIT_3C => X"7D568BEF080402000F7AAA8B55FFAABDFEFF7D16AA0008003FEBA55003DEBAA2",
INIT_3D => X"FFAAA8AAA080028BFF087BD54AA550402145550000010087FFFF45F78402145F",
INIT_3E => X"0000000000000000000000000000000000000F7D5555FFAAAAA8BFF002AAAA00",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_3,               -- Port A enable input
WEA      => wbe_a_hi_1024_3(1),               -- Port A write enable input
DIA(0)   => data_write_a(12),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_3(12),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_3,               -- Port B enable input
WEB      => wbe_b_hi_1024_3(1),               -- Port B write enable input
DIB(0)   => data_write_b(12),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_3(12),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_13_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10154A0441836CA2840512822007C18000E02700500030B31B300040081A042",
INIT_01 => X"00000804A000C04800020000000002404001000008220008A200100802110204",
INIT_02 => X"02200430000104000A4700804008000004100000000420918204D3033240400D",
INIT_03 => X"AA4003400008592400000590C40009141100000C6180C0000000C00001E14000",
INIT_04 => X"0800000102400120088054019000004160004190BAA0270000C8100000600206",
INIT_05 => X"21000012040610050040000227003AA0082400E94C1200000824424005220020",
INIT_06 => X"81963B180C001010580000080400000058000004109C00138000020024142581",
INIT_07 => X"002C8008000441600106400A9600010494020002B8AAA000EF003408000E2580",
INIT_08 => X"000000E48194408000A00A001210040441C80320040210000002ABF004102244",
INIT_09 => X"2A004009640040100400940412D4C4004000022000104200802D983000480120",
INIT_0A => X"8000202020401480000000000000080C90090881000145B0111A14004015080D",
INIT_0B => X"00000002004040AA08050400404040C11444000805200A402090024000008002",
INIT_0C => X"8410000A00280020020040800020040800020000801020000800010020400000",
INIT_0D => X"84A14250A055100050100490000500D00040080040290000084E4000B800610C",
INIT_0E => X"DCD13042BEDA36820228000000000000C000400081A08BC812A2092B02850942",
INIT_0F => X"89B9A260857DB400431969CA985D480949D32804A40AB137341C10B7D6A02EC0",
INIT_10 => X"E6ACA678001CE7D0296C213A460CA4271CA2168AEC1017606E6838216FAD4055",
INIT_11 => X"84AD4961C281B20213073C5FC0058008632D30D522CE80239DCC01AB013A4D20",
INIT_12 => X"2E6B13804A4B01D83461299900F6BD583A519104A0EEBD1A141010B2A4C8E116",
INIT_13 => X"89E5E40913419151EE0E94641828F72B5151EE0D184B321037AF5158BB02D085",
INIT_14 => X"562EC0B42162D68EE0073AE1C562EC13D521921A4170300B2B458B56B01C2280",
INIT_15 => X"00888A120240034000E6DC8285028014B82372011FC1E4F5E0A00929684EAF84",
INIT_16 => X"50942509425094250942509425094254940A1421420082020120908800480030",
INIT_17 => X"0942509425094250942509425094250942509425094250942509425094250942",
INIT_18 => X"9425094250942509425094250942509425094250942509425094250942509425",
INIT_19 => X"F7EFBBEEFF3F7DF7FF3E9F7DF7E2450228000000000000000000509425094250",
INIT_1A => X"BAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBF7DFDFDDD555555",
INIT_1B => X"EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAEBAE",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000000000F7EBF5FAFD7EBF5FAFD7",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"2ABEF00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0020105D557FEAA00557DE10AAD5554BA087FFFF55557BD54AAF7FBC01FFA280",
INIT_29 => X"7BD75EF087FFFFEF557BEAB45552E80155AA802AB45AA843FE0008557DFFF080",
INIT_2A => X"FAE820AA5D5557555082ABDF5508557DF45002ABDFFFF7803DE10AA80000AA08",
INIT_2B => X"0051555FFA2AA8200000557DFFFF7AA80000AAD1420AA087BD7555FFD168AAAF",
INIT_2C => X"5557FFDE10AAAEA8BFFA2FBD7545FFD157555085140010F7AEAABFFAAD542000",
INIT_2D => X"BA557BE8A10A284154BAFFAAAAB45007FC2155F7D155545AA80001EFAAFBEAB4",
INIT_2E => X"000A2D155410F7FFFFEBA08003FE00082AA8AAAAAFFC00BA00002AAAAF7D5574",
INIT_2F => X"0492E3F1C71C7BE8A2ABD7000000000000000000000000000000000000000000",
INIT_30 => X"3AE38145B78FD7000005010495B7AE921C517DE10A2DB50482147FFAF554971D",
INIT_31 => X"E3FE28B684070AA1C71D25D7007FFAFD7497BE8B5555208217DBE8A2AB45BE80",
INIT_32 => X"7FD257DFFD568A82FFA4870BA555F5056D002EBDF6D005B78F7D142ABDFC7F78",
INIT_33 => X"FAAAFBFFBED547038145B505FFB6A487000005F7AFD7F7A482038AADF4709214",
INIT_34 => X"AA8E071D7AAFBEFB455D71F8E00A2A0ADBC7A2FFD257DE3DF52555085142000F",
INIT_35 => X"21C002AA92FFDF574824171EAA10B680124BAFFAAAFB45007BC217DEBDB55555",
INIT_36 => X"00000000000000000000B6D550428FFF1FDE821C003FE001C2EAAAAAB6F5C208",
INIT_37 => X"0105D7BE8B55085142010AAD157545F7AEA8B550000000000000000000000000",
INIT_38 => X"01EFF7AAA8B55F7802AABA5D7FEAB45080015410007FEAA0055517DE00A2FFC0",
INIT_39 => X"E8BFF5D2ABDF55F7AABDEAAF784154BA5D5140145007BE8B55087BEAB555D040",
INIT_3A => X"0020BAA2FFD54105D7FC21EFFFD16AA10FF80174AA557FC21EF082EBFFEF007B",
INIT_3B => X"FBC0155085540000FFAEBFFEFF7D1554BA5D7BC01FFFF8015410007FEAB45F78",
INIT_3C => X"87FC01EFA2FFD7545AAAE97555A2FBFDF455D556AA00A2803FF45AAFFC21EFAA",
INIT_3D => X"552EAAAAAFFD1400005D042AA00F7FBD5410085568A10FF80020AAFFAABFF550",
INIT_3E => X"0000000000000000000000000000000000000F7D1400BAFFD57FE005D043FE10",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_3,               -- Port A enable input
WEA      => wbe_a_hi_1024_3(1),               -- Port A write enable input
DIA(0)   => data_write_a(13),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_3(13),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_3,               -- Port B enable input
WEB      => wbe_b_hi_1024_3(1),               -- Port B write enable input
DIB(0)   => data_write_b(13),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_3(13),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_14_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10020A000180000284008280000281800000030000000033022000000580002",
INIT_01 => X"000008020000204D006800000030824840000000084000084200090008510200",
INIT_02 => X"0220043170010A600A4D008040080000041000000028009002000F333240800C",
INIT_03 => X"111813400008002400000000C400090011000000610200001104D83000F14000",
INIT_04 => X"0801800100A000000000540084000040000040000800200000C8100000000748",
INIT_05 => X"0100000000001000000000002000080008000000001000000024024001200020",
INIT_06 => X"819EB84028001010000000080400000000000004108000100000020020040081",
INIT_07 => X"92040608000440100102400A94810206844200021DA2A0002000340800062C80",
INIT_08 => X"000000000084400008800A001214040441481500040000000000A7F408002244",
INIT_09 => X"0A0040090002008420401004104444004000020400214A208001000002400120",
INIT_0A => X"0400002020000000000000000000080C8008088100004590111B480040120000",
INIT_0B => X"1000000200404800000504016000002114000008020000020080024000000000",
INIT_0C => X"0410000010000000000040001000000000000040000000000001000000000000",
INIT_0D => X"04810244825010004010000000000000000000000000000000080000B8002104",
INIT_0E => X"0002C38280001202020800000000001000004000000000401022000002040902",
INIT_0F => X"20000587050001404E8084341CBA3404800828805200008000E0E0A000080002",
INIT_10 => X"4D18178E012010C00224004091C3514072C000444A0400080001C1C140001000",
INIT_11 => X"51709A07424142084458476001003809D0104B01C5710044020C4006010500C5",
INIT_12 => X"C26EE3803180C18006519462A00005001460E4730000050A1011004001060049",
INIT_13 => X"01F9E00660318000000538318740000140000001B4600CE80001400000002B62",
INIT_14 => X"0000000AD89857B0E0684411800000003799EB764D000330C300000000E3554B",
INIT_15 => X"0000021002002C000024008284001A0902000422E3F5960080480A0216A07240",
INIT_16 => X"4090240902409024090240902409024090081021020080015134920800480010",
INIT_17 => X"0902409024090240902409024090240902409024090240902409024090240902",
INIT_18 => X"9024090240902409024090240902409024090240902409024090240902409024",
INIT_19 => X"F5579B4E5C8FF0F7BE9D5F7DF650400200000000000000000000409024090240",
INIT_1A => X"9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7BF7DDDDDFCF3CF3D",
INIT_1B => X"F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE79E7",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000003FFF03F9FCFE7F3F9FCFE7F3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"420BA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"BD54AAF7FBC01FFA2802ABEFA2FBE8B55A2AE80000F7D5555555D2AAAABAAAD1",
INIT_29 => X"AA801FFA28402000AAAE955455500155EF0804155EFAAD5554BA087FFFF55557",
INIT_2A => X"7AEA8B45080417400AA843FE0008557DFFF0800020105D557FEAA00557DE10A2",
INIT_2B => X"087FFFFEF557BEAB45552E80155AA802AB4500516AA00A2AE800BAFFFFC20BAF",
INIT_2C => X"0AA80000AA005568ABAA28402010A2843FEBAFFFBD7410A2D168BFF087BD75EF",
INIT_2D => X"005D7FFDF4555517DFEF00043FEAA082ABDF5508557DF45002ABDFFFF7803DE1",
INIT_2E => X"000AAD1420AA087BD7555FFD168AAAFFAE820AA5D5557555002E80155A280000",
INIT_2F => X"0555412AA8ABAAADB40092000000000000000000000000000000000000000000",
INIT_30 => X"50482147FFAF554971D0492E3F1C71C7BE8A2ABD7A2FFEDB55B6A080038E3DB5",
INIT_31 => X"B7AE921C517DE10A2AE851FFB68402038AAAA955554900105FF0800175D7A2DB",
INIT_32 => X"A0800BAE3F1C0092EBAAADB6D080A12410BE803AE38145B78FD7000005010495",
INIT_33 => X"2D568BC71C71D25D7007FFAFD7497BE8B5555208217DBE8A2AB451C556FA00A2",
INIT_34 => X"142ABDFC7F78E3FE28B684070AA00516DABAA28402038B6803DE82F7F5D5410A",
INIT_35 => X"D002A80155B680000105D7FF8F455D5F78FD7000E3FEAA002EBDF6D005B78F7D",
INIT_36 => X"00000000000000000000AADF47092147FD257DFFD568A82FFA4870BA555F5056",
INIT_37 => X"F55FF84000AAAAFBC0145002AA8AAAAAFFC20000000000000000000000000000",
INIT_38 => X"01EF080417555A2FFC00105D7BE8B55085142010AAD157545F7AEA8B55A2FBFF",
INIT_39 => X"EAB45080015410007FEAA0055517DE00A2AA955FFFF80020BAAAAA9754508000",
INIT_3A => X"AA8B555D557FE00A280020BAAAD140000A2AEBFFEF082A82010F7802AABA5D7F",
INIT_3B => X"803DE00FFD557400AAD56AB455D5140145007BE8B55087BEAB555D04001EFF7A",
INIT_3C => X"82EBFFEF007BE8BFF5D2ABDF55F7AABDEAAF784154BA08557FEAAA284000AAFF",
INIT_3D => X"FF80174AA557FC21EF082A80145F780020105D7BEAB45557BE8B45082EBFEBA0",
INIT_3E => X"0000000000000000000000000000000000000A2FFD54105D7FC21EFFFD16AA10",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_3,               -- Port A enable input
WEA      => wbe_a_hi_1024_3(1),               -- Port A write enable input
DIA(0)   => data_write_a(14),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_3(14),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_3,               -- Port B enable input
WEB      => wbe_b_hi_1024_3(1),               -- Port B write enable input
DIB(0)   => data_write_b(14),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_3(14),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_15_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000A000000000284000280000001800020030000000033022000000180002",
INIT_01 => X"8000080000000048000000000000026040000000080000080200000000110200",
INIT_02 => X"0020042004010E60004C0080000800000410000000020090020000300245E005",
INIT_03 => X"0000010000080400000000408400480111000000610008000000C00000E54400",
INIT_04 => X"980000010000000088C2550080000040000040000008A00028C8100000120000",
INIT_05 => X"020004012E025000000001322000000A28008000011000000220004D41000000",
INIT_06 => X"819588000800101000011008040000100001060418800510000A620000000092",
INIT_07 => X"0000000800044004010C20008440810284020002102220002000340800062480",
INIT_08 => X"0000000001140800002C0A001214050540C800400406180000002DF004000244",
INIT_09 => X"1E00400900000000000016041044400440000000000042008001000000000022",
INIT_0A => X"0000000000000220000000000000080C00000081000045901118000040000000",
INIT_0B => X"0000000200404000010500004000000114000009000000000000004200000000",
INIT_0C => X"0000000000000000000040001000040001000000000000000001000020000800",
INIT_0D => X"000000000000001001208000180800000000030200000180800C400030002000",
INIT_0E => X"0000000000002600020800000000001080004000000000000002000000000000",
INIT_0F => X"A400000000000000000008000000000000000000000014800000000000000052",
INIT_10 => X"0000000000000000000000010240000000000000000000290000000000000000",
INIT_11 => X"2001C05838120800000000000000000000010000000000000000000000001804",
INIT_12 => X"081004000000000000A010000000000000902000000000180010002020000000",
INIT_13 => X"6600000000000000000024080000000000000000280400000000000000000000",
INIT_14 => X"0000000000200801000000000000000000501001920000000000000000000A40",
INIT_15 => X"0000020000000000000000003000000000000000000A101C3614000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000080000120980000000010",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000400200000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"28BEF00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"5555555D2AAAABAAAD1420BAFF8000010082A954BA00003DFEF085155400F784",
INIT_29 => X"AE95555A2FBE8BEFA2843DE00AA8015400FF84001EFA2FBE8B55A2AE80000F7D",
INIT_2A => X"2FBEAB45F7D56AABAAAD5554BA087FFFF55557BD54AAF7FBC01FFA2802ABEFF7",
INIT_2B => X"A28402000AAAE955455500155EF0804155EFFFFBE8BFF0800174AA557BFDE10A",
INIT_2C => X"A00557DE10F7D1574AAA2D16AB55FFD568BEF087FE8A1055003FE00A2AA801FF",
INIT_2D => X"00AA802AA00AAAE800BA5D0015545AA843FE0008557DFFF0800020105D557FEA",
INIT_2E => X"00000516AA00A2AE800BAFFFFC20BAF7AEA8B45080417400FFFFC21450800154",
INIT_2F => X"8FD7005150438F78A2DBFF000000000000000000000000000000000000000000",
INIT_30 => X"EDB55B6A080038E3DB50555412AA8ABAAADB40092E38E070280024904AA1C043",
INIT_31 => X"1C71C7BE8A2ABD7E3AA9257DA2FFE8BC7BE8E38E10A28017400E38A051FFA2FF",
INIT_32 => X"00124AA557FFDE10A2FBEDB6DF7D16AABAA2DB50482147FFAF554971D0492E3F",
INIT_33 => X"10038E38A2AE851FFB68402038AAAA955554900105FF0800175D7E3FFEFBD700",
INIT_34 => X"000005010495B7AE921C517DE10FFDF50482A2DB6AB45FFD56DBD7087BEAA384",
INIT_35 => X"0FFF1C017D140410400BE8E28A10AAA085082550A1057DBE803AE38145B78FD7",
INIT_36 => X"000000000000000000001C556FA00A2A0800BAE3F1C0092EBAAADB6D080A1241",
INIT_37 => X"4AA0800020BA550028B550855400AAF7AEBDFEF0000000000000000000000000",
INIT_38 => X"7400AAAE975EFA2FBFFF55FF84000AAAAFBC0145002AA8AAAAAFFC2000AAAA97",
INIT_39 => X"E8B55085142010AAD157545F7AEA8B55AAAE821EFAAFBEAB55F7AAA8A00AA841",
INIT_3A => X"417555AAFFFDF450804020AA557BFFE10A2FFFFFEFF7D568ABAA2FFC00105D7B",
INIT_3B => X"D17DF45007FE8AAA08002AAAAA2AA955FFFF80020BAAAAA975450800001EF080",
INIT_3C => X"7802AABA5D7FEAB45080015410007FEAA0055517DE00FFFBC2000AAFBE8B55F7",
INIT_3D => X"A2AEBFFEF082A82010FFD5421EF5D0000010F7AAA8A10AA8017400552A801EFF",
INIT_3E => X"00000000000000000000000000000000000005D557FE00A280020BAAAD140000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_3,               -- Port A enable input
WEA      => wbe_a_hi_1024_3(1),               -- Port A write enable input
DIA(0)   => data_write_a(15),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_3(15),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_3,               -- Port B enable input
WEB      => wbe_b_hi_1024_3(1),               -- Port B write enable input
DIB(0)   => data_write_b(15),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_3(15),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_16_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"DA22C618B1000482B688B186588884862A400438255FC38381441205BA803003",
INIT_01 => X"7045A80028404C211203A952A90341080B173340412000E1005D628000820484",
INIT_02 => X"428406A4000850848330118D0AAC55001349B108818005460229044001C01784",
INIT_03 => X"092C4020000500020000500986812C405000001A48202050000A214AC0650115",
INIT_04 => X"4804A55440256F504025E003A054F46415A4E62B6FE3307943965A00001A1152",
INIT_05 => X"0000001C40A5B950ADB8EA097057ECE14C86D2B7F85AAD17F4B100000B88148C",
INIT_06 => X"415401DCDCF2C0A8030140BCB0820A200342A1C641C1E8782F508F2B00003584",
INIT_07 => X"002701881A3202080AE00480A2002840BE1480FA004342AA6F12000054004867",
INIT_08 => X"08C54828091002000002B32A8C19064E486A8001510000014140C1E2A14891E0",
INIT_09 => X"015452B103020814004088B64102680B6596594800400413CAC0208944800000",
INIT_0A => X"96AA000484094C000000000000012C9000A0000D0A80000BF8028E87C1B99270",
INIT_0B => X"014808A02004200E540480212000A448C0082024AE50064B44000000000002A2",
INIT_0C => X"0004000D5846256AAEA811150445411150445411150445411150422A088A8200",
INIT_0D => X"00000004010042A204A0C5817D00005034052E40000817D00440004004AD3240",
INIT_0E => X"632B2673FA4587978A2004102800809225545155121740000004900090000000",
INIT_0F => X"00C6564CE7F4EA4B940076D296D003030800462CBD320018CAAAACFE9164C800",
INIT_10 => X"28834ADB1440A114793A4A30A40839AA14910D08DCB2640031955559FD3AC990",
INIT_11 => X"594AB0B1A025371CA0E034E8443C097A800EB090D4AAC91208ED2FA0CE5E09B1",
INIT_12 => X"7B50446083001B94BB38C540EBE61284BB304880E3E4579EDC00992980D58033",
INIT_13 => X"5511121840E7A2CD952ECC12ABC3E6ACB3DFB12ECE315000F61FF1727A85FDBC",
INIT_14 => X"75DEB07F6F2E7084517F126F8395CB2BEFBAB8BA8AF698228CC5E2F08ECA5159",
INIT_15 => X"5580A840A8009F8B108C80A1021B080AFC0DF6422C6077F4A77F20D0C0E21084",
INIT_16 => X"0000000000000000000000000000000000044000102A0001148442A110810359",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"558D11544C690DA64C1C4F68A360400000000000000000000000000000000000",
INIT_1A => X"14D14D14D14D14D14D14D14D14D14D14D14514514514514529E5F87869E79E78",
INIT_1B => X"D1E8F47A3D1E8F47A7D3E9F4FA7D3E9F4FA7D3E9F47A7D1E9F47A7D1E9F4D14D",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000007D3E9F4FA7D3E8F47A3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"C00AA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"03DFEF085155400F78428BEF087FFFFEFF7D168B55AAD17FFFF552EBFE00007F",
INIT_29 => X"2E975EFF7D568BFFFF80175EF0004000BA552A821FFFF8000010082A954BA000",
INIT_2A => X"55540000082EAABFFA2FBE8B55A2AE80000F7D5555555D2AAAABAAAD1420BA5D",
INIT_2B => X"A2FBE8BEFA2843DE00AA8015400FF84001EF0000020AA5D00154005D043FF455",
INIT_2C => X"FA2802ABEF557BEABEF5D0415410087FD74BAAAAEBFFEF557FC00AAF7AE95555",
INIT_2D => X"FFFFAABFEAAFF84001FF002A821FFAAD5554BA087FFFF55557BD54AAF7FBC01F",
INIT_2E => X"000FFFBE8BFF0800174AA557BFDE10A2FBEAB45F7D56AABA082A97545F7D16AB",
INIT_2F => X"FFEF552AB8E38087FC2092000000000000000000000000000000000000000000",
INIT_30 => X"070280024904AA1C0438FD7005150438F78A2DBFF0871F8FC7E3D56AB6DBEDB7",
INIT_31 => X"AA8ABAAADB400924920925EFF7D16ABFFE38E175EF1400000BA412E871FFE38E",
INIT_32 => X"0A1240055003FF6D5551420101C2EAFBD7A2FFEDB55B6A080038E3DB50555412",
INIT_33 => X"57FC00BAE3AA9257DA2FFE8BC7BE8E38E10A28017400E38A051FF0804050BA41",
INIT_34 => X"4971D0492E3F1C71C7BE8A2ABD74975EDBC7550E12410087FD74AAB6AABFFC75",
INIT_35 => X"A08249756DF7D168BC7F7AABAEAAF780051C70824851D7A2DB50482147FFAF55",
INIT_36 => X"00000000000000000000E3FFEFBD70000124AA557FFDE10A2FBEDB6DF7D16AAB",
INIT_37 => X"B55A2D16ABEFFFFBFDFFF552AAAAAA007BC00000000000000000000000000000",
INIT_38 => X"20AA002A955EFAAAA974AA0800020BA550028B550855400AAF7AEBDFEF08516A",
INIT_39 => X"000AAAAFBC0145002AA8AAAAAFFC20000000021EFF7D568BFFA2AA955FF5D040",
INIT_3A => X"E975EF0800174BA002E820105D003DFEF5D51420005D2ABFF45A2FBFFF55FF84",
INIT_3B => X"7BD74AAF7AEBDF455D7BC20BAAAAE821EFAAFBEAB55F7AAA8A00AA8417400AAA",
INIT_3C => X"2FFC00105D7BE8B55085142010AAD157545F7AEA8B5500557DF45552A8200000",
INIT_3D => X"A2FFFFFEFF7D568ABA0804155FFF7D568B55FFAAAAABAFF8415545000015555A",
INIT_3E => X"0000000000000000000000000000000000000AAFFFDF450804020AA557BFFE10",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_3,               -- Port A enable input
WEA      => wbe_a_hi_1024_3(2),               -- Port A write enable input
DIA(0)   => data_write_a(16),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_3(16),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_3,               -- Port B enable input
WEB      => wbe_b_hi_1024_3(2),               -- Port B write enable input
DIB(0)   => data_write_b(16),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_3(16),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_17_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"5284CE4FB7BD2C8994A13392DBD02E14006B82AC7E800D44D3DD2FD5F9B961C0",
INIT_01 => X"2EACD01F7E03FC6793F2199B39FC233C11D93AE6F3BB92B32091DBC339B24542",
INIT_02 => X"E63CCCC00A82C08092A2AFAE667033DB50853379C10BFDC5C6F4044443C817C6",
INIT_03 => X"7FF183635AEF9E3635AEF9E18E237040404446965C0607EE6DB7854AC4DE060C",
INIT_04 => X"D78AC33FB604488B000892EF17BE6D84196482236FE100294152E294350FB697",
INIT_05 => X"081B5F9B409420D0CDB47A05403F6CE0C08A4AB7F840EDB6F48100DFC8081081",
INIT_06 => X"768465354781CBC30316367077B4BDB50646E8D87100A8201ED01C19C020F71A",
INIT_07 => X"4002A110C922480A82D0841147162C48EBB9537A0022DC67987042EE976ABEA7",
INIT_08 => X"DB931BFEF91C00002CC0E019C0C82A4E4820C15A2330E004401891181168C4D1",
INIT_09 => X"09F3A1BC11EFBC66DB65307071477FF1030C397C060B4254064302042F803A69",
INIT_0A => X"3F330802162F3B7EE3F3EC7C7DEF207000F00059D2ED56D7EED2ED3C9A867DC0",
INIT_0B => X"185C44B91BC1740B7605040BE0018CFC7429F326B9E822FFC00074D5A0AB033A",
INIT_0C => X"00367A28FC1B7F7FEFFCFBFF3EFFCFBFF3EFFCFBFF3EFFCFBFF3EFFE7DFF9E00",
INIT_0D => X"0000000008004BA78428C7AD7FC94B533F5B4FFBD2FAD7FCCA786D43FE67C218",
INIT_0E => X"BA494CEBFD4F2667ABB6F68B29760593F33FA0CF170F40006001B1A05C000000",
INIT_0F => X"7F749299D7FAEB237DFE5865B6D2BF23265CBACE542A6FEE92333AFF33E0A9BF",
INIT_10 => X"F6C24B6D18C3C9F8E2881F3F787D776B5DB94A09955054DFDD246675FE7AC153",
INIT_11 => X"BFB349E08FF9A27EDE9FA8AEFD9E7467BFCB195CFEB56A1A70D34D1706FFFA3E",
INIT_12 => X"6FE219CA80725B875EED723FF7FCB2875EDAAFEAF7FD929BFD55BBC71D79F639",
INIT_13 => X"546670D018E7A6E581D7B6AB75FDFCECA6E581D7BB5DDFC6FF0EB7D7E859FDB5",
INIT_14 => X"B978177F6D6AF5ECDB5FB76A5F5FA165B456E0FB308710C49FCFB741598B9C7E",
INIT_15 => X"CFDAAB00AC00A8BBFC8B501CF7A0FED9A540EA1952586CEB54D143ACFF9A3BA9",
INIT_16 => X"000000000000000000000000000000000026E100002F382DBD9ECFE117805F20",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"4372003009EDCC4052E917114F981800C0000000000000000000000000000000",
INIT_1A => X"BA69A69AEBA69AEBA69A69AEBA69AEBA69A69A69A69A69A68698686981D75D74",
INIT_1B => X"6A351A8D46A351A8D068341A0D068341A0D068341A0D46A341A0D46A341A69AE",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000000000046A351A8D46A351A8D4",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"7FEAA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"17FFFF552EBFE00007FC00AA087FFFFFFFFFFFFFEFF7FBEAB450804001EFAAD5",
INIT_29 => X"D168A000004020AA5D7BE8B450051401EF087FD74AA087FFFFEFF7D168B55AAD",
INIT_2A => X"D7FEAB55FF80175EFFF8000010082A954BA00003DFEF085155400F78428BEFAA",
INIT_2B => X"F7D568BFFFF80175EF0004000BA552A821FF5D00020BA552A82000552A821555",
INIT_2C => X"AAAD1420BAFFFFFDF45AAD17FFFFAAFBC01EF5D0015555557BFDEBA5D2E975EF",
INIT_2D => X"BA007FEABEF005555555A2D1554BAA2FBE8B55A2AE80000F7D5555555D2AAAAB",
INIT_2E => X"0000000020AA5D00154005D043FF45555540000082EAABFF00516AA10552E820",
INIT_2F => X"8B550000071EFB6DF7AE92000000000000000000000000000000000000000000",
INIT_30 => X"F8FC7E3D56AB6DBEDB7FFEF552AB8E38087FC2092147FFFFFFFFFBFDFC7EBF5E",
INIT_31 => X"150438F78A2DBFFBED16AA381C0A07082497FEFB6D1451471EF007BD04920871",
INIT_32 => X"2A850105D2A80155417BEFB6DEB8E175FFE38E070280024904AA1C0438FD7005",
INIT_33 => X"D7BFAEBA4920925EFF7D16ABFFE38E175EF1400000BA412E871FF550A0009249",
INIT_34 => X"E3DB50555412AA8ABAAADB40092FFF5FFF6DAADF7FFD7B6F1C71EF55001756D5",
INIT_35 => X"7145B6AA28492487082007FEDBD700515556DA2DF50492A2FFEDB55B6A080038",
INIT_36 => X"000000000000000000000804050BA410A1240055003FF6D5551420101C2EAFBD",
INIT_37 => X"FEFF7FBFFF55A2D16AB550000175EFFFFBEAA000000000000000000000000000",
INIT_38 => X"55EF087FC200008516AB55A2D16ABEFFFFBFDFFF552AAAAAA007BC0000557FFD",
INIT_39 => X"020BA550028B550855400AAF7AEBDFEFF7D568AAA5D2A97410007BFFFFF55515",
INIT_3A => X"A955EF5D2E80010002A954005D2A82155087FFFFEFAAAA975EFAAAA974AA0800",
INIT_3B => X"D1575FF5504175EF5D7FEAAAA0000021EFF7D568BFFA2AA955FF5D04020AA002",
INIT_3C => X"2FBFFF55FF84000AAAAFBC0145002AA8AAAAAFFC2000FFD57DFFFAAFFFDF55FF",
INIT_3D => X"5D51420005D2ABFF45557FE8AAA000415410007BFFF450051555EFA2FBC0000A",
INIT_3E => X"00000000000000000000000000000000000000800174BA002E820105D003DFEF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_3,               -- Port A enable input
WEA      => wbe_a_hi_1024_3(2),               -- Port A write enable input
DIA(0)   => data_write_a(17),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_3(17),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_3,               -- Port B enable input
WEB      => wbe_b_hi_1024_3(2),               -- Port B write enable input
DIB(0)   => data_write_b(17),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_3(17),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_18_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"69844019080000A21A611406840014122A641074155FC28A2024001001801003",
INIT_01 => X"7443D920034004180005E9E3C90360C0041C0181002001602025800008440084",
INIT_02 => X"E2DCCCE61D5C008103F2000781FC0FEDEAC2161B0B8FB0008620044443006010",
INIT_03 => X"884E300802006900802006995C896D605200000856E24A040000640052141103",
INIT_04 => X"480520FC026125AC0025C9122644E3E40EC8E2001001302281841A009038A86A",
INIT_05 => X"432000040089983070019400F01010004C8DB841405A80A100B586200FAC24AE",
INIT_06 => X"09044359DC7040000000002C109B0E0A00A1104641C0803804000707284600E1",
INIT_07 => X"400D10100400481D5EB08501620000007500CE801241021FE78E404860140060",
INIT_08 => X"00880C0106A0528020019307CC082A0A4A6A01ED725021400040D028000A9729",
INIT_09 => X"00117063038000282081402E4106400B6186128040600C10C1C0200950508110",
INIT_0A => X"C0C30C2E21580C874004008080003C32A10A19090C02010E1022944061688000",
INIT_0B => X"0180A8062026000DC425C0301311324AA2373088479105D044A1022000001835",
INIT_0C => X"0D89844703649000000200000000000000000000000000000000000000000010",
INIT_0D => X"0D8306C182701404C1973010802020404084001E00010802046092B5001FB365",
INIT_0E => X"528EB314068AB8B803DB00002900800400FC503F08180050942E4200020C1B06",
INIT_0F => X"40A51D66280D6032C5F96D3C51555D5D7D5AA87285820814A3CCC501C2A60820",
INIT_10 => X"8B35A3FEBF1FEDFD9C2B30E0468AAAD5D48F37E8FC1304102947998A03984C10",
INIT_11 => X"440FE1DD772D37A0A321BC6968F32658BF2D4F2A80BF8FE3F9FE3AC362080529",
INIT_12 => X"5487910D7E5A6D961A28456A1832E5161A100DD5182BC54020EA67A189C6ED36",
INIT_13 => X"AA444CAF91EDD1B725868403BE06323551B725868A100ABD119753B70964122B",
INIT_14 => X"EDC259048ACD868EE3803D65CEDC258A8F80D55E007C3F8EBB56F4C5362C978F",
INIT_15 => X"3F240014BE84370001B6922070440556B15F7FABBC0031BCF2257C41634B14D4",
INIT_16 => X"C1B06C1B06C1B06C1B06C1B06C1B06C1B0491069068000004060300A005A0118",
INIT_17 => X"1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06",
INIT_18 => X"B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C",
INIT_19 => X"B28BBECEB80EE173C2300F7DF16000000000000000000000000041B06C1B06C1",
INIT_1A => X"8A28A28AAAAAAA28A28A28AAAAAAA28A28A28A28A28A28A2910591505C104104",
INIT_1B => X"28944A25128944A25128944A25128944A25128944A2552A954AA5128944AAAA2",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000128944A25128944A251",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"9540000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"BEAB450804001EFAAD57FEAA087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974BA082E",
INIT_29 => X"7FFFFFFFFFBFDF45AAD568B55080028B55002E82000087FFFFFFFFFFFFFEFF7F",
INIT_2A => X"0043DE10AA843DE00087FFFFEFF7D168B55AAD17FFFF552EBFE00007FC00AA08",
INIT_2B => X"0004020AA5D7BE8B450051401EF087FD74AAAAFFFDF45A2D16AB55F7FFFFFFF0",
INIT_2C => X"0F78428BEFAA80000000804154BA55042ABEF5D7FD75FFAAD540145AAD168A00",
INIT_2D => X"00082E95555085168A10557FD7545FF8000010082A954BA00003DFEF08515540",
INIT_2E => X"0005D00020BA552A82000552A821555D7FEAB55FF80175EF5D00020105D2A974",
INIT_2F => X"DFFF5D2A954AA082A92428000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFBFDFC7EBF5E8B550000071EFB6DF7AE921C7FFFFFFFFFFFFFFFF7FBF",
INIT_31 => X"AB8E38087FC2092087FFDFC7E3F1FAF55A2DF6DB7D1C002AB7D002A82028147F",
INIT_32 => X"DF6DB7DE3F5FAFC708003DE28B68E38E280871F8FC7E3D56AB6DBEDB7FFEF552",
INIT_33 => X"ADF4516DBED16AA381C0A07082497FEFB6D1451471EF007BD0492B6F1F8F55AA",
INIT_34 => X"1C0438FD7005150438F78A2DBFFA28407038140410492550A2ABC7497BD25FFA",
INIT_35 => X"F5D0E05000492097428002E9557D1C516FA28417BD5545E38E070280024904AA",
INIT_36 => X"00000000000000000000550A00092492A850105D2A80155417BEFB6DEB8E175F",
INIT_37 => X"FFFFFFFFDFEFF7FBFFFEF552E974AA082A820AA0000000000000000000000000",
INIT_38 => X"ABEF002A800AA557FFDFEFF7FBFFF55A2D16AB550000175EFFFFBEAA00557FFF",
INIT_39 => X"6ABEFFFFBFDFFF552AAAAAA007BC0000087BFDF45AAD568B55AAFBFDFEF55042",
INIT_3A => X"FC2000FFD56AB45A2FFFDFFFAAD16AB4500043DEAAFFAEAAAAA08516AB55A2D1",
INIT_3B => X"2AA8B45087FC01EFA2FFD55EFF7D568AAA5D2A97410007BFFFFF5551555EF087",
INIT_3C => X"AAA974AA0800020BA550028B550855400AAF7AEBDFEFA280154BA55040000055",
INIT_3D => X"087FFFFEFAAAA975EF5D2E974000804154BA082A975EF5D517DEAA007BD5545A",
INIT_3E => X"00000000000000000000000000000000000005D2E80010002A954005D2A82155",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_3,               -- Port A enable input
WEA      => wbe_a_hi_1024_3(2),               -- Port A write enable input
DIA(0)   => data_write_a(18),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_3(18),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_3,               -- Port B enable input
WEB      => wbe_b_hi_1024_3(2),               -- Port B write enable input
DIB(0)   => data_write_b(18),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_3(18),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_19_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"042200000000000041088001001AA00000000000000000000000500802000003",
INIT_01 => X"040048000024000000000404000000000A22000800000800004A200000000001",
INIT_02 => X"200C8840085EB00480060000001C008002489E0F000405EA0004040404000000",
INIT_03 => X"24004000000000000000000900002C4050000000000069500208400002E14100",
INIT_04 => X"4800200C0000000044002000C80020E40000E200000130200188000000800100",
INIT_05 => X"000000000080181000000000701000004C8000000058800000B1000009880480",
INIT_06 => X"80500081081040000000002C100040400000004641C080380400070100000000",
INIT_07 => X"4020109801A4CE005C00048380142810010564C4100114012002402028044808",
INIT_08 => X"0070700000000000000083004C3902420062000020E0000100004082A140102B",
INIT_09 => X"001150200000000000000026400000016186100000000010C04002C000000000",
INIT_0A => X"007C00008082C0002000000000002C3000000004050001030102040000000000",
INIT_0B => X"0000000000000000000000000000010000800011000000000000000000000BC0",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"000000000000000000000000000000042000760000000000000000010004B200",
INIT_0E => X"0D74002280300F0002FB069040000060000C5003000800000000000000000000",
INIT_0F => X"C01AE8004500744C780687DBA828008080A5FC0D385598035D0008A00C015660",
INIT_10 => X"39D8140040201BF861F0E7D693E6170022408116DFE0AB3006BA0011401D02AC",
INIT_11 => X"5412E4997F5249FD005043B8680CC98F00D0F2DD0140100406FE053A98F6ECC7",
INIT_12 => X"7418663001858040E153888000010840E165D0000000285C246A181C03FE4662",
INIT_13 => X"8199830066F0020858385974000001260208583854E2200000660208D6B1423F",
INIT_14 => X"8235AC508FCE8811042040F008235AE04420C040CF00C031C80009B8F224978B",
INIT_15 => X"030004E00000C220010808C10D9A92A74CD7CF4A09051110AD5A3C9200B7F280",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000118",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"07208BBA3F0C7010C660C7441920000000000000000000000000000000000000",
INIT_1A => X"861869A61861861861869A61861861861861861861861861A8208C4C1534D34C",
INIT_1B => X"984C26130984C26130984C26130984C26130984D26930984C26130984C261861",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000984C26130984C26130",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"174BA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFDFEF5D2A974BA082E95400F7FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0004",
INIT_29 => X"FFFFFFFFFFFFFFFFF7FBFDFFF552E974BAA2FFFFE10087FFFFFFFFFFFFFFFFFF",
INIT_2A => X"004001EFAAAEA8ABA087FFFFFFFFFFFFFEFF7FBEAB450804001EFAAD57FEAAF7",
INIT_2B => X"FFFBFDF45AAD568B55080028B55002E82000F7FFFFFFFFFFFFDFEFA2D568B550",
INIT_2C => X"0007FC00AAF7FFFFFFFF7FBE8B55AAD16ABEF5D2ABFF55080402010087FFFFFF",
INIT_2D => X"55A2FFFDFEF5D2EBFE00AAFFFFEBA087FFFFEFF7D168B55AAD17FFFF552EBFE0",
INIT_2E => X"000AAFFFDF45A2D16AB55F7FFFFFFF00043DE10AA843DE00557FFDFEFA2D16AB",
INIT_2F => X"FFEF552A974AA0000104AA000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFF7FBFDFFF5D2A954AA082A92428E3FFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"0071EFB6DF7AE92EBFFFFFFFFFFFFDFEFF7F5FAFC7492A974AAB6F5F8E101C7F",
INIT_32 => X"F1F8FD7AAD16AB450000001FFBEA4A8AAA147FFFFFFFFFBFDFC7EBF5E8B55000",
INIT_33 => X"00000010087FFDFC7E3F1FAF55A2DF6DB7D1C002AB7D002A82028FFFFFFFEFF7",
INIT_34 => X"BEDB7FFEF552AB8E38087FC2092F7FBF8FC7E3F5EAB45B6DF6FBEF5D2AB8F7D0",
INIT_35 => X"84971F8FC7AAD56DB6DBEF5F8FD7412ABFE28B6F5F8E820871F8FC7E3D56AB6D",
INIT_36 => X"00000000000000000000B6F1F8F55AADF6DB7DE3F5FAFC708003DE28B68E38E2",
INIT_37 => X"FFFFFFFFFFFFFFFFFDFEF552E954AA0004000AA0000000000000000000000000",
INIT_38 => X"54AAF7D568A00557FFFFFFFFFFFDFEFF7FBFFFEF552E974AA082A820AAA2FFFF",
INIT_39 => X"FFF55A2D16AB550000175EFFFFBEAA00A2FFFFFFFF7FBFDFFFFFD568B55002A9",
INIT_3A => X"A800AAF7FBFDFEFF7D56AB45AAD56AB450004001EFFF842AAAA557FFDFEFF7FB",
INIT_3B => X"FFFFFFF552AA8BEF080402000087BFDF45AAD568B55AAFBFDFEF55042ABEF002",
INIT_3C => X"8516AB55A2D16ABEFFFFBFDFFF552AAAAAA007BC0000FFFBE8B55AAD168B55F7",
INIT_3D => X"00043DEAAFFAEAAAAA08556AB55A2D57FFFFF7D568B45002ABDEAAFFD16AA000",
INIT_3E => X"0000000000000000000000000000000000000FFD56AB45A2FFFDFFFAAD16AB45",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_3,               -- Port A enable input
WEA      => wbe_a_hi_1024_3(2),               -- Port A write enable input
DIA(0)   => data_write_a(19),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_3(19),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_3,               -- Port B enable input
WEB      => wbe_b_hi_1024_3(2),               -- Port B write enable input
DIB(0)   => data_write_b(19),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_3(19),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_20_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000003",
INIT_01 => X"F55FF80000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"E05022020800008400F655001FFCFF80018FA804400000000000004400000001",
INIT_03 => X"00000000000000000000000900002CC07000000000000000000000000000013F",
INIT_04 => X"68002FFE40900010000180000001FFEC0012EE0C001370F40780000000000000",
INIT_05 => X"0840000880FCBBF0100E204DF0F88311DD8005080679800000F3000029980580",
INIT_06 => X"001000030817C8E8840155FDF9001001050023F6C3C3D0F87FA19F7F011000E4",
INIT_07 => X"000000090492260800008000EE00000000000000002101FF2002C00000004018",
INIT_08 => X"2A040001071004000013FF7FCA302C0C0008214800002101554031F800000000",
INIT_09 => X"801F57F200000090000489FEC0000001EFBEF0040008023FDFC0000000004006",
INIT_0A => X"0000000008000000000000000000ADF000000200000008000008028300110230",
INIT_0B => X"0000000000000800080000000000000000000000000000000800800A40000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"000000040900005C848538000020000000800000080000020000800101FFB600",
INIT_0E => X"00800000003A010003000000000000600FFC53FF001800000002004080000000",
INIT_0F => X"0001000000007408040000004000000004E9000008020000200000000E800800",
INIT_10 => X"00200000000313100010002000008000000000129600040000400000001D0010",
INIT_11 => X"81C012060000000000218F7840000100800004000000000066C0000080080000",
INIT_12 => X"800000000017C000100000000001A800080000000001A8040000002840008185",
INIT_13 => X"0000000006F00000100200000000012600001004000000000066000000801040",
INIT_14 => X"0000200410100000000005F00000020080090A0000000085C800002000586000",
INIT_15 => X"FF00400000000000020020020001000040283024E4F2860400008000030ED080",
INIT_16 => X"00000000000000000000000000000004010201001003020200000000000127DB",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"A0700030038200010089120104D2040020000000000000000000000000000000",
INIT_1A => X"2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2C30C30C30C30C306982121A1E79E79",
INIT_1B => X"32190C86432190C86432190C86432190C86432190C86432190C86432190CB2CB",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000432190C86432190C864",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0201000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF552A974AA0004174BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA0804",
INIT_29 => X"7FFFFFFFFFFFFFFFFFFFFFFEF552E954AA000400000F7FFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E954BA007FC00BA087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974BA082E9540000",
INIT_2B => X"FFFFFFFFFF7FBFDFFF552E974BAA2FFFFE10FFFFFFFFFFFFFFFFFFFFFBFDFFF5",
INIT_2C => X"FAAD57FEAA007FFFFFFFFFFFFFEFF7FBFFF550800020BAAAD56AAAAF7FFFFFFF",
INIT_2D => X"EFF7D56AB450000021EFA2D57DE10087FFFFFFFFFFFFFEFF7FBEAB450804001E",
INIT_2E => X"000F7FFFFFFFFFFFFDFEFA2D568B550004001EFAAAEA8ABA5D7FFFFFFFFFFFDF",
INIT_2F => X"FFFF5D2E954AA080005000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFEF552A974AA0000104AAFFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"A954AA082A92428087FFFFFFFFFFFFFFFFFFBFDFEF5D2E974AA000A07000E3FF",
INIT_32 => X"FFFFFEFF7FBFFFFF552E974AA0071C50BA1C7FFFFFFFFFFFFFFFF7FBFDFFF5D2",
INIT_33 => X"EDF6FABAEBFFFFFFFFFFFFDFEFF7F5FAFC7492A974AAB6F5F8E10E3FFFFFFFFF",
INIT_34 => X"EBF5E8B550000071EFB6DF7AE921C7FFFFFFFFFBFDFEFE3F5F8F450004050AAB",
INIT_35 => X"A497FFFFFFF7FBF8FC7EBD168B450804021FFB6D57DE28147FFFFFFFFFBFDFC7",
INIT_36 => X"00000000000000000000FFFFFFFEFF7F1F8FD7AAD16AB450000001FFBEA4A8AA",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2A954AA0800174100000000000000000000000000",
INIT_38 => X"74AA002E95410A2FFFFFFFFFFFFFFFFFFFFFDFEF552E954AA0004000AAFFFFFF",
INIT_39 => X"FDFEFF7FBFFFEF552E974AA082A820AA087FFFFFFFFFFFFFEFF7FBFDFFF5D2A9",
INIT_3A => X"568A00AAFFFFFFFFFFBFDFEFFFFFFDFEF5D2E954AA0051554BA557FFFFFFFFFF",
INIT_3B => X"D16AB450804174AAFFFFFFEBAA2FFFFFFFF7FBFDFFFFFD568B55002A954AAF7D",
INIT_3C => X"57FFDFEFF7FBFFF55A2D16AB550000175EFFFFBEAA005D7FFFFEFF7FBFDFFFAA",
INIT_3D => X"0004001EFFF842AAAA087BFDFEFF7FFEAB45A2D568B550804001EFF7D57DEBA5",
INIT_3E => X"0000000000000000000000000000000000000F7FBFDFEFF7D56AB45AAD56AB45",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_3,               -- Port A enable input
WEA      => wbe_a_hi_1024_3(2),               -- Port A write enable input
DIA(0)   => data_write_a(20),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_3(20),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_3,               -- Port B enable input
WEB      => wbe_b_hi_1024_3(2),               -- Port B write enable input
DIB(0)   => data_write_b(20),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_3(20),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_21_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"4A302428B824900A128C090A5C1800261500213C005FE812D10420054085A202",
INIT_01 => X"001FFE3440B609703B0427F801A40B8115BC4F655300340288A40D30040E4DD8",
INIT_02 => X"E00424256888D8819801000F9FFFFFFFF149FF1FCA448046C60A0D2437C517F9",
INIT_03 => X"20030640003250640003250F06002CC1740002019824E001CD357832440001FF",
INIT_04 => X"EA2C3FFD400006E04401A8837001FFFC004AEF00080B70E08FB5789421007C5C",
INIT_05 => X"00011A0C40F9FFF80920954FF0F00809DF84A0202879800000F3000029980780",
INIT_06 => X"0805984B7A1FC0A0000101FFF0480080002281F7C3C381F87C03DFFF00009004",
INIT_07 => X"B424068086A205481A60A19000908204A855B000A08A61FF20C3D004D331D340",
INIT_08 => X"1BFA0001600802000023F7FFC08D234B40C2028253000040114200000D0226C0",
INIT_09 => X"EF1F5FF054096C6ADBA169FFC202B1C1FFBEF0440021083DFFCE22DC2880E24D",
INIT_0A => X"45FF0C004041D84862A28C54518DBFF00020004C0A6044901112A0908AA0A300",
INIT_0B => X"018C241102068006C620C03882019480E63180855A492712CC01C49C20201BFE",
INIT_0C => X"08A9464116544302C02D92236488D92236488D92236488D922366446C911B210",
INIT_0D => X"08800444021048034004001890000806002804A0822189000900D80621FFBE00",
INIT_0E => X"060580261013813A2CC396506102C4053FFD5BFF00A04A00200602CA52001100",
INIT_0F => X"080C0B004C202621A85C09411500135844C196D3606941018150098404C1A304",
INIT_10 => X"B02901013416181C96C2C9C600890A2028172192C460D1820302A0130809834A",
INIT_11 => X"9C5E803408250180AC268D185DB3F4350B811068C00049A0A4AA68F05C96A001",
INIT_12 => X"002C006560138F032B1804101244C883052208209040CC849063A747512B7678",
INIT_13 => X"41401E240665750440C9488280254530314080C2C601040420352148A00501B1",
INIT_14 => X"500811204D000700114204A70422016149916011008CAA8858850B00C32591C0",
INIT_15 => X"FFC06E60AC0496022300233104663040808E991765205000070121D41D18D098",
INIT_16 => X"40100401004010040100401004010040102090010008000001C0E010020007DF",
INIT_17 => X"0100401004010040100401004010040100401004010040100401004010040100",
INIT_18 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_19 => X"FFEF9FEEFF7FFDF7FF3E3DFDF7E0000000000000000000000000401004010040",
INIT_1A => X"BEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBFFDFDFFFCF3CF3F",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFEFF7FBFDFEFF7FBFDFEFBEF",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000FFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0001000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E954AA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0004",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA0004154BAFFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"52E974BA0804000AAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0004174BAFF",
INIT_2B => X"FFFFFFFFFFFFFFFFEF552E954AA000400000007FFFFFFFFFFFFFFFFFFFFFFEF5",
INIT_2C => X"A082E95400007FFFFFFFFFFFFFFFFFFFFDFEF5D2E974BA002E97400007FFFFFF",
INIT_2D => X"FFFFFBFDFEF5D2A954AA002E974BA087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFBFDFFF5D2E954BA007FC00BA5D7FFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA000002000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080005000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"A974AA0000104AAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974BA0000174AAFFFF",
INIT_32 => X"FFFFFFFFFFFFDFEF552E954BA080A000AAE3FFFFFFFFFFFFFFFFFFFFFFFEF552",
INIT_33 => X"02A95400087FFFFFFFFFFFFFFFFFFBFDFEF5D2E974AA000A07000007FFFFFFFF",
INIT_34 => X"F7FBFDFFF5D2A954AA082A924281C7FFFFFFFFFFFFFFFFFFBFDFEF5D2A974BA0",
INIT_35 => X"A557FFFFFFFFFFFFFFFF7FBFDFFF552E974BA0020924BA1C7FFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000E3FFFFFFFFFFFFFFEFF7FBFFFFF552E974AA0071C50B",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0000020000000000000000000000000000",
INIT_38 => X"74BA0000174BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954AA080017410FFFFFF",
INIT_39 => X"FFFFFFFFFFDFEF552E954AA0004000AAF7FFFFFFFFFFFFFFFFFFFFFFFEF552A9",
INIT_3A => X"E95410087FFFFFFFFFFFFFFFF7FBFDFEF5D2A954BA082E800AAA2FFFFFFFFFFF",
INIT_3B => X"FBFFFFF552E954BA002E97410087FFFFFFFFFFFFFEFF7FBFDFFF5D2A974AA002",
INIT_3C => X"57FFFFFFFFFFFDFEFF7FBFFFEF552E974AA082A820AA557FFFFFFFFFFFFFEFF7",
INIT_3D => X"5D2E954AA0051554BA5D7FFFFFFFFFBFDFEFF7FFFFFEF5D2A974BA0000020AA5",
INIT_3E => X"0000000000000000000000000000000000000AAFFFFFFFFFFBFDFEFFFFFFDFEF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_3,               -- Port A enable input
WEA      => wbe_a_hi_1024_3(2),               -- Port A write enable input
DIA(0)   => data_write_a(21),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_3(21),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_3,               -- Port B enable input
WEB      => wbe_b_hi_1024_3(2),               -- Port B write enable input
DIB(0)   => data_write_b(21),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_3(21),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_22_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"5290F4CDE914905A14A43D33F488243E17122300F55FEB189B343A1140548380",
INIT_01 => X"A54007B259F6A975386262000C344BA9573C6FF57B18A5FB0ABFCD3C2C5F4F0C",
INIT_02 => X"021DFF8C38B3C009D203551040030071869D0040180AA2DC53DB89BEA8204001",
INIT_03 => X"2603475A969D0475A969D0460EAA401005111011BD506954EDB40F5EF41434C0",
INIT_04 => X"922D9002100ED69E443D988B0D5400103E48003D0800011E803B06B5B9125A15",
INIT_05 => X"281B5A0C06000408F4DF9422010D8802022F2124A8022492580040440002021C",
INIT_06 => X"F780C4C052881ADA0E05440205DA50930FA182010004700083E220800440B588",
INIT_07 => X"049D028B93FB561833D8094A02F5EA92FD7247E10305C40040D136E6A023F7FC",
INIT_08 => X"00028241680A0E002A9400803A884B5B5206B7C2E53CA25144009007A64EBD64",
INIT_09 => X"41008810240240C6694008010392354010000560141801002028A83D2A08E06D",
INIT_0A => X"34000000848BCA6902A29C54539C020E11810098D4067EFF9FF284D483E2AB41",
INIT_0B => X"500001840000C80B410014088040F4A944B1AA313C0022AA0011C0DC00028001",
INIT_0C => X"80B14004D158C8CA24A1C2A870AA1C2A870AA1C2A870AA1C2A872550E1543800",
INIT_0D => X"80A14050A01509E050854498B5281A1C34E506A2C6898B52A154DAC6B6000850",
INIT_0E => X"0B03001A483A4146603050080410089180008800143D83888281A2034A850142",
INIT_0F => X"A4160600349075238473F1210006133835E92273612B3482C090068A0E84AC56",
INIT_10 => X"30060181BA1B13959DC08DA902458870201970B29602562B0581200D141D0959",
INIT_11 => X"E042021C040D0152C8058B3840F044708E7E1C20A0106EA166C13AFC14AA3804",
INIT_12 => X"080E004B0C17C1439A9838301DC1A8438EA32C009DC1A8255300650458A1D588",
INIT_13 => X"018010E186F110A908E3A8CB0026C9A610A908E6A60F0807626610E160589C4C",
INIT_14 => X"2A701667334005800B1605F043858125E0D04110408D2485CA034681E43A1E40",
INIT_15 => X"00646002304244A91102C93A2D608D2A258DF8034188200C050171A41108F084",
INIT_16 => X"110441104411044110441104411044110466C440446CA06951D4EA8010009804",
INIT_17 => X"0040100401004411044110441104411044110441104411044110441104411044",
INIT_18 => X"0401004010040100401004010040100401004010040100401004010040100401",
INIT_19 => X"F7DFBFDEFE8FF1F7DEBDDF7DF7D05122890000000003FFFFFFFF900401004010",
INIT_1A => X"9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7BFFDFD7DDDF7DF7D",
INIT_1B => X"F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE79E7",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000003F9FCFE7F3F9FCFE7F3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA000400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0800",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000002000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2A954BA000015400FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080402010FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2A954BA0004154BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A0004174BAFFFFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0800154AAFFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF552A974AA0000174BAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974A",
INIT_2E => X"000007FFFFFFFFFFFFFFFFFFFFFFEF552E974BA0804000AAA2FFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080400010000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E954AA080005000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000402010FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2A954BA000417410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"804154BAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974BA0000174AAFFFFFFFFFFF",
INIT_34 => X"FFFFFFFEF552A974AA0000104AAE3FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0",
INIT_35 => X"AA2FFFFFFFFFFFFFFFFFFFFFFFEF552E954BA000E124BAE3FFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000007FFFFFFFFFFFFFFFFFFFFDFEF552E954BA080A000A",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804000100000000000000000000000000",
INIT_38 => X"54AA000400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2A954AA080017410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"0174BAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A954BA000415400FFFFFFFFFFFFF",
INIT_3B => X"FFFDFEF552E974AA0804174AAF7FFFFFFFFFFFFFFFFFFFFFFFEF552A974BA000",
INIT_3C => X"2FFFFFFFFFFFFFFFFFFFFFDFEF552E954AA0004000AAA2FFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2A954BA082E800AAAAFFFFFFFFFFFFFFFFFFFBFDFEF5D2E954BA002A820BAA",
INIT_3E => X"0000000000000000000000000000000000000087FFFFFFFFFFFFFFFF7FBFDFEF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_3,               -- Port A enable input
WEA      => wbe_a_hi_1024_3(2),               -- Port A write enable input
DIA(0)   => data_write_a(22),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_3(22),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_3,               -- Port B enable input
WEB      => wbe_b_hi_1024_3(2),               -- Port B write enable input
DIB(0)   => data_write_b(22),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_3(22),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_23_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"EF20906D902424807BC8241BC81801B97D38AD3C0800103362A6741C80A12A02",
INIT_01 => X"001FFF8409F089003B4422000D80C80106804A7951C5B9D1C828043EA28838F9",
INIT_02 => X"E01CEE21649C82C40800000F9FFEFF8E72CA7F5FC2E22809925A0D3611C877F8",
INIT_03 => X"24000400402670400402670D48222DC1764446838624000080007460C40001BF",
INIT_04 => X"68403FFC020560E0443E21037C01FFFC0002EE00628BF0E02FAD781014085014",
INIT_05 => X"0112000202FBFFF00920017FF0F0628BFF8488890979800002F702002BB807A0",
INIT_06 => X"EF85788B681FC000000001FFF0010000000001F7CBC385F87C0BFFFF20040001",
INIT_07 => X"F6E200000000C1440E3AE408009120071070FA07A1CB23FFA403F0C4D23BF7C0",
INIT_08 => X"0BF87CA400804000003FF7FFD8880A034AC09662305AB10555421006891A1089",
INIT_09 => X"BE1F5FEA10092C0896A243FFC0008087FFBEF2000000001DFFC612C0C0400100",
INIT_0A => X"41FF0C2060501000600000000001BFFA800808189A657EF81DD0C00079CC8001",
INIT_0B => X"018C24110A860006C620C0312241C482B20400CC52492710CC80060020A81BFE",
INIT_0C => X"0C08866907048320C20C10030400C10030400C10030400C10030400608018210",
INIT_0D => X"040002000041500300100040000500C000801000C02400000952800001FFBF04",
INIT_0E => X"FC850015385380380CDB86106502C5043FFD5FFF00A04BC010A7724B10000800",
INIT_0F => X"89F90A002A70A710A51C01C05904014861433602A1CAF13F2110055614C72FC0",
INIT_10 => X"E02D02001C1E14981B43253EE50C8220180F1082E06397E07E42200AAC298E57",
INIT_11 => X"8421802400A90022B0070FAE18019214A380344920080B21A58B02AC60BACDF0",
INIT_12 => X"0A2A000C480B0704B54028101AC49C84BB4100009AC49C80857A82D20CE8CB22",
INIT_13 => X"01E00C8103416445C12ED0400027C5292445C12D500B0005A62D344CB241D095",
INIT_14 => X"132C907425604680038706A35132C94BDD011010404428886AC91B11311C8280",
INIT_15 => X"FF000470BE0692020328CA0028042054A92771C50FC070110001C1680809591D",
INIT_16 => X"00802008020080200802008020080200800800200200000000000008004807DF",
INIT_17 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_18 => X"8020080200802008020080200802008020080200802008020080200802008020",
INIT_19 => X"0000000000000000000000000000000000000000000000000000008020080200",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080002010FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974AA000400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000400010FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974AA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080000010FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E954AA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954A",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA000015400FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080002010FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974AA000400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000402010FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E954AA080005000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA080407000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA00041741",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080000010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000402010FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2A954AA080002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954AA080017410FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"552A954BA000415400F7FFFFFFFFFFFFFFFFFFFFFFFFF552A954BA080015410F",
INIT_3E => X"0000000000000000000000000000000000000F7FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_3,               -- Port A enable input
WEA      => wbe_a_hi_1024_3(2),               -- Port A write enable input
DIA(0)   => data_write_a(23),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_3(23),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_3,               -- Port B enable input
WEB      => wbe_b_hi_1024_3(2),               -- Port B write enable input
DIB(0)   => data_write_b(23),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_3(23),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_24_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100600007FFF000080108004000800020000840041000080808",
INIT_02 => X"FC5CA803400EB8209000000F9FFEFF8E7240FF1FC22409EA04018E50074017F0",
INIT_03 => X"11100400000000400000000D00002CC07400000090C080019001010A000001BF",
INIT_04 => X"68003FFC00040000000000008001FFFC0002EE00000370E007A100000000E468",
INIT_05 => X"0000000000F8BFF00920004DF0F00001DF8000000079800000F3000029980780",
INIT_06 => X"6E461803081FC000000001FFF0000000000001F7C3C380F87C019FFF00000000",
INIT_07 => X"600C2400013649609C8000980040814210254000A00B21FF2003F2A80D500000",
INIT_08 => X"0BF80000000000000003F7FFD88D2B4A02C0940062EC2804001610020408178B",
INIT_09 => X"8E1F5FE010092C0892A041FFC0000001FFBEF0000000001DFFC002C000000000",
INIT_0A => X"41FF0C0000000000600000000001BFFA0000005501AA00000CE2000009400000",
INIT_0B => X"018C0411020600048620C030020502000200000400490510CC00040020201BF4",
INIT_0C => X"0808064106040300C00C10030400C10030400C10030400C10030400608018210",
INIT_0D => X"0000000000004003000000000000001200580000000000000000000001FFBE00",
INIT_0E => X"0086C022005381380FDB96516140C6043FFD5BFF000041000000004110000000",
INIT_0F => X"80010D804400A7240C840C201D0210840043B4804012500021E0088014C04940",
INIT_10 => X"4109038041021C980200D06410C1924030008142E06024A00043C01100298092",
INIT_11 => X"587CC200002100C14428090A1D02348190814C09C010104025AA40041A0D8005",
INIT_12 => X"022E0030300B0E46177004208000D8C61D7004300000D884817B00011306B2D9",
INIT_13 => X"01E003060344710009875C018100013831000985DC000C20003C310006143B70",
INIT_14 => X"4001850EDC004780144806A64400186CBF8961104000C3807884000846EB9500",
INIT_15 => X"FF0006E08C063C0220002201490418082010A57263E0100008000290161E711C",
INIT_16 => X"00000000000000000000000000000000000000000000000000000000000007DF",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"F2D0AEEAF6E7CC1132CDB4441990000000000000000000000000000000000000",
INIT_1A => X"BEFBE79E79E79E79E79EFBEFBEFBEFBEFBEF9EF9EF9EF9EFA69861219575D75F",
INIT_1B => X"783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1EFBEF",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000783C1E0F0783C1E0F0",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0201000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A000400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA000400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000400000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402010000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"00002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080002010FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000400010FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA00040000",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020100000000000000000000000000",
INIT_38 => X"74BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"000010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA000002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974AA000402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000002010F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_3,               -- Port A enable input
WEA      => wbe_a_hi_1024_3(3),               -- Port A write enable input
DIA(0)   => data_write_a(24),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_3(24),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_3,               -- Port B enable input
WEB      => wbe_b_hi_1024_3(3),               -- Port B write enable input
DIB(0)   => data_write_b(24),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_3(24),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_25_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100200002000000080100004000000020000800041000080808",
INIT_02 => X"FC400086000000800000000F9FFEFF8E738FFF1FC204010000000111568DD7F8",
INIT_03 => X"00000400000000400000000D00002CC4740000008000000080000000000001BF",
INIT_04 => X"68003FFF64A564AC000000000001FFFE0082EF00010370E007A1000000004000",
INIT_05 => X"0A00040148F8BFF80920804DF0F00101DFC040000079C92484F30499299837C1",
INIT_06 => X"66041803081FC0E0801101FFFD000E41002299F7E3C380F87C019FFF81200096",
INIT_07 => X"000000080480AE00000080000000000000000000A00B21FF2003E00000000000",
INIT_08 => X"1BF80000400A02000003F7FFFA0008000200A0400008A0000014100200081000",
INIT_09 => X"8E1F5FFA53EFBCACB2E369FFE0010001FFBEF80C40630C7DFFEEBAF000800202",
INIT_0A => X"41FF0C0600000000600000000001BFFE00301000000000000CC020000140000C",
INIT_0B => X"01DCCC31222730A49620C030020100000200000400490D10EC00040220201BF4",
INIT_0C => X"0808064106240300C00C10030400C10030400C10030400C10030400608018210",
INIT_0D => X"0883044582114013412080000000000000000000000000000012800001FFBE00",
INIT_0E => X"00040020000180380FC386106140C6043FFD5BFF00A04B80608003CB120C1106",
INIT_0F => X"0000080040000200040400000100000000009480000240000100080000400900",
INIT_10 => X"0001000000000808000000240000020000000100006004800002001000008012",
INIT_11 => X"0001001808220000002004001900000080800008000000000022400000088000",
INIT_12 => X"0010000000000E00110000000000408009000000000040808063004000008200",
INIT_13 => X"6000000000046100000240000000001021000004400000000010210000001010",
INIT_14 => X"4000000404000800000000060400000088000001800000001084000000088000",
INIT_15 => X"FF800C608C041002000002000006100000002100000000180600000000100018",
INIT_16 => X"4110441104411044110441104411044510629041040D180400000010028047DF",
INIT_17 => X"1104411044110441104411044110441104411044110441104411044110441104",
INIT_18 => X"1044110441104411044110441104411044110441104411044110441104411044",
INIT_19 => X"FBA2894A196A8C5A2932EC15DA080800002FFFFFFFFFFFFFFFFFC11044110441",
INIT_1A => X"2492492492492492492410410410410410410492410492412000531215A69A6B",
INIT_1B => X"158AC562B158AC562B158AC562B158AC562B1588C46231188C46231188C49249",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000B158AC562B158AC562B",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080000010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000010FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08000000",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_3,               -- Port A enable input
WEA      => wbe_a_hi_1024_3(3),               -- Port A write enable input
DIA(0)   => data_write_a(25),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_3(25),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_3,               -- Port B enable input
WEB      => wbe_b_hi_1024_3(3),               -- Port B write enable input
DIB(0)   => data_write_b(25),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_3(25),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_26_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"E9264EAB20190CA3BA4997AA9002AE9C001006B0778015CFA17E0811039879C7",
INIT_01 => X"2FFFF9BB1F773C7F9BB07DFFFDD863FC5FFF3FEFFBBF9FFB22FFFBC7B9F30686",
INIT_02 => X"E06CCC62052E708180F6FFBFFFFCFFFFF9C7FF7FC24332E642090000074037F6",
INIT_03 => X"428003739CD9863739CD9869FE2B7DEAF300029E4E300DFE69A6E644E6FF473F",
INIT_04 => X"7C2FEFFFF5BA124F003DD31EAFFFFFEE9FF7EE6F4C0770FFD7DC7CA53997B2B1",
INIT_05 => X"DFFB5421C1F8BBFAFDBFFACDF0FFCC05DDDBFF3690F9EDB7F5F7AFF639BD7DE3",
INIT_06 => X"EFD044ABC817C3E3A74667FDFFB6FF5727CC3BFEF7C3FAF87FF59F7FFBFEF69F",
INIT_07 => X"00003002132462052E708180EF060C18E5BEFB051225CDFF7002C4EEDE77F6E0",
INIT_08 => X"3FFF7D5000EC75088ED3FF7FC8790E46426CE06CB1F8E041051831FA3068D77E",
INIT_09 => X"C05FD7FF9BEFBDCEFBEE59FEF44F6603EFBEFAFCC2E35E7FDFD147CCF3F583FA",
INIT_0A => X"67FF1C7FBFADEB31E35768E8ED6BFDF3EB3EBF9DDBCE7FDC1DF8A760F3EACC02",
INIT_0B => X"5BDDCC3B336F7C548667D47B7737AF3FD62601EDC25B3533DCEB07F262213FFC",
INIT_0C => X"5F9A06E19F4D93A0EA0F78C35E30D78C35E30D78C35E30D78C35E986BC61AE31",
INIT_0D => X"5FD7AFEFDFFAF59B6FF28FE1D80D73D840607307DCFE1D80EF69A004DFFFF7FF",
INIT_0E => X"0004001F8041897B2FFFC6D86D70CE04FFFFF3FF1F5F5475BD7F72E4D75EBFAF",
INIT_0F => X"F60008003F008237B0040A00010003E020023E0201F45EC0010007E01047D17B",
INIT_10 => X"00010001DC0004C81003DE050A700200001DC0006863E8BD8002000FC0208FA2",
INIT_11 => X"2200E400002801E1A00004C21C0206F60081800800007B00010F02007EC09A0E",
INIT_12 => X"0880007E000807C7C1A612001E0015C7C19C22001E0015C59DFE82011A311AA0",
INIT_13 => X"00001BC00101F60409F0670840070809760409F06984800780097604067D0010",
INIT_14 => X"81019F40042100001F800203D81019EC085614000085C80023D81009CF008A74",
INIT_15 => X"FF802FFDFFAFD082003B032FB987E04021D481D4000819060801E0D00001231D",
INIT_16 => X"EBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEFFBFBFBFBBFCFBB0FFDFEFFEF2DFFFFFB",
INIT_17 => X"BFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAF",
INIT_18 => X"FAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFE",
INIT_19 => X"475B15BCF491E166CC8553F86EDB5C88646FFFFFFFFFFFFFFFFFEBFAFEBFAFEB",
INIT_1A => X"861861861861861861861861861861861861869A69A61861AFBD54D5F871C71D",
INIT_1B => X"984C26130984C26130984C26130984C26130984C26130984C26130984C261861",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000984C26130984C26130",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040201",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_3,               -- Port A enable input
WEA      => wbe_a_hi_1024_3(3),               -- Port A write enable input
DIA(0)   => data_write_a(26),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_3(26),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_3,               -- Port B enable input
WEB      => wbe_b_hi_1024_3(3),               -- Port B write enable input
DIB(0)   => data_write_b(26),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_3(26),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_27_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"00080A40000A41248002029000050A088000008242A0004404480002000A1155",
INIT_01 => X"2FFFF1C11F781C129C107DFFFE0860941E81258CA2B71C2220EC1B86E1A00002",
INIT_02 => X"E1000000810000014400FF6FFFF0FFFFF8007F1FC21110005080200000221FF0",
INIT_03 => X"4080026318C18226318C1821302232EAE00002BE001115FE48620040840A863F",
INIT_04 => X"643D4FFC2530000F003D821C0BFFFF8E9EF79E6D440748FED70060842105B0B0",
INIT_05 => X"D6F39020D1F8A3FAFDBFBACDC8FDC405D1DB7F1490E5EDB7D5CBADB2385D79C3",
INIT_06 => X"6FE000A38007C3032646EFF1F0B6FF46A78C39F8E723F2E47FE59C7F9ADA2612",
INIT_07 => X"00002820000000810000014401060C180190310540118DFF1000C0849673F6C0",
INIT_08 => X"3FF779100062B12A8EC3F47FC80208808210880C00082050000110023068D030",
INIT_09 => X"005F07E09BFFBD07FBAC09F8E42922038F7DF8BEC2E39C5F1FD047CEF1B582D8",
INIT_0A => X"63FF5D5F9FADE911E81C09818109E1F16B16B71092CE7ED81CF403601228C402",
INIT_0B => X"1BFDCC39732F3554866AD57C37BEAF1C152201A4C05B7531D56B05B06A213FF8",
INIT_0C => X"5BCA06F18FC59380F00E34430D10C34430D10C34430D10C34430F0861A2186B5",
INIT_0D => X"5B56ADAB5FAAE58B2F628EA0C80FA3F04040510768EA0C80CC61A0044DFFC6EB",
INIT_0E => X"0004001D800188792CE79715710AE4047FFD23FF315D54358D593474955AB6AD",
INIT_0F => X"520008003B000297B0040200010003E020001F0201E44A400100076000579129",
INIT_10 => X"00010001DC00004A10035E0408300200001DC000086BC8948002000EC000AF22",
INIT_11 => X"02002400002801E1A00000C01E0202F60080800800007B00000782006EC0820A",
INIT_12 => X"0080007E000006A7C10602001E0001A7C10C02001E0001C18DE282010A311AA0",
INIT_13 => X"00001BC00000FE0401F04300400708007E0401F04180800780007E04047D0010",
INIT_14 => X"81011F40040100001F800002F81011EC080604000085C80001F810094F008034",
INIT_15 => X"FF800C6DDDAFD082001B03249887E04001D481D4000009020801E0D00001021F",
INIT_16 => X"AB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6BF1EBDABD8E270BF84A25C6ACB777E3",
INIT_17 => X"B6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6AD",
INIT_18 => X"6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADA",
INIT_19 => X"490E2168100481CA860402104A471688747FFFFFFFFFFFFFFFFFAB6ADAB6ADAB",
INIT_1A => X"000000000000000000000000000000000008200000000000200072F210000001",
INIT_1B => X"05028140A05028140A05028140A05028140A0500804020100804020100800000",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000A05028140A05028140A",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040201",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_3,               -- Port A enable input
WEA      => wbe_a_hi_1024_3(3),               -- Port A write enable input
DIA(0)   => data_write_a(27),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_3(27),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_3,               -- Port B enable input
WEB      => wbe_b_hi_1024_3(3),               -- Port B write enable input
DIB(0)   => data_write_b(27),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_3(27),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_28_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"02200AA400180030808802A900002A08001280A08A801044104A1000001818C3",
INIT_01 => X"0AA00011460214428114180000882214413D0A71592A01D92213D28005210202",
INIT_02 => X"0451110A012100884000AA30200000000C100040104112101100008888200000",
INIT_03 => X"448000318C52A20318C52A20148810200111100C211004AA00034204200A2200",
INIT_04 => X"04004001001A90110000121402AA0000003C00000500000040080421080D0080",
INIT_05 => X"4060000C8001000000002E000000050000001610300000010000802202040012",
INIT_06 => X"1000002080001111001222000425A1040026A008000000000000000009328280",
INIT_07 => X"2491008A00491201210088400122448908A20402000408001000040820000000",
INIT_08 => X"20058310402A160026500000028040101004200C840082115554000112244814",
INIT_09 => X"4140000800000060000720000102028000000490160801020002200011100010",
INIT_0A => X"020000081B34211082B694D4D294000020020381040000000200032040004400",
INIT_0B => X"4800210C19808400500010009110091500020B408810000100200020408B0000",
INIT_0C => X"01028000080118020023604858121604858121604858121604858090B0242C00",
INIT_0D => X"010000800920040804020A6058003108402043058C460580653020005A004039",
INIT_0E => X"00000002800008014004104104420A00C000200005000010040A0020CC000200",
INIT_0F => X"520000000500000010000200000000000000280000040A40000000A000001029",
INIT_10 => X"00000000000000C0000002000830000000000000480008148000000140000020",
INIT_11 => X"020024000000000000000440000000020000800000000000000C00000040020A",
INIT_12 => X"00800000000001804006020000000500400C0200000005400A90000000100000",
INIT_13 => X"0000000000018200001003004000000142000010018080000001420000200000",
INIT_14 => X"8000080000010000000000018800008000060400000000000310000008000034",
INIT_15 => X"000002040080000000110006B081400000400000000009020000000000002200",
INIT_16 => X"802008020080200802008020080200802101210810C39A66A90A85420413A820",
INIT_17 => X"0200802008020080200802008020080200802008020080200802008020080200",
INIT_18 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_19 => X"DE21102C110A00246972BD89A40A0C22E1000000000000000000002008020080",
INIT_1A => X"2082082082082082082082082082082082082082082082080D35050758C30C31",
INIT_1B => X"0582C160B0582C160B0582C160B0582C160B0580C06030180C06030180C08208",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000B0582C160B0582C160B",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_3,               -- Port A enable input
WEA      => wbe_a_hi_1024_3(3),               -- Port A write enable input
DIA(0)   => data_write_a(28),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_3(28),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_3,               -- Port B enable input
WEB      => wbe_b_hi_1024_3(3),               -- Port B write enable input
DIB(0)   => data_write_b(28),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_3(28),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_29_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"79964E4BA01DACAB9E659792D00AAE160002829C7FDFEFCEE97C2815039D70C3",
INIT_01 => X"0ABFF9AB0775343F9AB01DF80D5821FC0FFF3FEFD1AF9FF1207FFBC7B9720586",
INIT_02 => X"002CCC60050E700080F6AAA7BFFC007189C7FF2FC00330E602800000074037F6",
INIT_03 => X"468003210868A63210868A68DA017D207200021C4E200CAA6186A40042FF4300",
INIT_04 => X"7C2FE002F0900001003C5316A6ABFFE21F36E02F0D03701F47D41800109FB281",
INIT_05 => X"4979440580F9B808F49F6A4DF00F8D01DC4B97369078249370F482E62BA41462",
INIT_06 => X"B250442BC81001E1870223FC0BF7F11507C423FE33C078F803F19F00E936721D",
INIT_07 => X"00011080012460050E700080EF020408EC8CFA01122149FF700200665A35D260",
INIT_08 => X"2BFD055040A452000443FF00007906464068406C31F84000000831FA1028575A",
INIT_09 => X"805FD017102690AA694551FE30444681E0820AD40201423FC00122C493500172",
INIT_0A => X"0600002AFFBE2330815568A8AD6ABC02A02A0B0CCB463B4C0748A720B1EA4C00",
INIT_0B => X"0850400A11414C005005000B51158936D20601A98A10200308A002E240010BFC",
INIT_0C => X"05928020194918A22A2268C81A32068C81A32068C81A32068C81A99034640C00",
INIT_0D => X"058102C48970541944B20FA1580561D040406305587A158046282000DBFFF13D",
INIT_0E => X"000000028040890327DCD28928324400DFFFF0001F1F0050342D42A086040B02",
INIT_0F => X"F60000000500802010000A000000000000022A0000141EC0000000A01000507B",
INIT_10 => X"00000000000004C0000082010A700000000000006800283D80000001402000A0",
INIT_11 => X"2200E4000000000000000442040004020001800000000000010D000010401A0E",
INIT_12 => X"08800000000801C040A6120000001540409C2200000015441DAC800010100000",
INIT_13 => X"0000000001019600081027084000000956000810298480000009560002200000",
INIT_14 => X"800088000021000000000201D800088000561400000000002358000088000A74",
INIT_15 => X"00802594A282C0000033010FB181E00020400000000819060000000000002305",
INIT_16 => X"C0B02C0B02C0B02C0B02C0B02C0B02C4B12B312912831A27FCFE7FFB175B6FF8",
INIT_17 => X"0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02",
INIT_18 => X"B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C",
INIT_19 => X"BBCF9F96EE7FFDF7FE783FFDFFEA0C00602FFFFFFFFFFFFFFFFFC0B02C0B02C0",
INIT_1A => X"EFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEEBAEBAEBAEBAEBBFFDF9FBEFFFFFFE",
INIT_1B => X"BFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFBEFB",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000FBFDFEFF7FBFDFEFF7F",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_3,               -- Port A enable input
WEA      => wbe_a_hi_1024_3(3),               -- Port A write enable input
DIA(0)   => data_write_a(29),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_3(29),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_3,               -- Port B enable input
WEB      => wbe_b_hi_1024_3(3),               -- Port B write enable input
DIB(0)   => data_write_b(29),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_3(29),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_30_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"F7FFBFFEFF9FE1F7FFBFFFFDFFD0000000000000000000000000000000000000",
INIT_1A => X"9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7AFBD75F5FDF7DF7F",
INIT_1B => X"F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE79E7",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000003F9FCFE7F3F9FCFE7F3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_3,               -- Port A enable input
WEA      => wbe_a_hi_1024_3(3),               -- Port A write enable input
DIA(0)   => data_write_a(30),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_3(30),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_3,               -- Port B enable input
WEB      => wbe_b_hi_1024_3(3),               -- Port B write enable input
DIB(0)   => data_write_b(30),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_3(30),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_31_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"129000008004A00804A40000400800020000000C005FEA005800200400050100",
INIT_01 => X"255FF18019700810180065FFFC0040801E80258CA2951C2200EC0906A0804140",
INIT_02 => X"E0000000000000011000550FDFF0FFFFF0007F1FC200000044000000000817F0",
INIT_03 => X"0000024210A30024210A3001002220C06044469200040154482000408400043F",
INIT_04 => X"602D0FFC2420000E003D80080955FF8E1ECA8E2D400340FE870060842100B030",
INIT_05 => X"0213100040F8A3F8FDBF944DC0FDC001D1CB6904A061EDB6D4C30490281831C1",
INIT_06 => X"6FC000830007C202060445F1F0D25E4207A099F0E303F0E07FE19C7F80402412",
INIT_07 => X"0000200000000000000001100004081001103107000185FF0000C0849673F6C0",
INIT_08 => X"1BF27A00000000000883F47FC800080002008000000820440000100220489020",
INIT_09 => X"011F07E013EFBC06FBA009F8E00120038F3CF82C44630C5D1FC002CCE0808248",
INIT_0A => X"61FF0C06C48BC801600000000001A1F00110101092CE7ED81CF0004012288000",
INIT_0B => X"11DCCC31222730048620C4382204A608142002A440492530C401049020221BF8",
INIT_0C => X"0888066187448380E00C10030400C10030400C10030400C10030600608018210",
INIT_0D => X"080204010200418301208480800D02D00040100240A808008840800405FF8640",
INIT_0E => X"0004001D000180780CE386106100C4043FFD03FF101D40008001304018081004",
INIT_0F => X"000008003A000217A0040000010003E02000160201E040000100074000478100",
INIT_10 => X"00010001DC00000810035C0400000200001DC0000063C0800002000E80008F02",
INIT_11 => X"00000000002801E1A00000801C0202F40080000800007B00000302006E808000",
INIT_12 => X"0000007E00000607810000001E000087810000001E000081846282010A211AA0",
INIT_13 => X"00001BC00000740401E0400000070800340401E04000000780003404045D0010",
INIT_14 => X"01011740040000001F8000025010116C080000000085C80000C8100947008000",
INIT_15 => X"FF800C609C06D082000A03200806A040019481D4000000000801E0D00001001D",
INIT_16 => X"010040100401004010040100401004010060C040040C200950402090128057C3",
INIT_17 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_18 => X"0040100401004010040100401004010040100401004010040100401004010040",
INIT_19 => X"00000000000000000000000000001000802FFFFFFFFFFFFFFFFF810040100401",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_3,               -- Port A enable input
WEA      => wbe_a_hi_1024_3(3),               -- Port A write enable input
DIA(0)   => data_write_a(31),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_3(31),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_3,               -- Port B enable input
WEB      => wbe_b_hi_1024_3(3),               -- Port B write enable input
DIB(0)   => data_write_b(31),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_3(31),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_0_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"ED39BA795990D275FB4A6E96ACC4731DEA4598B0AFB54867F6EE4618C3749803",
INIT_01 => X"8AA0047D8607944AC7DA180001ECA2444042106208408208C20022E9173734B3",
INIT_02 => X"1A7DDD79F9A73E6CCA7DAAF00001000008478020113D98E382FEDF333027C80F",
INIT_03 => X"75D341110C58F31110C58F32A208921F8051500147A0E4AB3493FB3A01EBE240",
INIT_04 => X"86424001531009B100425A97B2AA0001E03501D0A39C8F0078420001106D0C4C",
INIT_05 => X"BCC8CA2EBF03400700402BB20F00239E20341699198600000B08694B16434804",
INIT_06 => X"103FB860B2800161F8432200012DA185F80F24081C3C0707800E600056881308",
INIT_07 => X"B24197ABCDA467F9A73E6CCAFDC3870EEEEC44E2BDFE220094D03022210C011C",
INIT_08 => X"240581B5695EAA80262C080032BF07C7C1FC3F8E94F65B11555EAFFC1C306758",
INIT_09 => X"7E40000BEC004170040DB60017FED1CC0001045002984202003DB931192D60A5",
INIT_0A => X"120071411A74315881A28C141118000C5A85A60444210123820B43B40804674D",
INIT_0B => X"0820008E514045BB514F0106D1D8599581D3A958BC104A89215AC14C48898403",
INIT_0C => X"C261C01C48B1584A0CA3E2687A9A1E2687A9A1E2687A9A1E26870CD061343885",
INIT_0D => X"D274E93A758FA8683AC54B287522E10A74AF4AA59C568752662F5AC218000002",
INIT_0E => X"FF83C002783A0904231C70470C7E0B92800224008AE09FAD4BD48D1FC5D3A4E9",
INIT_0F => X"5BFF078004F075885DFBF7E15C06101C55E921F1F80FAB7FE0F0009E0E903EAD",
INIT_10 => X"F12E0380231F13978FF023FAFDBD9870380230F2D6081F56FFC1E0013C1D207D",
INIT_11 => X"DE7F263C0C8700125C0F8F3C43F1F10BBF7EFC61E01804E1E6C8F8FE807F67FB",
INIT_12 => X"02BE00017C17C1007E5E2E3081C5AC007E6F0E3081C5AC44418D65FE45DEE55B",
INIT_13 => X"61E0042786F103E9F01F9BC3C120C5A703E9F01F978B8C20666703E9F8A0FFED",
INIT_14 => X"FA7E283FFB414F80005F05F10FA7E283F78F6511C048278DCA174FF038FF15B4",
INIT_15 => X"0066A20B61692F293185D8D724E15D3FCC6B7C236FE0691B0700132C1F0EF880",
INIT_16 => X"3A4E93A4E93A4E93A4E93A4E93A4E93A4F942F92E9628540AD2A91442525A000",
INIT_17 => X"A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E9",
INIT_18 => X"4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93",
INIT_19 => X"55F3898E09B56C74DAB15D1CF13501AA495000000000000000003A4E93A4E93A",
INIT_1A => X"082082082082082082082082082082082082082082082082082084E41DC71C71",
INIT_1B => X"E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F82082",
INIT_1C => X"FFFFFFFFFFFFFFF94A5294A5294A5294A5294A52800003E1F0F87C3E1F0F87C3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"3060C183060C187FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"BDEBA0000000000000000000000000000000000000000000003060C183060C18",
INIT_28 => X"168ABA002E82145085155545F7AA975EFFFAABDE00FFAEBDFFF5D2EAAAAAF7AE",
INIT_29 => X"7FFFE10005542145557FD5545FF8000155087FC0155F7D168B55007BFDF45085",
INIT_2A => X"7FFC0010080017555555568AAAFFFFD7545AA8028A00A2802AABAFF8028BEF5D",
INIT_2B => X"FF842AABAA2AE95545FFD168ABAF7AEAAAAAA2FFFDF4500043FE105D2E954BAF",
INIT_2C => X"5007FD7400550415410002E974BA5D5168A00A2D142155005142010FFAE820AA",
INIT_2D => X"FFF780000BA007FE8AAAFF803FFFF5D2A821550000000BA007FD55FF5D7FC014",
INIT_2E => X"000AAFBEAA00007BFDFFF082EBDF455D5142000082E82145FFD17DFEFFFD168B",
INIT_2F => X"DFD75D2AA8A80EA8E2FE3F000000000000000000000000000000000000000000",
INIT_30 => X"68B551475FAF6D1C556F0AA1C24AABEA495FC716F002A975FFE3AA95E00EBAEB",
INIT_31 => X"42A0070071C50BAFEF1FAE0016D56A16D557BC257D415E0216FA3F1E8FC0145B",
INIT_32 => X"8010E004924874825D7FEAA85487FD24AFE3D02DAAAE12BD5545A2803AA00005",
INIT_33 => X"120155EA568E870BAEB8A05A2AEA8B50F55A2F150005A3A438BD04AFAB8F550A",
INIT_34 => X"545E055FFBE81D0BE8EA8A3AA05A2A5504001C74BA42A1571E8028E3DB7816D0",
INIT_35 => X"A5C7E3DFFFE90B45B47ABA497A82FFAFD2A82485FD2415A105C21451ED42A002",
INIT_36 => X"00000000000000000000B55EAAA100AA1D0F6F480B6A555A2A57A002A3D5FDB6",
INIT_37 => X"5EFAAAAB5E1AF3AABFF45592E88A0AFE80A8B0A0000000000000000000000000",
INIT_38 => X"65F520EBE9EF67D7BEA1FD5D556ABEF5D557FEBA55022A3F70C6B405F4D2AE97",
INIT_39 => X"C114728007521170821CE0FDE69411A8DED57CE1055555E5F58EFFC01FE2CACB",
INIT_3A => X"42341D5DEEBEF55080034E0A592A4AD0079C75D6070CC5CBB0280C029ABAA3EB",
INIT_3B => X"7F353AAF6C77F7F20D968BF57812A95E02A2AAB5EB0F280800EFAEE9F5D18F31",
INIT_3C => X"C91565455C141E41887D58AC448B69C30E02116220415A9540AA854140A0A204",
INIT_3D => X"DE6BE93172D7D625B556EEAB157ABEBE1B4D792A4AD1183454180DD3FDCAAAB7",
INIT_3E => X"F0000001FF0000001FF0000001FF0000001FF01EABC4B8014174FF7DA80F52FE",
INIT_3F => X"FF0000001FF0000001FF0000001FF0000001FF0000001FF0000001FF0000001F")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_4,               -- Port A enable input
WEA      => wbe_a_lo_1024_4(0),               -- Port A write enable input
DIA(0)   => data_write_a(0),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_4(0),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_4,               -- Port B enable input
WEB      => wbe_b_lo_1024_4(0),               -- Port B write enable input
DIB(0)   => data_write_b(0),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_4(0),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_1_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"212C001411984004084D000508C53810A03D1450E839B003342114428A000803",
INIT_01 => X"00000019400B100A8196000000CC004400400002000000000000028001340000",
INIT_02 => X"052137AE8031800C0044009000000000061800001CD4019802AD04CCCFC20004",
INIT_03 => X"04514108C60C21008C6042108400000201440020505100000043C30E10E9F000",
INIT_04 => X"02104001011DEFE088805681920000008000004001900800004002108C280008",
INIT_05 => X"040002340105000200000000080001900010000108040000000008411600401C",
INIT_06 => X"1034001042800808201000000001000820020000102000040000000000800180",
INIT_07 => X"64BF81A15EDFDE8031800C00843060C19E030022103600000450020800040004",
INIT_08 => X"00008004691687AA840008000090248CC84E000046000311555521F183060AC5",
INIT_09 => X"0820800D08100171000DB000154440C800400500000852020011200201012021",
INIT_0A => X"02000040001000880A2A04445004000102002041000001008208001440004140",
INIT_0B => X"4820018A1140440078050040511000102000A008183000010002404400000000",
INIT_0C => X"1000C80008000C030030880C2A030A00C28030A80C2A030A00C28018D4061401",
INIT_0D => X"10040802050080200284401C0022880F009E08008205C0020118088018000000",
INIT_0E => X"0F03C00280000000420860C60C0C0B92C0000000004000010042000040102008",
INIT_0F => X"001E078005000108400005E11C0610000000288058000003C0F000A000100000",
INIT_10 => X"F10E0380000000C202300000008D187038000000480800000781E00140002000",
INIT_11 => X"806302380C870010000004400100110800007861E0180000000C400680000001",
INIT_12 => X"023E00000000018000580C308000050000610C30800005000215006800000101",
INIT_13 => X"61E0000000018100B0001843812000014100B00016030C20000141002880026D",
INIT_14 => X"400A20009B404F80000000018400A20044096111C04000000304026000501580",
INIT_15 => X"0046820040082300218450C2800010094000482141E060190700100000002200",
INIT_16 => X"020080200802008020080200802008020080008008600500A82A1100A8000000",
INIT_17 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_18 => X"0080200802008020080200802008020080200802008020080200802008020080",
INIT_19 => X"81328A46BABEFC54A0810C7452B4428A14000000000000000000020080200802",
INIT_1A => X"AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA28A28A28A28A2A8218D2C0C924925",
INIT_1B => X"E974BA5D2E974BA5D2E974BA5D2E974BA5D2E975BADD6EB75BADD6EB75BAAAAA",
INIT_1C => X"FFFFFFFFFFFFFFFD8C6318C6318C6318C6318C63000002E974BA5D2E974BA5D2",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"70E1C3870E1C387FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"5555500000000000000000000000000000000000000000000070E1C3870E1C38",
INIT_28 => X"EBDF455D2EAABEFF7FFE8BFF5D0002155557FFFFFF007FC21EFA2FFD74AAAAD5",
INIT_29 => X"AA95400552AAAABAFFD1574105D7FD75FFAAAA800AAF7AA974BAFFFBE8B45F7A",
INIT_2A => X"0517DF555D2EAAA1055000015500557DF45AAD1400BAA2AE801550051555EFF7",
INIT_2B => X"FFD540155557FD5400F78028BFFFFFBEAB55F780020AAAA80020AA082EAAB550",
INIT_2C => X"AFF842ABEF5D517DF55552A974AAF7AE820AA0851574BAA2D1574AA5D7BFDEBA",
INIT_2D => X"EFAAD1575EF557FFFE10557FFFFFFFFD56AAAAFFFFD7555AAD168B45AAAEAAAB",
INIT_2E => X"0005D7FFDF4500043FE105D2E954BAF7AE80010082A97410557FEABFFAAFBE8B",
INIT_2F => X"51C7A2FBD5490BFD1C056A000000000000000000000000000000000000000000",
INIT_30 => X"974BAF7FFEFB45FFAABDF55492AA8BC2EBDFEAF7F1F840017D4975D2FEF147FC",
INIT_31 => X"080BEF495FC71D54124924385FAAA8AAAE3D145410F7F1D55D71C002DABAEBAA",
INIT_32 => X"002D082082AB8B6DBEDB7DF7F540E2AE85028B40155145F7AF6DBED5450AA1C2",
INIT_33 => X"78E021FF1471FDEAAFFD56F16D5571D2E28E38E0216FA2D1E8E80140F45082B4",
INIT_34 => X"A2DA3FB7DAAD4AAAAF487BC70BFA97F7AF6D417E92482BF84020BA495557E3FF",
INIT_35 => X"55554ADBD7A2FFC7BEFF6FFD7FC7002FD74951D71EDFFABFD16FAAAE92BD5545",
INIT_36 => X"00000000000000000000547AB8F550A8010E00492487482FFFE82A85EBAE2FFC",
INIT_37 => X"1EF005162BEF047FD5545AAFBF7400FBF9424F70000000000000000000000000",
INIT_38 => X"714F8338AAAA1D0AE974AAF7FFFDF55F7AABFF55082CA8B4DF6C1E8F5E540002",
INIT_39 => X"EABEF75550ACBB7582225FF5843404547184164AA5D2EBEEB0A2D555410D3555",
INIT_3A => X"FEAAEB083BC1000FF8409000512AEABFFDF79DCBF755962010BDCBBC21455D7F",
INIT_3B => X"801F8BA0C57740BDAA0688E5405D57D412F7D55F5E50C7F401BAAE8403CF5A3F",
INIT_3C => X"5D16BABAA3EBC3157ABD5FFE55F2AA9FEAFDF7F431A9F7FFE81FF013A8001AFF",
INIT_3D => X"FB863550229BCABEB7DA403FFFDA2FBF7FED2C7F955445079E280A00C56145EF",
INIT_3E => X"0000000000000000000000000000000000000596EBEF55080034E0A592A4AD00",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_4,               -- Port A enable input
WEA      => wbe_a_lo_1024_4(0),               -- Port A write enable input
DIA(0)   => data_write_a(1),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_4(1),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_4,               -- Port B enable input
WEB      => wbe_b_lo_1024_4(0),               -- Port B write enable input
DIB(0)   => data_write_b(1),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_4(1),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_2_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10E006600180111284380310006289800480032283E000A34301002001A0817",
INIT_01 => X"0005A00810790848048044A54E404350404000720885800802000906E4910200",
INIT_02 => X"407004208400408044C600C50AA055254010541A110222841200000002402544",
INIT_03 => X"0600011004182401004102408C28414043101000408118000145840440F5C415",
INIT_04 => X"5035855703A2900A000CD3088400F40688C9844409060850925E58A4081A0221",
INIT_05 => X"0200840D1021A15AC50494894850890540D1E12020C6E510818500440A280090",
INIT_06 => X"113044094002801020440090A8011A1224AB9380552102442884882A20004097",
INIT_07 => X"000100880004428400408044860000008C022402102100AA40004404B5075460",
INIT_08 => X"15C23440408C862A2A12382A8A5244145048C06085008010141521F000001240",
INIT_09 => X"400582B9033AA0E7AA4110B0506744810554542450694E710A836188C2C00222",
INIT_0A => X"443518360012C2210B020414109130A28038188096A06B8C120CA440A9C00802",
INIT_0B => X"1345E53300EC68005605002964AF222A5704004D080211121C80024200821780",
INIT_0C => X"181080C1110C882202211488452213C88472213C88472213488441109A442231",
INIT_0D => X"008204440210091341208041000810C00000300220201800A908000038AD0284",
INIT_0E => X"00040002804180300E88D28D206A40000554815500481440300000C44A081100",
INIT_0F => X"000008000500828700000000010000000002380000A00000010000A010050000",
INIT_10 => X"00010000000004CA000214000000020000000000684280000002000140200500",
INIT_11 => X"000000000020000000000442100002840000000800000000010C000026000000",
INIT_12 => X"00000000000805A4800000000000152300000000000015801272000100210020",
INIT_13 => X"000000000101C00000C000000000000940000120000000000009600004050000",
INIT_14 => X"0000130000000000000002018000106000000000000000002380000141000000",
INIT_15 => X"55000190000000000002000280000000011080C0000000000000000000002310",
INIT_16 => X"40902409064190641906419024090244902A9003004800415120D4A190804241",
INIT_17 => X"0900409004090641906419064190240902409024090641906419064190240902",
INIT_18 => X"9044090040900409004190441904419044090040900409004190441904419044",
INIT_19 => X"75960040138D70C030B51C50C7D100A2052F81F81F83F03F03F0419044190441",
INIT_1A => X"0410410410410410410410410410410410410410410410410248602081659659",
INIT_1B => X"5128944A25128944A25128944A25128944A25128944A25128944A25128941041",
INIT_1C => X"FFFFFFFFFFFFFFFE1084210842108421084210843FFF825128944A25128944A2",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"7FD5FF555815607FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"2AA000000000000000000000000000000000000000000000007FD5FF55581560",
INIT_28 => X"FC21EFA2FFD75EFAA8415410AA8415555087BFFF55A2AA800BAFFAE954000800",
INIT_29 => X"84155EFA2AEBDEAAA2FBEAABA5D7FE8B555551421455D0002145552EBFEBA007",
INIT_2A => X"2AEBDF555D2E954BAA2AA974BAFFFFE8B45552EBDF45FFAEAABFFF7FFE8B55F7",
INIT_2B => X"AAAAAAAAAFFD1574105D7FFFF555D2AAAAAA5D2E820BAA2FBEAB5555557DF55A",
INIT_2C => X"50055575EFFF84021555D043DEAA5D04021EF557FC21FFAA8428BFFAAAA954AA",
INIT_2D => X"10085568A00FF80175FFA2D17DFEFF7800215500557DF55AA80001FFAA800015",
INIT_2E => X"0005D00020AAAA80020AA082EAAB5500517DF555D042AA10A284154005D00154",
INIT_2F => X"00AAFFAA9543A080038A2A000000000000000000000000000000000000000000",
INIT_30 => X"0017D5D20B8EAA007FC51C7A2FBD55D2BE800042AFE8E1557D0075D2F45BEAA8",
INIT_31 => X"AA8BC7EBDFEAFEFFD00105FFBC20BDEAAA2FBF8AAA557BE8B6D5D5FFABEF4904",
INIT_32 => X"FFEFB6D555578F7DB6A0BDF7D480E174BFA02A974BAF7F5EFB455D2ABDF55492",
INIT_33 => X"ED1FDE90E3A497492B6AAADAAAE3D155E105571D55D71C002DABA5524820BAB6",
INIT_34 => X"BE8F401D7B6A0001470155C51D0092A071555D5E3AE821D00001FF0871C016DB",
INIT_35 => X"5BE8555400550A38428007FED000E3DA3DFD5E3DFFFBD5A38A021551C5F7AF6D",
INIT_36 => X"00000000000000000000410F45082B4002D082082AB8B6D1C5B7DF7FF78E075C",
INIT_37 => X"5EF005560B55F7AA800AAF7AA954AA00042AAA20000000000000000000000000",
INIT_38 => X"ABEF057D68F5F5A00021EF55042AAAA007FD5555AAFBD7545FBB8020A3F7AE97",
INIT_39 => X"7DF55D7AABFF5428ACA8F45A6C1E8F5EFF84165EFF7802BAB0A2FFEAABA557BE",
INIT_3A => X"CA8AA80800020AAF7FBFFFEF04552ABFFFF841FFE75CA882108202E974AAF7D5",
INIT_3B => X"00151FF0C57401E5F3D1E00A1A884174A8FFAEBFEB0A2D55541051555694F002",
INIT_3C => X"2AA801455D7FE8BFFF680800FFF7AAA155F595542455512A975455D3AA8A0055",
INIT_3D => X"5D79FCAF774AE005BE7895554005D2A8A0B882FFFFE10AAAAAB755A66B6AF56A",
INIT_3E => X"00000000000000000000000000000000000000C3BC1000FF8409000512AEABFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_4,               -- Port A enable input
WEA      => wbe_a_lo_1024_4(0),               -- Port A write enable input
DIA(0)   => data_write_a(2),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_4(2),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_4,               -- Port B enable input
WEB      => wbe_b_lo_1024_4(0),               -- Port B write enable input
DIB(0)   => data_write_b(2),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_4(2),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_3_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"210C00A20020000108430020001600B8156021104940741B3530400E02B92203",
INIT_01 => X"014C9BCA58B1296D24A402C992500B69404040028804A0080A000416A8D90A08",
INIT_02 => X"C12026A484318004404405C9C66E331352180D468B8203980300204442E02B34",
INIT_03 => X"04000748D60D24648D60524C88804D0215011020D15018148040C10A70E1D58C",
INIT_04 => X"18283333240FE41244187308C9104D70944852640901083801750EB0A418C220",
INIT_05 => X"0613142D01912CC2A1B4140528348900C612A104201C689044340ED413A07649",
INIT_06 => X"119000034019881822104C5E68035250A222829710A0A02C18C01A9920842413",
INIT_07 => X"402F00AB0016CA0431800444841020509D038B021230C1990001C644C8273200",
INIT_08 => X"16905000408482088290E8E64010248C4A5AA840C2000110001521F0810A92E7",
INIT_09 => X"0003CE6581BD016342A951AB146C4480530C3B2A8088D3542651670200C1826A",
INIT_0A => X"00735D36209A8A20020894004284B660821030C8990467401218004041020002",
INIT_0B => X"512445B740457154562F957CC08B00093700080D0A4851001D8302D20A0A1530",
INIT_0C => X"00508650008008021021A40861021840869021A408610218C0869810D6043095",
INIT_0D => X"1C8508438450801043A08090380A8834207007022209038080190000999C8F84",
INIT_0E => X"000400200000C0002A48A206204C4205F3304B33004C0041006240140A1C310A",
INIT_0F => X"0000080040000083800400000100000000008400018040000100080000510100",
INIT_10 => X"0001000000000800000244040000020000000100002A0080000200100000A702",
INIT_11 => X"000000000020000000200000080002C000800008000000000022000006808000",
INIT_12 => X"0000000000000A2281000000000040A3810000000000402001400000022002A0",
INIT_13 => X"000000000004200001C0400000000010200001C0400000000010000004490010",
INIT_14 => X"0001070004000000000000060000104C08000000000000001000000903008000",
INIT_15 => X"CC004050CA0C00020220200070040000010401C4000000000000000000100008",
INIT_16 => X"4310E4310A4210A4210A4210A4210A4210A8D0830A68010001B4DA881048061C",
INIT_17 => X"21084290A4210A4210A4210A4210A4210A4210A4210E4310E4310E4310E4310E",
INIT_18 => X"90A421084290A421084390E4310C4390E4310C4390E4310C4290A421084290A4",
INIT_19 => X"015303C0C78C706428A14C586291000A044001FFE000003FFC004290A4210842",
INIT_1A => X"2492492492492492492492492492492492410410410410412821600001249249",
INIT_1B => X"51A8D46A351A8D46A351A8D46A351A8D46A351A9D4EA753A9D4EA753A9D49249",
INIT_1C => X"FFFFFFFFFFFFFFFC00000000000000000000000038F56351A8D46A351A8D46A3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"55AB02055AB0207FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"420000000000000000000000000000000000000000000000007FFFAB57FFFAB5",
INIT_28 => X"A800BAFFAE9554508002AA00AA843DF55FFAA955EFA2D168B55557BEAA000055",
INIT_29 => X"002AB55AAAA955EF005568A00087BE8BFFA2D155410AA8415555087BFFF55A2A",
INIT_2A => X"AAABFF5508003FF555D0002145552ABFEBA007FC21EF007FD75FFAA841541008",
INIT_2B => X"082EBDEAAA2FBEAABA5D7FC0155005168B455D042AB45F7FFD741000042AA10A",
INIT_2C => X"FF7FBEAB55F7AABDEBA5D7FC2010A2D1575FFF7AA975555D2E80145F78415545",
INIT_2D => X"EF5555554AA087BC01FFFFAAAAB55552A954BAFFFFE8B55552EBDE00F7AEAABF",
INIT_2E => X"000082E820BAA2FBEAB5555557DF55A2AEBDF555D2E954BA002EAAABA002A821",
INIT_2F => X"FB7D5D7FEAA3808554203A000000000000000000000000000000000000000000",
INIT_30 => X"1557D1475FAF45BEAA800AAFFAA95578080038A2AA28E3AF55E3A0BA5D7AADB6",
INIT_31 => X"BD55D7BE80004AA1E8E2AB55B6A0925D7085F6AA10087FEABD7AAD57AEBAB68E",
INIT_32 => X"F5D0438140E2FA38B6AEBFF6D1D04AAFFA41040017D5D20B8EAA007FC51C7A2F",
INIT_33 => X"D0A901FFFF801557D1C20B8EAAA2FBE80AA557BE8B6D5D5FFABEF49002FB55FF",
INIT_34 => X"5D20BDE00EBAAA8BC7EBDFEAFEFAB8ABAE925D21C7010EADB525D7FFAE975C75",
INIT_35 => X"F002EADA921420871D74971D24820875C21D5EB8AA8FFF012A954BAFFF5EFB45",
INIT_36 => X"000000000000000000001C24820BAB6FFEFB6D555578F7DB6A0BDF7DEB8E125F",
INIT_37 => X"B55A28408145AAFFFFFFF5D7FEAABA0051400A20000000000000000000000000",
INIT_38 => X"AB55FAD568AA2AFAE975EF555168B55F7AA800BAF7AA955EF00042AAA2A2AEAA",
INIT_39 => X"2AAAA007FD55558A7BD7145FBB8020A35D2ABEF55F7800015F087FEAA00007FE",
INIT_3A => X"968F575D003FF55F7D5420BA5D2ABFEAAF7AE9DFF759A82AEF70800021EF5504",
INIT_3B => X"FFD5145FBAC9755F05040255FFD84175EF55002AAB0A2FFEAABA557BEA3EF057",
INIT_3C => X"82E974AAF7D57DF45552A3FF10AA8429F45A7D5EAF5FFBAEAAA10554155400AA",
INIT_3D => X"FF843FFE77C80825BC052ABFE10550415557085540000005156155FE90A8F5C0",
INIT_3E => X"00000000000000000000000000000000000005500020AAF7FBFFFEF04552ABFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_4,               -- Port A enable input
WEA      => wbe_a_lo_1024_4(0),               -- Port A write enable input
DIA(0)   => data_write_a(3),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_4(3),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_4,               -- Port B enable input
WEB      => wbe_b_lo_1024_4(0),               -- Port B write enable input
DIB(0)   => data_write_b(3),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_4(3),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_4_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A108400020612C80284210081034849800A00030300004833522C82D04A16002",
INIT_01 => X"2043998A1839284D1CA0650E1E504368403008418984014902030806A0D10200",
INIT_02 => X"C120042200000000044441CE01E80F00A49043118680008002000000026208E4",
INIT_03 => X"040001020019200020011209CC0164C060000000690111040144800042F5C403",
INIT_04 => X"7029AF0F81A00010CCA47700CC513CAC0D0B8E02010740E19754080108988021",
INIT_05 => X"02139405007133C0712244CD20F20105D583000020E9892201D304D42A9835E1",
INIT_06 => X"9190440300078002014405D9EE814C0284A883B6D7038AE079059B7800048092",
INIT_07 => X"000100AA0004408000000004840400008D200102503000782000C00C8025C000",
INIT_08 => X"00728A00408403220811991E02120C044058080004000001101121F220000260",
INIT_09 => X"811001E1185B38AD23C3707AD46440818F3CF80EC423CA7D01D123C80200816A",
INIT_0A => X"45810810A01B40216361056D6150F41200280001900439001FD8A00041400000",
INIT_0B => X"11FC88076266E800D605402962A820211500024808010512C40106D222223B14",
INIT_0C => X"0408804116040B02C02C500B0C02C100B0C02C100B0402C300B0401618058611",
INIT_0D => X"040200050200501301208482200D00D0A0408402C4282200A84800009B878680",
INIT_0E => X"00000020000100024AC88300300060090F0D830F00025400300204D018000804",
INIT_0F => X"8000000040000206A2000800000000000000950002E010000000080000588040",
INIT_10 => X"0000000000000808000554000200000000000100006D0020000000100000BB00",
INIT_11 => X"0000400000000000002000001A0002504001000000000000002280000D800800",
INIT_12 => X"0800000000000E2C802000000000408D801000000000408012440000200110A0",
INIT_13 => X"000000000004680003A0040000000010280003800800000000102800000B0000",
INIT_14 => X"000005C0002000000000000620000158000010000000000010A0000B00000200",
INIT_15 => X"C30146200400104002602600400000000294004000000004000000000010001A",
INIT_16 => X"0080200000008020000000802000000080080000004090014134DA101288C6DB",
INIT_17 => X"0802000000000401806010040180601004018060100000802000000080200000",
INIT_18 => X"8060180601004010040080200802000000000000802008020000000000008020",
INIT_19 => X"C0A28A063807E0500014063450404882846FFE000003FFC00000010040100401",
INIT_1A => X"AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA28A28A28A28A2934C8D0CCD145144",
INIT_1B => X"68341A0D068341A0D068341A0D068341A0D068351A8D46A351A8D46A351AAAAA",
INIT_1C => X"FFFFFFFFFFFFFFFC0000000000000000000000001FE32068341A0D068341A0D0",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"408102040810207FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"800AA00000000000000000000000000000000000000000000040810204081020",
INIT_28 => X"168B55557BEAB4500554200000557FE10FFFBEAA10007FD7410FFAA97555082A",
INIT_29 => X"55574105D2A800AA00043FEBA5D7FEAA00007BE8AAAAA843DF55FFAA955EFA2D",
INIT_2A => X"57BC00AAA2FFEAAAAAA8415555087BFFF55A2AA800BAFFAE9555508002AA0000",
INIT_2B => X"A2AA955EF005568A00087BE8BFFA2D17DE1000517FE10AAAAA8AAA002E975455",
INIT_2C => X"FAA8417410A2D140000F7FBC2010A2D157400AAAE974AAAAAA974BA08002AB55",
INIT_2D => X"EFA2AABDEAA087BEAAAAA2FBD54BA080002145552ABFEAA007FC21EF007FD75F",
INIT_2E => X"00055042AB45F7FFD741000042AA10AAAABFF5508003FF55F7D568A00552EA8B",
INIT_2F => X"5400F7A49057D0824850B8000000000000000000000000000000000000000000",
INIT_30 => X"3AF55F7A0925D7AADB6FB7D5D7FEAB7808554203A145178E00FFFBE8A101475D",
INIT_31 => X"A9557D080038AAA145157428492E8008200043FE925571EFA380871C7028A28E",
INIT_32 => X"AEA8A9200249056D4175C5092AAF5FDA38BE8E1557D1475FAF45BEAA800AAFFA",
INIT_33 => X"AA4954281C0E2FB55B6A0925D7085F6AA10087FEABD7AAD57AEBA08517DE00AA",
INIT_34 => X"007FC51C7007BD55D7BE80004AAFEDB42028EBFBC2028BED152438AAA092492A",
INIT_35 => X"AF7DF6AA00412EAABFFAA803DEBA0875EDA80BEF1C743840040017D5520B8EAA",
INIT_36 => X"0000000000000000000041002FB55FFF5D0438140E2FA38B6AEBFF6DBE84AAEB",
INIT_37 => X"A00FFFFEAA105D5155410FF84021EF0800154B20000000000000000000000000",
INIT_38 => X"DEBA0851574B2AAAEAAB55F78400145AAFFFFFEF5D7FEABFF0051400A25D5568",
INIT_39 => X"68B55F7AA800BAF7AA955EF00042AAA25555410BA082E8201000043FE005D517",
INIT_3A => X"568AA200557DE00AAAAAAA000804001FF005575408AA557FEB2FFAE975EF5551",
INIT_3B => X"D1550AAAA8002010F2AC154B25F2ABFF55F7800015F087FEAA00007FEAB55FAD",
INIT_3C => X"800021EF55042AAAA007FD5555087BD6145FAAC000A2A6FBC00BAAAFBC00BAF7",
INIT_3D => X"F7AEBDFF779A82AA43F7FBE8A00082EA8BFFAA843FEBA08517DE00F3F9574B30",
INIT_3E => X"000000000000000000000000000000000000008003FF55F7D5420BA5D2ABFEAA",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_4,               -- Port A enable input
WEA      => wbe_a_lo_1024_4(0),               -- Port A write enable input
DIA(0)   => data_write_a(4),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_4(4),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_4,               -- Port B enable input
WEB      => wbe_b_lo_1024_4(0),               -- Port B write enable input
DIB(0)   => data_write_b(4),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_4(4),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_5_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50DF4A0791B3FCB694379283C81FD996A091832102004A336A20E03C040C002",
INIT_01 => X"805FBDC69830A84D5C6A60000C34C26841280A00084000C8C212892EEAD53235",
INIT_02 => X"3B2026B578918E640A4F01CF8011FF0002080000082CA9998276DF7772C7C80D",
INIT_03 => X"37134108420D700084205702A4008A1D9100002171C0E0051554D93A11F5D140",
INIT_04 => X"8A41A0FC03A56DA000425A819410E3816C086198A388B702A8CA1210844A0C4C",
INIT_05 => X"B1808A062E8BC835F5E84532D708238A282F00A9291224800A2861490343082C",
INIT_06 => X"903FB8483A90581859050424100940825C6184401CDC451B860A6507160C4100",
INIT_07 => X"D26F068BCC96CDF8918E640E96D1A3469D6300E2FFEA27F8E4D23248130E259C",
INIT_08 => X"0BFA82E568442B2A082C0A7E3014250D49DA37A2420619000002AFF48D1222E5",
INIT_09 => X"3F005001E40969289429360416DCD1C46083030604B1CA20C03DF83B0A2C60A5",
INIT_0A => X"14613C71005A10492B888120288F480D58858449026145B3830F449449062B4F",
INIT_0B => X"11AC04934AC648BFD727C031E64170A137D5AA5C3E4B0F8A3C58C34C002290E3",
INIT_0C => X"CA29C6CC50384B6AC6AC86AB31AACA6AB39AAC86AB39AACA6AB3055643559C31",
INIT_0D => X"C673E33CF28F38603855401985228A0614BD30A0A2819852011E5AC2B87F9182",
INIT_0E => X"FF87C002F87A803E460B2516510CA594FF0044FFA4B08BAC4BB2CD0F09CF84E3",
INIT_0F => X"0DFF0F8005F0F5100DFFF5E15D06101C55EB29F1E00BE53FE1F000BE1E802F94",
INIT_10 => X"F12F0380231F17D78FC029FFF58D9A70380230F2FE0017C37FC3E0017C3D005F",
INIT_11 => X"FC7F023C0CA700125C0F8F7E43F1F001BFFE7C69E01804E1E7CCF8FC003FF5F1",
INIT_12 => X"023E00017C1FC1A4BFD82C3081C5BD27BFE30C3081C5BD00C02365D645CEEF5B",
INIT_13 => X"61E0042787F181E9C1EFD8CB8120C5AF41E9C18FD60F0C20666F41E9F009FFFD",
INIT_14 => X"7A7C077FFF404F80005F07F187A7D14BFFC96111C048278DEB074F9930FF9D80",
INIT_15 => X"C064014B8B652E2B3120C81284641D3E8DBF7D636FE860190700132C1F0EFB80",
INIT_16 => X"38CE1384E3384E338CE138CE1384E33C4E3ECE32E128882551349A1CBAA44103",
INIT_17 => X"84E3384E3384E3384E338CE138CE1384E3384E338CE138CE1384E3384E338CE1",
INIT_18 => X"CE138CE138CE138CE1384E3384E3384E3384E338CE138CE138CE138CE1384E33",
INIT_19 => X"F5E5BB4E7F7B9DB7FF3A1B6DB7E8410A8C000000000000000000384E3384E338",
INIT_1A => X"BEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEF9F7CFDFDDCF3CF3D",
INIT_1B => X"BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEFBEF",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000001711C7BBDDEEF77BBDDEEF77",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"FDFFF00000000000000000000000000000000000000000000080000000000000",
INIT_28 => X"FD7410FFAA97410082A800AAAAAE955450055421FFFFFBC0010AAD5574BA557F",
INIT_29 => X"7FD74000055574BA5D7FD7555A2D5575EF55517FF5500557FE10FFFBEAA10007",
INIT_2A => X"0002AABA5D2ABFFFFAA843DF55FFAA955EFA2D168B55557BEAB5500554200000",
INIT_2B => X"5D2A800AA00043FEBA5D7FEAA00007BC00AAAAAEBDF45A28428B45FFD168BFF0",
INIT_2C => X"5080028A00A2FFFDE00F7D57FEBAFF80174BAAAD1555EF555555555005557410",
INIT_2D => X"BA5D2E821FFA2D5554BA557BD75FFAA8415555087BFFF55A2AA800BAFFAE9555",
INIT_2E => X"00000517FE10AAAAA8AAA002E97545557BC00AAA2FFEAAAA082A97545F7D5420",
INIT_2F => X"7010BEDF524AA5571FDFEF000000000000000000000000000000000000000000",
INIT_30 => X"78E00EBFBE8A101475D5400F7A49043D0824850B8A2AE9756D145B401FFFFFFC",
INIT_31 => X"FEAB7D0855420BA1471D74380851524BA5571D757DB6D5525EF555178F6D1451",
INIT_32 => X"8A28B6DEBDF6DBEF1C0A28AAA5524BFFFFA28E3AF55F7A0925D7AADB6FB7D5D7",
INIT_33 => X"5555057D145152428492E8008200043FE925571EFA380871C7028B6AEBDF45B6",
INIT_34 => X"BEAA800AAFFAA9557D080038AAAA2FBF8E10EBD578EAAFF8415482BED1555EF5",
INIT_35 => X"81C209256DFFDF420BA552A821FFB6DF574A85575C55EFBE8E1557D1475FAF45",
INIT_36 => X"0000000000000000000008517DE00AAAEA8A9200249056D4175C50920875FDA3",
INIT_37 => X"5FF5D7BC21EFF7FBD7400F7FBC00BA55557DFF70000000000000000000000000",
INIT_38 => X"01FF5D5568BE7555568A00AAFFEAA105D5155410FF84020AA0800154B2AAAA97",
INIT_39 => X"00145AAFFFFFEF5D7FEABFF0051400A25551554BA0051400BA5551575EFF7D14",
INIT_3A => X"1574B2FFAABFF45FFAAAABFFAAFFFDFFF552EA8AAA55043DFF7AAAEAAB55F784",
INIT_3B => X"8002410FFD5575EF5555421E75555400BA082E8201000043FE005D517DEBA085",
INIT_3C => X"FAE975EF555168B55F7AA800BAF7AA955EF00002AAA2A2FBE8A00A2D16AAAAFF",
INIT_3D => X"0055554088A557FEB25D00021FFFFFFC00BA552A821EFFFFFD74BA5D51575F7F",
INIT_3E => X"000000000000000000000000000000000000000557DE00AAAAAAA000804001FF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_4,               -- Port A enable input
WEA      => wbe_a_lo_1024_4(0),               -- Port A write enable input
DIA(0)   => data_write_a(5),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_4(5),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_4,               -- Port B enable input
WEB      => wbe_b_lo_1024_4(0),               -- Port B write enable input
DIB(0)   => data_write_b(5),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_4(5),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_6_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10800B0061A01002840002C03002818000402322520070B313301C4389B2082",
INIT_01 => X"250041CA3839684D18A160000C52426841000000090800090210080008110200",
INIT_02 => X"0020042080010000044654C0000C008010000000001020900200200002620814",
INIT_03 => X"060881021088200021080200E4000A0891000020610111500104C00000F14400",
INIT_04 => X"0880000100000002000052288144004281C050400100280000C8100000080001",
INIT_05 => X"928080840001100A08009000280201000850E022401400002028214043410820",
INIT_06 => X"10100518090012122100C808049310002040000410A0001400000200120840D2",
INIT_07 => X"000100800004400001000000860408108C22000A502010074120044800040001",
INIT_08 => X"50000040D0C4E2088003FD01C01004044058082004000000000121F020408244",
INIT_09 => X"00BF17E9001205A5204911F814444080400100020000D200DFD16400C2A40AA0",
INIT_0A => X"04611C17849000022862A1596C8B5DF04834948900000100220C244840000880",
INIT_0B => X"03AD0413424E4044D665C070C22602291504400D084915020448114080201000",
INIT_0C => X"5E08864011088B22D22C008B0022C408B1022C208B0822C608B1111600458010",
INIT_0D => X"4251A12CD28A300429688001000800000020280204001000A00804309A002182",
INIT_0E => X"0000000280402400420800000000006200FC10002442042429324294014E8CA7",
INIT_0F => X"A40000000500800840000800000000000002280018001480000000A010100052",
INIT_10 => X"00000000000004C2003000010240000000000000680800290000000140202000",
INIT_11 => X"2000C0000000000000000442000001080001000000000000010C000280001804",
INIT_12 => X"08000000000801C300A010000000156000902000000015101200002800000000",
INIT_13 => X"000000000101800038002408000000094000386028040000000940000ED40000",
INIT_14 => X"0003B000002000000000020180002A24005010000000000023000060C7000A40",
INIT_15 => X"3F0280090321000040A410C28108000160008094000810040000000000002300",
INIT_16 => X"284A5284A728CA5284A528CA728CA52C4A5A0A32A300940101349A0408240818",
INIT_17 => X"9CA1294A329CA5284A728CA7284A5284A728CA5284A528CA728CA5284A728CA7",
INIT_18 => X"CA3294A129CA3294A129CA1294A329CA1294A3294A129CA3294A129CA3294A32",
INIT_19 => X"F5F78BCE7F8FF0F4FA955F7CF7F40A80145D55555556AAAAAAAAA94A329CA129",
INIT_1A => X"8E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E39B6CEDECDDF7DF7D",
INIT_1B => X"F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE38E3",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000001A1A33F9FCFE7F3F9FCFE7F3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"555FF00000000000000000000000000000000000000000000080000000000000",
INIT_28 => X"BC0010AAD5574BA557FFDFFF087BFDF45F7AA974AAAAAA97555F784174BAF7D5",
INIT_29 => X"515555508043FE00F7AA97555A2FBD7410AA8428AAAAAAE955450055421FFFFF",
INIT_2A => X"7D1575EFFFAA9555500557FE10FFFBEAA10007FD7410FFAA97400082A800AA08",
INIT_2B => X"0055574BA5D7FD7555A2D5575EF55517FF55A2AA97400552AAAB45082E80155F",
INIT_2C => X"500554200000003DE10FFD5401FFF7AAA8A10082EAAB45A2FFC2000007FD7400",
INIT_2D => X"10AA803FE105D516AABAFF843FFFFAA843DF55FFAA955EFA2D168B55557BEAB5",
INIT_2E => X"000AAAEBDF45A28428B45FFD168BFF00002AABA5D2ABFFFF087BD5545007BFDE",
INIT_2F => X"256DEB84104BAFFD1525FF000000000000000000000000000000000000000000",
INIT_30 => X"9756D145B401FFFFFFC7010BEDF524AA5571FDFEF1C7BFFF55FFA095482B6A49",
INIT_31 => X"4904380824850381C5B5057D1C003DE28F7A49057DAAF5D2428A2842AAAAA2AE",
INIT_32 => X"2AAFB451C2A8017DE3DF525FFFFA49756D145178E00EBFBE8A101475D5400F7A",
INIT_33 => X"2F1C50381471D74380851524BA5571D757DB6D5525EF555178F6DAAA49542841",
INIT_34 => X"AADB6FB7D5D7FEAB7D0855420BA1C0E3FE00E3DB471EFE3AAAAA00082EA8B6DA",
INIT_35 => X"F1C7BD057D1C71FFE10A28038E1049516AAB8FF8428FEFA28E3AF55F7A0925D7",
INIT_36 => X"00000000000000000000B6AEBDF45B68A28B6DEBDF6DBEF1C0A28AAA5524BFFF",
INIT_37 => X"F55F78017400F780001FFAA84000AAFFD1401E70000000000000000000000000",
INIT_38 => X"20BAAA8428AA2AAAA975FF5D7BC21EFF7FBD7400F7FBC00BA55557DFF7557BFD",
INIT_39 => X"EAA105D5155410FF84020AA0800154B2557FC01EF55043FEAAFF80021EFA2D14",
INIT_3A => X"568BE7AA80174AA082ABDF555D2A821EFAAFBC01FFF780155F7555568A00AAFF",
INIT_3B => X"AEA8A10082EA8BEFAAD5554B25551554BA0051400BA5551575EFF7D1401FF5D5",
INIT_3C => X"AAEAAB55F78400145AAFFFFFEF5D7FEABFF0051400A25D2EBFE10AAFFD55EFA2",
INIT_3D => X"552EA8AAA55043DFF7557BC01EF55557DE00AA842AA0000516AABAFF8428BE7A",
INIT_3E => X"0000000000000000000000000000000000000FFAABFF45FFAAAABFFAAFFFDFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_4,               -- Port A enable input
WEA      => wbe_a_lo_1024_4(0),               -- Port A write enable input
DIA(0)   => data_write_a(6),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_4(6),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_4,               -- Port B enable input
WEB      => wbe_b_lo_1024_4(0),               -- Port B write enable input
DIB(0)   => data_write_b(6),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_4(6),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_7_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10844B00482258A2842112C02450418800002300500030B313300C418992002",
INIT_01 => X"000009CA3839684D1CA0E0000E51424840000000080000080200080008510204",
INIT_02 => X"0120042086010000044600C00008000004100000000260900200000002402004",
INIT_03 => X"8628A10000082400000002408400080011000000610008000208C00000E14400",
INIT_04 => X"0911800100A000000000524084000040000050001140200100C8100000080102",
INIT_05 => X"0300812401011000000000002000114008008060441000000020024093000000",
INIT_06 => X"9190431C0D4010100000880804010010800000041080081000000200010424B2",
INIT_07 => X"000100AA0004408601000004860000008C02000A103010006928040800062481",
INIT_08 => X"84000048D484C20888000A0002120484C048007004000000000021F000000244",
INIT_09 => X"00A06009881201A520491004106C48A04040002400A15A208001650004001020",
INIT_0A => X"C99E1060201002044809C1040140A001004808810000459033189C0A400118A0",
INIT_0B => X"102000024040484050050041648A0041140C500B08821054C000264120000400",
INIT_0C => X"0404A083260E0832132011880462011880462051881462051881D31018C40620",
INIT_0D => X"0001000080001000813094801A8F80F00A600B52602801A88848011118003700",
INIT_0E => X"000003C007C002808228010410082042C000C000000004001002000400040002",
INIT_0F => X"A4000007800F80C840000800009864038A1200081C0014800000F001F0200052",
INIT_10 => X"00002C0E00E0E4004038000102400002C0E00E0D20100029000001E003E04000",
INIT_11 => X"2000C04031100E0403D0700300080908000100000661801E1900040380001804",
INIT_12 => X"0840878083E8003780A01043203A101780902043203A10082410082880000000",
INIT_13 => X"0601E0187900181035E0240806483248181035E0280410C8198818100DDD0000",
INIT_14 => X"0403774000201021E020FA006040376C00501022131210722060806D47000A40",
INIT_15 => X"00928A0002000110888600C032128201519480D40009902430160403E0E00506",
INIT_16 => X"01000000020080601802000000000405000A0020020081014134928820480010",
INIT_17 => X"0802018040000000006018020080200804010000000000806018020080000004",
INIT_18 => X"0000000001806008020000001006008020080001004008020080201004000020",
INIT_19 => X"0000000000000000000000000000400A004618618618C30C30C3000020180600",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000000B0840000000000000000000",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"1555500000000000000000000000000000000000000000000080000000000000",
INIT_28 => X"A97555F784174BAF7D5555FFF780155EFAAAEA8ABAAAFBFDE0055556AA005D04",
INIT_29 => X"55555EFAAFFFDFEFAAAAAAB455D556AA00FFAE95555087BFDF45F7AA974AAAAA",
INIT_2A => X"02EAAAAA082EA8A00AAAE955450055421FFFFFBC0010AAD5574BA557FFDFFF55",
INIT_2B => X"08043FE00F7AA97555A2FBD7410AA8428AAA557BFDFFF55003DFFFF7FBEAA000",
INIT_2C => X"0082A800AAF7AE975FFA28000010552EBDE00007BEAAAAA2D140000085155555",
INIT_2D => X"45087FEAB455D516AB55557BD55FF00557FE10FFFBEAA10007FD7410FFAA9740",
INIT_2E => X"000A2AA97400552AAAB45082E80155F7D1575EFFFAA955555D51574AAAAFFD55",
INIT_2F => X"AE105D556AA10410E17555000000000000000000000000000000000000000000",
INIT_30 => X"FFF55FFA095482B6A49256DEB84104BAFFD1525FFFF8E175C7A2AAAAA82A2F1F",
INIT_31 => X"F524AA5571FDFEF415B575D7AAF1FFFD7AAAAAFB7D495F6AA10E3AE905551C7B",
INIT_32 => X"003AFEFEBFBEAA001C2EA8A821C2EAAA00A2AE9756D145B401FFFFFFC7010BED",
INIT_33 => X"EDB470101C5B5057D1C003DE28F7A49057DAAF5D2428A2842AAAA497BFAFFF49",
INIT_34 => X"1475D5400F7A490438082485038F7A4905C7A28A070384120BDE100075EAA82B",
INIT_35 => X"D495150492BEF1D2555087BE8B7D555F6AB57417BC05D7145178E00EBFBE8A10",
INIT_36 => X"00000000000000000000AAA495428412AAFB451C2A8017DE3DF525FFFFA49756",
INIT_37 => X"555A2AEA8A10AAD568A00555168A10002E9754D0000000000000000000000000",
INIT_38 => X"8A10AAAE8215D557BFDF55F78017400F780001FFAA84000AAFFD1401E7FFAA97",
INIT_39 => X"C21EFF7FBD7400F7FBC00BA55557DFF7007BD5555AAD57DF55AAAEBDFEF007BE",
INIT_3A => X"428AA2007FE8BFF080028BFFAAFFEAA105D2EAAA005D2AAAA18AAAA975FF5D7B",
INIT_3B => X"043DE0000516AA10F7FBD7408557FC01EF55043FEAAFF80021EFA2D1420BAAA8",
INIT_3C => X"55568A00AAFFEAA105D5155410FF84020AA0800154B2FF8402145A2AA954AA00",
INIT_3D => X"AAFBC01FFF780155F7005140000FFD140145007FE8BEF557BEAB55087FC215D5",
INIT_3E => X"0000000000000000000000000000000000000AA80174AA082ABDF555D2A821EF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_4,               -- Port A enable input
WEA      => wbe_a_lo_1024_4(0),               -- Port A write enable input
DIA(0)   => data_write_a(7),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_4(7),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_4,               -- Port B enable input
WEB      => wbe_b_lo_1024_4(0),               -- Port B write enable input
DIB(0)   => data_write_b(7),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_4(7),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_8_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00000648E2840112C00000418000002700500030B3132000400812082",
INIT_01 => X"100008480009004C04A100000252024840000000180800080200010040110204",
INIT_02 => X"0020042000490000004600804008000005100000000024900200000002400004",
INIT_03 => X"0A0C33400008082400000080A4004B0891000020610112000040C00000E5C000",
INIT_04 => X"18800001000000000000512080000040800150400824280110C8100000120200",
INIT_05 => X"908084A10100100200004080280008240810802206940000012C214451610800",
INIT_06 => X"81B000080860109021400008040000202048020414A0021400040200322824C1",
INIT_07 => X"000000080004408049000004860000008402001A50208000630C040800062483",
INIT_08 => X"440000428644212280800A00021004044048002124000000000021F000000244",
INIT_09 => X"00004009001001010008100414644410400102228000D20080114502006409A2",
INIT_0A => X"000051312000042200294429148A4801C80C8C81000045907118040340020832",
INIT_0B => X"4020000240404140004D0544C4AA0001150410090302500011C813428A000400",
INIT_0C => X"46501090008820240240409000240009000240009000240009000120204808A5",
INIT_0D => X"42D1A168D09A301468402480004780F00140080860280004085904309A002196",
INIT_0E => X"00783FC00044340242280000000000020000C0000442106419120004034685A3",
INIT_0F => X"8000F07F800088A80000081EA2F9EC0000064004081010001E0FF00011104040",
INIT_10 => X"0ED0FC7E00000422201080000202658FC7E0000021882020003C1FE000222080",
INIT_11 => X"018059C3F350FE0C00000002A0040500000103961FE780000110010090000800",
INIT_12 => X"FD41FF80000830200021C1CF600012200010D1CF600012121600100810000004",
INIT_13 => X"9E1FE000010A1802100004343ED8000898021000087073D80008980200800002",
INIT_14 => X"0080200000BEB07FE00002086008020000209AEE3F300000246020200000620B",
INIT_15 => X"0088881903210000440610C8000A808040000208901786E4F0FE0C0000000166",
INIT_16 => X"685A1685A769DA368DA368DA769DA36CDA121A11A141800011309284002C0810",
INIT_17 => X"95A5685A1685A5695A368DA368DA769DA368DA368DA7695A1685A1685A5695A1",
INIT_18 => X"5A1695A568DA368DA369DA768DA1685A1695A5685A168DA369DA768DA368DA16",
INIT_19 => X"A4028A0A543EBC57A10A1E75D64108080468618618630C30C30C69DA5685A168",
INIT_1A => X"9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7BF3CCD8DF5B2DB2C",
INIT_1B => X"F87D3E1F4F87D3E1F4F87D3E1F4F87D3E1F4F87C3E1F0F87C3E1F0F87C3E79E7",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000006A6D4F87D3E1F4F87D3E1F4",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"155FF00000000000000000000000000000000000000000000080000000000000",
INIT_28 => X"BFDE0055556AA005D0415555080000000087BEAA10F7803DE00FFAEBFFFF0800",
INIT_29 => X"2AA8AAA557FC0010F780154105D7FC2145005155555F780155EFAAAEA8ABAAAF",
INIT_2A => X"7FFFFF55AA80155FF087BFDF45F7AA974AAAAAA97555F784174BAF7D5555FF55",
INIT_2B => X"AAFFFDFEFAAAAAAB455D556AA00FFAE95555AAFFE8A00552EBFE00F7D17FF45F",
INIT_2C => X"A557FFDFFF5504000AAAAAAA8B55F7D140010552E821EFAAAABDF555555555EF",
INIT_2D => X"55AA8028A00A2D57FF45557BE8A00AAAE955450055421FFFFFBC0010AAD5574B",
INIT_2E => X"000557BFDFFF55003DFFFF7FBEAA00002EAAAAA082EA8A00002AA8A10F784021",
INIT_2F => X"FE10F7AEBAFFF080A175D7000000000000000000000000000000000000000000",
INIT_30 => X"175C7A2AAAAA82A2F1FAE105D556AA10410E17555080E000280071E8A00EB8E3",
INIT_31 => X"4104BAFFD1525FF492EA8AAA5571C2000FF8A17400557FC015514555757DFF8E",
INIT_32 => X"2ABDE10EBDF7AF6DE3FFF8F7DB68A105D71C7BFFF55FFA095482B6A49256DEB8",
INIT_33 => X"AA0BDF6D415B575D7AAF1FFFD7AAAAAFB7D495F6AA10E3AE90555A2FBE8A3849",
INIT_34 => X"FFFFC7010BEDF524AA5571FDFEF550E00082B6A0AFB55F7D1420104124821D7A",
INIT_35 => X"01C2EA8A00F7800017DA2842FA00B6D578F6D557FFDA00A2AE9756D145B401FF",
INIT_36 => X"00000000000000000000497BFAFFF49003AFEFEBFBEAA001C2EA8A821C2EAAA0",
INIT_37 => X"0BA08556AA00AAAABFE00F7AEAABEF082E955450000000000000000000000000",
INIT_38 => X"21555D51575EFFFAA97555A2AEA8A10AAD568A00555168A10002E9754D082E82",
INIT_39 => X"17400F780001FFAA84000AAFFD1401E7082EAAABA5D5140010F7AE974105D7BC",
INIT_3A => X"E8215DA2FFE8ABA082ABFE00AAFBEABFFAAFBEABFFF7AA80145557BFDF55F780",
INIT_3B => X"D540000000402145AA843FFFF007BD5555AAD57DF55AAAEBDFEF007BE8A10AAA",
INIT_3C => X"AAA975FF5D7BC21EFF7FBD7400F7FBC00BA55557DFF75D2E82010F7843DF45FF",
INIT_3D => X"5D2EAAA005D2AAAA185D2AAAA10F780021FFA2803DE10FFD16ABFF5D7BFDE10A",
INIT_3E => X"0000000000000000000000000000000000000007FE8BFF080028BFFAAFFEAA10",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_4,               -- Port A enable input
WEA      => wbe_a_lo_1024_4(1),               -- Port A write enable input
DIA(0)   => data_write_a(8),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_4(8),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_4,               -- Port B enable input
WEB      => wbe_b_lo_1024_4(1),               -- Port B write enable input
DIB(0)   => data_write_b(8),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_4(8),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_9_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00018248A2840112C00002C18000002300500030B3132000400812006",
INIT_01 => X"400008000000004C0020000000100248413C0A61590001D90213C10008110204",
INIT_02 => X"01A0042080010000054600C04008000004100000001020900200200002420804",
INIT_03 => X"024003400008012400000010E4004B0891000020610310000144C00000F5C000",
INIT_04 => X"1801800100E000000000510084000040010050020810200000C8900000320200",
INIT_05 => X"918004311104100000000000200008100800002000100000002C234415610820",
INIT_06 => X"81B00008080010100000980804000008800042041080001000100200322C2481",
INIT_07 => X"0000811800044080010000058600000086020002502080006000040800062C80",
INIT_08 => X"0000004001D4618008800A00061004044048002004000000000061F000000244",
INIT_09 => X"000040090802009420409004104444084001022400214A2080014400026401A2",
INIT_0A => X"04000071200000A003CA294140200800C80C8C8100004590111C040040120800",
INIT_0B => X"12210002404848502847040164880021150400080222000200C8034200000000",
INIT_0C => X"4610088010080421021040841021000841021000841021000841010800420820",
INIT_0D => X"42D0A16C529A321068500484000500D10042080040284000084900001A002196",
INIT_0E => X"00000002804000004228010410082002C000C0002400046419120410034285A1",
INIT_0F => X"A00000000500800800000800000000000002290008001080000000A010100042",
INIT_10 => X"00000000000004C2001000000240000000000000680800280000000140202000",
INIT_11 => X"0000C0000000000000000442020001000001000000000000010C800080000804",
INIT_12 => X"08000000000801A7802010000000152780102000000015000600000800000000",
INIT_13 => X"000000000101900011E0240000000009500011E0280000000009500004DD0000",
INIT_14 => X"000137400020000000000201C000136C00101000000000002340002947000240",
INIT_15 => X"0080881901210000000600C280028000419480D4000010040000000000002304",
INIT_16 => X"68DA368DA1685A1685A1685A1685A16C5A121A13A141950051309284A82C0010",
INIT_17 => X"85A1685A1685A1685A368DA368DA368DA368DA368DA368DA368DA368DA368DA3",
INIT_18 => X"5A1685A168DA368DA368DA368DA368DA368DA368DA3685A1685A1685A1685A16",
INIT_19 => X"0157344CCCF48DE68A895C38E2540A8010100000000000000000685A1685A168",
INIT_1A => X"14514514514514514514514514514514514D34D34D34D34D28E1004039248209",
INIT_1B => X"D268341A4D268341A0D069349A0D069349A0D068341A0D068341A0D068345145",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000014D490D069349A0D068341A4",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"EAABA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"03DE00FFAEBFFFF0800155FFAAFBE8B45002A974AAAA803DFFFAA843DF45FFFF",
INIT_29 => X"7BFDE00A2FBD7400F7FBFDFFFA2AEBDE00AAFBEAABA080000000087BEAA10F78",
INIT_2A => X"055401FFF7AEAAA10F780155EFAAAEA8ABAAAFBFDE0055556AA005D041555508",
INIT_2B => X"557FC0010F780154105D7FC2145005155555557BE8BEF007FFDEAAAAD1555EF0",
INIT_2C => X"AF7D5555FFF780154AA5D2AA8A10F7AA974AA082E80010A2AAAAA10552AA8AAA",
INIT_2D => X"BAF7D17FEBAA2AEBDF45002EAAABA087BFDF45F7AA974AAAAAA97555F784174B",
INIT_2E => X"000AAFFE8A00552EBFE00F7D17FF45F7FFFFF55AA80155FF080400145FFFBEAA",
INIT_2F => X"8FC7BE8A3DF7DF7F5E8A92000000000000000000000000000000000000000000",
INIT_30 => X"000280071E8A00EB8E3FE10F7AEBAFFF080A175D7BEF1E8B6D002090482B68E3",
INIT_31 => X"56AA10410E175550871FFE00A2FBD0400FFF5FDFC7B6A0BDE38B6F5E8A92080E",
INIT_32 => X"7BFAE82A2DB555C71C5B451D7FFAAA8A38FF8E175C7A2AAAAA82A2F1FAE105D5",
INIT_33 => X"2AEADA38492EA8AAA5571C2000FF8A17400557FC015514555757D5D71E8BEF14",
INIT_34 => X"B6A49256DEB84104BAFFD1525FFFF84174BA5D20AAA00E3AA904BA142A87010A",
INIT_35 => X"7000400155FFFBEDA82FFD57DEBAAAA0BFF7D0024ADA921C7BFFF55FFA095482",
INIT_36 => X"00000000000000000000A2FBE8A38492ABDE10EBDF7AF6DE3FFF8F7DB68A105D",
INIT_37 => X"BEF080402000F7AAA8B55FFAABDFEFF7D16AA000000000000000000000000000",
INIT_38 => X"FEAAFFD16AA00082E820BA08556AA00AAAABFE00F7AEAABEF082E95545F7D568",
INIT_39 => X"A8A10AAD568A00555168A10002E9754D00517DE00A2FFC2000F7D17FF55FF803",
INIT_3A => X"1575EF555568BEF5D7FE8A10AAFFD55555D7FD5555FFAAA8AAAFFAA97555A2AE",
INIT_3B => X"AE800AA552A97400A2AEBDEAA082EAAABA5D5140010F7AE974105D7BC21555D5",
INIT_3C => X"57BFDF55F78017400F780001FFAA84000AAFFD1401E7FF80174AA5D0028A00AA",
INIT_3D => X"AAFBEABFFF7AA80145080002145F7FBFFE00FFD17FEAAA2803DFEF08043FE005",
INIT_3E => X"0000000000000000000000000000000000000A2FFE8ABA082ABFE00AAFBEABFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_4,               -- Port A enable input
WEA      => wbe_a_lo_1024_4(1),               -- Port A write enable input
DIA(0)   => data_write_a(9),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_4(9),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_4,               -- Port B enable input
WEB      => wbe_b_lo_1024_4(1),               -- Port B write enable input
DIB(0)   => data_write_b(9),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_4(9),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_10_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00018248A2840112C00002C18000202300500030B3132000400992006",
INIT_01 => X"254008000000004C002000000010026840000000080000080200010008110204",
INIT_02 => X"0020042000010000004455800008000004100000000000900200000002400004",
INIT_03 => X"020001021089000021081000C400090011000000610001540104C00000F14400",
INIT_04 => X"0811800101A00002000050088554004200C840000000200080C8100000000001",
INIT_05 => X"030080001000100800009400200000000840E020201000000024024001200020",
INIT_06 => X"81B00008080012120004CC080492500280208004148000100000020020042493",
INIT_07 => X"0000000800044080010000048404081085020002502000006000040800062480",
INIT_08 => X"100202400084410808000A00021004044048000004000000000021F020408264",
INIT_09 => X"010040090002008420401004144440004040022484214A2080110108C2C00320",
INIT_0A => X"04004166A48A0001080000000000080080181881000045901118044040020800",
INIT_0B => X"1201000200484910000F0105602622291404020902005002018002400A022000",
INIT_0C => X"0440001011808020120004801120044800120004801120044800110002400884",
INIT_0D => X"008000440210100041308480800F82F00040180260A808008848000018002104",
INIT_0E => X"000000028040000002280104100820020000400020000440100204100A000100",
INIT_0F => X"040000000500800800000000000000000002280008000400000000A010100010",
INIT_10 => X"00000000000004C2001000010000000000000000680800010000000140202000",
INIT_11 => X"200000000000000000000442000001000000000000000000010C000080001000",
INIT_12 => X"00000000000801C0008000000000154000800000000015000410000800000000",
INIT_13 => X"0000000001019800180000080000000958001800000400000009580002800000",
INIT_14 => X"0000A0000000000000000201E0000A0000400000000000002360002080000800",
INIT_15 => X"0080881000000000000600C28102800060000000000800000000000000002306",
INIT_16 => X"401004010040100401004010040100441020D0030008840051309A90BA884010",
INIT_17 => X"0902409024090240900401004010040100401004010040100401004010040100",
INIT_18 => X"1004010040902409024090240902409024090240902409024090240902409024",
INIT_19 => X"F546890A940FE0D3971243555205428290100000000000000000401004010040",
INIT_1A => X"8A28A28A28A28A28A28A28A28A28A28A28A28A28A28A28A29554199854514514",
INIT_1B => X"2B95CAE532994CA6532995CAE572B94CA6532994CA6532994CA6532994CA28A2",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000002718E72B94CA6532994CA657",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"FDE1000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"03DFFFAA843DF45FFFFEAABA007FC2155F7D155545AA80001EFAAFBEAB45557F",
INIT_29 => X"042AB55FFD168B55AA8000010FFFBE8BFFF78402155AAFBE8B45002A974AAAA8",
INIT_2A => X"AD16AABA002ABDE10080000000087BEAA10F7803DE00FFAEBFFFF0800155FF00",
INIT_2B => X"A2FBD7400F7FBFDFFFA2AEBDE00AAFBEAABAA2FFD741055003DFEFF7AA801FFA",
INIT_2C => X"05D0415555007FD74105555555EFF7FBC0145F78028A00A2D142155087BFDE00",
INIT_2D => X"55AAD168ABA002A975FFF7AEBDEBAF780155EFAAAEA8ABAAAFBFDE0055556AA0",
INIT_2E => X"000557BE8BEF007FFDEAAAAD1555EF0055401FFF7AEAAA105D042ABFF5D556AB",
INIT_2F => X"71D7AAFBEFB455D71F8E00000000000000000000000000000000000000000000",
INIT_30 => X"E8B6D002090482B68E38FC7BE8A3DF7DF7F5E8A92007BC217DEBDB55555AA8E0",
INIT_31 => X"EBAFFF080A175D700042AB7DEBDB6DB55BE8E05000EBFFE8BC7E38E07145BEF1",
INIT_32 => X"0A3DFD7F7A4821D7A2D16FA82142EB8E00080E000280071E8A00EB8E3FE10F7A",
INIT_33 => X"ED1421450871FFE00A2FBD0400FFF5FDFC7B6A0BDE38B6F5E8A92B6FBD541049",
INIT_34 => X"A2F1FAE105D556AA10410E175550071D54104951555D7EBF5C5155E3842AA00B",
INIT_35 => X"8410E2ABD749516FB55BED16FA820820955EFE3AEBDEAAFF8E175C7A2AAAAA82",
INIT_36 => X"000000000000000000005D71E8BEF147BFAE82A2DB555C71C5B451D7FFAAA8A3",
INIT_37 => X"1EFA2FFD7545AAAE97555A2FBFDF455D556AA000000000000000000000000000",
INIT_38 => X"8B45AAAA95545F7D568BEF080402000F7AAA8B55FFAABDFEFF7D16AA00087FC0",
INIT_39 => X"6AA00AAAABFE00F7AEAABEF082E9554500042ABFFA2FFFFF45F7AE97400AAFFE",
INIT_3A => X"16AA00FFFBD5400082EBFF45F78400155A2D57FE00552EA8A00082E820BA0855",
INIT_3B => X"D557555A2802AA10FFD54214500517DE00A2FFC2000F7D17FF55FF803FEAAFFD",
INIT_3C => X"FAA97555A2AEA8A10AAD568A00555168A10002E9754D085155410085557555AA",
INIT_3D => X"5D7FD5555FFAAA8AAA002AAAB4508557DF55F7D17FE000804155FFAAAABDEAAF",
INIT_3E => X"0000000000000000000000000000000000000555568BEF5D7FE8A10AAFFD5555",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_4,               -- Port A enable input
WEA      => wbe_a_lo_1024_4(1),               -- Port A write enable input
DIA(0)   => data_write_a(10),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_4(10),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_4,               -- Port B enable input
WEB      => wbe_b_lo_1024_4(1),               -- Port B write enable input
DIB(0)   => data_write_b(10),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_4(10),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_11_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A101C4B05A0034CA2840712C2D001419000002300500030B31B20084EC992002",
INIT_01 => X"90000986B83028491800E0000C26426040000000080000088200080802512224",
INIT_02 => X"1A2004205E010640024D00800008000004100000040EC090820018003241A00C",
INIT_03 => X"28639100000C5C00000045C08400C8001100000061806A001618C03001E54400",
INIT_04 => X"1A800001000009A0804059A190000040400040008058220008C8100000120D4E",
INIT_05 => X"02000E81080250010000002022000058080400000E1200000020004401000004",
INIT_06 => X"819435143F20101010001008040800B8100102041088011100022200000024B2",
INIT_07 => X"90640D280884453E01064002944180008402001295BA100022E4340800062D82",
INIT_08 => X"400000093204802200280A0012160585C1D808D004000000000323F40C102244",
INIT_09 => X"380040098010001100009204107C5950400000220080C200800900020C006827",
INIT_0A => X"80007100004016EA080801010000080D00200081000045B0511D289940103399",
INIT_0B => X"002000024040410A000D0104408810C115D9C008050042400100D04E88000002",
INIT_0C => X"00655010009264201200C7B421ED0C7B421ED0C7B431ED087B43176843DA1085",
INIT_0D => X"0401020080400A10012494881A4F80F209500BB2602881A488485C1318002000",
INIT_0E => X"6619A540124814800228010410082022C00040002020090020220C9600040802",
INIT_0F => X"ACCC334A802491600C587949B6D0141B4CC600D5761B1599865A500490B86A56",
INIT_10 => X"BAC845542056A61686EC81E3A6CB68AA2C622C9A251C352B330CB4A0092170D8",
INIT_11 => X"BCCAD0B5A81536080CC6B21A21B1FC09CB0F1076D4A200B2AD4068F4101639B5",
INIT_12 => X"4D2CC281E31AA0103AB8D5514066380804B268A2E060901204112566F10AC418",
INIT_13 => X"D551443C47281002540B2C9AAAA8662A1152B202AE3554403028115AA88201A1",
INIT_14 => X"548A20A0492A2724A0621620402A020141F172FB182A32AB6845AB6200251BC9",
INIT_15 => X"00C00A000200074044E6801832728080D00A380B753952C4877E0104DDE4D124",
INIT_16 => X"0080200802008020080200802008020480080022020081010124988800400010",
INIT_17 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_18 => X"0000000000802008020080200802008020080200802008020080200802008020",
INIT_19 => X"55062608804180C0B10A42104201400204000000000000000000000000000000",
INIT_1A => X"00000000000000000000000000000000000820820820820801C4149470000000",
INIT_1B => X"0000000000000000040200000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000007E0F0000000000000100800",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"000AA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0001EFAAFBEAB45557FFDE10082ABDF5508557DF45002ABDFFFF7803DE10AA80",
INIT_29 => X"AEBFF45FFAEBFEAA002A801FFF7FFE8A10A28000000007FC2155F7D155545AA8",
INIT_2A => X"2AABFE10082ABFFEFAAFBE8B45002A974AAAA803DFFFAA843DF45FFFFEAABAA2",
INIT_2B => X"FFD168B55AA8000010FFFBE8BFFF78402155AAD155555A28428BFF002ABDE00A",
INIT_2C => X"F0800155FF00557FF45557FC2010002A80010A2842AAAA007BFFF4500042AB55",
INIT_2D => X"FF5D00154BAF7FBE8BEFFFD540000080000000087BEAA10F7803DE00FFAEBFFF",
INIT_2E => X"000A2FFD741055003DFEFF7AA801FFAAD16AABA002ABDE10A2D168A10A284021",
INIT_2F => X"DFC7F78E3FE28B684070AA000000000000000000000000000000000000000000",
INIT_30 => X"C217DEBDB55555AA8E071D7AAFBEFB455D71F8E00002EBDF6D005B78F7D142AB",
INIT_31 => X"A3DF7DF7F5E8A92BEAEBFF7DEBA0BDEAA1C2A801C7E3FFEFA10B68407038007B",
INIT_32 => X"8A28BFF082ABAE10B6AAB8E280820B8FEFBEF1E8B6D002090482B68E38FC7BE8",
INIT_33 => X"07FF8F7D00042AB7DEBDB6DB55BE8E05000EBFFE8BC7E38E07145B6D15756DA2",
INIT_34 => X"EB8E3FE10F7AEBAFFF080A175D708517DF7D497BC5028142A87000A28A2AA920",
INIT_35 => X"0B6DB6AA28A280001FF5D0A10482FFFFEFBC7E3DF42028080E000280071E8A00",
INIT_36 => X"00000000000000000000B6FBD5410490A3DFD7F7A4821D7A2D16FA82142EB8E0",
INIT_37 => X"FEF007BE8BFF5D2ABDF55F7AABDEAAF784154BA0000000000000000000000000",
INIT_38 => X"DE00FF84154BA087FC01EFA2FFD7545AAAE97555A2FBFDF455D556AA00082EBF",
INIT_39 => X"02000F7AAA8B55FFAABDFEFF7D16AA00FFAEBFFEFAA803DEBA5D2E82155A2FBF",
INIT_3A => X"A95545F7D5555FFAAAAA8BFF002AAAA00FFAAA8AAA080028BFFF7D568BEF0804",
INIT_3B => X"2E95400A2AEA8A00007FEABFF00042ABFFA2FFFFF45F7AE97400AAFFE8B45AAA",
INIT_3C => X"82E820BA08556AA00AAAABFE00F7AEAABEF082E9554508557DFFF007BD54BA5D",
INIT_3D => X"A2D57FE00552EA8A00FFFFE8AAAAA80001FF5D2E82000F7FFFFF45AAFFC20BA0",
INIT_3E => X"0000000000000000000000000000000000000FFFBD5400082EBFF45F78400155",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_4,               -- Port A enable input
WEA      => wbe_a_lo_1024_4(1),               -- Port A write enable input
DIA(0)   => data_write_a(11),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_4(11),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_4,               -- Port B enable input
WEB      => wbe_b_lo_1024_4(1),               -- Port B write enable input
DIB(0)   => data_write_b(11),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_4(11),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_12_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50080B01BC002006940202C0DE041196A83183000000023322287E0FC000006",
INIT_01 => X"75400D849830C84C5823E0000C17424840000000080000088200002802153231",
INIT_02 => X"18A026B43ED180040147558040090000061800000C06ED9802768F4472C52005",
INIT_03 => X"2A67E34A528D0524A52850528400C8001100000171C02B550618C91A10E55440",
INIT_04 => X"1BC0000100056C8280825DE98154004300C840800850240080CA921084520A07",
INIT_05 => X"02000F832000500C0000941024000852084060202E100001002000448100000C",
INIT_06 => X"819A1D1C3FE01A1A40045408049A50BA4020C6041090001200006200000000F2",
INIT_07 => X"C26A0719CC96CC6ED18A64019695A854870300FA3968B20068FC06080106249F",
INIT_08 => X"D002024B3E040800008C0A002610240D494A06F3460409000000E3F0AD5282E5",
INIT_09 => X"27A06009200040000400120412445D78400001000410420080218029CC807A27",
INIT_0A => X"18000006848A026F000000000000080000F010C100204593F11A6CDF48003BF8",
INIT_0B => X"000000820040402B28050400400432C9349DF21A31A00ACC0000F04F80020001",
INIT_0C => X"00357804611AE45D05D0833430CD0833420CD0C33420CD0833430668619A1000",
INIT_0D => X"0000000000000A74812DF00E87E80A079F9F90FA0280E87E800C7FF3B8002000",
INIT_0E => X"3B6B0E404D26160682082002000401EA0000C40000800A006002818808000000",
INIT_0F => X"A476D61C809A4DA84272592D6246FC1B17B541F97E1B348EDA93900B2B286C56",
INIT_10 => X"30C669E622DBC325CFD881A962454CFBE5403AB99594362B1DB52720165650D9",
INIT_11 => X"F8D2D39A3745261E4A95A110A3F855000E4B1D32BAB504BB7490FCFF912A3834",
INIT_12 => X"B90E9B018C7530200AB8F8BF41F9A22006B37DC8E1F9A21A70116D4C5080651C",
INIT_13 => X"118780319CCA08AB1001ACDF34B8F1C688AB1002AE3F7B807B6289F368828C4C",
INIT_14 => X"2AF020233376A5ECC016B1A827CDA21160F051DE610A34C50427E6E220323E4A",
INIT_15 => X"0077020000000439FDC05C5806781FAB46095A0B5199B0AC55521524F1864022",
INIT_16 => X"000000000000000000000000000000000026C000002884000130921092804010",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"8020080200000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0051B946088881360A95090CB054420290100000000000000000008020080200",
INIT_1A => X"041041041041041041041041041041041049249249249249200100002D451451",
INIT_1B => X"92C964B2592C964B2592C964B2592C964B2592C86432190C86432190C8641041",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000003800F592C964B2592C964B25",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"7DE1000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"ABDFFFF7803DE10AA80000AAAA843FE0008557DFFF0800020105D557FEAA0055",
INIT_29 => X"D5420000051555FFA2AA8200000557DFFFF7AA80000082ABDF5508557DF45002",
INIT_2A => X"82AA8AAAAAFFC00BA007FC2155F7D155545AA80001EFAAFBEAB45557FFDE10AA",
INIT_2B => X"FFAEBFEAA002A801FFF7FFE8A10A28000000A2D155410F7FFFFEBA08003FE000",
INIT_2C => X"5FFFFEAABA000028A105D2ABFE10A2AABFE1055516ABEF5D517DEAAA2AEBFF45",
INIT_2D => X"55002A820AA08557DFFFF7AA82155AAFBE8B45002A974AAAA803DFFFAA843DF4",
INIT_2E => X"000AAD155555A28428BFF002ABDE00A2AABFE10082ABFFEF0855420000004175",
INIT_2F => X"5010495B7AE921C517DE10000000000000000000000000000000000000000000",
INIT_30 => X"BDF6D005B78F7D142ABDFC7F78E3FE28B684070AABE803AE38145B78FD700000",
INIT_31 => X"BEFB455D71F8E00BED547038145B505FFB6A487000005F7AFD7F7A482038002E",
INIT_32 => X"F1FDE821C003FE001C2EAAAAAB6F5C2082007BC217DEBDB55555AA8E071D7AAF",
INIT_33 => X"D517DEAABEAEBFF7DEBA0BDEAA1C2A801C7E3FFEFA10B68407038B6D550428FF",
INIT_34 => X"B68E38FC7BE8A3DF7DF7F5E8A9200002FA285D20BDE28A2A4B8E10555B68BEF5",
INIT_35 => X"F085F47038140010555142082082005F7DFD7F7A482155BEF1E8B6D002090482",
INIT_36 => X"00000000000000000000B6D15756DA28A28BFF082ABAE10B6AAB8E280820B8FE",
INIT_37 => X"ABA5D7FEAB45080015410007FEAA0055517DE000000000000000000000000000",
INIT_38 => X"AB45F780020BA082EBFFEF007BE8BFF5D2ABDF55F7AABDEAAF784154BAF7802A",
INIT_39 => X"D7545AAAE97555A2FBFDF455D556AA00F7D1554BA5D7BC01FFFF8015410007FE",
INIT_3A => X"4154BAF7D1400BAFFD57FE005D043FE10552EAAAAAFFD140000087FC01EFA2FF",
INIT_3B => X"8428A105D7FEABEF55557DEBAFFAEBFFEFAA803DEBA5D2E82155A2FBFDE00FF8",
INIT_3C => X"7D568BEF080402000F7AAA8B55FFAABDFEFF7D16AA0008003FEBA55003DEBAA2",
INIT_3D => X"FFAAA8AAA080028BFF087BD54AA550402145550000010087FFFF45F78402145F",
INIT_3E => X"0000000000000000000000000000000000000F7D5555FFAAAAA8BFF002AAAA00",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_4,               -- Port A enable input
WEA      => wbe_a_lo_1024_4(1),               -- Port A write enable input
DIA(0)   => data_write_a(12),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_4(12),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_4,               -- Port B enable input
WEB      => wbe_b_lo_1024_4(1),               -- Port B write enable input
DIB(0)   => data_write_b(12),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_4(12),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_13_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10154A0441836CA2840512822007C18000E02700500030B31B300040081A042",
INIT_01 => X"00000804A000C04800020000000002404001000008220008A200100802110204",
INIT_02 => X"02200430000104000A4700804008000004100000000420918204D3033240400D",
INIT_03 => X"AA4003400008592400000590C40009141100000C6180C0000000C00001E14000",
INIT_04 => X"0800000102400120088054019000004160004190BAA0270000C8100000600206",
INIT_05 => X"21000012040610050040000227003AA0082400E94C1200000824424005220020",
INIT_06 => X"81963B180C001010580000080400000058000004109C00138000020024142581",
INIT_07 => X"002C8008000441600106400A9600010494020002B8AAA000EF003408000E2580",
INIT_08 => X"000000E48194408000A00A001210040441C80320040210000002ABF004102244",
INIT_09 => X"2A004009640040100400940412D4C4004000022000104200802D983000480120",
INIT_0A => X"8000202020401480000000000000080C90090881000145B0111A14004015080D",
INIT_0B => X"00000002004040AA08050400404040C11444000805200A402090024000008002",
INIT_0C => X"8410000A00280020020040800020040800020000801020000800010020400000",
INIT_0D => X"84A14250A055100050100490000500D00040080040290000084E4000B800610C",
INIT_0E => X"DCD13042BEDA36820228000000000000C000400081A08BC812A2092B02850942",
INIT_0F => X"89B9A260857DB400431969CA985D480949D32804A40AB137341C10B7D6A02EC0",
INIT_10 => X"E6ACA678001CE7D0296C213A460CA4271CA2168AEC1017606E6838216FAD4055",
INIT_11 => X"84AD4961C281B20213073C5FC0058008632D30D522CE80239DCC01AB013A4D20",
INIT_12 => X"2E6B13804A4B01D83461299900F6BD583A519104A0EEBD1A141010B2A4C8E116",
INIT_13 => X"89E5E40913419151EE0E94641828F72B5151EE0D184B321037AF5158BB02D085",
INIT_14 => X"562EC0B42162D68EE0073AE1C562EC13D521921A4170300B2B458B56B01C2280",
INIT_15 => X"00888A120240034000E6DC8285028014B82372011FC1E4F5E0A00929684EAF84",
INIT_16 => X"50942509425094250942509425094254940A1421420082020120908800480030",
INIT_17 => X"0942509425094250942509425094250942509425094250942509425094250942",
INIT_18 => X"9425094250942509425094250942509425094250942509425094250942509425",
INIT_19 => X"F7EFBBEEFF3F7DF7FF3E9F7DF7E2450228000000000000000000509425094250",
INIT_1A => X"BAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBF7DFDFDDD555555",
INIT_1B => X"EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAEBAE",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000000000F7EBF5FAFD7EBF5FAFD7",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"2ABEF00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0020105D557FEAA00557DE10AAD5554BA087FFFF55557BD54AAF7FBC01FFA280",
INIT_29 => X"7BD75EF087FFFFEF557BEAB45552E80155AA802AB45AA843FE0008557DFFF080",
INIT_2A => X"FAE820AA5D5557555082ABDF5508557DF45002ABDFFFF7803DE10AA80000AA08",
INIT_2B => X"0051555FFA2AA8200000557DFFFF7AA80000AAD1420AA087BD7555FFD168AAAF",
INIT_2C => X"5557FFDE10AAAEA8BFFA2FBD7545FFD157555085140010F7AEAABFFAAD542000",
INIT_2D => X"BA557BE8A10A284154BAFFAAAAB45007FC2155F7D155545AA80001EFAAFBEAB4",
INIT_2E => X"000A2D155410F7FFFFEBA08003FE00082AA8AAAAAFFC00BA00002AAAAF7D5574",
INIT_2F => X"0492E3F1C71C7BE8A2ABD7000000000000000000000000000000000000000000",
INIT_30 => X"3AE38145B78FD7000005010495B7AE921C517DE10A2DB50482147FFAF554971D",
INIT_31 => X"E3FE28B684070AA1C71D25D7007FFAFD7497BE8B5555208217DBE8A2AB45BE80",
INIT_32 => X"7FD257DFFD568A82FFA4870BA555F5056D002EBDF6D005B78F7D142ABDFC7F78",
INIT_33 => X"FAAAFBFFBED547038145B505FFB6A487000005F7AFD7F7A482038AADF4709214",
INIT_34 => X"AA8E071D7AAFBEFB455D71F8E00A2A0ADBC7A2FFD257DE3DF52555085142000F",
INIT_35 => X"21C002AA92FFDF574824171EAA10B680124BAFFAAAFB45007BC217DEBDB55555",
INIT_36 => X"00000000000000000000B6D550428FFF1FDE821C003FE001C2EAAAAAB6F5C208",
INIT_37 => X"0105D7BE8B55085142010AAD157545F7AEA8B550000000000000000000000000",
INIT_38 => X"01EFF7AAA8B55F7802AABA5D7FEAB45080015410007FEAA0055517DE00A2FFC0",
INIT_39 => X"E8BFF5D2ABDF55F7AABDEAAF784154BA5D5140145007BE8B55087BEAB555D040",
INIT_3A => X"0020BAA2FFD54105D7FC21EFFFD16AA10FF80174AA557FC21EF082EBFFEF007B",
INIT_3B => X"FBC0155085540000FFAEBFFEFF7D1554BA5D7BC01FFFF8015410007FEAB45F78",
INIT_3C => X"87FC01EFA2FFD7545AAAE97555A2FBFDF455D556AA00A2803FF45AAFFC21EFAA",
INIT_3D => X"552EAAAAAFFD1400005D042AA00F7FBD5410085568A10FF80020AAFFAABFF550",
INIT_3E => X"0000000000000000000000000000000000000F7D1400BAFFD57FE005D043FE10",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_4,               -- Port A enable input
WEA      => wbe_a_lo_1024_4(1),               -- Port A write enable input
DIA(0)   => data_write_a(13),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_4(13),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_4,               -- Port B enable input
WEB      => wbe_b_lo_1024_4(1),               -- Port B write enable input
DIB(0)   => data_write_b(13),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_4(13),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_14_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10020A000180000284008280000281800000030000000033022000000580002",
INIT_01 => X"000008020000204D006800000030824840000000084000084200090008510200",
INIT_02 => X"0220043170010A600A4D008040080000041000000028009002000F333240800C",
INIT_03 => X"111813400008002400000000C400090011000000610200001104D83000F14000",
INIT_04 => X"0801800100A000000000540084000040000040000800200000C8100000000748",
INIT_05 => X"0100000000001000000000002000080008000000001000000024024001200020",
INIT_06 => X"819EB84028001010000000080400000000000004108000100000020020040081",
INIT_07 => X"92040608000440100102400A94810206844200021DA2A0002000340800062C80",
INIT_08 => X"000000000084400008800A001214040441481500040000000000A7F408002244",
INIT_09 => X"0A0040090002008420401004104444004000020400214A208001000002400120",
INIT_0A => X"0400002020000000000000000000080C8008088100004590111B480040120000",
INIT_0B => X"1000000200404800000504016000002114000008020000020080024000000000",
INIT_0C => X"0410000010000000000040001000000000000040000000000001000000000000",
INIT_0D => X"04810244825010004010000000000000000000000000000000080000B8002104",
INIT_0E => X"0002C38280001202020800000000001000004000000000401022000002040902",
INIT_0F => X"20000587050001404E8084341CBA3404800828805200008000E0E0A000080002",
INIT_10 => X"4D18178E012010C00224004091C3514072C000444A0400080001C1C140001000",
INIT_11 => X"51709A07424142084458476001003809D0104B01C5710044020C4006010500C5",
INIT_12 => X"C26EE3803180C18006519462A00005001460E4730000050A1011004001060049",
INIT_13 => X"01F9E00660318000000538318740000140000001B4600CE80001400000002B62",
INIT_14 => X"0000000AD89857B0E0684411800000003799EB764D000330C300000000E3554B",
INIT_15 => X"0000021002002C000024008284001A0902000422E3F5960080480A0216A07240",
INIT_16 => X"4090240902409024090240902409024090081021020080015134920800480010",
INIT_17 => X"0902409024090240902409024090240902409024090240902409024090240902",
INIT_18 => X"9024090240902409024090240902409024090240902409024090240902409024",
INIT_19 => X"F5579B4E5C8FF0F7BE9D5F7DF650400200000000000000000000409024090240",
INIT_1A => X"9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7BF7DDDDDFCF3CF3D",
INIT_1B => X"F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE79E7",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000003FFF03F9FCFE7F3F9FCFE7F3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"420BA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"BD54AAF7FBC01FFA2802ABEFA2FBE8B55A2AE80000F7D5555555D2AAAABAAAD1",
INIT_29 => X"AA801FFA28402000AAAE955455500155EF0804155EFAAD5554BA087FFFF55557",
INIT_2A => X"7AEA8B45080417400AA843FE0008557DFFF0800020105D557FEAA00557DE10A2",
INIT_2B => X"087FFFFEF557BEAB45552E80155AA802AB4500516AA00A2AE800BAFFFFC20BAF",
INIT_2C => X"0AA80000AA005568ABAA28402010A2843FEBAFFFBD7410A2D168BFF087BD75EF",
INIT_2D => X"005D7FFDF4555517DFEF00043FEAA082ABDF5508557DF45002ABDFFFF7803DE1",
INIT_2E => X"000AAD1420AA087BD7555FFD168AAAFFAE820AA5D5557555002E80155A280000",
INIT_2F => X"0555412AA8ABAAADB40092000000000000000000000000000000000000000000",
INIT_30 => X"50482147FFAF554971D0492E3F1C71C7BE8A2ABD7A2FFEDB55B6A080038E3DB5",
INIT_31 => X"B7AE921C517DE10A2AE851FFB68402038AAAA955554900105FF0800175D7A2DB",
INIT_32 => X"A0800BAE3F1C0092EBAAADB6D080A12410BE803AE38145B78FD7000005010495",
INIT_33 => X"2D568BC71C71D25D7007FFAFD7497BE8B5555208217DBE8A2AB451C556FA00A2",
INIT_34 => X"142ABDFC7F78E3FE28B684070AA00516DABAA28402038B6803DE82F7F5D5410A",
INIT_35 => X"D002A80155B680000105D7FF8F455D5F78FD7000E3FEAA002EBDF6D005B78F7D",
INIT_36 => X"00000000000000000000AADF47092147FD257DFFD568A82FFA4870BA555F5056",
INIT_37 => X"F55FF84000AAAAFBC0145002AA8AAAAAFFC20000000000000000000000000000",
INIT_38 => X"01EF080417555A2FFC00105D7BE8B55085142010AAD157545F7AEA8B55A2FBFF",
INIT_39 => X"EAB45080015410007FEAA0055517DE00A2AA955FFFF80020BAAAAA9754508000",
INIT_3A => X"AA8B555D557FE00A280020BAAAD140000A2AEBFFEF082A82010F7802AABA5D7F",
INIT_3B => X"803DE00FFD557400AAD56AB455D5140145007BE8B55087BEAB555D04001EFF7A",
INIT_3C => X"82EBFFEF007BE8BFF5D2ABDF55F7AABDEAAF784154BA08557FEAAA284000AAFF",
INIT_3D => X"FF80174AA557FC21EF082A80145F780020105D7BEAB45557BE8B45082EBFEBA0",
INIT_3E => X"0000000000000000000000000000000000000A2FFD54105D7FC21EFFFD16AA10",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_4,               -- Port A enable input
WEA      => wbe_a_lo_1024_4(1),               -- Port A write enable input
DIA(0)   => data_write_a(14),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_4(14),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_4,               -- Port B enable input
WEB      => wbe_b_lo_1024_4(1),               -- Port B write enable input
DIB(0)   => data_write_b(14),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_4(14),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_15_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000A000000000284000280000001800020030000000033022000000180002",
INIT_01 => X"8000080000000048000000000000026040000000080000080200000000110200",
INIT_02 => X"0020042004010E60004C0080000800000410000000020090020000300245E005",
INIT_03 => X"0000010000080400000000408400480111000000610008000000C00000E54400",
INIT_04 => X"980000010000000088C2550080000040000040000008A00028C8100000120000",
INIT_05 => X"020004012E025000000001322000000A28008000011000000220004D41000000",
INIT_06 => X"819588000800101000011008040000100001060418800510000A620000000092",
INIT_07 => X"0000000800044004010C20008440810284020002102220002000340800062480",
INIT_08 => X"0000000001140800002C0A001214050540C800400406180000002DF004000244",
INIT_09 => X"1E00400900000000000016041044400440000000000042008001000000000022",
INIT_0A => X"0000000000000220000000000000080C00000081000045901118000040000000",
INIT_0B => X"0000000200404000010500004000000114000009000000000000004200000000",
INIT_0C => X"0000000000000000000040001000040001000000000000000001000020000800",
INIT_0D => X"000000000000001001208000180800000000030200000180800C400030002000",
INIT_0E => X"0000000000002600020800000000001080004000000000000002000000000000",
INIT_0F => X"A400000000000000000008000000000000000000000014800000000000000052",
INIT_10 => X"0000000000000000000000010240000000000000000000290000000000000000",
INIT_11 => X"2001C05838120800000000000000000000010000000000000000000000001804",
INIT_12 => X"081004000000000000A010000000000000902000000000180010002020000000",
INIT_13 => X"6600000000000000000024080000000000000000280400000000000000000000",
INIT_14 => X"0000000000200801000000000000000000501001920000000000000000000A40",
INIT_15 => X"0000020000000000000000003000000000000000000A101C3614000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000080000120980000000010",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000400200000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"28BEF00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"5555555D2AAAABAAAD1420BAFF8000010082A954BA00003DFEF085155400F784",
INIT_29 => X"AE95555A2FBE8BEFA2843DE00AA8015400FF84001EFA2FBE8B55A2AE80000F7D",
INIT_2A => X"2FBEAB45F7D56AABAAAD5554BA087FFFF55557BD54AAF7FBC01FFA2802ABEFF7",
INIT_2B => X"A28402000AAAE955455500155EF0804155EFFFFBE8BFF0800174AA557BFDE10A",
INIT_2C => X"A00557DE10F7D1574AAA2D16AB55FFD568BEF087FE8A1055003FE00A2AA801FF",
INIT_2D => X"00AA802AA00AAAE800BA5D0015545AA843FE0008557DFFF0800020105D557FEA",
INIT_2E => X"00000516AA00A2AE800BAFFFFC20BAF7AEA8B45080417400FFFFC21450800154",
INIT_2F => X"8FD7005150438F78A2DBFF000000000000000000000000000000000000000000",
INIT_30 => X"EDB55B6A080038E3DB50555412AA8ABAAADB40092E38E070280024904AA1C043",
INIT_31 => X"1C71C7BE8A2ABD7E3AA9257DA2FFE8BC7BE8E38E10A28017400E38A051FFA2FF",
INIT_32 => X"00124AA557FFDE10A2FBEDB6DF7D16AABAA2DB50482147FFAF554971D0492E3F",
INIT_33 => X"10038E38A2AE851FFB68402038AAAA955554900105FF0800175D7E3FFEFBD700",
INIT_34 => X"000005010495B7AE921C517DE10FFDF50482A2DB6AB45FFD56DBD7087BEAA384",
INIT_35 => X"0FFF1C017D140410400BE8E28A10AAA085082550A1057DBE803AE38145B78FD7",
INIT_36 => X"000000000000000000001C556FA00A2A0800BAE3F1C0092EBAAADB6D080A1241",
INIT_37 => X"4AA0800020BA550028B550855400AAF7AEBDFEF0000000000000000000000000",
INIT_38 => X"7400AAAE975EFA2FBFFF55FF84000AAAAFBC0145002AA8AAAAAFFC2000AAAA97",
INIT_39 => X"E8B55085142010AAD157545F7AEA8B55AAAE821EFAAFBEAB55F7AAA8A00AA841",
INIT_3A => X"417555AAFFFDF450804020AA557BFFE10A2FFFFFEFF7D568ABAA2FFC00105D7B",
INIT_3B => X"D17DF45007FE8AAA08002AAAAA2AA955FFFF80020BAAAAA975450800001EF080",
INIT_3C => X"7802AABA5D7FEAB45080015410007FEAA0055517DE00FFFBC2000AAFBE8B55F7",
INIT_3D => X"A2AEBFFEF082A82010FFD5421EF5D0000010F7AAA8A10AA8017400552A801EFF",
INIT_3E => X"00000000000000000000000000000000000005D557FE00A280020BAAAD140000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_4,               -- Port A enable input
WEA      => wbe_a_lo_1024_4(1),               -- Port A write enable input
DIA(0)   => data_write_a(15),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_4(15),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_4,               -- Port B enable input
WEB      => wbe_b_lo_1024_4(1),               -- Port B write enable input
DIB(0)   => data_write_b(15),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_4(15),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_16_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"DA22C618B1000482B688B186588884862A400438255FC38381441205BA803003",
INIT_01 => X"7045A80028404C211203A952A90341080B173340412000E1005D628000820484",
INIT_02 => X"428406A4000850848330118D0AAC55001349B108818005460229044001C01784",
INIT_03 => X"092C4020000500020000500986812C405000001A48202050000A214AC0650115",
INIT_04 => X"4804A55440256F504025E003A054F46415A4E62B6FE3307943965A00001A1152",
INIT_05 => X"0000001C40A5B950ADB8EA097057ECE14C86D2B7F85AAD17F4B100000B88148C",
INIT_06 => X"415401DCDCF2C0A8030140BCB0820A200342A1C641C1E8782F508F2B00003584",
INIT_07 => X"002701881A3202080AE00480A2002840BE1480FA004342AA6F12000054004867",
INIT_08 => X"08C54828091002000002B32A8C19064E486A8001510000014140C1E2A14891E0",
INIT_09 => X"015452B103020814004088B64102680B6596594800400413CAC0208944800000",
INIT_0A => X"96AA000484094C000000000000012C9000A0000D0A80000BF8028E87C1B99270",
INIT_0B => X"014808A02004200E540480212000A448C0082024AE50064B44000000000002A2",
INIT_0C => X"0004000D5846256AAEA811150445411150445411150445411150422A088A8200",
INIT_0D => X"00000004010042A204A0C5817D00005034052E40000817D00440004004AD3240",
INIT_0E => X"632B2673FA4587978A2004102800809225545155121740000004900090000000",
INIT_0F => X"00C6564CE7F4EA4B940076D296D003030800462CBD320018CAAAACFE9164C800",
INIT_10 => X"28834ADB1440A114793A4A30A40839AA14910D08DCB2640031955559FD3AC990",
INIT_11 => X"594AB0B1A025371CA0E034E8443C097A800EB090D4AAC91208ED2FA0CE5E09B1",
INIT_12 => X"7B50446083001B94BB38C540EBE61284BB304880E3E4579EDC00992980D58033",
INIT_13 => X"5511121840E7A2CD952ECC12ABC3E6ACB3DFB12ECE315000F61FF1727A85FDBC",
INIT_14 => X"75DEB07F6F2E7084517F126F8395CB2BEFBAB8BA8AF698228CC5E2F08ECA5159",
INIT_15 => X"5580A840A8009F8B108C80A1021B080AFC0DF6422C6077F4A77F20D0C0E21084",
INIT_16 => X"0000000000000000000000000000000000044000102A0001148442A110810359",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"558D11544C690DA64C1C4F68A360400000000000000000000000000000000000",
INIT_1A => X"14D14D14D14D14D14D14D14D14D14D14D14514514514514529E5F87869E79E78",
INIT_1B => X"D1E8F47A3D1E8F47A7D3E9F4FA7D3E9F4FA7D3E9F47A7D1E9F47A7D1E9F4D14D",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000007D3E9F4FA7D3E8F47A3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"C00AA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"03DFEF085155400F78428BEF087FFFFEFF7D168B55AAD17FFFF552EBFE00007F",
INIT_29 => X"2E975EFF7D568BFFFF80175EF0004000BA552A821FFFF8000010082A954BA000",
INIT_2A => X"55540000082EAABFFA2FBE8B55A2AE80000F7D5555555D2AAAABAAAD1420BA5D",
INIT_2B => X"A2FBE8BEFA2843DE00AA8015400FF84001EF0000020AA5D00154005D043FF455",
INIT_2C => X"FA2802ABEF557BEABEF5D0415410087FD74BAAAAEBFFEF557FC00AAF7AE95555",
INIT_2D => X"FFFFAABFEAAFF84001FF002A821FFAAD5554BA087FFFF55557BD54AAF7FBC01F",
INIT_2E => X"000FFFBE8BFF0800174AA557BFDE10A2FBEAB45F7D56AABA082A97545F7D16AB",
INIT_2F => X"FFEF552AB8E38087FC2092000000000000000000000000000000000000000000",
INIT_30 => X"070280024904AA1C0438FD7005150438F78A2DBFF0871F8FC7E3D56AB6DBEDB7",
INIT_31 => X"AA8ABAAADB400924920925EFF7D16ABFFE38E175EF1400000BA412E871FFE38E",
INIT_32 => X"0A1240055003FF6D5551420101C2EAFBD7A2FFEDB55B6A080038E3DB50555412",
INIT_33 => X"57FC00BAE3AA9257DA2FFE8BC7BE8E38E10A28017400E38A051FF0804050BA41",
INIT_34 => X"4971D0492E3F1C71C7BE8A2ABD74975EDBC7550E12410087FD74AAB6AABFFC75",
INIT_35 => X"A08249756DF7D168BC7F7AABAEAAF780051C70824851D7A2DB50482147FFAF55",
INIT_36 => X"00000000000000000000E3FFEFBD70000124AA557FFDE10A2FBEDB6DF7D16AAB",
INIT_37 => X"B55A2D16ABEFFFFBFDFFF552AAAAAA007BC00000000000000000000000000000",
INIT_38 => X"20AA002A955EFAAAA974AA0800020BA550028B550855400AAF7AEBDFEF08516A",
INIT_39 => X"000AAAAFBC0145002AA8AAAAAFFC20000000021EFF7D568BFFA2AA955FF5D040",
INIT_3A => X"E975EF0800174BA002E820105D003DFEF5D51420005D2ABFF45A2FBFFF55FF84",
INIT_3B => X"7BD74AAF7AEBDF455D7BC20BAAAAE821EFAAFBEAB55F7AAA8A00AA8417400AAA",
INIT_3C => X"2FFC00105D7BE8B55085142010AAD157545F7AEA8B5500557DF45552A8200000",
INIT_3D => X"A2FFFFFEFF7D568ABA0804155FFF7D568B55FFAAAAABAFF8415545000015555A",
INIT_3E => X"0000000000000000000000000000000000000AAFFFDF450804020AA557BFFE10",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_4,               -- Port A enable input
WEA      => wbe_a_lo_1024_4(2),               -- Port A write enable input
DIA(0)   => data_write_a(16),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_4(16),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_4,               -- Port B enable input
WEB      => wbe_b_lo_1024_4(2),               -- Port B write enable input
DIB(0)   => data_write_b(16),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_4(16),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_17_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"5284CE4FB7BD2C8994A13392DBD02E14006B82AC7E800D44D3DD2FD5F9B961C0",
INIT_01 => X"2EACD01F7E03FC6793F2199B39FC233C11D93AE6F3BB92B32091DBC339B24542",
INIT_02 => X"E63CCCC00A82C08092A2AFAE667033DB50853379C10BFDC5C6F4044443C817C6",
INIT_03 => X"7FF183635AEF9E3635AEF9E18E237040404446965C0607EE6DB7854AC4DE060C",
INIT_04 => X"D78AC33FB604488B000892EF17BE6D84196482236FE100294152E294350FB697",
INIT_05 => X"081B5F9B409420D0CDB47A05403F6CE0C08A4AB7F840EDB6F48100DFC8081081",
INIT_06 => X"768465354781CBC30316367077B4BDB50646E8D87100A8201ED01C19C020F71A",
INIT_07 => X"4002A110C922480A82D0841147162C48EBB9537A0022DC67987042EE976ABEA7",
INIT_08 => X"DB931BFEF91C00002CC0E019C0C82A4E4820C15A2330E004401891181168C4D1",
INIT_09 => X"09F3A1BC11EFBC66DB65307071477FF1030C397C060B4254064302042F803A69",
INIT_0A => X"3F330802162F3B7EE3F3EC7C7DEF207000F00059D2ED56D7EED2ED3C9A867DC0",
INIT_0B => X"185C44B91BC1740B7605040BE0018CFC7429F326B9E822FFC00074D5A0AB033A",
INIT_0C => X"00367A28FC1B7F7FEFFCFBFF3EFFCFBFF3EFFCFBFF3EFFCFBFF3EFFE7DFF9E00",
INIT_0D => X"0000000008004BA78428C7AD7FC94B533F5B4FFBD2FAD7FCCA786D43FE67C218",
INIT_0E => X"BA494CEBFD4F2667ABB6F68B29760593F33FA0CF170F40006001B1A05C000000",
INIT_0F => X"7F749299D7FAEB237DFE5865B6D2BF23265CBACE542A6FEE92333AFF33E0A9BF",
INIT_10 => X"F6C24B6D18C3C9F8E2881F3F787D776B5DB94A09955054DFDD246675FE7AC153",
INIT_11 => X"BFB349E08FF9A27EDE9FA8AEFD9E7467BFCB195CFEB56A1A70D34D1706FFFA3E",
INIT_12 => X"6FE219CA80725B875EED723FF7FCB2875EDAAFEAF7FD929BFD55BBC71D79F639",
INIT_13 => X"546670D018E7A6E581D7B6AB75FDFCECA6E581D7BB5DDFC6FF0EB7D7E859FDB5",
INIT_14 => X"B978177F6D6AF5ECDB5FB76A5F5FA165B456E0FB308710C49FCFB741598B9C7E",
INIT_15 => X"CFDAAB00AC00A8BBFC8B501CF7A0FED9A540EA1952586CEB54D143ACFF9A3BA9",
INIT_16 => X"000000000000000000000000000000000026E100002F382DBD9ECFE117805F20",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"4372003009EDCC4052E917114F981800C0000000000000000000000000000000",
INIT_1A => X"BA69A69AEBA69AEBA69A69AEBA69AEBA69A69A69A69A69A68698686981D75D74",
INIT_1B => X"6A351A8D46A351A8D068341A0D068341A0D068341A0D46A341A0D46A341A69AE",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000000000046A351A8D46A351A8D4",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"7FEAA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"17FFFF552EBFE00007FC00AA087FFFFFFFFFFFFFEFF7FBEAB450804001EFAAD5",
INIT_29 => X"D168A000004020AA5D7BE8B450051401EF087FD74AA087FFFFEFF7D168B55AAD",
INIT_2A => X"D7FEAB55FF80175EFFF8000010082A954BA00003DFEF085155400F78428BEFAA",
INIT_2B => X"F7D568BFFFF80175EF0004000BA552A821FF5D00020BA552A82000552A821555",
INIT_2C => X"AAAD1420BAFFFFFDF45AAD17FFFFAAFBC01EF5D0015555557BFDEBA5D2E975EF",
INIT_2D => X"BA007FEABEF005555555A2D1554BAA2FBE8B55A2AE80000F7D5555555D2AAAAB",
INIT_2E => X"0000000020AA5D00154005D043FF45555540000082EAABFF00516AA10552E820",
INIT_2F => X"8B550000071EFB6DF7AE92000000000000000000000000000000000000000000",
INIT_30 => X"F8FC7E3D56AB6DBEDB7FFEF552AB8E38087FC2092147FFFFFFFFFBFDFC7EBF5E",
INIT_31 => X"150438F78A2DBFFBED16AA381C0A07082497FEFB6D1451471EF007BD04920871",
INIT_32 => X"2A850105D2A80155417BEFB6DEB8E175FFE38E070280024904AA1C0438FD7005",
INIT_33 => X"D7BFAEBA4920925EFF7D16ABFFE38E175EF1400000BA412E871FF550A0009249",
INIT_34 => X"E3DB50555412AA8ABAAADB40092FFF5FFF6DAADF7FFD7B6F1C71EF55001756D5",
INIT_35 => X"7145B6AA28492487082007FEDBD700515556DA2DF50492A2FFEDB55B6A080038",
INIT_36 => X"000000000000000000000804050BA410A1240055003FF6D5551420101C2EAFBD",
INIT_37 => X"FEFF7FBFFF55A2D16AB550000175EFFFFBEAA000000000000000000000000000",
INIT_38 => X"55EF087FC200008516AB55A2D16ABEFFFFBFDFFF552AAAAAA007BC0000557FFD",
INIT_39 => X"020BA550028B550855400AAF7AEBDFEFF7D568AAA5D2A97410007BFFFFF55515",
INIT_3A => X"A955EF5D2E80010002A954005D2A82155087FFFFEFAAAA975EFAAAA974AA0800",
INIT_3B => X"D1575FF5504175EF5D7FEAAAA0000021EFF7D568BFFA2AA955FF5D04020AA002",
INIT_3C => X"2FBFFF55FF84000AAAAFBC0145002AA8AAAAAFFC2000FFD57DFFFAAFFFDF55FF",
INIT_3D => X"5D51420005D2ABFF45557FE8AAA000415410007BFFF450051555EFA2FBC0000A",
INIT_3E => X"00000000000000000000000000000000000000800174BA002E820105D003DFEF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_4,               -- Port A enable input
WEA      => wbe_a_lo_1024_4(2),               -- Port A write enable input
DIA(0)   => data_write_a(17),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_4(17),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_4,               -- Port B enable input
WEB      => wbe_b_lo_1024_4(2),               -- Port B write enable input
DIB(0)   => data_write_b(17),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_4(17),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_18_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"69844019080000A21A611406840014122A641074155FC28A2024001001801003",
INIT_01 => X"7443D920034004180005E9E3C90360C0041C0181002001602025800008440084",
INIT_02 => X"E2DCCCE61D5C008103F2000781FC0FEDEAC2161B0B8FB0008620044443006010",
INIT_03 => X"884E300802006900802006995C896D605200000856E24A040000640052141103",
INIT_04 => X"480520FC026125AC0025C9122644E3E40EC8E2001001302281841A009038A86A",
INIT_05 => X"432000040089983070019400F01010004C8DB841405A80A100B586200FAC24AE",
INIT_06 => X"09044359DC7040000000002C109B0E0A00A1104641C0803804000707284600E1",
INIT_07 => X"400D10100400481D5EB08501620000007500CE801241021FE78E404860140060",
INIT_08 => X"00880C0106A0528020019307CC082A0A4A6A01ED725021400040D028000A9729",
INIT_09 => X"00117063038000282081402E4106400B6186128040600C10C1C0200950508110",
INIT_0A => X"C0C30C2E21580C874004008080003C32A10A19090C02010E1022944061688000",
INIT_0B => X"0180A8062026000DC425C0301311324AA2373088479105D044A1022000001835",
INIT_0C => X"0D89844703649000000200000000000000000000000000000000000000000010",
INIT_0D => X"0D8306C182701404C1973010802020404084001E00010802046092B5001FB365",
INIT_0E => X"528EB314068AB8B803DB00002900800400FC503F08180050942E4200020C1B06",
INIT_0F => X"40A51D66280D6032C5F96D3C51555D5D7D5AA87285820814A3CCC501C2A60820",
INIT_10 => X"8B35A3FEBF1FEDFD9C2B30E0468AAAD5D48F37E8FC1304102947998A03984C10",
INIT_11 => X"440FE1DD772D37A0A321BC6968F32658BF2D4F2A80BF8FE3F9FE3AC362080529",
INIT_12 => X"5487910D7E5A6D961A28456A1832E5161A100DD5182BC54020EA67A189C6ED36",
INIT_13 => X"AA444CAF91EDD1B725868403BE06323551B725868A100ABD119753B70964122B",
INIT_14 => X"EDC259048ACD868EE3803D65CEDC258A8F80D55E007C3F8EBB56F4C5362C978F",
INIT_15 => X"3F240014BE84370001B6922070440556B15F7FABBC0031BCF2257C41634B14D4",
INIT_16 => X"C1B06C1B06C1B06C1B06C1B06C1B06C1B0491069068000004060300A005A0118",
INIT_17 => X"1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06",
INIT_18 => X"B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C",
INIT_19 => X"B28BBECEB80EE173C2300F7DF16000000000000000000000000041B06C1B06C1",
INIT_1A => X"8A28A28AAAAAAA28A28A28AAAAAAA28A28A28A28A28A28A2910591505C104104",
INIT_1B => X"28944A25128944A25128944A25128944A25128944A2552A954AA5128944AAAA2",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000128944A25128944A251",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"9540000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"BEAB450804001EFAAD57FEAA087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974BA082E",
INIT_29 => X"7FFFFFFFFFBFDF45AAD568B55080028B55002E82000087FFFFFFFFFFFFFEFF7F",
INIT_2A => X"0043DE10AA843DE00087FFFFEFF7D168B55AAD17FFFF552EBFE00007FC00AA08",
INIT_2B => X"0004020AA5D7BE8B450051401EF087FD74AAAAFFFDF45A2D16AB55F7FFFFFFF0",
INIT_2C => X"0F78428BEFAA80000000804154BA55042ABEF5D7FD75FFAAD540145AAD168A00",
INIT_2D => X"00082E95555085168A10557FD7545FF8000010082A954BA00003DFEF08515540",
INIT_2E => X"0005D00020BA552A82000552A821555D7FEAB55FF80175EF5D00020105D2A974",
INIT_2F => X"DFFF5D2A954AA082A92428000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFBFDFC7EBF5E8B550000071EFB6DF7AE921C7FFFFFFFFFFFFFFFF7FBF",
INIT_31 => X"AB8E38087FC2092087FFDFC7E3F1FAF55A2DF6DB7D1C002AB7D002A82028147F",
INIT_32 => X"DF6DB7DE3F5FAFC708003DE28B68E38E280871F8FC7E3D56AB6DBEDB7FFEF552",
INIT_33 => X"ADF4516DBED16AA381C0A07082497FEFB6D1451471EF007BD0492B6F1F8F55AA",
INIT_34 => X"1C0438FD7005150438F78A2DBFFA28407038140410492550A2ABC7497BD25FFA",
INIT_35 => X"F5D0E05000492097428002E9557D1C516FA28417BD5545E38E070280024904AA",
INIT_36 => X"00000000000000000000550A00092492A850105D2A80155417BEFB6DEB8E175F",
INIT_37 => X"FFFFFFFFDFEFF7FBFFFEF552E974AA082A820AA0000000000000000000000000",
INIT_38 => X"ABEF002A800AA557FFDFEFF7FBFFF55A2D16AB550000175EFFFFBEAA00557FFF",
INIT_39 => X"6ABEFFFFBFDFFF552AAAAAA007BC0000087BFDF45AAD568B55AAFBFDFEF55042",
INIT_3A => X"FC2000FFD56AB45A2FFFDFFFAAD16AB4500043DEAAFFAEAAAAA08516AB55A2D1",
INIT_3B => X"2AA8B45087FC01EFA2FFD55EFF7D568AAA5D2A97410007BFFFFF5551555EF087",
INIT_3C => X"AAA974AA0800020BA550028B550855400AAF7AEBDFEFA280154BA55040000055",
INIT_3D => X"087FFFFEFAAAA975EF5D2E974000804154BA082A975EF5D517DEAA007BD5545A",
INIT_3E => X"00000000000000000000000000000000000005D2E80010002A954005D2A82155",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_4,               -- Port A enable input
WEA      => wbe_a_lo_1024_4(2),               -- Port A write enable input
DIA(0)   => data_write_a(18),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_4(18),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_4,               -- Port B enable input
WEB      => wbe_b_lo_1024_4(2),               -- Port B write enable input
DIB(0)   => data_write_b(18),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_4(18),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_19_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"042200000000000041088001001AA00000000000000000000000500802000003",
INIT_01 => X"040048000024000000000404000000000A22000800000800004A200000000001",
INIT_02 => X"200C8840085EB00480060000001C008002489E0F000405EA0004040404000000",
INIT_03 => X"24004000000000000000000900002C4050000000000069500208400002E14100",
INIT_04 => X"4800200C0000000044002000C80020E40000E200000130200188000000800100",
INIT_05 => X"000000000080181000000000701000004C8000000058800000B1000009880480",
INIT_06 => X"80500081081040000000002C100040400000004641C080380400070100000000",
INIT_07 => X"4020109801A4CE005C00048380142810010564C4100114012002402028044808",
INIT_08 => X"0070700000000000000083004C3902420062000020E0000100004082A140102B",
INIT_09 => X"001150200000000000000026400000016186100000000010C04002C000000000",
INIT_0A => X"007C00008082C0002000000000002C3000000004050001030102040000000000",
INIT_0B => X"0000000000000000000000000000010000800011000000000000000000000BC0",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"000000000000000000000000000000042000760000000000000000010004B200",
INIT_0E => X"0D74002280300F0002FB069040000060000C5003000800000000000000000000",
INIT_0F => X"C01AE8004500744C780687DBA828008080A5FC0D385598035D0008A00C015660",
INIT_10 => X"39D8140040201BF861F0E7D693E6170022408116DFE0AB3006BA0011401D02AC",
INIT_11 => X"5412E4997F5249FD005043B8680CC98F00D0F2DD0140100406FE053A98F6ECC7",
INIT_12 => X"7418663001858040E153888000010840E165D0000000285C246A181C03FE4662",
INIT_13 => X"8199830066F0020858385974000001260208583854E2200000660208D6B1423F",
INIT_14 => X"8235AC508FCE8811042040F008235AE04420C040CF00C031C80009B8F224978B",
INIT_15 => X"030004E00000C220010808C10D9A92A74CD7CF4A09051110AD5A3C9200B7F280",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000118",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"07208BBA3F0C7010C660C7441920000000000000000000000000000000000000",
INIT_1A => X"861869A61861861861869A61861861861861861861861861A8208C4C1534D34C",
INIT_1B => X"984C26130984C26130984C26130984C26130984D26930984C26130984C261861",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000984C26130984C26130",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"174BA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFDFEF5D2A974BA082E95400F7FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0004",
INIT_29 => X"FFFFFFFFFFFFFFFFF7FBFDFFF552E974BAA2FFFFE10087FFFFFFFFFFFFFFFFFF",
INIT_2A => X"004001EFAAAEA8ABA087FFFFFFFFFFFFFEFF7FBEAB450804001EFAAD57FEAAF7",
INIT_2B => X"FFFBFDF45AAD568B55080028B55002E82000F7FFFFFFFFFFFFDFEFA2D568B550",
INIT_2C => X"0007FC00AAF7FFFFFFFF7FBE8B55AAD16ABEF5D2ABFF55080402010087FFFFFF",
INIT_2D => X"55A2FFFDFEF5D2EBFE00AAFFFFEBA087FFFFEFF7D168B55AAD17FFFF552EBFE0",
INIT_2E => X"000AAFFFDF45A2D16AB55F7FFFFFFF00043DE10AA843DE00557FFDFEFA2D16AB",
INIT_2F => X"FFEF552A974AA0000104AA000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFF7FBFDFFF5D2A954AA082A92428E3FFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"0071EFB6DF7AE92EBFFFFFFFFFFFFDFEFF7F5FAFC7492A974AAB6F5F8E101C7F",
INIT_32 => X"F1F8FD7AAD16AB450000001FFBEA4A8AAA147FFFFFFFFFBFDFC7EBF5E8B55000",
INIT_33 => X"00000010087FFDFC7E3F1FAF55A2DF6DB7D1C002AB7D002A82028FFFFFFFEFF7",
INIT_34 => X"BEDB7FFEF552AB8E38087FC2092F7FBF8FC7E3F5EAB45B6DF6FBEF5D2AB8F7D0",
INIT_35 => X"84971F8FC7AAD56DB6DBEF5F8FD7412ABFE28B6F5F8E820871F8FC7E3D56AB6D",
INIT_36 => X"00000000000000000000B6F1F8F55AADF6DB7DE3F5FAFC708003DE28B68E38E2",
INIT_37 => X"FFFFFFFFFFFFFFFFFDFEF552E954AA0004000AA0000000000000000000000000",
INIT_38 => X"54AAF7D568A00557FFFFFFFFFFFDFEFF7FBFFFEF552E974AA082A820AAA2FFFF",
INIT_39 => X"FFF55A2D16AB550000175EFFFFBEAA00A2FFFFFFFF7FBFDFFFFFD568B55002A9",
INIT_3A => X"A800AAF7FBFDFEFF7D56AB45AAD56AB450004001EFFF842AAAA557FFDFEFF7FB",
INIT_3B => X"FFFFFFF552AA8BEF080402000087BFDF45AAD568B55AAFBFDFEF55042ABEF002",
INIT_3C => X"8516AB55A2D16ABEFFFFBFDFFF552AAAAAA007BC0000FFFBE8B55AAD168B55F7",
INIT_3D => X"00043DEAAFFAEAAAAA08556AB55A2D57FFFFF7D568B45002ABDEAAFFD16AA000",
INIT_3E => X"0000000000000000000000000000000000000FFD56AB45A2FFFDFFFAAD16AB45",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_4,               -- Port A enable input
WEA      => wbe_a_lo_1024_4(2),               -- Port A write enable input
DIA(0)   => data_write_a(19),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_4(19),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_4,               -- Port B enable input
WEB      => wbe_b_lo_1024_4(2),               -- Port B write enable input
DIB(0)   => data_write_b(19),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_4(19),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_20_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000003",
INIT_01 => X"F55FF80000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"E05022020800008400F655001FFCFF80018FA804400000000000004400000001",
INIT_03 => X"00000000000000000000000900002CC07000000000000000000000000000013F",
INIT_04 => X"68002FFE40900010000180000001FFEC0012EE0C001370F40780000000000000",
INIT_05 => X"0840000880FCBBF0100E204DF0F88311DD8005080679800000F3000029980580",
INIT_06 => X"001000030817C8E8840155FDF9001001050023F6C3C3D0F87FA19F7F011000E4",
INIT_07 => X"000000090492260800008000EE00000000000000002101FF2002C00000004018",
INIT_08 => X"2A040001071004000013FF7FCA302C0C0008214800002101554031F800000000",
INIT_09 => X"801F57F200000090000489FEC0000001EFBEF0040008023FDFC0000000004006",
INIT_0A => X"0000000008000000000000000000ADF000000200000008000008028300110230",
INIT_0B => X"0000000000000800080000000000000000000000000000000800800A40000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"000000040900005C848538000020000000800000080000020000800101FFB600",
INIT_0E => X"00800000003A010003000000000000600FFC53FF001800000002004080000000",
INIT_0F => X"0001000000007408040000004000000004E9000008020000200000000E800800",
INIT_10 => X"00200000000313100010002000008000000000129600040000400000001D0010",
INIT_11 => X"81C012060000000000218F7840000100800004000000000066C0000080080000",
INIT_12 => X"800000000017C000100000000001A800080000000001A8040000002840008185",
INIT_13 => X"0000000006F00000100200000000012600001004000000000066000000801040",
INIT_14 => X"0000200410100000000005F00000020080090A0000000085C800002000586000",
INIT_15 => X"FF00400000000000020020020001000040283024E4F2860400008000030ED080",
INIT_16 => X"00000000000000000000000000000004010201001003020200000000000127DB",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"A0700030038200010089120104D2040020000000000000000000000000000000",
INIT_1A => X"2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2C30C30C30C30C306982121A1E79E79",
INIT_1B => X"32190C86432190C86432190C86432190C86432190C86432190C86432190CB2CB",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000432190C86432190C864",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0201000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF552A974AA0004174BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA0804",
INIT_29 => X"7FFFFFFFFFFFFFFFFFFFFFFEF552E954AA000400000F7FFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E954BA007FC00BA087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974BA082E9540000",
INIT_2B => X"FFFFFFFFFF7FBFDFFF552E974BAA2FFFFE10FFFFFFFFFFFFFFFFFFFFFBFDFFF5",
INIT_2C => X"FAAD57FEAA007FFFFFFFFFFFFFEFF7FBFFF550800020BAAAD56AAAAF7FFFFFFF",
INIT_2D => X"EFF7D56AB450000021EFA2D57DE10087FFFFFFFFFFFFFEFF7FBEAB450804001E",
INIT_2E => X"000F7FFFFFFFFFFFFDFEFA2D568B550004001EFAAAEA8ABA5D7FFFFFFFFFFFDF",
INIT_2F => X"FFFF5D2E954AA080005000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFEF552A974AA0000104AAFFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"A954AA082A92428087FFFFFFFFFFFFFFFFFFBFDFEF5D2E974AA000A07000E3FF",
INIT_32 => X"FFFFFEFF7FBFFFFF552E974AA0071C50BA1C7FFFFFFFFFFFFFFFF7FBFDFFF5D2",
INIT_33 => X"EDF6FABAEBFFFFFFFFFFFFDFEFF7F5FAFC7492A974AAB6F5F8E10E3FFFFFFFFF",
INIT_34 => X"EBF5E8B550000071EFB6DF7AE921C7FFFFFFFFFBFDFEFE3F5F8F450004050AAB",
INIT_35 => X"A497FFFFFFF7FBF8FC7EBD168B450804021FFB6D57DE28147FFFFFFFFFBFDFC7",
INIT_36 => X"00000000000000000000FFFFFFFEFF7F1F8FD7AAD16AB450000001FFBEA4A8AA",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2A954AA0800174100000000000000000000000000",
INIT_38 => X"74AA002E95410A2FFFFFFFFFFFFFFFFFFFFFDFEF552E954AA0004000AAFFFFFF",
INIT_39 => X"FDFEFF7FBFFFEF552E974AA082A820AA087FFFFFFFFFFFFFEFF7FBFDFFF5D2A9",
INIT_3A => X"568A00AAFFFFFFFFFFBFDFEFFFFFFDFEF5D2E954AA0051554BA557FFFFFFFFFF",
INIT_3B => X"D16AB450804174AAFFFFFFEBAA2FFFFFFFF7FBFDFFFFFD568B55002A954AAF7D",
INIT_3C => X"57FFDFEFF7FBFFF55A2D16AB550000175EFFFFBEAA005D7FFFFEFF7FBFDFFFAA",
INIT_3D => X"0004001EFFF842AAAA087BFDFEFF7FFEAB45A2D568B550804001EFF7D57DEBA5",
INIT_3E => X"0000000000000000000000000000000000000F7FBFDFEFF7D56AB45AAD56AB45",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_4,               -- Port A enable input
WEA      => wbe_a_lo_1024_4(2),               -- Port A write enable input
DIA(0)   => data_write_a(20),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_4(20),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_4,               -- Port B enable input
WEB      => wbe_b_lo_1024_4(2),               -- Port B write enable input
DIB(0)   => data_write_b(20),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_4(20),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_21_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"4A302428B824900A128C090A5C1800261500213C005FE812D10420054085A202",
INIT_01 => X"001FFE3440B609703B0427F801A40B8115BC4F655300340288A40D30040E4DD8",
INIT_02 => X"E00424256888D8819801000F9FFFFFFFF149FF1FCA448046C60A0D2437C517F9",
INIT_03 => X"20030640003250640003250F06002CC1740002019824E001CD357832440001FF",
INIT_04 => X"EA2C3FFD400006E04401A8837001FFFC004AEF00080B70E08FB5789421007C5C",
INIT_05 => X"00011A0C40F9FFF80920954FF0F00809DF84A0202879800000F3000029980780",
INIT_06 => X"0805984B7A1FC0A0000101FFF0480080002281F7C3C381F87C03DFFF00009004",
INIT_07 => X"B424068086A205481A60A19000908204A855B000A08A61FF20C3D004D331D340",
INIT_08 => X"1BFA0001600802000023F7FFC08D234B40C2028253000040114200000D0226C0",
INIT_09 => X"EF1F5FF054096C6ADBA169FFC202B1C1FFBEF0440021083DFFCE22DC2880E24D",
INIT_0A => X"45FF0C004041D84862A28C54518DBFF00020004C0A6044901112A0908AA0A300",
INIT_0B => X"018C241102068006C620C03882019480E63180855A492712CC01C49C20201BFE",
INIT_0C => X"08A9464116544302C02D92236488D92236488D92236488D922366446C911B210",
INIT_0D => X"08800444021048034004001890000806002804A0822189000900D80621FFBE00",
INIT_0E => X"060580261013813A2CC396506102C4053FFD5BFF00A04A00200602CA52001100",
INIT_0F => X"080C0B004C202621A85C09411500135844C196D3606941018150098404C1A304",
INIT_10 => X"B02901013416181C96C2C9C600890A2028172192C460D1820302A0130809834A",
INIT_11 => X"9C5E803408250180AC268D185DB3F4350B811068C00049A0A4AA68F05C96A001",
INIT_12 => X"002C006560138F032B1804101244C883052208209040CC849063A747512B7678",
INIT_13 => X"41401E240665750440C9488280254530314080C2C601040420352148A00501B1",
INIT_14 => X"500811204D000700114204A70422016149916011008CAA8858850B00C32591C0",
INIT_15 => X"FFC06E60AC0496022300233104663040808E991765205000070121D41D18D098",
INIT_16 => X"40100401004010040100401004010040102090010008000001C0E010020007DF",
INIT_17 => X"0100401004010040100401004010040100401004010040100401004010040100",
INIT_18 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_19 => X"FFEF9FEEFF7FFDF7FF3E3DFDF7E0000000000000000000000000401004010040",
INIT_1A => X"BEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBFFDFDFFFCF3CF3F",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFEFF7FBFDFEFF7FBFDFEFBEF",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000FFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0001000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E954AA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0004",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA0004154BAFFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"52E974BA0804000AAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0004174BAFF",
INIT_2B => X"FFFFFFFFFFFFFFFFEF552E954AA000400000007FFFFFFFFFFFFFFFFFFFFFFEF5",
INIT_2C => X"A082E95400007FFFFFFFFFFFFFFFFFFFFDFEF5D2E974BA002E97400007FFFFFF",
INIT_2D => X"FFFFFBFDFEF5D2A954AA002E974BA087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFBFDFFF5D2E954BA007FC00BA5D7FFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA000002000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080005000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"A974AA0000104AAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974BA0000174AAFFFF",
INIT_32 => X"FFFFFFFFFFFFDFEF552E954BA080A000AAE3FFFFFFFFFFFFFFFFFFFFFFFEF552",
INIT_33 => X"02A95400087FFFFFFFFFFFFFFFFFFBFDFEF5D2E974AA000A07000007FFFFFFFF",
INIT_34 => X"F7FBFDFFF5D2A954AA082A924281C7FFFFFFFFFFFFFFFFFFBFDFEF5D2A974BA0",
INIT_35 => X"A557FFFFFFFFFFFFFFFF7FBFDFFF552E974BA0020924BA1C7FFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000E3FFFFFFFFFFFFFFEFF7FBFFFFF552E974AA0071C50B",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0000020000000000000000000000000000",
INIT_38 => X"74BA0000174BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954AA080017410FFFFFF",
INIT_39 => X"FFFFFFFFFFDFEF552E954AA0004000AAF7FFFFFFFFFFFFFFFFFFFFFFFEF552A9",
INIT_3A => X"E95410087FFFFFFFFFFFFFFFF7FBFDFEF5D2A954BA082E800AAA2FFFFFFFFFFF",
INIT_3B => X"FBFFFFF552E954BA002E97410087FFFFFFFFFFFFFEFF7FBFDFFF5D2A974AA002",
INIT_3C => X"57FFFFFFFFFFFDFEFF7FBFFFEF552E974AA082A820AA557FFFFFFFFFFFFFEFF7",
INIT_3D => X"5D2E954AA0051554BA5D7FFFFFFFFFBFDFEFF7FFFFFEF5D2A974BA0000020AA5",
INIT_3E => X"0000000000000000000000000000000000000AAFFFFFFFFFFBFDFEFFFFFFDFEF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_4,               -- Port A enable input
WEA      => wbe_a_lo_1024_4(2),               -- Port A write enable input
DIA(0)   => data_write_a(21),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_4(21),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_4,               -- Port B enable input
WEB      => wbe_b_lo_1024_4(2),               -- Port B write enable input
DIB(0)   => data_write_b(21),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_4(21),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_22_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"5290F4CDE914905A14A43D33F488243E17122300F55FEB189B343A1140548380",
INIT_01 => X"A54007B259F6A975386262000C344BA9573C6FF57B18A5FB0ABFCD3C2C5F4F0C",
INIT_02 => X"021DFF8C38B3C009D203551040030071869D0040180AA2DC53DB89BEA8204001",
INIT_03 => X"2603475A969D0475A969D0460EAA401005111011BD506954EDB40F5EF41434C0",
INIT_04 => X"922D9002100ED69E443D988B0D5400103E48003D0800011E803B06B5B9125A15",
INIT_05 => X"281B5A0C06000408F4DF9422010D8802022F2124A8022492580040440002021C",
INIT_06 => X"F780C4C052881ADA0E05440205DA50930FA182010004700083E220800440B588",
INIT_07 => X"049D028B93FB561833D8094A02F5EA92FD7247E10305C40040D136E6A023F7FC",
INIT_08 => X"00028241680A0E002A9400803A884B5B5206B7C2E53CA25144009007A64EBD64",
INIT_09 => X"41008810240240C6694008010392354010000560141801002028A83D2A08E06D",
INIT_0A => X"34000000848BCA6902A29C54539C020E11810098D4067EFF9FF284D483E2AB41",
INIT_0B => X"500001840000C80B410014088040F4A944B1AA313C0022AA0011C0DC00028001",
INIT_0C => X"80B14004D158C8CA24A1C2A870AA1C2A870AA1C2A870AA1C2A872550E1543800",
INIT_0D => X"80A14050A01509E050854498B5281A1C34E506A2C6898B52A154DAC6B6000850",
INIT_0E => X"0B03001A483A4146603050080410089180008800143D83888281A2034A850142",
INIT_0F => X"A4160600349075238473F1210006133835E92273612B3482C090068A0E84AC56",
INIT_10 => X"30060181BA1B13959DC08DA902458870201970B29602562B0581200D141D0959",
INIT_11 => X"E042021C040D0152C8058B3840F044708E7E1C20A0106EA166C13AFC14AA3804",
INIT_12 => X"080E004B0C17C1439A9838301DC1A8438EA32C009DC1A8255300650458A1D588",
INIT_13 => X"018010E186F110A908E3A8CB0026C9A610A908E6A60F0807626610E160589C4C",
INIT_14 => X"2A701667334005800B1605F043858125E0D04110408D2485CA034681E43A1E40",
INIT_15 => X"00646002304244A91102C93A2D608D2A258DF8034188200C050171A41108F084",
INIT_16 => X"110441104411044110441104411044110466C440446CA06951D4EA8010009804",
INIT_17 => X"0040100401004411044110441104411044110441104411044110441104411044",
INIT_18 => X"0401004010040100401004010040100401004010040100401004010040100401",
INIT_19 => X"F7DFBFDEFE8FF1F7DEBDDF7DF7D05122890000000003FFFFFFFF900401004010",
INIT_1A => X"9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7BFFDFD7DDDF7DF7D",
INIT_1B => X"F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE79E7",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000003F9FCFE7F3F9FCFE7F3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA000400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0800",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000002000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2A954BA000015400FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080402010FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2A954BA0004154BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A0004174BAFFFFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0800154AAFFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF552A974AA0000174BAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974A",
INIT_2E => X"000007FFFFFFFFFFFFFFFFFFFFFFEF552E974BA0804000AAA2FFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080400010000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E954AA080005000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000402010FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2A954BA000417410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"804154BAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974BA0000174AAFFFFFFFFFFF",
INIT_34 => X"FFFFFFFEF552A974AA0000104AAE3FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0",
INIT_35 => X"AA2FFFFFFFFFFFFFFFFFFFFFFFEF552E954BA000E124BAE3FFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000007FFFFFFFFFFFFFFFFFFFFDFEF552E954BA080A000A",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804000100000000000000000000000000",
INIT_38 => X"54AA000400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2A954AA080017410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"0174BAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A954BA000415400FFFFFFFFFFFFF",
INIT_3B => X"FFFDFEF552E974AA0804174AAF7FFFFFFFFFFFFFFFFFFFFFFFEF552A974BA000",
INIT_3C => X"2FFFFFFFFFFFFFFFFFFFFFDFEF552E954AA0004000AAA2FFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2A954BA082E800AAAAFFFFFFFFFFFFFFFFFFFBFDFEF5D2E954BA002A820BAA",
INIT_3E => X"0000000000000000000000000000000000000087FFFFFFFFFFFFFFFF7FBFDFEF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_4,               -- Port A enable input
WEA      => wbe_a_lo_1024_4(2),               -- Port A write enable input
DIA(0)   => data_write_a(22),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_4(22),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_4,               -- Port B enable input
WEB      => wbe_b_lo_1024_4(2),               -- Port B write enable input
DIB(0)   => data_write_b(22),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_4(22),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_23_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"EF20906D902424807BC8241BC81801B97D38AD3C0800103362A6741C80A12A02",
INIT_01 => X"001FFF8409F089003B4422000D80C80106804A7951C5B9D1C828043EA28838F9",
INIT_02 => X"E01CEE21649C82C40800000F9FFEFF8E72CA7F5FC2E22809925A0D3611C877F8",
INIT_03 => X"24000400402670400402670D48222DC1764446838624000080007460C40001BF",
INIT_04 => X"68403FFC020560E0443E21037C01FFFC0002EE00628BF0E02FAD781014085014",
INIT_05 => X"0112000202FBFFF00920017FF0F0628BFF8488890979800002F702002BB807A0",
INIT_06 => X"EF85788B681FC000000001FFF0010000000001F7CBC385F87C0BFFFF20040001",
INIT_07 => X"F6E200000000C1440E3AE408009120071070FA07A1CB23FFA403F0C4D23BF7C0",
INIT_08 => X"0BF87CA400804000003FF7FFD8880A034AC09662305AB10555421006891A1089",
INIT_09 => X"BE1F5FEA10092C0896A243FFC0008087FFBEF2000000001DFFC612C0C0400100",
INIT_0A => X"41FF0C2060501000600000000001BFFA800808189A657EF81DD0C00079CC8001",
INIT_0B => X"018C24110A860006C620C0312241C482B20400CC52492710CC80060020A81BFE",
INIT_0C => X"0C08866907048320C20C10030400C10030400C10030400C10030400608018210",
INIT_0D => X"040002000041500300100040000500C000801000C02400000952800001FFBF04",
INIT_0E => X"FC850015385380380CDB86106502C5043FFD5FFF00A04BC010A7724B10000800",
INIT_0F => X"89F90A002A70A710A51C01C05904014861433602A1CAF13F2110055614C72FC0",
INIT_10 => X"E02D02001C1E14981B43253EE50C8220180F1082E06397E07E42200AAC298E57",
INIT_11 => X"8421802400A90022B0070FAE18019214A380344920080B21A58B02AC60BACDF0",
INIT_12 => X"0A2A000C480B0704B54028101AC49C84BB4100009AC49C80857A82D20CE8CB22",
INIT_13 => X"01E00C8103416445C12ED0400027C5292445C12D500B0005A62D344CB241D095",
INIT_14 => X"132C907425604680038706A35132C94BDD011010404428886AC91B11311C8280",
INIT_15 => X"FF000470BE0692020328CA0028042054A92771C50FC070110001C1680809591D",
INIT_16 => X"00802008020080200802008020080200800800200200000000000008004807DF",
INIT_17 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_18 => X"8020080200802008020080200802008020080200802008020080200802008020",
INIT_19 => X"0000000000000000000000000000000000000000000000000000008020080200",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080002010FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974AA000400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000400010FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974AA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080000010FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E954AA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954A",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA000015400FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080002010FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974AA000400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000402010FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E954AA080005000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA080407000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA00041741",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080000010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000402010FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2A954AA080002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954AA080017410FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"552A954BA000415400F7FFFFFFFFFFFFFFFFFFFFFFFFF552A954BA080015410F",
INIT_3E => X"0000000000000000000000000000000000000F7FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_4,               -- Port A enable input
WEA      => wbe_a_lo_1024_4(2),               -- Port A write enable input
DIA(0)   => data_write_a(23),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_4(23),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_4,               -- Port B enable input
WEB      => wbe_b_lo_1024_4(2),               -- Port B write enable input
DIB(0)   => data_write_b(23),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_4(23),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_24_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100600007FFF000080108004000800020000840041000080808",
INIT_02 => X"FC5CA803400EB8209000000F9FFEFF8E7240FF1FC22409EA04018E50074017F0",
INIT_03 => X"11100400000000400000000D00002CC07400000090C080019001010A000001BF",
INIT_04 => X"68003FFC00040000000000008001FFFC0002EE00000370E007A100000000E468",
INIT_05 => X"0000000000F8BFF00920004DF0F00001DF8000000079800000F3000029980780",
INIT_06 => X"6E461803081FC000000001FFF0000000000001F7C3C380F87C019FFF00000000",
INIT_07 => X"600C2400013649609C8000980040814210254000A00B21FF2003F2A80D500000",
INIT_08 => X"0BF80000000000000003F7FFD88D2B4A02C0940062EC2804001610020408178B",
INIT_09 => X"8E1F5FE010092C0892A041FFC0000001FFBEF0000000001DFFC002C000000000",
INIT_0A => X"41FF0C0000000000600000000001BFFA0000005501AA00000CE2000009400000",
INIT_0B => X"018C0411020600048620C030020502000200000400490510CC00040020201BF4",
INIT_0C => X"0808064106040300C00C10030400C10030400C10030400C10030400608018210",
INIT_0D => X"0000000000004003000000000000001200580000000000000000000001FFBE00",
INIT_0E => X"0086C022005381380FDB96516140C6043FFD5BFF000041000000004110000000",
INIT_0F => X"80010D804400A7240C840C201D0210840043B4804012500021E0088014C04940",
INIT_10 => X"4109038041021C980200D06410C1924030008142E06024A00043C01100298092",
INIT_11 => X"587CC200002100C14428090A1D02348190814C09C010104025AA40041A0D8005",
INIT_12 => X"022E0030300B0E46177004208000D8C61D7004300000D884817B00011306B2D9",
INIT_13 => X"01E003060344710009875C018100013831000985DC000C20003C310006143B70",
INIT_14 => X"4001850EDC004780144806A64400186CBF8961104000C3807884000846EB9500",
INIT_15 => X"FF0006E08C063C0220002201490418082010A57263E0100008000290161E711C",
INIT_16 => X"00000000000000000000000000000000000000000000000000000000000007DF",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"F2D0AEEAF6E7CC1132CDB4441990000000000000000000000000000000000000",
INIT_1A => X"BEFBE79E79E79E79E79EFBEFBEFBEFBEFBEF9EF9EF9EF9EFA69861219575D75F",
INIT_1B => X"783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1EFBEF",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000783C1E0F0783C1E0F0",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0201000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A000400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA000400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000400000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402010000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"00002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080002010FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000400010FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA00040000",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020100000000000000000000000000",
INIT_38 => X"74BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"000010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA000002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974AA000402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000002010F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_4,               -- Port A enable input
WEA      => wbe_a_lo_1024_4(3),               -- Port A write enable input
DIA(0)   => data_write_a(24),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_4(24),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_4,               -- Port B enable input
WEB      => wbe_b_lo_1024_4(3),               -- Port B write enable input
DIB(0)   => data_write_b(24),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_4(24),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_25_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100200002000000080100004000000020000800041000080808",
INIT_02 => X"FC400086000000800000000F9FFEFF8E738FFF1FC204010000000111568DD7F8",
INIT_03 => X"00000400000000400000000D00002CC4740000008000000080000000000001BF",
INIT_04 => X"68003FFF64A564AC000000000001FFFE0082EF00010370E007A1000000004000",
INIT_05 => X"0A00040148F8BFF80920804DF0F00101DFC040000079C92484F30499299837C1",
INIT_06 => X"66041803081FC0E0801101FFFD000E41002299F7E3C380F87C019FFF81200096",
INIT_07 => X"000000080480AE00000080000000000000000000A00B21FF2003E00000000000",
INIT_08 => X"1BF80000400A02000003F7FFFA0008000200A0400008A0000014100200081000",
INIT_09 => X"8E1F5FFA53EFBCACB2E369FFE0010001FFBEF80C40630C7DFFEEBAF000800202",
INIT_0A => X"41FF0C0600000000600000000001BFFE00301000000000000CC020000140000C",
INIT_0B => X"01DCCC31222730A49620C030020100000200000400490D10EC00040220201BF4",
INIT_0C => X"0808064106240300C00C10030400C10030400C10030400C10030400608018210",
INIT_0D => X"0883044582114013412080000000000000000000000000000012800001FFBE00",
INIT_0E => X"00040020000180380FC386106140C6043FFD5BFF00A04B80608003CB120C1106",
INIT_0F => X"0000080040000200040400000100000000009480000240000100080000400900",
INIT_10 => X"0001000000000808000000240000020000000100006004800002001000008012",
INIT_11 => X"0001001808220000002004001900000080800008000000000022400000088000",
INIT_12 => X"0010000000000E00110000000000408009000000000040808063004000008200",
INIT_13 => X"6000000000046100000240000000001021000004400000000010210000001010",
INIT_14 => X"4000000404000800000000060400000088000001800000001084000000088000",
INIT_15 => X"FF800C608C041002000002000006100000002100000000180600000000100018",
INIT_16 => X"4110441104411044110441104411044510629041040D180400000010028047DF",
INIT_17 => X"1104411044110441104411044110441104411044110441104411044110441104",
INIT_18 => X"1044110441104411044110441104411044110441104411044110441104411044",
INIT_19 => X"FBA2894A196A8C5A2932EC15DA080800002FFFFFFFFFFFFFFFFFC11044110441",
INIT_1A => X"2492492492492492492410410410410410410492410492412000531215A69A6B",
INIT_1B => X"158AC562B158AC562B158AC562B158AC562B1588C46231188C46231188C49249",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000B158AC562B158AC562B",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080000010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000010FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08000000",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_4,               -- Port A enable input
WEA      => wbe_a_lo_1024_4(3),               -- Port A write enable input
DIA(0)   => data_write_a(25),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_4(25),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_4,               -- Port B enable input
WEB      => wbe_b_lo_1024_4(3),               -- Port B write enable input
DIB(0)   => data_write_b(25),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_4(25),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_26_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"E9264EAB20190CA3BA4997AA9002AE9C001006B0778015CFA17E0811039879C7",
INIT_01 => X"2FFFF9BB1F773C7F9BB07DFFFDD863FC5FFF3FEFFBBF9FFB22FFFBC7B9F30686",
INIT_02 => X"E06CCC62052E708180F6FFBFFFFCFFFFF9C7FF7FC24332E642090000074037F6",
INIT_03 => X"428003739CD9863739CD9869FE2B7DEAF300029E4E300DFE69A6E644E6FF473F",
INIT_04 => X"7C2FEFFFF5BA124F003DD31EAFFFFFEE9FF7EE6F4C0770FFD7DC7CA53997B2B1",
INIT_05 => X"DFFB5421C1F8BBFAFDBFFACDF0FFCC05DDDBFF3690F9EDB7F5F7AFF639BD7DE3",
INIT_06 => X"EFD044ABC817C3E3A74667FDFFB6FF5727CC3BFEF7C3FAF87FF59F7FFBFEF69F",
INIT_07 => X"00003002132462052E708180EF060C18E5BEFB051225CDFF7002C4EEDE77F6E0",
INIT_08 => X"3FFF7D5000EC75088ED3FF7FC8790E46426CE06CB1F8E041051831FA3068D77E",
INIT_09 => X"C05FD7FF9BEFBDCEFBEE59FEF44F6603EFBEFAFCC2E35E7FDFD147CCF3F583FA",
INIT_0A => X"67FF1C7FBFADEB31E35768E8ED6BFDF3EB3EBF9DDBCE7FDC1DF8A760F3EACC02",
INIT_0B => X"5BDDCC3B336F7C548667D47B7737AF3FD62601EDC25B3533DCEB07F262213FFC",
INIT_0C => X"5F9A06E19F4D93A0EA0F78C35E30D78C35E30D78C35E30D78C35E986BC61AE31",
INIT_0D => X"5FD7AFEFDFFAF59B6FF28FE1D80D73D840607307DCFE1D80EF69A004DFFFF7FF",
INIT_0E => X"0004001F8041897B2FFFC6D86D70CE04FFFFF3FF1F5F5475BD7F72E4D75EBFAF",
INIT_0F => X"F60008003F008237B0040A00010003E020023E0201F45EC0010007E01047D17B",
INIT_10 => X"00010001DC0004C81003DE050A700200001DC0006863E8BD8002000FC0208FA2",
INIT_11 => X"2200E400002801E1A00004C21C0206F60081800800007B00010F02007EC09A0E",
INIT_12 => X"0880007E000807C7C1A612001E0015C7C19C22001E0015C59DFE82011A311AA0",
INIT_13 => X"00001BC00101F60409F0670840070809760409F06984800780097604067D0010",
INIT_14 => X"81019F40042100001F800203D81019EC085614000085C80023D81009CF008A74",
INIT_15 => X"FF802FFDFFAFD082003B032FB987E04021D481D4000819060801E0D00001231D",
INIT_16 => X"EBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEFFBFBFBFBBFCFBB0FFDFEFFEF2DFFFFFB",
INIT_17 => X"BFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAF",
INIT_18 => X"FAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFE",
INIT_19 => X"475B15BCF491E166CC8553F86EDB5C88646FFFFFFFFFFFFFFFFFEBFAFEBFAFEB",
INIT_1A => X"861861861861861861861861861861861861869A69A61861AFBD54D5F871C71D",
INIT_1B => X"984C26130984C26130984C26130984C26130984C26130984C26130984C261861",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000984C26130984C26130",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040201",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_4,               -- Port A enable input
WEA      => wbe_a_lo_1024_4(3),               -- Port A write enable input
DIA(0)   => data_write_a(26),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_4(26),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_4,               -- Port B enable input
WEB      => wbe_b_lo_1024_4(3),               -- Port B write enable input
DIB(0)   => data_write_b(26),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_4(26),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_27_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"00080A40000A41248002029000050A088000008242A0004404480002000A1155",
INIT_01 => X"2FFFF1C11F781C129C107DFFFE0860941E81258CA2B71C2220EC1B86E1A00002",
INIT_02 => X"E1000000810000014400FF6FFFF0FFFFF8007F1FC21110005080200000221FF0",
INIT_03 => X"4080026318C18226318C1821302232EAE00002BE001115FE48620040840A863F",
INIT_04 => X"643D4FFC2530000F003D821C0BFFFF8E9EF79E6D440748FED70060842105B0B0",
INIT_05 => X"D6F39020D1F8A3FAFDBFBACDC8FDC405D1DB7F1490E5EDB7D5CBADB2385D79C3",
INIT_06 => X"6FE000A38007C3032646EFF1F0B6FF46A78C39F8E723F2E47FE59C7F9ADA2612",
INIT_07 => X"00002820000000810000014401060C180190310540118DFF1000C0849673F6C0",
INIT_08 => X"3FF779100062B12A8EC3F47FC80208808210880C00082050000110023068D030",
INIT_09 => X"005F07E09BFFBD07FBAC09F8E42922038F7DF8BEC2E39C5F1FD047CEF1B582D8",
INIT_0A => X"63FF5D5F9FADE911E81C09818109E1F16B16B71092CE7ED81CF403601228C402",
INIT_0B => X"1BFDCC39732F3554866AD57C37BEAF1C152201A4C05B7531D56B05B06A213FF8",
INIT_0C => X"5BCA06F18FC59380F00E34430D10C34430D10C34430D10C34430F0861A2186B5",
INIT_0D => X"5B56ADAB5FAAE58B2F628EA0C80FA3F04040510768EA0C80CC61A0044DFFC6EB",
INIT_0E => X"0004001D800188792CE79715710AE4047FFD23FF315D54358D593474955AB6AD",
INIT_0F => X"520008003B000297B0040200010003E020001F0201E44A400100076000579129",
INIT_10 => X"00010001DC00004A10035E0408300200001DC000086BC8948002000EC000AF22",
INIT_11 => X"02002400002801E1A00000C01E0202F60080800800007B00000782006EC0820A",
INIT_12 => X"0080007E000006A7C10602001E0001A7C10C02001E0001C18DE282010A311AA0",
INIT_13 => X"00001BC00000FE0401F04300400708007E0401F04180800780007E04047D0010",
INIT_14 => X"81011F40040100001F800002F81011EC080604000085C80001F810094F008034",
INIT_15 => X"FF800C6DDDAFD082001B03249887E04001D481D4000009020801E0D00001021F",
INIT_16 => X"AB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6BF1EBDABD8E270BF84A25C6ACB777E3",
INIT_17 => X"B6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6AD",
INIT_18 => X"6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADA",
INIT_19 => X"490E2168100481CA860402104A471688747FFFFFFFFFFFFFFFFFAB6ADAB6ADAB",
INIT_1A => X"000000000000000000000000000000000008200000000000200072F210000001",
INIT_1B => X"05028140A05028140A05028140A05028140A0500804020100804020100800000",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000A05028140A05028140A",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040201",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_4,               -- Port A enable input
WEA      => wbe_a_lo_1024_4(3),               -- Port A write enable input
DIA(0)   => data_write_a(27),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_4(27),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_4,               -- Port B enable input
WEB      => wbe_b_lo_1024_4(3),               -- Port B write enable input
DIB(0)   => data_write_b(27),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_4(27),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_28_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"02200AA400180030808802A900002A08001280A08A801044104A1000001818C3",
INIT_01 => X"0AA00011460214428114180000882214413D0A71592A01D92213D28005210202",
INIT_02 => X"0451110A012100884000AA30200000000C100040104112101100008888200000",
INIT_03 => X"448000318C52A20318C52A20148810200111100C211004AA00034204200A2200",
INIT_04 => X"04004001001A90110000121402AA0000003C00000500000040080421080D0080",
INIT_05 => X"4060000C8001000000002E000000050000001610300000010000802202040012",
INIT_06 => X"1000002080001111001222000425A1040026A008000000000000000009328280",
INIT_07 => X"2491008A00491201210088400122448908A20402000408001000040820000000",
INIT_08 => X"20058310402A160026500000028040101004200C840082115554000112244814",
INIT_09 => X"4140000800000060000720000102028000000490160801020002200011100010",
INIT_0A => X"020000081B34211082B694D4D294000020020381040000000200032040004400",
INIT_0B => X"4800210C19808400500010009110091500020B408810000100200020408B0000",
INIT_0C => X"01028000080118020023604858121604858121604858121604858090B0242C00",
INIT_0D => X"010000800920040804020A6058003108402043058C460580653020005A004039",
INIT_0E => X"00000002800008014004104104420A00C000200005000010040A0020CC000200",
INIT_0F => X"520000000500000010000200000000000000280000040A40000000A000001029",
INIT_10 => X"00000000000000C0000002000830000000000000480008148000000140000020",
INIT_11 => X"020024000000000000000440000000020000800000000000000C00000040020A",
INIT_12 => X"00800000000001804006020000000500400C0200000005400A90000000100000",
INIT_13 => X"0000000000018200001003004000000142000010018080000001420000200000",
INIT_14 => X"8000080000010000000000018800008000060400000000000310000008000034",
INIT_15 => X"000002040080000000110006B081400000400000000009020000000000002200",
INIT_16 => X"802008020080200802008020080200802101210810C39A66A90A85420413A820",
INIT_17 => X"0200802008020080200802008020080200802008020080200802008020080200",
INIT_18 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_19 => X"DE21102C110A00246972BD89A40A0C22E1000000000000000000002008020080",
INIT_1A => X"2082082082082082082082082082082082082082082082080D35050758C30C31",
INIT_1B => X"0582C160B0582C160B0582C160B0582C160B0580C06030180C06030180C08208",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000B0582C160B0582C160B",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_4,               -- Port A enable input
WEA      => wbe_a_lo_1024_4(3),               -- Port A write enable input
DIA(0)   => data_write_a(28),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_4(28),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_4,               -- Port B enable input
WEB      => wbe_b_lo_1024_4(3),               -- Port B write enable input
DIB(0)   => data_write_b(28),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_4(28),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_29_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"79964E4BA01DACAB9E659792D00AAE160002829C7FDFEFCEE97C2815039D70C3",
INIT_01 => X"0ABFF9AB0775343F9AB01DF80D5821FC0FFF3FEFD1AF9FF1207FFBC7B9720586",
INIT_02 => X"002CCC60050E700080F6AAA7BFFC007189C7FF2FC00330E602800000074037F6",
INIT_03 => X"468003210868A63210868A68DA017D207200021C4E200CAA6186A40042FF4300",
INIT_04 => X"7C2FE002F0900001003C5316A6ABFFE21F36E02F0D03701F47D41800109FB281",
INIT_05 => X"4979440580F9B808F49F6A4DF00F8D01DC4B97369078249370F482E62BA41462",
INIT_06 => X"B250442BC81001E1870223FC0BF7F11507C423FE33C078F803F19F00E936721D",
INIT_07 => X"00011080012460050E700080EF020408EC8CFA01122149FF700200665A35D260",
INIT_08 => X"2BFD055040A452000443FF00007906464068406C31F84000000831FA1028575A",
INIT_09 => X"805FD017102690AA694551FE30444681E0820AD40201423FC00122C493500172",
INIT_0A => X"0600002AFFBE2330815568A8AD6ABC02A02A0B0CCB463B4C0748A720B1EA4C00",
INIT_0B => X"0850400A11414C005005000B51158936D20601A98A10200308A002E240010BFC",
INIT_0C => X"05928020194918A22A2268C81A32068C81A32068C81A32068C81A99034640C00",
INIT_0D => X"058102C48970541944B20FA1580561D040406305587A158046282000DBFFF13D",
INIT_0E => X"000000028040890327DCD28928324400DFFFF0001F1F0050342D42A086040B02",
INIT_0F => X"F60000000500802010000A000000000000022A0000141EC0000000A01000507B",
INIT_10 => X"00000000000004C0000082010A700000000000006800283D80000001402000A0",
INIT_11 => X"2200E4000000000000000442040004020001800000000000010D000010401A0E",
INIT_12 => X"08800000000801C040A6120000001540409C2200000015441DAC800010100000",
INIT_13 => X"0000000001019600081027084000000956000810298480000009560002200000",
INIT_14 => X"800088000021000000000201D800088000561400000000002358000088000A74",
INIT_15 => X"00802594A282C0000033010FB181E00020400000000819060000000000002305",
INIT_16 => X"C0B02C0B02C0B02C0B02C0B02C0B02C4B12B312912831A27FCFE7FFB175B6FF8",
INIT_17 => X"0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02",
INIT_18 => X"B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C",
INIT_19 => X"BBCF9F96EE7FFDF7FE783FFDFFEA0C00602FFFFFFFFFFFFFFFFFC0B02C0B02C0",
INIT_1A => X"EFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEEBAEBAEBAEBAEBBFFDF9FBEFFFFFFE",
INIT_1B => X"BFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFBEFB",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000FBFDFEFF7FBFDFEFF7F",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_4,               -- Port A enable input
WEA      => wbe_a_lo_1024_4(3),               -- Port A write enable input
DIA(0)   => data_write_a(29),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_4(29),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_4,               -- Port B enable input
WEB      => wbe_b_lo_1024_4(3),               -- Port B write enable input
DIB(0)   => data_write_b(29),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_4(29),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_30_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"F7FFBFFEFF9FE1F7FFBFFFFDFFD0000000000000000000000000000000000000",
INIT_1A => X"9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7AFBD75F5FDF7DF7F",
INIT_1B => X"F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE79E7",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000003F9FCFE7F3F9FCFE7F3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_4,               -- Port A enable input
WEA      => wbe_a_lo_1024_4(3),               -- Port A write enable input
DIA(0)   => data_write_a(30),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_4(30),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_4,               -- Port B enable input
WEB      => wbe_b_lo_1024_4(3),               -- Port B write enable input
DIB(0)   => data_write_b(30),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_4(30),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_31_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"129000008004A00804A40000400800020000000C005FEA005800200400050100",
INIT_01 => X"255FF18019700810180065FFFC0040801E80258CA2951C2200EC0906A0804140",
INIT_02 => X"E0000000000000011000550FDFF0FFFFF0007F1FC200000044000000000817F0",
INIT_03 => X"0000024210A30024210A3001002220C06044469200040154482000408400043F",
INIT_04 => X"602D0FFC2420000E003D80080955FF8E1ECA8E2D400340FE870060842100B030",
INIT_05 => X"0213100040F8A3F8FDBF944DC0FDC001D1CB6904A061EDB6D4C30490281831C1",
INIT_06 => X"6FC000830007C202060445F1F0D25E4207A099F0E303F0E07FE19C7F80402412",
INIT_07 => X"0000200000000000000001100004081001103107000185FF0000C0849673F6C0",
INIT_08 => X"1BF27A00000000000883F47FC800080002008000000820440000100220489020",
INIT_09 => X"011F07E013EFBC06FBA009F8E00120038F3CF82C44630C5D1FC002CCE0808248",
INIT_0A => X"61FF0C06C48BC801600000000001A1F00110101092CE7ED81CF0004012288000",
INIT_0B => X"11DCCC31222730048620C4382204A608142002A440492530C401049020221BF8",
INIT_0C => X"0888066187448380E00C10030400C10030400C10030400C10030600608018210",
INIT_0D => X"080204010200418301208480800D02D00040100240A808008840800405FF8640",
INIT_0E => X"0004001D000180780CE386106100C4043FFD03FF101D40008001304018081004",
INIT_0F => X"000008003A000217A0040000010003E02000160201E040000100074000478100",
INIT_10 => X"00010001DC00000810035C0400000200001DC0000063C0800002000E80008F02",
INIT_11 => X"00000000002801E1A00000801C0202F40080000800007B00000302006E808000",
INIT_12 => X"0000007E00000607810000001E000087810000001E000081846282010A211AA0",
INIT_13 => X"00001BC00000740401E0400000070800340401E04000000780003404045D0010",
INIT_14 => X"01011740040000001F8000025010116C080000000085C80000C8100947008000",
INIT_15 => X"FF800C609C06D082000A03200806A040019481D4000000000801E0D00001001D",
INIT_16 => X"010040100401004010040100401004010060C040040C200950402090128057C3",
INIT_17 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_18 => X"0040100401004010040100401004010040100401004010040100401004010040",
INIT_19 => X"00000000000000000000000000001000802FFFFFFFFFFFFFFFFF810040100401",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_1024_4,               -- Port A enable input
WEA      => wbe_a_lo_1024_4(3),               -- Port A write enable input
DIA(0)   => data_write_a(31),        -- Port A data input
DOA(0)   => data_read_a_lo_1024_4(31),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_1024_4,               -- Port B enable input
WEB      => wbe_b_lo_1024_4(3),               -- Port B write enable input
DIB(0)   => data_write_b(31),        -- Port B data input
DOB(0)   => data_read_b_lo_1024_4(31),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_0_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"ED39BA795990D275FB4A6E96ACC4731DEA4598B0AFB54867F6EE4618C3749803",
INIT_01 => X"8AA0047D8607944AC7DA180001ECA2444042106208408208C20022E9173734B3",
INIT_02 => X"1A7DDD79F9A73E6CCA7DAAF00001000008478020113D98E382FEDF333027C80F",
INIT_03 => X"75D341110C58F31110C58F32A208921F8051500147A0E4AB3493FB3A01EBE240",
INIT_04 => X"86424001531009B100425A97B2AA0001E03501D0A39C8F0078420001106D0C4C",
INIT_05 => X"BCC8CA2EBF03400700402BB20F00239E20341699198600000B08694B16434804",
INIT_06 => X"103FB860B2800161F8432200012DA185F80F24081C3C0707800E600056881308",
INIT_07 => X"B24197ABCDA467F9A73E6CCAFDC3870EEEEC44E2BDFE220094D03022210C011C",
INIT_08 => X"240581B5695EAA80262C080032BF07C7C1FC3F8E94F65B11555EAFFC1C306758",
INIT_09 => X"7E40000BEC004170040DB60017FED1CC0001045002984202003DB931192D60A5",
INIT_0A => X"120071411A74315881A28C141118000C5A85A60444210123820B43B40804674D",
INIT_0B => X"0820008E514045BB514F0106D1D8599581D3A958BC104A89215AC14C48898403",
INIT_0C => X"C261C01C48B1584A0CA3E2687A9A1E2687A9A1E2687A9A1E26870CD061343885",
INIT_0D => X"D274E93A758FA8683AC54B287522E10A74AF4AA59C568752662F5AC218000002",
INIT_0E => X"FF83C002783A0904231C70470C7E0B92800224008AE09FAD4BD48D1FC5D3A4E9",
INIT_0F => X"5BFF078004F075885DFBF7E15C06101C55E921F1F80FAB7FE0F0009E0E903EAD",
INIT_10 => X"F12E0380231F13978FF023FAFDBD9870380230F2D6081F56FFC1E0013C1D207D",
INIT_11 => X"DE7F263C0C8700125C0F8F3C43F1F10BBF7EFC61E01804E1E6C8F8FE807F67FB",
INIT_12 => X"02BE00017C17C1007E5E2E3081C5AC007E6F0E3081C5AC44418D65FE45DEE55B",
INIT_13 => X"61E0042786F103E9F01F9BC3C120C5A703E9F01F978B8C20666703E9F8A0FFED",
INIT_14 => X"FA7E283FFB414F80005F05F10FA7E283F78F6511C048278DCA174FF038FF15B4",
INIT_15 => X"0066A20B61692F293185D8D724E15D3FCC6B7C236FE0691B0700132C1F0EF880",
INIT_16 => X"3A4E93A4E93A4E93A4E93A4E93A4E93A4F942F92E9628540AD2A91442525A000",
INIT_17 => X"A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E9",
INIT_18 => X"4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93",
INIT_19 => X"55F3898E09B56C74DAB15D1CF13501AA495000000000000000003A4E93A4E93A",
INIT_1A => X"082082082082082082082082082082082082082082082082082084E41DC71C71",
INIT_1B => X"E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F82082",
INIT_1C => X"FFFFFFFFFFFFFFF94A5294A5294A5294A5294A52800003E1F0F87C3E1F0F87C3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"3060C183060C187FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"BDEBA0000000000000000000000000000000000000000000003060C183060C18",
INIT_28 => X"168ABA002E82145085155545F7AA975EFFFAABDE00FFAEBDFFF5D2EAAAAAF7AE",
INIT_29 => X"7FFFE10005542145557FD5545FF8000155087FC0155F7D168B55007BFDF45085",
INIT_2A => X"7FFC0010080017555555568AAAFFFFD7545AA8028A00A2802AABAFF8028BEF5D",
INIT_2B => X"FF842AABAA2AE95545FFD168ABAF7AEAAAAAA2FFFDF4500043FE105D2E954BAF",
INIT_2C => X"5007FD7400550415410002E974BA5D5168A00A2D142155005142010FFAE820AA",
INIT_2D => X"FFF780000BA007FE8AAAFF803FFFF5D2A821550000000BA007FD55FF5D7FC014",
INIT_2E => X"000AAFBEAA00007BFDFFF082EBDF455D5142000082E82145FFD17DFEFFFD168B",
INIT_2F => X"DFD75D2AA8A80EA8E2FE3F000000000000000000000000000000000000000000",
INIT_30 => X"68B551475FAF6D1C556F0AA1C24AABEA495FC716F002A975FFE3AA95E00EBAEB",
INIT_31 => X"42A0070071C50BAFEF1FAE0016D56A16D557BC257D415E0216FA3F1E8FC0145B",
INIT_32 => X"8010E004924874825D7FEAA85487FD24AFE3D02DAAAE12BD5545A2803AA00005",
INIT_33 => X"120155EA568E870BAEB8A05A2AEA8B50F55A2F150005A3A438BD04AFAB8F550A",
INIT_34 => X"545E055FFBE81D0BE8EA8A3AA05A2A5504001C74BA42A1571E8028E3DB7816D0",
INIT_35 => X"A5C7E3DFFFE90B45B47ABA497A82FFAFD2A82485FD2415A105C21451ED42A002",
INIT_36 => X"00000000000000000000B55EAAA100AA1D0F6F480B6A555A2A57A002A3D5FDB6",
INIT_37 => X"5EFAAAAB5E1AF3AABFF45592E88A0AFE80A8B0A0000000000000000000000000",
INIT_38 => X"65F520EBE9EF67D7BEA1FD5D556ABEF5D557FEBA55022A3F70C6B405F4D2AE97",
INIT_39 => X"C114728007521170821CE0FDE69411A8DED57CE1055555E5F58EFFC01FE2CACB",
INIT_3A => X"42341D5DEEBEF55080034E0A592A4AD0079C75D6070CC5CBB0280C029ABAA3EB",
INIT_3B => X"7F353AAF6C77F7F20D968BF57812A95E02A2AAB5EB0F280800EFAEE9F5D18F31",
INIT_3C => X"C91565455C141E41887D58AC448B69C30E02116220415A9540AA854140A0A204",
INIT_3D => X"DE6BE93172D7D625B556EEAB157ABEBE1B4D792A4AD1183454180DD3FDCAAAB7",
INIT_3E => X"F0000001FF0000001FF0000001FF0000001FF01EABC4B8014174FF7DA80F52FE",
INIT_3F => X"FF0000001FF0000001FF0000001FF0000001FF0000001FF0000001FF0000001F")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_4,               -- Port A enable input
WEA      => wbe_a_hi_1024_4(0),               -- Port A write enable input
DIA(0)   => data_write_a(0),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_4(0),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_4,               -- Port B enable input
WEB      => wbe_b_hi_1024_4(0),               -- Port B write enable input
DIB(0)   => data_write_b(0),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_4(0),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_1_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"212C001411984004084D000508C53810A03D1450E839B003342114428A000803",
INIT_01 => X"00000019400B100A8196000000CC004400400002000000000000028001340000",
INIT_02 => X"052137AE8031800C0044009000000000061800001CD4019802AD04CCCFC20004",
INIT_03 => X"04514108C60C21008C6042108400000201440020505100000043C30E10E9F000",
INIT_04 => X"02104001011DEFE088805681920000008000004001900800004002108C280008",
INIT_05 => X"040002340105000200000000080001900010000108040000000008411600401C",
INIT_06 => X"1034001042800808201000000001000820020000102000040000000000800180",
INIT_07 => X"64BF81A15EDFDE8031800C00843060C19E030022103600000450020800040004",
INIT_08 => X"00008004691687AA840008000090248CC84E000046000311555521F183060AC5",
INIT_09 => X"0820800D08100171000DB000154440C800400500000852020011200201012021",
INIT_0A => X"02000040001000880A2A04445004000102002041000001008208001440004140",
INIT_0B => X"4820018A1140440078050040511000102000A008183000010002404400000000",
INIT_0C => X"1000C80008000C030030880C2A030A00C28030A80C2A030A00C28018D4061401",
INIT_0D => X"10040802050080200284401C0022880F009E08008205C0020118088018000000",
INIT_0E => X"0F03C00280000000420860C60C0C0B92C0000000004000010042000040102008",
INIT_0F => X"001E078005000108400005E11C0610000000288058000003C0F000A000100000",
INIT_10 => X"F10E0380000000C202300000008D187038000000480800000781E00140002000",
INIT_11 => X"806302380C870010000004400100110800007861E0180000000C400680000001",
INIT_12 => X"023E00000000018000580C308000050000610C30800005000215006800000101",
INIT_13 => X"61E0000000018100B0001843812000014100B00016030C20000141002880026D",
INIT_14 => X"400A20009B404F80000000018400A20044096111C04000000304026000501580",
INIT_15 => X"0046820040082300218450C2800010094000482141E060190700100000002200",
INIT_16 => X"020080200802008020080200802008020080008008600500A82A1100A8000000",
INIT_17 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_18 => X"0080200802008020080200802008020080200802008020080200802008020080",
INIT_19 => X"81328A46BABEFC54A0810C7452B4428A14000000000000000000020080200802",
INIT_1A => X"AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA28A28A28A28A2A8218D2C0C924925",
INIT_1B => X"E974BA5D2E974BA5D2E974BA5D2E974BA5D2E975BADD6EB75BADD6EB75BAAAAA",
INIT_1C => X"FFFFFFFFFFFFFFFD8C6318C6318C6318C6318C63000002E974BA5D2E974BA5D2",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"70E1C3870E1C387FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"5555500000000000000000000000000000000000000000000070E1C3870E1C38",
INIT_28 => X"EBDF455D2EAABEFF7FFE8BFF5D0002155557FFFFFF007FC21EFA2FFD74AAAAD5",
INIT_29 => X"AA95400552AAAABAFFD1574105D7FD75FFAAAA800AAF7AA974BAFFFBE8B45F7A",
INIT_2A => X"0517DF555D2EAAA1055000015500557DF45AAD1400BAA2AE801550051555EFF7",
INIT_2B => X"FFD540155557FD5400F78028BFFFFFBEAB55F780020AAAA80020AA082EAAB550",
INIT_2C => X"AFF842ABEF5D517DF55552A974AAF7AE820AA0851574BAA2D1574AA5D7BFDEBA",
INIT_2D => X"EFAAD1575EF557FFFE10557FFFFFFFFD56AAAAFFFFD7555AAD168B45AAAEAAAB",
INIT_2E => X"0005D7FFDF4500043FE105D2E954BAF7AE80010082A97410557FEABFFAAFBE8B",
INIT_2F => X"51C7A2FBD5490BFD1C056A000000000000000000000000000000000000000000",
INIT_30 => X"974BAF7FFEFB45FFAABDF55492AA8BC2EBDFEAF7F1F840017D4975D2FEF147FC",
INIT_31 => X"080BEF495FC71D54124924385FAAA8AAAE3D145410F7F1D55D71C002DABAEBAA",
INIT_32 => X"002D082082AB8B6DBEDB7DF7F540E2AE85028B40155145F7AF6DBED5450AA1C2",
INIT_33 => X"78E021FF1471FDEAAFFD56F16D5571D2E28E38E0216FA2D1E8E80140F45082B4",
INIT_34 => X"A2DA3FB7DAAD4AAAAF487BC70BFA97F7AF6D417E92482BF84020BA495557E3FF",
INIT_35 => X"55554ADBD7A2FFC7BEFF6FFD7FC7002FD74951D71EDFFABFD16FAAAE92BD5545",
INIT_36 => X"00000000000000000000547AB8F550A8010E00492487482FFFE82A85EBAE2FFC",
INIT_37 => X"1EF005162BEF047FD5545AAFBF7400FBF9424F70000000000000000000000000",
INIT_38 => X"714F8338AAAA1D0AE974AAF7FFFDF55F7AABFF55082CA8B4DF6C1E8F5E540002",
INIT_39 => X"EABEF75550ACBB7582225FF5843404547184164AA5D2EBEEB0A2D555410D3555",
INIT_3A => X"FEAAEB083BC1000FF8409000512AEABFFDF79DCBF755962010BDCBBC21455D7F",
INIT_3B => X"801F8BA0C57740BDAA0688E5405D57D412F7D55F5E50C7F401BAAE8403CF5A3F",
INIT_3C => X"5D16BABAA3EBC3157ABD5FFE55F2AA9FEAFDF7F431A9F7FFE81FF013A8001AFF",
INIT_3D => X"FB863550229BCABEB7DA403FFFDA2FBF7FED2C7F955445079E280A00C56145EF",
INIT_3E => X"0000000000000000000000000000000000000596EBEF55080034E0A592A4AD00",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_4,               -- Port A enable input
WEA      => wbe_a_hi_1024_4(0),               -- Port A write enable input
DIA(0)   => data_write_a(1),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_4(1),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_4,               -- Port B enable input
WEB      => wbe_b_hi_1024_4(0),               -- Port B write enable input
DIB(0)   => data_write_b(1),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_4(1),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_2_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10E006600180111284380310006289800480032283E000A34301002001A0817",
INIT_01 => X"0005A00810790848048044A54E404350404000720885800802000906E4910200",
INIT_02 => X"407004208400408044C600C50AA055254010541A110222841200000002402544",
INIT_03 => X"0600011004182401004102408C28414043101000408118000145840440F5C415",
INIT_04 => X"5035855703A2900A000CD3088400F40688C9844409060850925E58A4081A0221",
INIT_05 => X"0200840D1021A15AC50494894850890540D1E12020C6E510818500440A280090",
INIT_06 => X"113044094002801020440090A8011A1224AB9380552102442884882A20004097",
INIT_07 => X"000100880004428400408044860000008C022402102100AA40004404B5075460",
INIT_08 => X"15C23440408C862A2A12382A8A5244145048C06085008010141521F000001240",
INIT_09 => X"400582B9033AA0E7AA4110B0506744810554542450694E710A836188C2C00222",
INIT_0A => X"443518360012C2210B020414109130A28038188096A06B8C120CA440A9C00802",
INIT_0B => X"1345E53300EC68005605002964AF222A5704004D080211121C80024200821780",
INIT_0C => X"181080C1110C882202211488452213C88472213C88472213488441109A442231",
INIT_0D => X"008204440210091341208041000810C00000300220201800A908000038AD0284",
INIT_0E => X"00040002804180300E88D28D206A40000554815500481440300000C44A081100",
INIT_0F => X"000008000500828700000000010000000002380000A00000010000A010050000",
INIT_10 => X"00010000000004CA000214000000020000000000684280000002000140200500",
INIT_11 => X"000000000020000000000442100002840000000800000000010C000026000000",
INIT_12 => X"00000000000805A4800000000000152300000000000015801272000100210020",
INIT_13 => X"000000000101C00000C000000000000940000120000000000009600004050000",
INIT_14 => X"0000130000000000000002018000106000000000000000002380000141000000",
INIT_15 => X"55000190000000000002000280000000011080C0000000000000000000002310",
INIT_16 => X"40902409064190641906419024090244902A9003004800415120D4A190804241",
INIT_17 => X"0900409004090641906419064190240902409024090641906419064190240902",
INIT_18 => X"9044090040900409004190441904419044090040900409004190441904419044",
INIT_19 => X"75960040138D70C030B51C50C7D100A2052F81F81F83F03F03F0419044190441",
INIT_1A => X"0410410410410410410410410410410410410410410410410248602081659659",
INIT_1B => X"5128944A25128944A25128944A25128944A25128944A25128944A25128941041",
INIT_1C => X"FFFFFFFFFFFFFFFE1084210842108421084210843FFF825128944A25128944A2",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"7FD5FF555815607FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"2AA000000000000000000000000000000000000000000000007FD5FF55581560",
INIT_28 => X"FC21EFA2FFD75EFAA8415410AA8415555087BFFF55A2AA800BAFFAE954000800",
INIT_29 => X"84155EFA2AEBDEAAA2FBEAABA5D7FE8B555551421455D0002145552EBFEBA007",
INIT_2A => X"2AEBDF555D2E954BAA2AA974BAFFFFE8B45552EBDF45FFAEAABFFF7FFE8B55F7",
INIT_2B => X"AAAAAAAAAFFD1574105D7FFFF555D2AAAAAA5D2E820BAA2FBEAB5555557DF55A",
INIT_2C => X"50055575EFFF84021555D043DEAA5D04021EF557FC21FFAA8428BFFAAAA954AA",
INIT_2D => X"10085568A00FF80175FFA2D17DFEFF7800215500557DF55AA80001FFAA800015",
INIT_2E => X"0005D00020AAAA80020AA082EAAB5500517DF555D042AA10A284154005D00154",
INIT_2F => X"00AAFFAA9543A080038A2A000000000000000000000000000000000000000000",
INIT_30 => X"0017D5D20B8EAA007FC51C7A2FBD55D2BE800042AFE8E1557D0075D2F45BEAA8",
INIT_31 => X"AA8BC7EBDFEAFEFFD00105FFBC20BDEAAA2FBF8AAA557BE8B6D5D5FFABEF4904",
INIT_32 => X"FFEFB6D555578F7DB6A0BDF7D480E174BFA02A974BAF7F5EFB455D2ABDF55492",
INIT_33 => X"ED1FDE90E3A497492B6AAADAAAE3D155E105571D55D71C002DABA5524820BAB6",
INIT_34 => X"BE8F401D7B6A0001470155C51D0092A071555D5E3AE821D00001FF0871C016DB",
INIT_35 => X"5BE8555400550A38428007FED000E3DA3DFD5E3DFFFBD5A38A021551C5F7AF6D",
INIT_36 => X"00000000000000000000410F45082B4002D082082AB8B6D1C5B7DF7FF78E075C",
INIT_37 => X"5EF005560B55F7AA800AAF7AA954AA00042AAA20000000000000000000000000",
INIT_38 => X"ABEF057D68F5F5A00021EF55042AAAA007FD5555AAFBD7545FBB8020A3F7AE97",
INIT_39 => X"7DF55D7AABFF5428ACA8F45A6C1E8F5EFF84165EFF7802BAB0A2FFEAABA557BE",
INIT_3A => X"CA8AA80800020AAF7FBFFFEF04552ABFFFF841FFE75CA882108202E974AAF7D5",
INIT_3B => X"00151FF0C57401E5F3D1E00A1A884174A8FFAEBFEB0A2D55541051555694F002",
INIT_3C => X"2AA801455D7FE8BFFF680800FFF7AAA155F595542455512A975455D3AA8A0055",
INIT_3D => X"5D79FCAF774AE005BE7895554005D2A8A0B882FFFFE10AAAAAB755A66B6AF56A",
INIT_3E => X"00000000000000000000000000000000000000C3BC1000FF8409000512AEABFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_4,               -- Port A enable input
WEA      => wbe_a_hi_1024_4(0),               -- Port A write enable input
DIA(0)   => data_write_a(2),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_4(2),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_4,               -- Port B enable input
WEB      => wbe_b_hi_1024_4(0),               -- Port B write enable input
DIB(0)   => data_write_b(2),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_4(2),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_3_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"210C00A20020000108430020001600B8156021104940741B3530400E02B92203",
INIT_01 => X"014C9BCA58B1296D24A402C992500B69404040028804A0080A000416A8D90A08",
INIT_02 => X"C12026A484318004404405C9C66E331352180D468B8203980300204442E02B34",
INIT_03 => X"04000748D60D24648D60524C88804D0215011020D15018148040C10A70E1D58C",
INIT_04 => X"18283333240FE41244187308C9104D70944852640901083801750EB0A418C220",
INIT_05 => X"0613142D01912CC2A1B4140528348900C612A104201C689044340ED413A07649",
INIT_06 => X"119000034019881822104C5E68035250A222829710A0A02C18C01A9920842413",
INIT_07 => X"402F00AB0016CA0431800444841020509D038B021230C1990001C644C8273200",
INIT_08 => X"16905000408482088290E8E64010248C4A5AA840C2000110001521F0810A92E7",
INIT_09 => X"0003CE6581BD016342A951AB146C4480530C3B2A8088D3542651670200C1826A",
INIT_0A => X"00735D36209A8A20020894004284B660821030C8990467401218004041020002",
INIT_0B => X"512445B740457154562F957CC08B00093700080D0A4851001D8302D20A0A1530",
INIT_0C => X"00508650008008021021A40861021840869021A408610218C0869810D6043095",
INIT_0D => X"1C8508438450801043A08090380A8834207007022209038080190000999C8F84",
INIT_0E => X"000400200000C0002A48A206204C4205F3304B33004C0041006240140A1C310A",
INIT_0F => X"0000080040000083800400000100000000008400018040000100080000510100",
INIT_10 => X"0001000000000800000244040000020000000100002A0080000200100000A702",
INIT_11 => X"000000000020000000200000080002C000800008000000000022000006808000",
INIT_12 => X"0000000000000A2281000000000040A3810000000000402001400000022002A0",
INIT_13 => X"000000000004200001C0400000000010200001C0400000000010000004490010",
INIT_14 => X"0001070004000000000000060000104C08000000000000001000000903008000",
INIT_15 => X"CC004050CA0C00020220200070040000010401C4000000000000000000100008",
INIT_16 => X"4310E4310A4210A4210A4210A4210A4210A8D0830A68010001B4DA881048061C",
INIT_17 => X"21084290A4210A4210A4210A4210A4210A4210A4210E4310E4310E4310E4310E",
INIT_18 => X"90A421084290A421084390E4310C4390E4310C4390E4310C4290A421084290A4",
INIT_19 => X"015303C0C78C706428A14C586291000A044001FFE000003FFC004290A4210842",
INIT_1A => X"2492492492492492492492492492492492410410410410412821600001249249",
INIT_1B => X"51A8D46A351A8D46A351A8D46A351A8D46A351A9D4EA753A9D4EA753A9D49249",
INIT_1C => X"FFFFFFFFFFFFFFFC00000000000000000000000038F56351A8D46A351A8D46A3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"55AB02055AB0207FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"420000000000000000000000000000000000000000000000007FFFAB57FFFAB5",
INIT_28 => X"A800BAFFAE9554508002AA00AA843DF55FFAA955EFA2D168B55557BEAA000055",
INIT_29 => X"002AB55AAAA955EF005568A00087BE8BFFA2D155410AA8415555087BFFF55A2A",
INIT_2A => X"AAABFF5508003FF555D0002145552ABFEBA007FC21EF007FD75FFAA841541008",
INIT_2B => X"082EBDEAAA2FBEAABA5D7FC0155005168B455D042AB45F7FFD741000042AA10A",
INIT_2C => X"FF7FBEAB55F7AABDEBA5D7FC2010A2D1575FFF7AA975555D2E80145F78415545",
INIT_2D => X"EF5555554AA087BC01FFFFAAAAB55552A954BAFFFFE8B55552EBDE00F7AEAABF",
INIT_2E => X"000082E820BAA2FBEAB5555557DF55A2AEBDF555D2E954BA002EAAABA002A821",
INIT_2F => X"FB7D5D7FEAA3808554203A000000000000000000000000000000000000000000",
INIT_30 => X"1557D1475FAF45BEAA800AAFFAA95578080038A2AA28E3AF55E3A0BA5D7AADB6",
INIT_31 => X"BD55D7BE80004AA1E8E2AB55B6A0925D7085F6AA10087FEABD7AAD57AEBAB68E",
INIT_32 => X"F5D0438140E2FA38B6AEBFF6D1D04AAFFA41040017D5D20B8EAA007FC51C7A2F",
INIT_33 => X"D0A901FFFF801557D1C20B8EAAA2FBE80AA557BE8B6D5D5FFABEF49002FB55FF",
INIT_34 => X"5D20BDE00EBAAA8BC7EBDFEAFEFAB8ABAE925D21C7010EADB525D7FFAE975C75",
INIT_35 => X"F002EADA921420871D74971D24820875C21D5EB8AA8FFF012A954BAFFF5EFB45",
INIT_36 => X"000000000000000000001C24820BAB6FFEFB6D555578F7DB6A0BDF7DEB8E125F",
INIT_37 => X"B55A28408145AAFFFFFFF5D7FEAABA0051400A20000000000000000000000000",
INIT_38 => X"AB55FAD568AA2AFAE975EF555168B55F7AA800BAF7AA955EF00042AAA2A2AEAA",
INIT_39 => X"2AAAA007FD55558A7BD7145FBB8020A35D2ABEF55F7800015F087FEAA00007FE",
INIT_3A => X"968F575D003FF55F7D5420BA5D2ABFEAAF7AE9DFF759A82AEF70800021EF5504",
INIT_3B => X"FFD5145FBAC9755F05040255FFD84175EF55002AAB0A2FFEAABA557BEA3EF057",
INIT_3C => X"82E974AAF7D57DF45552A3FF10AA8429F45A7D5EAF5FFBAEAAA10554155400AA",
INIT_3D => X"FF843FFE77C80825BC052ABFE10550415557085540000005156155FE90A8F5C0",
INIT_3E => X"00000000000000000000000000000000000005500020AAF7FBFFFEF04552ABFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_4,               -- Port A enable input
WEA      => wbe_a_hi_1024_4(0),               -- Port A write enable input
DIA(0)   => data_write_a(3),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_4(3),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_4,               -- Port B enable input
WEB      => wbe_b_hi_1024_4(0),               -- Port B write enable input
DIB(0)   => data_write_b(3),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_4(3),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_4_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A108400020612C80284210081034849800A00030300004833522C82D04A16002",
INIT_01 => X"2043998A1839284D1CA0650E1E504368403008418984014902030806A0D10200",
INIT_02 => X"C120042200000000044441CE01E80F00A49043118680008002000000026208E4",
INIT_03 => X"040001020019200020011209CC0164C060000000690111040144800042F5C403",
INIT_04 => X"7029AF0F81A00010CCA47700CC513CAC0D0B8E02010740E19754080108988021",
INIT_05 => X"02139405007133C0712244CD20F20105D583000020E9892201D304D42A9835E1",
INIT_06 => X"9190440300078002014405D9EE814C0284A883B6D7038AE079059B7800048092",
INIT_07 => X"000100AA0004408000000004840400008D200102503000782000C00C8025C000",
INIT_08 => X"00728A00408403220811991E02120C044058080004000001101121F220000260",
INIT_09 => X"811001E1185B38AD23C3707AD46440818F3CF80EC423CA7D01D123C80200816A",
INIT_0A => X"45810810A01B40216361056D6150F41200280001900439001FD8A00041400000",
INIT_0B => X"11FC88076266E800D605402962A820211500024808010512C40106D222223B14",
INIT_0C => X"0408804116040B02C02C500B0C02C100B0C02C100B0402C300B0401618058611",
INIT_0D => X"040200050200501301208482200D00D0A0408402C4282200A84800009B878680",
INIT_0E => X"00000020000100024AC88300300060090F0D830F00025400300204D018000804",
INIT_0F => X"8000000040000206A2000800000000000000950002E010000000080000588040",
INIT_10 => X"0000000000000808000554000200000000000100006D0020000000100000BB00",
INIT_11 => X"0000400000000000002000001A0002504001000000000000002280000D800800",
INIT_12 => X"0800000000000E2C802000000000408D801000000000408012440000200110A0",
INIT_13 => X"000000000004680003A0040000000010280003800800000000102800000B0000",
INIT_14 => X"000005C0002000000000000620000158000010000000000010A0000B00000200",
INIT_15 => X"C30146200400104002602600400000000294004000000004000000000010001A",
INIT_16 => X"0080200000008020000000802000000080080000004090014134DA101288C6DB",
INIT_17 => X"0802000000000401806010040180601004018060100000802000000080200000",
INIT_18 => X"8060180601004010040080200802000000000000802008020000000000008020",
INIT_19 => X"C0A28A063807E0500014063450404882846FFE000003FFC00000010040100401",
INIT_1A => X"AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA28A28A28A28A2934C8D0CCD145144",
INIT_1B => X"68341A0D068341A0D068341A0D068341A0D068351A8D46A351A8D46A351AAAAA",
INIT_1C => X"FFFFFFFFFFFFFFFC0000000000000000000000001FE32068341A0D068341A0D0",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"408102040810207FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"800AA00000000000000000000000000000000000000000000040810204081020",
INIT_28 => X"168B55557BEAB4500554200000557FE10FFFBEAA10007FD7410FFAA97555082A",
INIT_29 => X"55574105D2A800AA00043FEBA5D7FEAA00007BE8AAAAA843DF55FFAA955EFA2D",
INIT_2A => X"57BC00AAA2FFEAAAAAA8415555087BFFF55A2AA800BAFFAE9555508002AA0000",
INIT_2B => X"A2AA955EF005568A00087BE8BFFA2D17DE1000517FE10AAAAA8AAA002E975455",
INIT_2C => X"FAA8417410A2D140000F7FBC2010A2D157400AAAE974AAAAAA974BA08002AB55",
INIT_2D => X"EFA2AABDEAA087BEAAAAA2FBD54BA080002145552ABFEAA007FC21EF007FD75F",
INIT_2E => X"00055042AB45F7FFD741000042AA10AAAABFF5508003FF55F7D568A00552EA8B",
INIT_2F => X"5400F7A49057D0824850B8000000000000000000000000000000000000000000",
INIT_30 => X"3AF55F7A0925D7AADB6FB7D5D7FEAB7808554203A145178E00FFFBE8A101475D",
INIT_31 => X"A9557D080038AAA145157428492E8008200043FE925571EFA380871C7028A28E",
INIT_32 => X"AEA8A9200249056D4175C5092AAF5FDA38BE8E1557D1475FAF45BEAA800AAFFA",
INIT_33 => X"AA4954281C0E2FB55B6A0925D7085F6AA10087FEABD7AAD57AEBA08517DE00AA",
INIT_34 => X"007FC51C7007BD55D7BE80004AAFEDB42028EBFBC2028BED152438AAA092492A",
INIT_35 => X"AF7DF6AA00412EAABFFAA803DEBA0875EDA80BEF1C743840040017D5520B8EAA",
INIT_36 => X"0000000000000000000041002FB55FFF5D0438140E2FA38B6AEBFF6DBE84AAEB",
INIT_37 => X"A00FFFFEAA105D5155410FF84021EF0800154B20000000000000000000000000",
INIT_38 => X"DEBA0851574B2AAAEAAB55F78400145AAFFFFFEF5D7FEABFF0051400A25D5568",
INIT_39 => X"68B55F7AA800BAF7AA955EF00042AAA25555410BA082E8201000043FE005D517",
INIT_3A => X"568AA200557DE00AAAAAAA000804001FF005575408AA557FEB2FFAE975EF5551",
INIT_3B => X"D1550AAAA8002010F2AC154B25F2ABFF55F7800015F087FEAA00007FEAB55FAD",
INIT_3C => X"800021EF55042AAAA007FD5555087BD6145FAAC000A2A6FBC00BAAAFBC00BAF7",
INIT_3D => X"F7AEBDFF779A82AA43F7FBE8A00082EA8BFFAA843FEBA08517DE00F3F9574B30",
INIT_3E => X"000000000000000000000000000000000000008003FF55F7D5420BA5D2ABFEAA",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_4,               -- Port A enable input
WEA      => wbe_a_hi_1024_4(0),               -- Port A write enable input
DIA(0)   => data_write_a(4),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_4(4),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_4,               -- Port B enable input
WEB      => wbe_b_hi_1024_4(0),               -- Port B write enable input
DIB(0)   => data_write_b(4),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_4(4),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_5_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50DF4A0791B3FCB694379283C81FD996A091832102004A336A20E03C040C002",
INIT_01 => X"805FBDC69830A84D5C6A60000C34C26841280A00084000C8C212892EEAD53235",
INIT_02 => X"3B2026B578918E640A4F01CF8011FF0002080000082CA9998276DF7772C7C80D",
INIT_03 => X"37134108420D700084205702A4008A1D9100002171C0E0051554D93A11F5D140",
INIT_04 => X"8A41A0FC03A56DA000425A819410E3816C086198A388B702A8CA1210844A0C4C",
INIT_05 => X"B1808A062E8BC835F5E84532D708238A282F00A9291224800A2861490343082C",
INIT_06 => X"903FB8483A90581859050424100940825C6184401CDC451B860A6507160C4100",
INIT_07 => X"D26F068BCC96CDF8918E640E96D1A3469D6300E2FFEA27F8E4D23248130E259C",
INIT_08 => X"0BFA82E568442B2A082C0A7E3014250D49DA37A2420619000002AFF48D1222E5",
INIT_09 => X"3F005001E40969289429360416DCD1C46083030604B1CA20C03DF83B0A2C60A5",
INIT_0A => X"14613C71005A10492B888120288F480D58858449026145B3830F449449062B4F",
INIT_0B => X"11AC04934AC648BFD727C031E64170A137D5AA5C3E4B0F8A3C58C34C002290E3",
INIT_0C => X"CA29C6CC50384B6AC6AC86AB31AACA6AB39AAC86AB39AACA6AB3055643559C31",
INIT_0D => X"C673E33CF28F38603855401985228A0614BD30A0A2819852011E5AC2B87F9182",
INIT_0E => X"FF87C002F87A803E460B2516510CA594FF0044FFA4B08BAC4BB2CD0F09CF84E3",
INIT_0F => X"0DFF0F8005F0F5100DFFF5E15D06101C55EB29F1E00BE53FE1F000BE1E802F94",
INIT_10 => X"F12F0380231F17D78FC029FFF58D9A70380230F2FE0017C37FC3E0017C3D005F",
INIT_11 => X"FC7F023C0CA700125C0F8F7E43F1F001BFFE7C69E01804E1E7CCF8FC003FF5F1",
INIT_12 => X"023E00017C1FC1A4BFD82C3081C5BD27BFE30C3081C5BD00C02365D645CEEF5B",
INIT_13 => X"61E0042787F181E9C1EFD8CB8120C5AF41E9C18FD60F0C20666F41E9F009FFFD",
INIT_14 => X"7A7C077FFF404F80005F07F187A7D14BFFC96111C048278DEB074F9930FF9D80",
INIT_15 => X"C064014B8B652E2B3120C81284641D3E8DBF7D636FE860190700132C1F0EFB80",
INIT_16 => X"38CE1384E3384E338CE138CE1384E33C4E3ECE32E128882551349A1CBAA44103",
INIT_17 => X"84E3384E3384E3384E338CE138CE1384E3384E338CE138CE1384E3384E338CE1",
INIT_18 => X"CE138CE138CE138CE1384E3384E3384E3384E338CE138CE138CE138CE1384E33",
INIT_19 => X"F5E5BB4E7F7B9DB7FF3A1B6DB7E8410A8C000000000000000000384E3384E338",
INIT_1A => X"BEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEF9F7CFDFDDCF3CF3D",
INIT_1B => X"BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEFBEF",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000001711C7BBDDEEF77BBDDEEF77",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"FDFFF00000000000000000000000000000000000000000000080000000000000",
INIT_28 => X"FD7410FFAA97410082A800AAAAAE955450055421FFFFFBC0010AAD5574BA557F",
INIT_29 => X"7FD74000055574BA5D7FD7555A2D5575EF55517FF5500557FE10FFFBEAA10007",
INIT_2A => X"0002AABA5D2ABFFFFAA843DF55FFAA955EFA2D168B55557BEAB5500554200000",
INIT_2B => X"5D2A800AA00043FEBA5D7FEAA00007BC00AAAAAEBDF45A28428B45FFD168BFF0",
INIT_2C => X"5080028A00A2FFFDE00F7D57FEBAFF80174BAAAD1555EF555555555005557410",
INIT_2D => X"BA5D2E821FFA2D5554BA557BD75FFAA8415555087BFFF55A2AA800BAFFAE9555",
INIT_2E => X"00000517FE10AAAAA8AAA002E97545557BC00AAA2FFEAAAA082A97545F7D5420",
INIT_2F => X"7010BEDF524AA5571FDFEF000000000000000000000000000000000000000000",
INIT_30 => X"78E00EBFBE8A101475D5400F7A49043D0824850B8A2AE9756D145B401FFFFFFC",
INIT_31 => X"FEAB7D0855420BA1471D74380851524BA5571D757DB6D5525EF555178F6D1451",
INIT_32 => X"8A28B6DEBDF6DBEF1C0A28AAA5524BFFFFA28E3AF55F7A0925D7AADB6FB7D5D7",
INIT_33 => X"5555057D145152428492E8008200043FE925571EFA380871C7028B6AEBDF45B6",
INIT_34 => X"BEAA800AAFFAA9557D080038AAAA2FBF8E10EBD578EAAFF8415482BED1555EF5",
INIT_35 => X"81C209256DFFDF420BA552A821FFB6DF574A85575C55EFBE8E1557D1475FAF45",
INIT_36 => X"0000000000000000000008517DE00AAAEA8A9200249056D4175C50920875FDA3",
INIT_37 => X"5FF5D7BC21EFF7FBD7400F7FBC00BA55557DFF70000000000000000000000000",
INIT_38 => X"01FF5D5568BE7555568A00AAFFEAA105D5155410FF84020AA0800154B2AAAA97",
INIT_39 => X"00145AAFFFFFEF5D7FEABFF0051400A25551554BA0051400BA5551575EFF7D14",
INIT_3A => X"1574B2FFAABFF45FFAAAABFFAAFFFDFFF552EA8AAA55043DFF7AAAEAAB55F784",
INIT_3B => X"8002410FFD5575EF5555421E75555400BA082E8201000043FE005D517DEBA085",
INIT_3C => X"FAE975EF555168B55F7AA800BAF7AA955EF00002AAA2A2FBE8A00A2D16AAAAFF",
INIT_3D => X"0055554088A557FEB25D00021FFFFFFC00BA552A821EFFFFFD74BA5D51575F7F",
INIT_3E => X"000000000000000000000000000000000000000557DE00AAAAAAA000804001FF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_4,               -- Port A enable input
WEA      => wbe_a_hi_1024_4(0),               -- Port A write enable input
DIA(0)   => data_write_a(5),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_4(5),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_4,               -- Port B enable input
WEB      => wbe_b_hi_1024_4(0),               -- Port B write enable input
DIB(0)   => data_write_b(5),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_4(5),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_6_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10800B0061A01002840002C03002818000402322520070B313301C4389B2082",
INIT_01 => X"250041CA3839684D18A160000C52426841000000090800090210080008110200",
INIT_02 => X"0020042080010000044654C0000C008010000000001020900200200002620814",
INIT_03 => X"060881021088200021080200E4000A0891000020610111500104C00000F14400",
INIT_04 => X"0880000100000002000052288144004281C050400100280000C8100000080001",
INIT_05 => X"928080840001100A08009000280201000850E022401400002028214043410820",
INIT_06 => X"10100518090012122100C808049310002040000410A0001400000200120840D2",
INIT_07 => X"000100800004400001000000860408108C22000A502010074120044800040001",
INIT_08 => X"50000040D0C4E2088003FD01C01004044058082004000000000121F020408244",
INIT_09 => X"00BF17E9001205A5204911F814444080400100020000D200DFD16400C2A40AA0",
INIT_0A => X"04611C17849000022862A1596C8B5DF04834948900000100220C244840000880",
INIT_0B => X"03AD0413424E4044D665C070C22602291504400D084915020448114080201000",
INIT_0C => X"5E08864011088B22D22C008B0022C408B1022C208B0822C608B1111600458010",
INIT_0D => X"4251A12CD28A300429688001000800000020280204001000A00804309A002182",
INIT_0E => X"0000000280402400420800000000006200FC10002442042429324294014E8CA7",
INIT_0F => X"A40000000500800840000800000000000002280018001480000000A010100052",
INIT_10 => X"00000000000004C2003000010240000000000000680800290000000140202000",
INIT_11 => X"2000C0000000000000000442000001080001000000000000010C000280001804",
INIT_12 => X"08000000000801C300A010000000156000902000000015101200002800000000",
INIT_13 => X"000000000101800038002408000000094000386028040000000940000ED40000",
INIT_14 => X"0003B000002000000000020180002A24005010000000000023000060C7000A40",
INIT_15 => X"3F0280090321000040A410C28108000160008094000810040000000000002300",
INIT_16 => X"284A5284A728CA5284A528CA728CA52C4A5A0A32A300940101349A0408240818",
INIT_17 => X"9CA1294A329CA5284A728CA7284A5284A728CA5284A528CA728CA5284A728CA7",
INIT_18 => X"CA3294A129CA3294A129CA1294A329CA1294A3294A129CA3294A129CA3294A32",
INIT_19 => X"F5F78BCE7F8FF0F4FA955F7CF7F40A80145D55555556AAAAAAAAA94A329CA129",
INIT_1A => X"8E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E39B6CEDECDDF7DF7D",
INIT_1B => X"F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE38E3",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000001A1A33F9FCFE7F3F9FCFE7F3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"555FF00000000000000000000000000000000000000000000080000000000000",
INIT_28 => X"BC0010AAD5574BA557FFDFFF087BFDF45F7AA974AAAAAA97555F784174BAF7D5",
INIT_29 => X"515555508043FE00F7AA97555A2FBD7410AA8428AAAAAAE955450055421FFFFF",
INIT_2A => X"7D1575EFFFAA9555500557FE10FFFBEAA10007FD7410FFAA97400082A800AA08",
INIT_2B => X"0055574BA5D7FD7555A2D5575EF55517FF55A2AA97400552AAAB45082E80155F",
INIT_2C => X"500554200000003DE10FFD5401FFF7AAA8A10082EAAB45A2FFC2000007FD7400",
INIT_2D => X"10AA803FE105D516AABAFF843FFFFAA843DF55FFAA955EFA2D168B55557BEAB5",
INIT_2E => X"000AAAEBDF45A28428B45FFD168BFF00002AABA5D2ABFFFF087BD5545007BFDE",
INIT_2F => X"256DEB84104BAFFD1525FF000000000000000000000000000000000000000000",
INIT_30 => X"9756D145B401FFFFFFC7010BEDF524AA5571FDFEF1C7BFFF55FFA095482B6A49",
INIT_31 => X"4904380824850381C5B5057D1C003DE28F7A49057DAAF5D2428A2842AAAAA2AE",
INIT_32 => X"2AAFB451C2A8017DE3DF525FFFFA49756D145178E00EBFBE8A101475D5400F7A",
INIT_33 => X"2F1C50381471D74380851524BA5571D757DB6D5525EF555178F6DAAA49542841",
INIT_34 => X"AADB6FB7D5D7FEAB7D0855420BA1C0E3FE00E3DB471EFE3AAAAA00082EA8B6DA",
INIT_35 => X"F1C7BD057D1C71FFE10A28038E1049516AAB8FF8428FEFA28E3AF55F7A0925D7",
INIT_36 => X"00000000000000000000B6AEBDF45B68A28B6DEBDF6DBEF1C0A28AAA5524BFFF",
INIT_37 => X"F55F78017400F780001FFAA84000AAFFD1401E70000000000000000000000000",
INIT_38 => X"20BAAA8428AA2AAAA975FF5D7BC21EFF7FBD7400F7FBC00BA55557DFF7557BFD",
INIT_39 => X"EAA105D5155410FF84020AA0800154B2557FC01EF55043FEAAFF80021EFA2D14",
INIT_3A => X"568BE7AA80174AA082ABDF555D2A821EFAAFBC01FFF780155F7555568A00AAFF",
INIT_3B => X"AEA8A10082EA8BEFAAD5554B25551554BA0051400BA5551575EFF7D1401FF5D5",
INIT_3C => X"AAEAAB55F78400145AAFFFFFEF5D7FEABFF0051400A25D2EBFE10AAFFD55EFA2",
INIT_3D => X"552EA8AAA55043DFF7557BC01EF55557DE00AA842AA0000516AABAFF8428BE7A",
INIT_3E => X"0000000000000000000000000000000000000FFAABFF45FFAAAABFFAAFFFDFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_4,               -- Port A enable input
WEA      => wbe_a_hi_1024_4(0),               -- Port A write enable input
DIA(0)   => data_write_a(6),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_4(6),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_4,               -- Port B enable input
WEB      => wbe_b_hi_1024_4(0),               -- Port B write enable input
DIB(0)   => data_write_b(6),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_4(6),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_7_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10844B00482258A2842112C02450418800002300500030B313300C418992002",
INIT_01 => X"000009CA3839684D1CA0E0000E51424840000000080000080200080008510204",
INIT_02 => X"0120042086010000044600C00008000004100000000260900200000002402004",
INIT_03 => X"8628A10000082400000002408400080011000000610008000208C00000E14400",
INIT_04 => X"0911800100A000000000524084000040000050001140200100C8100000080102",
INIT_05 => X"0300812401011000000000002000114008008060441000000020024093000000",
INIT_06 => X"9190431C0D4010100000880804010010800000041080081000000200010424B2",
INIT_07 => X"000100AA0004408601000004860000008C02000A103010006928040800062481",
INIT_08 => X"84000048D484C20888000A0002120484C048007004000000000021F000000244",
INIT_09 => X"00A06009881201A520491004106C48A04040002400A15A208001650004001020",
INIT_0A => X"C99E1060201002044809C1040140A001004808810000459033189C0A400118A0",
INIT_0B => X"102000024040484050050041648A0041140C500B08821054C000264120000400",
INIT_0C => X"0404A083260E0832132011880462011880462051881462051881D31018C40620",
INIT_0D => X"0001000080001000813094801A8F80F00A600B52602801A88848011118003700",
INIT_0E => X"000003C007C002808228010410082042C000C000000004001002000400040002",
INIT_0F => X"A4000007800F80C840000800009864038A1200081C0014800000F001F0200052",
INIT_10 => X"00002C0E00E0E4004038000102400002C0E00E0D20100029000001E003E04000",
INIT_11 => X"2000C04031100E0403D0700300080908000100000661801E1900040380001804",
INIT_12 => X"0840878083E8003780A01043203A101780902043203A10082410082880000000",
INIT_13 => X"0601E0187900181035E0240806483248181035E0280410C8198818100DDD0000",
INIT_14 => X"0403774000201021E020FA006040376C00501022131210722060806D47000A40",
INIT_15 => X"00928A0002000110888600C032128201519480D40009902430160403E0E00506",
INIT_16 => X"01000000020080601802000000000405000A0020020081014134928820480010",
INIT_17 => X"0802018040000000006018020080200804010000000000806018020080000004",
INIT_18 => X"0000000001806008020000001006008020080001004008020080201004000020",
INIT_19 => X"0000000000000000000000000000400A004618618618C30C30C3000020180600",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000000B0840000000000000000000",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"1555500000000000000000000000000000000000000000000080000000000000",
INIT_28 => X"A97555F784174BAF7D5555FFF780155EFAAAEA8ABAAAFBFDE0055556AA005D04",
INIT_29 => X"55555EFAAFFFDFEFAAAAAAB455D556AA00FFAE95555087BFDF45F7AA974AAAAA",
INIT_2A => X"02EAAAAA082EA8A00AAAE955450055421FFFFFBC0010AAD5574BA557FFDFFF55",
INIT_2B => X"08043FE00F7AA97555A2FBD7410AA8428AAA557BFDFFF55003DFFFF7FBEAA000",
INIT_2C => X"0082A800AAF7AE975FFA28000010552EBDE00007BEAAAAA2D140000085155555",
INIT_2D => X"45087FEAB455D516AB55557BD55FF00557FE10FFFBEAA10007FD7410FFAA9740",
INIT_2E => X"000A2AA97400552AAAB45082E80155F7D1575EFFFAA955555D51574AAAAFFD55",
INIT_2F => X"AE105D556AA10410E17555000000000000000000000000000000000000000000",
INIT_30 => X"FFF55FFA095482B6A49256DEB84104BAFFD1525FFFF8E175C7A2AAAAA82A2F1F",
INIT_31 => X"F524AA5571FDFEF415B575D7AAF1FFFD7AAAAAFB7D495F6AA10E3AE905551C7B",
INIT_32 => X"003AFEFEBFBEAA001C2EA8A821C2EAAA00A2AE9756D145B401FFFFFFC7010BED",
INIT_33 => X"EDB470101C5B5057D1C003DE28F7A49057DAAF5D2428A2842AAAA497BFAFFF49",
INIT_34 => X"1475D5400F7A490438082485038F7A4905C7A28A070384120BDE100075EAA82B",
INIT_35 => X"D495150492BEF1D2555087BE8B7D555F6AB57417BC05D7145178E00EBFBE8A10",
INIT_36 => X"00000000000000000000AAA495428412AAFB451C2A8017DE3DF525FFFFA49756",
INIT_37 => X"555A2AEA8A10AAD568A00555168A10002E9754D0000000000000000000000000",
INIT_38 => X"8A10AAAE8215D557BFDF55F78017400F780001FFAA84000AAFFD1401E7FFAA97",
INIT_39 => X"C21EFF7FBD7400F7FBC00BA55557DFF7007BD5555AAD57DF55AAAEBDFEF007BE",
INIT_3A => X"428AA2007FE8BFF080028BFFAAFFEAA105D2EAAA005D2AAAA18AAAA975FF5D7B",
INIT_3B => X"043DE0000516AA10F7FBD7408557FC01EF55043FEAAFF80021EFA2D1420BAAA8",
INIT_3C => X"55568A00AAFFEAA105D5155410FF84020AA0800154B2FF8402145A2AA954AA00",
INIT_3D => X"AAFBC01FFF780155F7005140000FFD140145007FE8BEF557BEAB55087FC215D5",
INIT_3E => X"0000000000000000000000000000000000000AA80174AA082ABDF555D2A821EF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_4,               -- Port A enable input
WEA      => wbe_a_hi_1024_4(0),               -- Port A write enable input
DIA(0)   => data_write_a(7),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_4(7),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_4,               -- Port B enable input
WEB      => wbe_b_hi_1024_4(0),               -- Port B write enable input
DIB(0)   => data_write_b(7),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_4(7),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_8_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00000648E2840112C00000418000002700500030B3132000400812082",
INIT_01 => X"100008480009004C04A100000252024840000000180800080200010040110204",
INIT_02 => X"0020042000490000004600804008000005100000000024900200000002400004",
INIT_03 => X"0A0C33400008082400000080A4004B0891000020610112000040C00000E5C000",
INIT_04 => X"18800001000000000000512080000040800150400824280110C8100000120200",
INIT_05 => X"908084A10100100200004080280008240810802206940000012C214451610800",
INIT_06 => X"81B000080860109021400008040000202048020414A0021400040200322824C1",
INIT_07 => X"000000080004408049000004860000008402001A50208000630C040800062483",
INIT_08 => X"440000428644212280800A00021004044048002124000000000021F000000244",
INIT_09 => X"00004009001001010008100414644410400102228000D20080114502006409A2",
INIT_0A => X"000051312000042200294429148A4801C80C8C81000045907118040340020832",
INIT_0B => X"4020000240404140004D0544C4AA0001150410090302500011C813428A000400",
INIT_0C => X"46501090008820240240409000240009000240009000240009000120204808A5",
INIT_0D => X"42D1A168D09A301468402480004780F00140080860280004085904309A002196",
INIT_0E => X"00783FC00044340242280000000000020000C0000442106419120004034685A3",
INIT_0F => X"8000F07F800088A80000081EA2F9EC0000064004081010001E0FF00011104040",
INIT_10 => X"0ED0FC7E00000422201080000202658FC7E0000021882020003C1FE000222080",
INIT_11 => X"018059C3F350FE0C00000002A0040500000103961FE780000110010090000800",
INIT_12 => X"FD41FF80000830200021C1CF600012200010D1CF600012121600100810000004",
INIT_13 => X"9E1FE000010A1802100004343ED8000898021000087073D80008980200800002",
INIT_14 => X"0080200000BEB07FE00002086008020000209AEE3F300000246020200000620B",
INIT_15 => X"0088881903210000440610C8000A808040000208901786E4F0FE0C0000000166",
INIT_16 => X"685A1685A769DA368DA368DA769DA36CDA121A11A141800011309284002C0810",
INIT_17 => X"95A5685A1685A5695A368DA368DA769DA368DA368DA7695A1685A1685A5695A1",
INIT_18 => X"5A1695A568DA368DA369DA768DA1685A1695A5685A168DA369DA768DA368DA16",
INIT_19 => X"A4028A0A543EBC57A10A1E75D64108080468618618630C30C30C69DA5685A168",
INIT_1A => X"9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7BF3CCD8DF5B2DB2C",
INIT_1B => X"F87D3E1F4F87D3E1F4F87D3E1F4F87D3E1F4F87C3E1F0F87C3E1F0F87C3E79E7",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000006A6D4F87D3E1F4F87D3E1F4",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"155FF00000000000000000000000000000000000000000000080000000000000",
INIT_28 => X"BFDE0055556AA005D0415555080000000087BEAA10F7803DE00FFAEBFFFF0800",
INIT_29 => X"2AA8AAA557FC0010F780154105D7FC2145005155555F780155EFAAAEA8ABAAAF",
INIT_2A => X"7FFFFF55AA80155FF087BFDF45F7AA974AAAAAA97555F784174BAF7D5555FF55",
INIT_2B => X"AAFFFDFEFAAAAAAB455D556AA00FFAE95555AAFFE8A00552EBFE00F7D17FF45F",
INIT_2C => X"A557FFDFFF5504000AAAAAAA8B55F7D140010552E821EFAAAABDF555555555EF",
INIT_2D => X"55AA8028A00A2D57FF45557BE8A00AAAE955450055421FFFFFBC0010AAD5574B",
INIT_2E => X"000557BFDFFF55003DFFFF7FBEAA00002EAAAAA082EA8A00002AA8A10F784021",
INIT_2F => X"FE10F7AEBAFFF080A175D7000000000000000000000000000000000000000000",
INIT_30 => X"175C7A2AAAAA82A2F1FAE105D556AA10410E17555080E000280071E8A00EB8E3",
INIT_31 => X"4104BAFFD1525FF492EA8AAA5571C2000FF8A17400557FC015514555757DFF8E",
INIT_32 => X"2ABDE10EBDF7AF6DE3FFF8F7DB68A105D71C7BFFF55FFA095482B6A49256DEB8",
INIT_33 => X"AA0BDF6D415B575D7AAF1FFFD7AAAAAFB7D495F6AA10E3AE90555A2FBE8A3849",
INIT_34 => X"FFFFC7010BEDF524AA5571FDFEF550E00082B6A0AFB55F7D1420104124821D7A",
INIT_35 => X"01C2EA8A00F7800017DA2842FA00B6D578F6D557FFDA00A2AE9756D145B401FF",
INIT_36 => X"00000000000000000000497BFAFFF49003AFEFEBFBEAA001C2EA8A821C2EAAA0",
INIT_37 => X"0BA08556AA00AAAABFE00F7AEAABEF082E955450000000000000000000000000",
INIT_38 => X"21555D51575EFFFAA97555A2AEA8A10AAD568A00555168A10002E9754D082E82",
INIT_39 => X"17400F780001FFAA84000AAFFD1401E7082EAAABA5D5140010F7AE974105D7BC",
INIT_3A => X"E8215DA2FFE8ABA082ABFE00AAFBEABFFAAFBEABFFF7AA80145557BFDF55F780",
INIT_3B => X"D540000000402145AA843FFFF007BD5555AAD57DF55AAAEBDFEF007BE8A10AAA",
INIT_3C => X"AAA975FF5D7BC21EFF7FBD7400F7FBC00BA55557DFF75D2E82010F7843DF45FF",
INIT_3D => X"5D2EAAA005D2AAAA185D2AAAA10F780021FFA2803DE10FFD16ABFF5D7BFDE10A",
INIT_3E => X"0000000000000000000000000000000000000007FE8BFF080028BFFAAFFEAA10",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_4,               -- Port A enable input
WEA      => wbe_a_hi_1024_4(1),               -- Port A write enable input
DIA(0)   => data_write_a(8),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_4(8),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_4,               -- Port B enable input
WEB      => wbe_b_hi_1024_4(1),               -- Port B write enable input
DIB(0)   => data_write_b(8),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_4(8),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_9_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00018248A2840112C00002C18000002300500030B3132000400812006",
INIT_01 => X"400008000000004C0020000000100248413C0A61590001D90213C10008110204",
INIT_02 => X"01A0042080010000054600C04008000004100000001020900200200002420804",
INIT_03 => X"024003400008012400000010E4004B0891000020610310000144C00000F5C000",
INIT_04 => X"1801800100E000000000510084000040010050020810200000C8900000320200",
INIT_05 => X"918004311104100000000000200008100800002000100000002C234415610820",
INIT_06 => X"81B00008080010100000980804000008800042041080001000100200322C2481",
INIT_07 => X"0000811800044080010000058600000086020002502080006000040800062C80",
INIT_08 => X"0000004001D4618008800A00061004044048002004000000000061F000000244",
INIT_09 => X"000040090802009420409004104444084001022400214A2080014400026401A2",
INIT_0A => X"04000071200000A003CA294140200800C80C8C8100004590111C040040120800",
INIT_0B => X"12210002404848502847040164880021150400080222000200C8034200000000",
INIT_0C => X"4610088010080421021040841021000841021000841021000841010800420820",
INIT_0D => X"42D0A16C529A321068500484000500D10042080040284000084900001A002196",
INIT_0E => X"00000002804000004228010410082002C000C0002400046419120410034285A1",
INIT_0F => X"A00000000500800800000800000000000002290008001080000000A010100042",
INIT_10 => X"00000000000004C2001000000240000000000000680800280000000140202000",
INIT_11 => X"0000C0000000000000000442020001000001000000000000010C800080000804",
INIT_12 => X"08000000000801A7802010000000152780102000000015000600000800000000",
INIT_13 => X"000000000101900011E0240000000009500011E0280000000009500004DD0000",
INIT_14 => X"000137400020000000000201C000136C00101000000000002340002947000240",
INIT_15 => X"0080881901210000000600C280028000419480D4000010040000000000002304",
INIT_16 => X"68DA368DA1685A1685A1685A1685A16C5A121A13A141950051309284A82C0010",
INIT_17 => X"85A1685A1685A1685A368DA368DA368DA368DA368DA368DA368DA368DA368DA3",
INIT_18 => X"5A1685A168DA368DA368DA368DA368DA368DA368DA3685A1685A1685A1685A16",
INIT_19 => X"0157344CCCF48DE68A895C38E2540A8010100000000000000000685A1685A168",
INIT_1A => X"14514514514514514514514514514514514D34D34D34D34D28E1004039248209",
INIT_1B => X"D268341A4D268341A0D069349A0D069349A0D068341A0D068341A0D068345145",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000014D490D069349A0D068341A4",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"EAABA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"03DE00FFAEBFFFF0800155FFAAFBE8B45002A974AAAA803DFFFAA843DF45FFFF",
INIT_29 => X"7BFDE00A2FBD7400F7FBFDFFFA2AEBDE00AAFBEAABA080000000087BEAA10F78",
INIT_2A => X"055401FFF7AEAAA10F780155EFAAAEA8ABAAAFBFDE0055556AA005D041555508",
INIT_2B => X"557FC0010F780154105D7FC2145005155555557BE8BEF007FFDEAAAAD1555EF0",
INIT_2C => X"AF7D5555FFF780154AA5D2AA8A10F7AA974AA082E80010A2AAAAA10552AA8AAA",
INIT_2D => X"BAF7D17FEBAA2AEBDF45002EAAABA087BFDF45F7AA974AAAAAA97555F784174B",
INIT_2E => X"000AAFFE8A00552EBFE00F7D17FF45F7FFFFF55AA80155FF080400145FFFBEAA",
INIT_2F => X"8FC7BE8A3DF7DF7F5E8A92000000000000000000000000000000000000000000",
INIT_30 => X"000280071E8A00EB8E3FE10F7AEBAFFF080A175D7BEF1E8B6D002090482B68E3",
INIT_31 => X"56AA10410E175550871FFE00A2FBD0400FFF5FDFC7B6A0BDE38B6F5E8A92080E",
INIT_32 => X"7BFAE82A2DB555C71C5B451D7FFAAA8A38FF8E175C7A2AAAAA82A2F1FAE105D5",
INIT_33 => X"2AEADA38492EA8AAA5571C2000FF8A17400557FC015514555757D5D71E8BEF14",
INIT_34 => X"B6A49256DEB84104BAFFD1525FFFF84174BA5D20AAA00E3AA904BA142A87010A",
INIT_35 => X"7000400155FFFBEDA82FFD57DEBAAAA0BFF7D0024ADA921C7BFFF55FFA095482",
INIT_36 => X"00000000000000000000A2FBE8A38492ABDE10EBDF7AF6DE3FFF8F7DB68A105D",
INIT_37 => X"BEF080402000F7AAA8B55FFAABDFEFF7D16AA000000000000000000000000000",
INIT_38 => X"FEAAFFD16AA00082E820BA08556AA00AAAABFE00F7AEAABEF082E95545F7D568",
INIT_39 => X"A8A10AAD568A00555168A10002E9754D00517DE00A2FFC2000F7D17FF55FF803",
INIT_3A => X"1575EF555568BEF5D7FE8A10AAFFD55555D7FD5555FFAAA8AAAFFAA97555A2AE",
INIT_3B => X"AE800AA552A97400A2AEBDEAA082EAAABA5D5140010F7AE974105D7BC21555D5",
INIT_3C => X"57BFDF55F78017400F780001FFAA84000AAFFD1401E7FF80174AA5D0028A00AA",
INIT_3D => X"AAFBEABFFF7AA80145080002145F7FBFFE00FFD17FEAAA2803DFEF08043FE005",
INIT_3E => X"0000000000000000000000000000000000000A2FFE8ABA082ABFE00AAFBEABFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_4,               -- Port A enable input
WEA      => wbe_a_hi_1024_4(1),               -- Port A write enable input
DIA(0)   => data_write_a(9),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_4(9),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_4,               -- Port B enable input
WEB      => wbe_b_hi_1024_4(1),               -- Port B write enable input
DIB(0)   => data_write_b(9),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_4(9),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_10_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00018248A2840112C00002C18000202300500030B3132000400992006",
INIT_01 => X"254008000000004C002000000010026840000000080000080200010008110204",
INIT_02 => X"0020042000010000004455800008000004100000000000900200000002400004",
INIT_03 => X"020001021089000021081000C400090011000000610001540104C00000F14400",
INIT_04 => X"0811800101A00002000050088554004200C840000000200080C8100000000001",
INIT_05 => X"030080001000100800009400200000000840E020201000000024024001200020",
INIT_06 => X"81B00008080012120004CC080492500280208004148000100000020020042493",
INIT_07 => X"0000000800044080010000048404081085020002502000006000040800062480",
INIT_08 => X"100202400084410808000A00021004044048000004000000000021F020408264",
INIT_09 => X"010040090002008420401004144440004040022484214A2080110108C2C00320",
INIT_0A => X"04004166A48A0001080000000000080080181881000045901118044040020800",
INIT_0B => X"1201000200484910000F0105602622291404020902005002018002400A022000",
INIT_0C => X"0440001011808020120004801120044800120004801120044800110002400884",
INIT_0D => X"008000440210100041308480800F82F00040180260A808008848000018002104",
INIT_0E => X"000000028040000002280104100820020000400020000440100204100A000100",
INIT_0F => X"040000000500800800000000000000000002280008000400000000A010100010",
INIT_10 => X"00000000000004C2001000010000000000000000680800010000000140202000",
INIT_11 => X"200000000000000000000442000001000000000000000000010C000080001000",
INIT_12 => X"00000000000801C0008000000000154000800000000015000410000800000000",
INIT_13 => X"0000000001019800180000080000000958001800000400000009580002800000",
INIT_14 => X"0000A0000000000000000201E0000A0000400000000000002360002080000800",
INIT_15 => X"0080881000000000000600C28102800060000000000800000000000000002306",
INIT_16 => X"401004010040100401004010040100441020D0030008840051309A90BA884010",
INIT_17 => X"0902409024090240900401004010040100401004010040100401004010040100",
INIT_18 => X"1004010040902409024090240902409024090240902409024090240902409024",
INIT_19 => X"F546890A940FE0D3971243555205428290100000000000000000401004010040",
INIT_1A => X"8A28A28A28A28A28A28A28A28A28A28A28A28A28A28A28A29554199854514514",
INIT_1B => X"2B95CAE532994CA6532995CAE572B94CA6532994CA6532994CA6532994CA28A2",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000002718E72B94CA6532994CA657",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"FDE1000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"03DFFFAA843DF45FFFFEAABA007FC2155F7D155545AA80001EFAAFBEAB45557F",
INIT_29 => X"042AB55FFD168B55AA8000010FFFBE8BFFF78402155AAFBE8B45002A974AAAA8",
INIT_2A => X"AD16AABA002ABDE10080000000087BEAA10F7803DE00FFAEBFFFF0800155FF00",
INIT_2B => X"A2FBD7400F7FBFDFFFA2AEBDE00AAFBEAABAA2FFD741055003DFEFF7AA801FFA",
INIT_2C => X"05D0415555007FD74105555555EFF7FBC0145F78028A00A2D142155087BFDE00",
INIT_2D => X"55AAD168ABA002A975FFF7AEBDEBAF780155EFAAAEA8ABAAAFBFDE0055556AA0",
INIT_2E => X"000557BE8BEF007FFDEAAAAD1555EF0055401FFF7AEAAA105D042ABFF5D556AB",
INIT_2F => X"71D7AAFBEFB455D71F8E00000000000000000000000000000000000000000000",
INIT_30 => X"E8B6D002090482B68E38FC7BE8A3DF7DF7F5E8A92007BC217DEBDB55555AA8E0",
INIT_31 => X"EBAFFF080A175D700042AB7DEBDB6DB55BE8E05000EBFFE8BC7E38E07145BEF1",
INIT_32 => X"0A3DFD7F7A4821D7A2D16FA82142EB8E00080E000280071E8A00EB8E3FE10F7A",
INIT_33 => X"ED1421450871FFE00A2FBD0400FFF5FDFC7B6A0BDE38B6F5E8A92B6FBD541049",
INIT_34 => X"A2F1FAE105D556AA10410E175550071D54104951555D7EBF5C5155E3842AA00B",
INIT_35 => X"8410E2ABD749516FB55BED16FA820820955EFE3AEBDEAAFF8E175C7A2AAAAA82",
INIT_36 => X"000000000000000000005D71E8BEF147BFAE82A2DB555C71C5B451D7FFAAA8A3",
INIT_37 => X"1EFA2FFD7545AAAE97555A2FBFDF455D556AA000000000000000000000000000",
INIT_38 => X"8B45AAAA95545F7D568BEF080402000F7AAA8B55FFAABDFEFF7D16AA00087FC0",
INIT_39 => X"6AA00AAAABFE00F7AEAABEF082E9554500042ABFFA2FFFFF45F7AE97400AAFFE",
INIT_3A => X"16AA00FFFBD5400082EBFF45F78400155A2D57FE00552EA8A00082E820BA0855",
INIT_3B => X"D557555A2802AA10FFD54214500517DE00A2FFC2000F7D17FF55FF803FEAAFFD",
INIT_3C => X"FAA97555A2AEA8A10AAD568A00555168A10002E9754D085155410085557555AA",
INIT_3D => X"5D7FD5555FFAAA8AAA002AAAB4508557DF55F7D17FE000804155FFAAAABDEAAF",
INIT_3E => X"0000000000000000000000000000000000000555568BEF5D7FE8A10AAFFD5555",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_4,               -- Port A enable input
WEA      => wbe_a_hi_1024_4(1),               -- Port A write enable input
DIA(0)   => data_write_a(10),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_4(10),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_4,               -- Port B enable input
WEB      => wbe_b_hi_1024_4(1),               -- Port B write enable input
DIB(0)   => data_write_b(10),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_4(10),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_11_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A101C4B05A0034CA2840712C2D001419000002300500030B31B20084EC992002",
INIT_01 => X"90000986B83028491800E0000C26426040000000080000088200080802512224",
INIT_02 => X"1A2004205E010640024D00800008000004100000040EC090820018003241A00C",
INIT_03 => X"28639100000C5C00000045C08400C8001100000061806A001618C03001E54400",
INIT_04 => X"1A800001000009A0804059A190000040400040008058220008C8100000120D4E",
INIT_05 => X"02000E81080250010000002022000058080400000E1200000020004401000004",
INIT_06 => X"819435143F20101010001008040800B8100102041088011100022200000024B2",
INIT_07 => X"90640D280884453E01064002944180008402001295BA100022E4340800062D82",
INIT_08 => X"400000093204802200280A0012160585C1D808D004000000000323F40C102244",
INIT_09 => X"380040098010001100009204107C5950400000220080C200800900020C006827",
INIT_0A => X"80007100004016EA080801010000080D00200081000045B0511D289940103399",
INIT_0B => X"002000024040410A000D0104408810C115D9C008050042400100D04E88000002",
INIT_0C => X"00655010009264201200C7B421ED0C7B421ED0C7B431ED087B43176843DA1085",
INIT_0D => X"0401020080400A10012494881A4F80F209500BB2602881A488485C1318002000",
INIT_0E => X"6619A540124814800228010410082022C00040002020090020220C9600040802",
INIT_0F => X"ACCC334A802491600C587949B6D0141B4CC600D5761B1599865A500490B86A56",
INIT_10 => X"BAC845542056A61686EC81E3A6CB68AA2C622C9A251C352B330CB4A0092170D8",
INIT_11 => X"BCCAD0B5A81536080CC6B21A21B1FC09CB0F1076D4A200B2AD4068F4101639B5",
INIT_12 => X"4D2CC281E31AA0103AB8D5514066380804B268A2E060901204112566F10AC418",
INIT_13 => X"D551443C47281002540B2C9AAAA8662A1152B202AE3554403028115AA88201A1",
INIT_14 => X"548A20A0492A2724A0621620402A020141F172FB182A32AB6845AB6200251BC9",
INIT_15 => X"00C00A000200074044E6801832728080D00A380B753952C4877E0104DDE4D124",
INIT_16 => X"0080200802008020080200802008020480080022020081010124988800400010",
INIT_17 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_18 => X"0000000000802008020080200802008020080200802008020080200802008020",
INIT_19 => X"55062608804180C0B10A42104201400204000000000000000000000000000000",
INIT_1A => X"00000000000000000000000000000000000820820820820801C4149470000000",
INIT_1B => X"0000000000000000040200000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000007E0F0000000000000100800",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"000AA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0001EFAAFBEAB45557FFDE10082ABDF5508557DF45002ABDFFFF7803DE10AA80",
INIT_29 => X"AEBFF45FFAEBFEAA002A801FFF7FFE8A10A28000000007FC2155F7D155545AA8",
INIT_2A => X"2AABFE10082ABFFEFAAFBE8B45002A974AAAA803DFFFAA843DF45FFFFEAABAA2",
INIT_2B => X"FFD168B55AA8000010FFFBE8BFFF78402155AAD155555A28428BFF002ABDE00A",
INIT_2C => X"F0800155FF00557FF45557FC2010002A80010A2842AAAA007BFFF4500042AB55",
INIT_2D => X"FF5D00154BAF7FBE8BEFFFD540000080000000087BEAA10F7803DE00FFAEBFFF",
INIT_2E => X"000A2FFD741055003DFEFF7AA801FFAAD16AABA002ABDE10A2D168A10A284021",
INIT_2F => X"DFC7F78E3FE28B684070AA000000000000000000000000000000000000000000",
INIT_30 => X"C217DEBDB55555AA8E071D7AAFBEFB455D71F8E00002EBDF6D005B78F7D142AB",
INIT_31 => X"A3DF7DF7F5E8A92BEAEBFF7DEBA0BDEAA1C2A801C7E3FFEFA10B68407038007B",
INIT_32 => X"8A28BFF082ABAE10B6AAB8E280820B8FEFBEF1E8B6D002090482B68E38FC7BE8",
INIT_33 => X"07FF8F7D00042AB7DEBDB6DB55BE8E05000EBFFE8BC7E38E07145B6D15756DA2",
INIT_34 => X"EB8E3FE10F7AEBAFFF080A175D708517DF7D497BC5028142A87000A28A2AA920",
INIT_35 => X"0B6DB6AA28A280001FF5D0A10482FFFFEFBC7E3DF42028080E000280071E8A00",
INIT_36 => X"00000000000000000000B6FBD5410490A3DFD7F7A4821D7A2D16FA82142EB8E0",
INIT_37 => X"FEF007BE8BFF5D2ABDF55F7AABDEAAF784154BA0000000000000000000000000",
INIT_38 => X"DE00FF84154BA087FC01EFA2FFD7545AAAE97555A2FBFDF455D556AA00082EBF",
INIT_39 => X"02000F7AAA8B55FFAABDFEFF7D16AA00FFAEBFFEFAA803DEBA5D2E82155A2FBF",
INIT_3A => X"A95545F7D5555FFAAAAA8BFF002AAAA00FFAAA8AAA080028BFFF7D568BEF0804",
INIT_3B => X"2E95400A2AEA8A00007FEABFF00042ABFFA2FFFFF45F7AE97400AAFFE8B45AAA",
INIT_3C => X"82E820BA08556AA00AAAABFE00F7AEAABEF082E9554508557DFFF007BD54BA5D",
INIT_3D => X"A2D57FE00552EA8A00FFFFE8AAAAA80001FF5D2E82000F7FFFFF45AAFFC20BA0",
INIT_3E => X"0000000000000000000000000000000000000FFFBD5400082EBFF45F78400155",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_4,               -- Port A enable input
WEA      => wbe_a_hi_1024_4(1),               -- Port A write enable input
DIA(0)   => data_write_a(11),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_4(11),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_4,               -- Port B enable input
WEB      => wbe_b_hi_1024_4(1),               -- Port B write enable input
DIB(0)   => data_write_b(11),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_4(11),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_12_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50080B01BC002006940202C0DE041196A83183000000023322287E0FC000006",
INIT_01 => X"75400D849830C84C5823E0000C17424840000000080000088200002802153231",
INIT_02 => X"18A026B43ED180040147558040090000061800000C06ED9802768F4472C52005",
INIT_03 => X"2A67E34A528D0524A52850528400C8001100000171C02B550618C91A10E55440",
INIT_04 => X"1BC0000100056C8280825DE98154004300C840800850240080CA921084520A07",
INIT_05 => X"02000F832000500C0000941024000852084060202E100001002000448100000C",
INIT_06 => X"819A1D1C3FE01A1A40045408049A50BA4020C6041090001200006200000000F2",
INIT_07 => X"C26A0719CC96CC6ED18A64019695A854870300FA3968B20068FC06080106249F",
INIT_08 => X"D002024B3E040800008C0A002610240D494A06F3460409000000E3F0AD5282E5",
INIT_09 => X"27A06009200040000400120412445D78400001000410420080218029CC807A27",
INIT_0A => X"18000006848A026F000000000000080000F010C100204593F11A6CDF48003BF8",
INIT_0B => X"000000820040402B28050400400432C9349DF21A31A00ACC0000F04F80020001",
INIT_0C => X"00357804611AE45D05D0833430CD0833420CD0C33420CD0833430668619A1000",
INIT_0D => X"0000000000000A74812DF00E87E80A079F9F90FA0280E87E800C7FF3B8002000",
INIT_0E => X"3B6B0E404D26160682082002000401EA0000C40000800A006002818808000000",
INIT_0F => X"A476D61C809A4DA84272592D6246FC1B17B541F97E1B348EDA93900B2B286C56",
INIT_10 => X"30C669E622DBC325CFD881A962454CFBE5403AB99594362B1DB52720165650D9",
INIT_11 => X"F8D2D39A3745261E4A95A110A3F855000E4B1D32BAB504BB7490FCFF912A3834",
INIT_12 => X"B90E9B018C7530200AB8F8BF41F9A22006B37DC8E1F9A21A70116D4C5080651C",
INIT_13 => X"118780319CCA08AB1001ACDF34B8F1C688AB1002AE3F7B807B6289F368828C4C",
INIT_14 => X"2AF020233376A5ECC016B1A827CDA21160F051DE610A34C50427E6E220323E4A",
INIT_15 => X"0077020000000439FDC05C5806781FAB46095A0B5199B0AC55521524F1864022",
INIT_16 => X"000000000000000000000000000000000026C000002884000130921092804010",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"8020080200000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0051B946088881360A95090CB054420290100000000000000000008020080200",
INIT_1A => X"041041041041041041041041041041041049249249249249200100002D451451",
INIT_1B => X"92C964B2592C964B2592C964B2592C964B2592C86432190C86432190C8641041",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000003800F592C964B2592C964B25",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"7DE1000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"ABDFFFF7803DE10AA80000AAAA843FE0008557DFFF0800020105D557FEAA0055",
INIT_29 => X"D5420000051555FFA2AA8200000557DFFFF7AA80000082ABDF5508557DF45002",
INIT_2A => X"82AA8AAAAAFFC00BA007FC2155F7D155545AA80001EFAAFBEAB45557FFDE10AA",
INIT_2B => X"FFAEBFEAA002A801FFF7FFE8A10A28000000A2D155410F7FFFFEBA08003FE000",
INIT_2C => X"5FFFFEAABA000028A105D2ABFE10A2AABFE1055516ABEF5D517DEAAA2AEBFF45",
INIT_2D => X"55002A820AA08557DFFFF7AA82155AAFBE8B45002A974AAAA803DFFFAA843DF4",
INIT_2E => X"000AAD155555A28428BFF002ABDE00A2AABFE10082ABFFEF0855420000004175",
INIT_2F => X"5010495B7AE921C517DE10000000000000000000000000000000000000000000",
INIT_30 => X"BDF6D005B78F7D142ABDFC7F78E3FE28B684070AABE803AE38145B78FD700000",
INIT_31 => X"BEFB455D71F8E00BED547038145B505FFB6A487000005F7AFD7F7A482038002E",
INIT_32 => X"F1FDE821C003FE001C2EAAAAAB6F5C2082007BC217DEBDB55555AA8E071D7AAF",
INIT_33 => X"D517DEAABEAEBFF7DEBA0BDEAA1C2A801C7E3FFEFA10B68407038B6D550428FF",
INIT_34 => X"B68E38FC7BE8A3DF7DF7F5E8A9200002FA285D20BDE28A2A4B8E10555B68BEF5",
INIT_35 => X"F085F47038140010555142082082005F7DFD7F7A482155BEF1E8B6D002090482",
INIT_36 => X"00000000000000000000B6D15756DA28A28BFF082ABAE10B6AAB8E280820B8FE",
INIT_37 => X"ABA5D7FEAB45080015410007FEAA0055517DE000000000000000000000000000",
INIT_38 => X"AB45F780020BA082EBFFEF007BE8BFF5D2ABDF55F7AABDEAAF784154BAF7802A",
INIT_39 => X"D7545AAAE97555A2FBFDF455D556AA00F7D1554BA5D7BC01FFFF8015410007FE",
INIT_3A => X"4154BAF7D1400BAFFD57FE005D043FE10552EAAAAAFFD140000087FC01EFA2FF",
INIT_3B => X"8428A105D7FEABEF55557DEBAFFAEBFFEFAA803DEBA5D2E82155A2FBFDE00FF8",
INIT_3C => X"7D568BEF080402000F7AAA8B55FFAABDFEFF7D16AA0008003FEBA55003DEBAA2",
INIT_3D => X"FFAAA8AAA080028BFF087BD54AA550402145550000010087FFFF45F78402145F",
INIT_3E => X"0000000000000000000000000000000000000F7D5555FFAAAAA8BFF002AAAA00",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_4,               -- Port A enable input
WEA      => wbe_a_hi_1024_4(1),               -- Port A write enable input
DIA(0)   => data_write_a(12),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_4(12),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_4,               -- Port B enable input
WEB      => wbe_b_hi_1024_4(1),               -- Port B write enable input
DIB(0)   => data_write_b(12),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_4(12),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_13_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10154A0441836CA2840512822007C18000E02700500030B31B300040081A042",
INIT_01 => X"00000804A000C04800020000000002404001000008220008A200100802110204",
INIT_02 => X"02200430000104000A4700804008000004100000000420918204D3033240400D",
INIT_03 => X"AA4003400008592400000590C40009141100000C6180C0000000C00001E14000",
INIT_04 => X"0800000102400120088054019000004160004190BAA0270000C8100000600206",
INIT_05 => X"21000012040610050040000227003AA0082400E94C1200000824424005220020",
INIT_06 => X"81963B180C001010580000080400000058000004109C00138000020024142581",
INIT_07 => X"002C8008000441600106400A9600010494020002B8AAA000EF003408000E2580",
INIT_08 => X"000000E48194408000A00A001210040441C80320040210000002ABF004102244",
INIT_09 => X"2A004009640040100400940412D4C4004000022000104200802D983000480120",
INIT_0A => X"8000202020401480000000000000080C90090881000145B0111A14004015080D",
INIT_0B => X"00000002004040AA08050400404040C11444000805200A402090024000008002",
INIT_0C => X"8410000A00280020020040800020040800020000801020000800010020400000",
INIT_0D => X"84A14250A055100050100490000500D00040080040290000084E4000B800610C",
INIT_0E => X"DCD13042BEDA36820228000000000000C000400081A08BC812A2092B02850942",
INIT_0F => X"89B9A260857DB400431969CA985D480949D32804A40AB137341C10B7D6A02EC0",
INIT_10 => X"E6ACA678001CE7D0296C213A460CA4271CA2168AEC1017606E6838216FAD4055",
INIT_11 => X"84AD4961C281B20213073C5FC0058008632D30D522CE80239DCC01AB013A4D20",
INIT_12 => X"2E6B13804A4B01D83461299900F6BD583A519104A0EEBD1A141010B2A4C8E116",
INIT_13 => X"89E5E40913419151EE0E94641828F72B5151EE0D184B321037AF5158BB02D085",
INIT_14 => X"562EC0B42162D68EE0073AE1C562EC13D521921A4170300B2B458B56B01C2280",
INIT_15 => X"00888A120240034000E6DC8285028014B82372011FC1E4F5E0A00929684EAF84",
INIT_16 => X"50942509425094250942509425094254940A1421420082020120908800480030",
INIT_17 => X"0942509425094250942509425094250942509425094250942509425094250942",
INIT_18 => X"9425094250942509425094250942509425094250942509425094250942509425",
INIT_19 => X"F7EFBBEEFF3F7DF7FF3E9F7DF7E2450228000000000000000000509425094250",
INIT_1A => X"BAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBF7DFDFDDD555555",
INIT_1B => X"EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAEBAE",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000000000F7EBF5FAFD7EBF5FAFD7",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"2ABEF00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0020105D557FEAA00557DE10AAD5554BA087FFFF55557BD54AAF7FBC01FFA280",
INIT_29 => X"7BD75EF087FFFFEF557BEAB45552E80155AA802AB45AA843FE0008557DFFF080",
INIT_2A => X"FAE820AA5D5557555082ABDF5508557DF45002ABDFFFF7803DE10AA80000AA08",
INIT_2B => X"0051555FFA2AA8200000557DFFFF7AA80000AAD1420AA087BD7555FFD168AAAF",
INIT_2C => X"5557FFDE10AAAEA8BFFA2FBD7545FFD157555085140010F7AEAABFFAAD542000",
INIT_2D => X"BA557BE8A10A284154BAFFAAAAB45007FC2155F7D155545AA80001EFAAFBEAB4",
INIT_2E => X"000A2D155410F7FFFFEBA08003FE00082AA8AAAAAFFC00BA00002AAAAF7D5574",
INIT_2F => X"0492E3F1C71C7BE8A2ABD7000000000000000000000000000000000000000000",
INIT_30 => X"3AE38145B78FD7000005010495B7AE921C517DE10A2DB50482147FFAF554971D",
INIT_31 => X"E3FE28B684070AA1C71D25D7007FFAFD7497BE8B5555208217DBE8A2AB45BE80",
INIT_32 => X"7FD257DFFD568A82FFA4870BA555F5056D002EBDF6D005B78F7D142ABDFC7F78",
INIT_33 => X"FAAAFBFFBED547038145B505FFB6A487000005F7AFD7F7A482038AADF4709214",
INIT_34 => X"AA8E071D7AAFBEFB455D71F8E00A2A0ADBC7A2FFD257DE3DF52555085142000F",
INIT_35 => X"21C002AA92FFDF574824171EAA10B680124BAFFAAAFB45007BC217DEBDB55555",
INIT_36 => X"00000000000000000000B6D550428FFF1FDE821C003FE001C2EAAAAAB6F5C208",
INIT_37 => X"0105D7BE8B55085142010AAD157545F7AEA8B550000000000000000000000000",
INIT_38 => X"01EFF7AAA8B55F7802AABA5D7FEAB45080015410007FEAA0055517DE00A2FFC0",
INIT_39 => X"E8BFF5D2ABDF55F7AABDEAAF784154BA5D5140145007BE8B55087BEAB555D040",
INIT_3A => X"0020BAA2FFD54105D7FC21EFFFD16AA10FF80174AA557FC21EF082EBFFEF007B",
INIT_3B => X"FBC0155085540000FFAEBFFEFF7D1554BA5D7BC01FFFF8015410007FEAB45F78",
INIT_3C => X"87FC01EFA2FFD7545AAAE97555A2FBFDF455D556AA00A2803FF45AAFFC21EFAA",
INIT_3D => X"552EAAAAAFFD1400005D042AA00F7FBD5410085568A10FF80020AAFFAABFF550",
INIT_3E => X"0000000000000000000000000000000000000F7D1400BAFFD57FE005D043FE10",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_4,               -- Port A enable input
WEA      => wbe_a_hi_1024_4(1),               -- Port A write enable input
DIA(0)   => data_write_a(13),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_4(13),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_4,               -- Port B enable input
WEB      => wbe_b_hi_1024_4(1),               -- Port B write enable input
DIB(0)   => data_write_b(13),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_4(13),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_14_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10020A000180000284008280000281800000030000000033022000000580002",
INIT_01 => X"000008020000204D006800000030824840000000084000084200090008510200",
INIT_02 => X"0220043170010A600A4D008040080000041000000028009002000F333240800C",
INIT_03 => X"111813400008002400000000C400090011000000610200001104D83000F14000",
INIT_04 => X"0801800100A000000000540084000040000040000800200000C8100000000748",
INIT_05 => X"0100000000001000000000002000080008000000001000000024024001200020",
INIT_06 => X"819EB84028001010000000080400000000000004108000100000020020040081",
INIT_07 => X"92040608000440100102400A94810206844200021DA2A0002000340800062C80",
INIT_08 => X"000000000084400008800A001214040441481500040000000000A7F408002244",
INIT_09 => X"0A0040090002008420401004104444004000020400214A208001000002400120",
INIT_0A => X"0400002020000000000000000000080C8008088100004590111B480040120000",
INIT_0B => X"1000000200404800000504016000002114000008020000020080024000000000",
INIT_0C => X"0410000010000000000040001000000000000040000000000001000000000000",
INIT_0D => X"04810244825010004010000000000000000000000000000000080000B8002104",
INIT_0E => X"0002C38280001202020800000000001000004000000000401022000002040902",
INIT_0F => X"20000587050001404E8084341CBA3404800828805200008000E0E0A000080002",
INIT_10 => X"4D18178E012010C00224004091C3514072C000444A0400080001C1C140001000",
INIT_11 => X"51709A07424142084458476001003809D0104B01C5710044020C4006010500C5",
INIT_12 => X"C26EE3803180C18006519462A00005001460E4730000050A1011004001060049",
INIT_13 => X"01F9E00660318000000538318740000140000001B4600CE80001400000002B62",
INIT_14 => X"0000000AD89857B0E0684411800000003799EB764D000330C300000000E3554B",
INIT_15 => X"0000021002002C000024008284001A0902000422E3F5960080480A0216A07240",
INIT_16 => X"4090240902409024090240902409024090081021020080015134920800480010",
INIT_17 => X"0902409024090240902409024090240902409024090240902409024090240902",
INIT_18 => X"9024090240902409024090240902409024090240902409024090240902409024",
INIT_19 => X"F5579B4E5C8FF0F7BE9D5F7DF650400200000000000000000000409024090240",
INIT_1A => X"9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7BF7DDDDDFCF3CF3D",
INIT_1B => X"F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE79E7",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000003FFF03F9FCFE7F3F9FCFE7F3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"420BA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"BD54AAF7FBC01FFA2802ABEFA2FBE8B55A2AE80000F7D5555555D2AAAABAAAD1",
INIT_29 => X"AA801FFA28402000AAAE955455500155EF0804155EFAAD5554BA087FFFF55557",
INIT_2A => X"7AEA8B45080417400AA843FE0008557DFFF0800020105D557FEAA00557DE10A2",
INIT_2B => X"087FFFFEF557BEAB45552E80155AA802AB4500516AA00A2AE800BAFFFFC20BAF",
INIT_2C => X"0AA80000AA005568ABAA28402010A2843FEBAFFFBD7410A2D168BFF087BD75EF",
INIT_2D => X"005D7FFDF4555517DFEF00043FEAA082ABDF5508557DF45002ABDFFFF7803DE1",
INIT_2E => X"000AAD1420AA087BD7555FFD168AAAFFAE820AA5D5557555002E80155A280000",
INIT_2F => X"0555412AA8ABAAADB40092000000000000000000000000000000000000000000",
INIT_30 => X"50482147FFAF554971D0492E3F1C71C7BE8A2ABD7A2FFEDB55B6A080038E3DB5",
INIT_31 => X"B7AE921C517DE10A2AE851FFB68402038AAAA955554900105FF0800175D7A2DB",
INIT_32 => X"A0800BAE3F1C0092EBAAADB6D080A12410BE803AE38145B78FD7000005010495",
INIT_33 => X"2D568BC71C71D25D7007FFAFD7497BE8B5555208217DBE8A2AB451C556FA00A2",
INIT_34 => X"142ABDFC7F78E3FE28B684070AA00516DABAA28402038B6803DE82F7F5D5410A",
INIT_35 => X"D002A80155B680000105D7FF8F455D5F78FD7000E3FEAA002EBDF6D005B78F7D",
INIT_36 => X"00000000000000000000AADF47092147FD257DFFD568A82FFA4870BA555F5056",
INIT_37 => X"F55FF84000AAAAFBC0145002AA8AAAAAFFC20000000000000000000000000000",
INIT_38 => X"01EF080417555A2FFC00105D7BE8B55085142010AAD157545F7AEA8B55A2FBFF",
INIT_39 => X"EAB45080015410007FEAA0055517DE00A2AA955FFFF80020BAAAAA9754508000",
INIT_3A => X"AA8B555D557FE00A280020BAAAD140000A2AEBFFEF082A82010F7802AABA5D7F",
INIT_3B => X"803DE00FFD557400AAD56AB455D5140145007BE8B55087BEAB555D04001EFF7A",
INIT_3C => X"82EBFFEF007BE8BFF5D2ABDF55F7AABDEAAF784154BA08557FEAAA284000AAFF",
INIT_3D => X"FF80174AA557FC21EF082A80145F780020105D7BEAB45557BE8B45082EBFEBA0",
INIT_3E => X"0000000000000000000000000000000000000A2FFD54105D7FC21EFFFD16AA10",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_4,               -- Port A enable input
WEA      => wbe_a_hi_1024_4(1),               -- Port A write enable input
DIA(0)   => data_write_a(14),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_4(14),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_4,               -- Port B enable input
WEB      => wbe_b_hi_1024_4(1),               -- Port B write enable input
DIB(0)   => data_write_b(14),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_4(14),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_15_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000A000000000284000280000001800020030000000033022000000180002",
INIT_01 => X"8000080000000048000000000000026040000000080000080200000000110200",
INIT_02 => X"0020042004010E60004C0080000800000410000000020090020000300245E005",
INIT_03 => X"0000010000080400000000408400480111000000610008000000C00000E54400",
INIT_04 => X"980000010000000088C2550080000040000040000008A00028C8100000120000",
INIT_05 => X"020004012E025000000001322000000A28008000011000000220004D41000000",
INIT_06 => X"819588000800101000011008040000100001060418800510000A620000000092",
INIT_07 => X"0000000800044004010C20008440810284020002102220002000340800062480",
INIT_08 => X"0000000001140800002C0A001214050540C800400406180000002DF004000244",
INIT_09 => X"1E00400900000000000016041044400440000000000042008001000000000022",
INIT_0A => X"0000000000000220000000000000080C00000081000045901118000040000000",
INIT_0B => X"0000000200404000010500004000000114000009000000000000004200000000",
INIT_0C => X"0000000000000000000040001000040001000000000000000001000020000800",
INIT_0D => X"000000000000001001208000180800000000030200000180800C400030002000",
INIT_0E => X"0000000000002600020800000000001080004000000000000002000000000000",
INIT_0F => X"A400000000000000000008000000000000000000000014800000000000000052",
INIT_10 => X"0000000000000000000000010240000000000000000000290000000000000000",
INIT_11 => X"2001C05838120800000000000000000000010000000000000000000000001804",
INIT_12 => X"081004000000000000A010000000000000902000000000180010002020000000",
INIT_13 => X"6600000000000000000024080000000000000000280400000000000000000000",
INIT_14 => X"0000000000200801000000000000000000501001920000000000000000000A40",
INIT_15 => X"0000020000000000000000003000000000000000000A101C3614000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000080000120980000000010",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000400200000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"28BEF00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"5555555D2AAAABAAAD1420BAFF8000010082A954BA00003DFEF085155400F784",
INIT_29 => X"AE95555A2FBE8BEFA2843DE00AA8015400FF84001EFA2FBE8B55A2AE80000F7D",
INIT_2A => X"2FBEAB45F7D56AABAAAD5554BA087FFFF55557BD54AAF7FBC01FFA2802ABEFF7",
INIT_2B => X"A28402000AAAE955455500155EF0804155EFFFFBE8BFF0800174AA557BFDE10A",
INIT_2C => X"A00557DE10F7D1574AAA2D16AB55FFD568BEF087FE8A1055003FE00A2AA801FF",
INIT_2D => X"00AA802AA00AAAE800BA5D0015545AA843FE0008557DFFF0800020105D557FEA",
INIT_2E => X"00000516AA00A2AE800BAFFFFC20BAF7AEA8B45080417400FFFFC21450800154",
INIT_2F => X"8FD7005150438F78A2DBFF000000000000000000000000000000000000000000",
INIT_30 => X"EDB55B6A080038E3DB50555412AA8ABAAADB40092E38E070280024904AA1C043",
INIT_31 => X"1C71C7BE8A2ABD7E3AA9257DA2FFE8BC7BE8E38E10A28017400E38A051FFA2FF",
INIT_32 => X"00124AA557FFDE10A2FBEDB6DF7D16AABAA2DB50482147FFAF554971D0492E3F",
INIT_33 => X"10038E38A2AE851FFB68402038AAAA955554900105FF0800175D7E3FFEFBD700",
INIT_34 => X"000005010495B7AE921C517DE10FFDF50482A2DB6AB45FFD56DBD7087BEAA384",
INIT_35 => X"0FFF1C017D140410400BE8E28A10AAA085082550A1057DBE803AE38145B78FD7",
INIT_36 => X"000000000000000000001C556FA00A2A0800BAE3F1C0092EBAAADB6D080A1241",
INIT_37 => X"4AA0800020BA550028B550855400AAF7AEBDFEF0000000000000000000000000",
INIT_38 => X"7400AAAE975EFA2FBFFF55FF84000AAAAFBC0145002AA8AAAAAFFC2000AAAA97",
INIT_39 => X"E8B55085142010AAD157545F7AEA8B55AAAE821EFAAFBEAB55F7AAA8A00AA841",
INIT_3A => X"417555AAFFFDF450804020AA557BFFE10A2FFFFFEFF7D568ABAA2FFC00105D7B",
INIT_3B => X"D17DF45007FE8AAA08002AAAAA2AA955FFFF80020BAAAAA975450800001EF080",
INIT_3C => X"7802AABA5D7FEAB45080015410007FEAA0055517DE00FFFBC2000AAFBE8B55F7",
INIT_3D => X"A2AEBFFEF082A82010FFD5421EF5D0000010F7AAA8A10AA8017400552A801EFF",
INIT_3E => X"00000000000000000000000000000000000005D557FE00A280020BAAAD140000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_4,               -- Port A enable input
WEA      => wbe_a_hi_1024_4(1),               -- Port A write enable input
DIA(0)   => data_write_a(15),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_4(15),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_4,               -- Port B enable input
WEB      => wbe_b_hi_1024_4(1),               -- Port B write enable input
DIB(0)   => data_write_b(15),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_4(15),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_16_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"DA22C618B1000482B688B186588884862A400438255FC38381441205BA803003",
INIT_01 => X"7045A80028404C211203A952A90341080B173340412000E1005D628000820484",
INIT_02 => X"428406A4000850848330118D0AAC55001349B108818005460229044001C01784",
INIT_03 => X"092C4020000500020000500986812C405000001A48202050000A214AC0650115",
INIT_04 => X"4804A55440256F504025E003A054F46415A4E62B6FE3307943965A00001A1152",
INIT_05 => X"0000001C40A5B950ADB8EA097057ECE14C86D2B7F85AAD17F4B100000B88148C",
INIT_06 => X"415401DCDCF2C0A8030140BCB0820A200342A1C641C1E8782F508F2B00003584",
INIT_07 => X"002701881A3202080AE00480A2002840BE1480FA004342AA6F12000054004867",
INIT_08 => X"08C54828091002000002B32A8C19064E486A8001510000014140C1E2A14891E0",
INIT_09 => X"015452B103020814004088B64102680B6596594800400413CAC0208944800000",
INIT_0A => X"96AA000484094C000000000000012C9000A0000D0A80000BF8028E87C1B99270",
INIT_0B => X"014808A02004200E540480212000A448C0082024AE50064B44000000000002A2",
INIT_0C => X"0004000D5846256AAEA811150445411150445411150445411150422A088A8200",
INIT_0D => X"00000004010042A204A0C5817D00005034052E40000817D00440004004AD3240",
INIT_0E => X"632B2673FA4587978A2004102800809225545155121740000004900090000000",
INIT_0F => X"00C6564CE7F4EA4B940076D296D003030800462CBD320018CAAAACFE9164C800",
INIT_10 => X"28834ADB1440A114793A4A30A40839AA14910D08DCB2640031955559FD3AC990",
INIT_11 => X"594AB0B1A025371CA0E034E8443C097A800EB090D4AAC91208ED2FA0CE5E09B1",
INIT_12 => X"7B50446083001B94BB38C540EBE61284BB304880E3E4579EDC00992980D58033",
INIT_13 => X"5511121840E7A2CD952ECC12ABC3E6ACB3DFB12ECE315000F61FF1727A85FDBC",
INIT_14 => X"75DEB07F6F2E7084517F126F8395CB2BEFBAB8BA8AF698228CC5E2F08ECA5159",
INIT_15 => X"5580A840A8009F8B108C80A1021B080AFC0DF6422C6077F4A77F20D0C0E21084",
INIT_16 => X"0000000000000000000000000000000000044000102A0001148442A110810359",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"558D11544C690DA64C1C4F68A360400000000000000000000000000000000000",
INIT_1A => X"14D14D14D14D14D14D14D14D14D14D14D14514514514514529E5F87869E79E78",
INIT_1B => X"D1E8F47A3D1E8F47A7D3E9F4FA7D3E9F4FA7D3E9F47A7D1E9F47A7D1E9F4D14D",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000007D3E9F4FA7D3E8F47A3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"C00AA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"03DFEF085155400F78428BEF087FFFFEFF7D168B55AAD17FFFF552EBFE00007F",
INIT_29 => X"2E975EFF7D568BFFFF80175EF0004000BA552A821FFFF8000010082A954BA000",
INIT_2A => X"55540000082EAABFFA2FBE8B55A2AE80000F7D5555555D2AAAABAAAD1420BA5D",
INIT_2B => X"A2FBE8BEFA2843DE00AA8015400FF84001EF0000020AA5D00154005D043FF455",
INIT_2C => X"FA2802ABEF557BEABEF5D0415410087FD74BAAAAEBFFEF557FC00AAF7AE95555",
INIT_2D => X"FFFFAABFEAAFF84001FF002A821FFAAD5554BA087FFFF55557BD54AAF7FBC01F",
INIT_2E => X"000FFFBE8BFF0800174AA557BFDE10A2FBEAB45F7D56AABA082A97545F7D16AB",
INIT_2F => X"FFEF552AB8E38087FC2092000000000000000000000000000000000000000000",
INIT_30 => X"070280024904AA1C0438FD7005150438F78A2DBFF0871F8FC7E3D56AB6DBEDB7",
INIT_31 => X"AA8ABAAADB400924920925EFF7D16ABFFE38E175EF1400000BA412E871FFE38E",
INIT_32 => X"0A1240055003FF6D5551420101C2EAFBD7A2FFEDB55B6A080038E3DB50555412",
INIT_33 => X"57FC00BAE3AA9257DA2FFE8BC7BE8E38E10A28017400E38A051FF0804050BA41",
INIT_34 => X"4971D0492E3F1C71C7BE8A2ABD74975EDBC7550E12410087FD74AAB6AABFFC75",
INIT_35 => X"A08249756DF7D168BC7F7AABAEAAF780051C70824851D7A2DB50482147FFAF55",
INIT_36 => X"00000000000000000000E3FFEFBD70000124AA557FFDE10A2FBEDB6DF7D16AAB",
INIT_37 => X"B55A2D16ABEFFFFBFDFFF552AAAAAA007BC00000000000000000000000000000",
INIT_38 => X"20AA002A955EFAAAA974AA0800020BA550028B550855400AAF7AEBDFEF08516A",
INIT_39 => X"000AAAAFBC0145002AA8AAAAAFFC20000000021EFF7D568BFFA2AA955FF5D040",
INIT_3A => X"E975EF0800174BA002E820105D003DFEF5D51420005D2ABFF45A2FBFFF55FF84",
INIT_3B => X"7BD74AAF7AEBDF455D7BC20BAAAAE821EFAAFBEAB55F7AAA8A00AA8417400AAA",
INIT_3C => X"2FFC00105D7BE8B55085142010AAD157545F7AEA8B5500557DF45552A8200000",
INIT_3D => X"A2FFFFFEFF7D568ABA0804155FFF7D568B55FFAAAAABAFF8415545000015555A",
INIT_3E => X"0000000000000000000000000000000000000AAFFFDF450804020AA557BFFE10",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_4,               -- Port A enable input
WEA      => wbe_a_hi_1024_4(2),               -- Port A write enable input
DIA(0)   => data_write_a(16),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_4(16),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_4,               -- Port B enable input
WEB      => wbe_b_hi_1024_4(2),               -- Port B write enable input
DIB(0)   => data_write_b(16),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_4(16),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_17_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"5284CE4FB7BD2C8994A13392DBD02E14006B82AC7E800D44D3DD2FD5F9B961C0",
INIT_01 => X"2EACD01F7E03FC6793F2199B39FC233C11D93AE6F3BB92B32091DBC339B24542",
INIT_02 => X"E63CCCC00A82C08092A2AFAE667033DB50853379C10BFDC5C6F4044443C817C6",
INIT_03 => X"7FF183635AEF9E3635AEF9E18E237040404446965C0607EE6DB7854AC4DE060C",
INIT_04 => X"D78AC33FB604488B000892EF17BE6D84196482236FE100294152E294350FB697",
INIT_05 => X"081B5F9B409420D0CDB47A05403F6CE0C08A4AB7F840EDB6F48100DFC8081081",
INIT_06 => X"768465354781CBC30316367077B4BDB50646E8D87100A8201ED01C19C020F71A",
INIT_07 => X"4002A110C922480A82D0841147162C48EBB9537A0022DC67987042EE976ABEA7",
INIT_08 => X"DB931BFEF91C00002CC0E019C0C82A4E4820C15A2330E004401891181168C4D1",
INIT_09 => X"09F3A1BC11EFBC66DB65307071477FF1030C397C060B4254064302042F803A69",
INIT_0A => X"3F330802162F3B7EE3F3EC7C7DEF207000F00059D2ED56D7EED2ED3C9A867DC0",
INIT_0B => X"185C44B91BC1740B7605040BE0018CFC7429F326B9E822FFC00074D5A0AB033A",
INIT_0C => X"00367A28FC1B7F7FEFFCFBFF3EFFCFBFF3EFFCFBFF3EFFCFBFF3EFFE7DFF9E00",
INIT_0D => X"0000000008004BA78428C7AD7FC94B533F5B4FFBD2FAD7FCCA786D43FE67C218",
INIT_0E => X"BA494CEBFD4F2667ABB6F68B29760593F33FA0CF170F40006001B1A05C000000",
INIT_0F => X"7F749299D7FAEB237DFE5865B6D2BF23265CBACE542A6FEE92333AFF33E0A9BF",
INIT_10 => X"F6C24B6D18C3C9F8E2881F3F787D776B5DB94A09955054DFDD246675FE7AC153",
INIT_11 => X"BFB349E08FF9A27EDE9FA8AEFD9E7467BFCB195CFEB56A1A70D34D1706FFFA3E",
INIT_12 => X"6FE219CA80725B875EED723FF7FCB2875EDAAFEAF7FD929BFD55BBC71D79F639",
INIT_13 => X"546670D018E7A6E581D7B6AB75FDFCECA6E581D7BB5DDFC6FF0EB7D7E859FDB5",
INIT_14 => X"B978177F6D6AF5ECDB5FB76A5F5FA165B456E0FB308710C49FCFB741598B9C7E",
INIT_15 => X"CFDAAB00AC00A8BBFC8B501CF7A0FED9A540EA1952586CEB54D143ACFF9A3BA9",
INIT_16 => X"000000000000000000000000000000000026E100002F382DBD9ECFE117805F20",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"4372003009EDCC4052E917114F981800C0000000000000000000000000000000",
INIT_1A => X"BA69A69AEBA69AEBA69A69AEBA69AEBA69A69A69A69A69A68698686981D75D74",
INIT_1B => X"6A351A8D46A351A8D068341A0D068341A0D068341A0D46A341A0D46A341A69AE",
INIT_1C => X"FFFFFFFFFFFFFFF80000000000000000000000000000046A351A8D46A351A8D4",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"7FEAA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"17FFFF552EBFE00007FC00AA087FFFFFFFFFFFFFEFF7FBEAB450804001EFAAD5",
INIT_29 => X"D168A000004020AA5D7BE8B450051401EF087FD74AA087FFFFEFF7D168B55AAD",
INIT_2A => X"D7FEAB55FF80175EFFF8000010082A954BA00003DFEF085155400F78428BEFAA",
INIT_2B => X"F7D568BFFFF80175EF0004000BA552A821FF5D00020BA552A82000552A821555",
INIT_2C => X"AAAD1420BAFFFFFDF45AAD17FFFFAAFBC01EF5D0015555557BFDEBA5D2E975EF",
INIT_2D => X"BA007FEABEF005555555A2D1554BAA2FBE8B55A2AE80000F7D5555555D2AAAAB",
INIT_2E => X"0000000020AA5D00154005D043FF45555540000082EAABFF00516AA10552E820",
INIT_2F => X"8B550000071EFB6DF7AE92000000000000000000000000000000000000000000",
INIT_30 => X"F8FC7E3D56AB6DBEDB7FFEF552AB8E38087FC2092147FFFFFFFFFBFDFC7EBF5E",
INIT_31 => X"150438F78A2DBFFBED16AA381C0A07082497FEFB6D1451471EF007BD04920871",
INIT_32 => X"2A850105D2A80155417BEFB6DEB8E175FFE38E070280024904AA1C0438FD7005",
INIT_33 => X"D7BFAEBA4920925EFF7D16ABFFE38E175EF1400000BA412E871FF550A0009249",
INIT_34 => X"E3DB50555412AA8ABAAADB40092FFF5FFF6DAADF7FFD7B6F1C71EF55001756D5",
INIT_35 => X"7145B6AA28492487082007FEDBD700515556DA2DF50492A2FFEDB55B6A080038",
INIT_36 => X"000000000000000000000804050BA410A1240055003FF6D5551420101C2EAFBD",
INIT_37 => X"FEFF7FBFFF55A2D16AB550000175EFFFFBEAA000000000000000000000000000",
INIT_38 => X"55EF087FC200008516AB55A2D16ABEFFFFBFDFFF552AAAAAA007BC0000557FFD",
INIT_39 => X"020BA550028B550855400AAF7AEBDFEFF7D568AAA5D2A97410007BFFFFF55515",
INIT_3A => X"A955EF5D2E80010002A954005D2A82155087FFFFEFAAAA975EFAAAA974AA0800",
INIT_3B => X"D1575FF5504175EF5D7FEAAAA0000021EFF7D568BFFA2AA955FF5D04020AA002",
INIT_3C => X"2FBFFF55FF84000AAAAFBC0145002AA8AAAAAFFC2000FFD57DFFFAAFFFDF55FF",
INIT_3D => X"5D51420005D2ABFF45557FE8AAA000415410007BFFF450051555EFA2FBC0000A",
INIT_3E => X"00000000000000000000000000000000000000800174BA002E820105D003DFEF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_4,               -- Port A enable input
WEA      => wbe_a_hi_1024_4(2),               -- Port A write enable input
DIA(0)   => data_write_a(17),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_4(17),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_4,               -- Port B enable input
WEB      => wbe_b_hi_1024_4(2),               -- Port B write enable input
DIB(0)   => data_write_b(17),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_4(17),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_18_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"69844019080000A21A611406840014122A641074155FC28A2024001001801003",
INIT_01 => X"7443D920034004180005E9E3C90360C0041C0181002001602025800008440084",
INIT_02 => X"E2DCCCE61D5C008103F2000781FC0FEDEAC2161B0B8FB0008620044443006010",
INIT_03 => X"884E300802006900802006995C896D605200000856E24A040000640052141103",
INIT_04 => X"480520FC026125AC0025C9122644E3E40EC8E2001001302281841A009038A86A",
INIT_05 => X"432000040089983070019400F01010004C8DB841405A80A100B586200FAC24AE",
INIT_06 => X"09044359DC7040000000002C109B0E0A00A1104641C0803804000707284600E1",
INIT_07 => X"400D10100400481D5EB08501620000007500CE801241021FE78E404860140060",
INIT_08 => X"00880C0106A0528020019307CC082A0A4A6A01ED725021400040D028000A9729",
INIT_09 => X"00117063038000282081402E4106400B6186128040600C10C1C0200950508110",
INIT_0A => X"C0C30C2E21580C874004008080003C32A10A19090C02010E1022944061688000",
INIT_0B => X"0180A8062026000DC425C0301311324AA2373088479105D044A1022000001835",
INIT_0C => X"0D89844703649000000200000000000000000000000000000000000000000010",
INIT_0D => X"0D8306C182701404C1973010802020404084001E00010802046092B5001FB365",
INIT_0E => X"528EB314068AB8B803DB00002900800400FC503F08180050942E4200020C1B06",
INIT_0F => X"40A51D66280D6032C5F96D3C51555D5D7D5AA87285820814A3CCC501C2A60820",
INIT_10 => X"8B35A3FEBF1FEDFD9C2B30E0468AAAD5D48F37E8FC1304102947998A03984C10",
INIT_11 => X"440FE1DD772D37A0A321BC6968F32658BF2D4F2A80BF8FE3F9FE3AC362080529",
INIT_12 => X"5487910D7E5A6D961A28456A1832E5161A100DD5182BC54020EA67A189C6ED36",
INIT_13 => X"AA444CAF91EDD1B725868403BE06323551B725868A100ABD119753B70964122B",
INIT_14 => X"EDC259048ACD868EE3803D65CEDC258A8F80D55E007C3F8EBB56F4C5362C978F",
INIT_15 => X"3F240014BE84370001B6922070440556B15F7FABBC0031BCF2257C41634B14D4",
INIT_16 => X"C1B06C1B06C1B06C1B06C1B06C1B06C1B0491069068000004060300A005A0118",
INIT_17 => X"1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06",
INIT_18 => X"B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C",
INIT_19 => X"B28BBECEB80EE173C2300F7DF16000000000000000000000000041B06C1B06C1",
INIT_1A => X"8A28A28AAAAAAA28A28A28AAAAAAA28A28A28A28A28A28A2910591505C104104",
INIT_1B => X"28944A25128944A25128944A25128944A25128944A2552A954AA5128944AAAA2",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000128944A25128944A251",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"9540000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"BEAB450804001EFAAD57FEAA087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974BA082E",
INIT_29 => X"7FFFFFFFFFBFDF45AAD568B55080028B55002E82000087FFFFFFFFFFFFFEFF7F",
INIT_2A => X"0043DE10AA843DE00087FFFFEFF7D168B55AAD17FFFF552EBFE00007FC00AA08",
INIT_2B => X"0004020AA5D7BE8B450051401EF087FD74AAAAFFFDF45A2D16AB55F7FFFFFFF0",
INIT_2C => X"0F78428BEFAA80000000804154BA55042ABEF5D7FD75FFAAD540145AAD168A00",
INIT_2D => X"00082E95555085168A10557FD7545FF8000010082A954BA00003DFEF08515540",
INIT_2E => X"0005D00020BA552A82000552A821555D7FEAB55FF80175EF5D00020105D2A974",
INIT_2F => X"DFFF5D2A954AA082A92428000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFBFDFC7EBF5E8B550000071EFB6DF7AE921C7FFFFFFFFFFFFFFFF7FBF",
INIT_31 => X"AB8E38087FC2092087FFDFC7E3F1FAF55A2DF6DB7D1C002AB7D002A82028147F",
INIT_32 => X"DF6DB7DE3F5FAFC708003DE28B68E38E280871F8FC7E3D56AB6DBEDB7FFEF552",
INIT_33 => X"ADF4516DBED16AA381C0A07082497FEFB6D1451471EF007BD0492B6F1F8F55AA",
INIT_34 => X"1C0438FD7005150438F78A2DBFFA28407038140410492550A2ABC7497BD25FFA",
INIT_35 => X"F5D0E05000492097428002E9557D1C516FA28417BD5545E38E070280024904AA",
INIT_36 => X"00000000000000000000550A00092492A850105D2A80155417BEFB6DEB8E175F",
INIT_37 => X"FFFFFFFFDFEFF7FBFFFEF552E974AA082A820AA0000000000000000000000000",
INIT_38 => X"ABEF002A800AA557FFDFEFF7FBFFF55A2D16AB550000175EFFFFBEAA00557FFF",
INIT_39 => X"6ABEFFFFBFDFFF552AAAAAA007BC0000087BFDF45AAD568B55AAFBFDFEF55042",
INIT_3A => X"FC2000FFD56AB45A2FFFDFFFAAD16AB4500043DEAAFFAEAAAAA08516AB55A2D1",
INIT_3B => X"2AA8B45087FC01EFA2FFD55EFF7D568AAA5D2A97410007BFFFFF5551555EF087",
INIT_3C => X"AAA974AA0800020BA550028B550855400AAF7AEBDFEFA280154BA55040000055",
INIT_3D => X"087FFFFEFAAAA975EF5D2E974000804154BA082A975EF5D517DEAA007BD5545A",
INIT_3E => X"00000000000000000000000000000000000005D2E80010002A954005D2A82155",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_4,               -- Port A enable input
WEA      => wbe_a_hi_1024_4(2),               -- Port A write enable input
DIA(0)   => data_write_a(18),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_4(18),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_4,               -- Port B enable input
WEB      => wbe_b_hi_1024_4(2),               -- Port B write enable input
DIB(0)   => data_write_b(18),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_4(18),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_19_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"042200000000000041088001001AA00000000000000000000000500802000003",
INIT_01 => X"040048000024000000000404000000000A22000800000800004A200000000001",
INIT_02 => X"200C8840085EB00480060000001C008002489E0F000405EA0004040404000000",
INIT_03 => X"24004000000000000000000900002C4050000000000069500208400002E14100",
INIT_04 => X"4800200C0000000044002000C80020E40000E200000130200188000000800100",
INIT_05 => X"000000000080181000000000701000004C8000000058800000B1000009880480",
INIT_06 => X"80500081081040000000002C100040400000004641C080380400070100000000",
INIT_07 => X"4020109801A4CE005C00048380142810010564C4100114012002402028044808",
INIT_08 => X"0070700000000000000083004C3902420062000020E0000100004082A140102B",
INIT_09 => X"001150200000000000000026400000016186100000000010C04002C000000000",
INIT_0A => X"007C00008082C0002000000000002C3000000004050001030102040000000000",
INIT_0B => X"0000000000000000000000000000010000800011000000000000000000000BC0",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"000000000000000000000000000000042000760000000000000000010004B200",
INIT_0E => X"0D74002280300F0002FB069040000060000C5003000800000000000000000000",
INIT_0F => X"C01AE8004500744C780687DBA828008080A5FC0D385598035D0008A00C015660",
INIT_10 => X"39D8140040201BF861F0E7D693E6170022408116DFE0AB3006BA0011401D02AC",
INIT_11 => X"5412E4997F5249FD005043B8680CC98F00D0F2DD0140100406FE053A98F6ECC7",
INIT_12 => X"7418663001858040E153888000010840E165D0000000285C246A181C03FE4662",
INIT_13 => X"8199830066F0020858385974000001260208583854E2200000660208D6B1423F",
INIT_14 => X"8235AC508FCE8811042040F008235AE04420C040CF00C031C80009B8F224978B",
INIT_15 => X"030004E00000C220010808C10D9A92A74CD7CF4A09051110AD5A3C9200B7F280",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000118",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"07208BBA3F0C7010C660C7441920000000000000000000000000000000000000",
INIT_1A => X"861869A61861861861869A61861861861861861861861861A8208C4C1534D34C",
INIT_1B => X"984C26130984C26130984C26130984C26130984D26930984C26130984C261861",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000984C26130984C26130",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"174BA00000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFDFEF5D2A974BA082E95400F7FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0004",
INIT_29 => X"FFFFFFFFFFFFFFFFF7FBFDFFF552E974BAA2FFFFE10087FFFFFFFFFFFFFFFFFF",
INIT_2A => X"004001EFAAAEA8ABA087FFFFFFFFFFFFFEFF7FBEAB450804001EFAAD57FEAAF7",
INIT_2B => X"FFFBFDF45AAD568B55080028B55002E82000F7FFFFFFFFFFFFDFEFA2D568B550",
INIT_2C => X"0007FC00AAF7FFFFFFFF7FBE8B55AAD16ABEF5D2ABFF55080402010087FFFFFF",
INIT_2D => X"55A2FFFDFEF5D2EBFE00AAFFFFEBA087FFFFEFF7D168B55AAD17FFFF552EBFE0",
INIT_2E => X"000AAFFFDF45A2D16AB55F7FFFFFFF00043DE10AA843DE00557FFDFEFA2D16AB",
INIT_2F => X"FFEF552A974AA0000104AA000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFF7FBFDFFF5D2A954AA082A92428E3FFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"0071EFB6DF7AE92EBFFFFFFFFFFFFDFEFF7F5FAFC7492A974AAB6F5F8E101C7F",
INIT_32 => X"F1F8FD7AAD16AB450000001FFBEA4A8AAA147FFFFFFFFFBFDFC7EBF5E8B55000",
INIT_33 => X"00000010087FFDFC7E3F1FAF55A2DF6DB7D1C002AB7D002A82028FFFFFFFEFF7",
INIT_34 => X"BEDB7FFEF552AB8E38087FC2092F7FBF8FC7E3F5EAB45B6DF6FBEF5D2AB8F7D0",
INIT_35 => X"84971F8FC7AAD56DB6DBEF5F8FD7412ABFE28B6F5F8E820871F8FC7E3D56AB6D",
INIT_36 => X"00000000000000000000B6F1F8F55AADF6DB7DE3F5FAFC708003DE28B68E38E2",
INIT_37 => X"FFFFFFFFFFFFFFFFFDFEF552E954AA0004000AA0000000000000000000000000",
INIT_38 => X"54AAF7D568A00557FFFFFFFFFFFDFEFF7FBFFFEF552E974AA082A820AAA2FFFF",
INIT_39 => X"FFF55A2D16AB550000175EFFFFBEAA00A2FFFFFFFF7FBFDFFFFFD568B55002A9",
INIT_3A => X"A800AAF7FBFDFEFF7D56AB45AAD56AB450004001EFFF842AAAA557FFDFEFF7FB",
INIT_3B => X"FFFFFFF552AA8BEF080402000087BFDF45AAD568B55AAFBFDFEF55042ABEF002",
INIT_3C => X"8516AB55A2D16ABEFFFFBFDFFF552AAAAAA007BC0000FFFBE8B55AAD168B55F7",
INIT_3D => X"00043DEAAFFAEAAAAA08556AB55A2D57FFFFF7D568B45002ABDEAAFFD16AA000",
INIT_3E => X"0000000000000000000000000000000000000FFD56AB45A2FFFDFFFAAD16AB45",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_4,               -- Port A enable input
WEA      => wbe_a_hi_1024_4(2),               -- Port A write enable input
DIA(0)   => data_write_a(19),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_4(19),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_4,               -- Port B enable input
WEB      => wbe_b_hi_1024_4(2),               -- Port B write enable input
DIB(0)   => data_write_b(19),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_4(19),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_20_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000003",
INIT_01 => X"F55FF80000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"E05022020800008400F655001FFCFF80018FA804400000000000004400000001",
INIT_03 => X"00000000000000000000000900002CC07000000000000000000000000000013F",
INIT_04 => X"68002FFE40900010000180000001FFEC0012EE0C001370F40780000000000000",
INIT_05 => X"0840000880FCBBF0100E204DF0F88311DD8005080679800000F3000029980580",
INIT_06 => X"001000030817C8E8840155FDF9001001050023F6C3C3D0F87FA19F7F011000E4",
INIT_07 => X"000000090492260800008000EE00000000000000002101FF2002C00000004018",
INIT_08 => X"2A040001071004000013FF7FCA302C0C0008214800002101554031F800000000",
INIT_09 => X"801F57F200000090000489FEC0000001EFBEF0040008023FDFC0000000004006",
INIT_0A => X"0000000008000000000000000000ADF000000200000008000008028300110230",
INIT_0B => X"0000000000000800080000000000000000000000000000000800800A40000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"000000040900005C848538000020000000800000080000020000800101FFB600",
INIT_0E => X"00800000003A010003000000000000600FFC53FF001800000002004080000000",
INIT_0F => X"0001000000007408040000004000000004E9000008020000200000000E800800",
INIT_10 => X"00200000000313100010002000008000000000129600040000400000001D0010",
INIT_11 => X"81C012060000000000218F7840000100800004000000000066C0000080080000",
INIT_12 => X"800000000017C000100000000001A800080000000001A8040000002840008185",
INIT_13 => X"0000000006F00000100200000000012600001004000000000066000000801040",
INIT_14 => X"0000200410100000000005F00000020080090A0000000085C800002000586000",
INIT_15 => X"FF00400000000000020020020001000040283024E4F2860400008000030ED080",
INIT_16 => X"00000000000000000000000000000004010201001003020200000000000127DB",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"A0700030038200010089120104D2040020000000000000000000000000000000",
INIT_1A => X"2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2C30C30C30C30C306982121A1E79E79",
INIT_1B => X"32190C86432190C86432190C86432190C86432190C86432190C86432190CB2CB",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000432190C86432190C864",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0201000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF552A974AA0004174BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA0804",
INIT_29 => X"7FFFFFFFFFFFFFFFFFFFFFFEF552E954AA000400000F7FFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E954BA007FC00BA087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974BA082E9540000",
INIT_2B => X"FFFFFFFFFF7FBFDFFF552E974BAA2FFFFE10FFFFFFFFFFFFFFFFFFFFFBFDFFF5",
INIT_2C => X"FAAD57FEAA007FFFFFFFFFFFFFEFF7FBFFF550800020BAAAD56AAAAF7FFFFFFF",
INIT_2D => X"EFF7D56AB450000021EFA2D57DE10087FFFFFFFFFFFFFEFF7FBEAB450804001E",
INIT_2E => X"000F7FFFFFFFFFFFFDFEFA2D568B550004001EFAAAEA8ABA5D7FFFFFFFFFFFDF",
INIT_2F => X"FFFF5D2E954AA080005000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFEF552A974AA0000104AAFFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"A954AA082A92428087FFFFFFFFFFFFFFFFFFBFDFEF5D2E974AA000A07000E3FF",
INIT_32 => X"FFFFFEFF7FBFFFFF552E974AA0071C50BA1C7FFFFFFFFFFFFFFFF7FBFDFFF5D2",
INIT_33 => X"EDF6FABAEBFFFFFFFFFFFFDFEFF7F5FAFC7492A974AAB6F5F8E10E3FFFFFFFFF",
INIT_34 => X"EBF5E8B550000071EFB6DF7AE921C7FFFFFFFFFBFDFEFE3F5F8F450004050AAB",
INIT_35 => X"A497FFFFFFF7FBF8FC7EBD168B450804021FFB6D57DE28147FFFFFFFFFBFDFC7",
INIT_36 => X"00000000000000000000FFFFFFFEFF7F1F8FD7AAD16AB450000001FFBEA4A8AA",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2A954AA0800174100000000000000000000000000",
INIT_38 => X"74AA002E95410A2FFFFFFFFFFFFFFFFFFFFFDFEF552E954AA0004000AAFFFFFF",
INIT_39 => X"FDFEFF7FBFFFEF552E974AA082A820AA087FFFFFFFFFFFFFEFF7FBFDFFF5D2A9",
INIT_3A => X"568A00AAFFFFFFFFFFBFDFEFFFFFFDFEF5D2E954AA0051554BA557FFFFFFFFFF",
INIT_3B => X"D16AB450804174AAFFFFFFEBAA2FFFFFFFF7FBFDFFFFFD568B55002A954AAF7D",
INIT_3C => X"57FFDFEFF7FBFFF55A2D16AB550000175EFFFFBEAA005D7FFFFEFF7FBFDFFFAA",
INIT_3D => X"0004001EFFF842AAAA087BFDFEFF7FFEAB45A2D568B550804001EFF7D57DEBA5",
INIT_3E => X"0000000000000000000000000000000000000F7FBFDFEFF7D56AB45AAD56AB45",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_4,               -- Port A enable input
WEA      => wbe_a_hi_1024_4(2),               -- Port A write enable input
DIA(0)   => data_write_a(20),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_4(20),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_4,               -- Port B enable input
WEB      => wbe_b_hi_1024_4(2),               -- Port B write enable input
DIB(0)   => data_write_b(20),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_4(20),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_21_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"4A302428B824900A128C090A5C1800261500213C005FE812D10420054085A202",
INIT_01 => X"001FFE3440B609703B0427F801A40B8115BC4F655300340288A40D30040E4DD8",
INIT_02 => X"E00424256888D8819801000F9FFFFFFFF149FF1FCA448046C60A0D2437C517F9",
INIT_03 => X"20030640003250640003250F06002CC1740002019824E001CD357832440001FF",
INIT_04 => X"EA2C3FFD400006E04401A8837001FFFC004AEF00080B70E08FB5789421007C5C",
INIT_05 => X"00011A0C40F9FFF80920954FF0F00809DF84A0202879800000F3000029980780",
INIT_06 => X"0805984B7A1FC0A0000101FFF0480080002281F7C3C381F87C03DFFF00009004",
INIT_07 => X"B424068086A205481A60A19000908204A855B000A08A61FF20C3D004D331D340",
INIT_08 => X"1BFA0001600802000023F7FFC08D234B40C2028253000040114200000D0226C0",
INIT_09 => X"EF1F5FF054096C6ADBA169FFC202B1C1FFBEF0440021083DFFCE22DC2880E24D",
INIT_0A => X"45FF0C004041D84862A28C54518DBFF00020004C0A6044901112A0908AA0A300",
INIT_0B => X"018C241102068006C620C03882019480E63180855A492712CC01C49C20201BFE",
INIT_0C => X"08A9464116544302C02D92236488D92236488D92236488D922366446C911B210",
INIT_0D => X"08800444021048034004001890000806002804A0822189000900D80621FFBE00",
INIT_0E => X"060580261013813A2CC396506102C4053FFD5BFF00A04A00200602CA52001100",
INIT_0F => X"080C0B004C202621A85C09411500135844C196D3606941018150098404C1A304",
INIT_10 => X"B02901013416181C96C2C9C600890A2028172192C460D1820302A0130809834A",
INIT_11 => X"9C5E803408250180AC268D185DB3F4350B811068C00049A0A4AA68F05C96A001",
INIT_12 => X"002C006560138F032B1804101244C883052208209040CC849063A747512B7678",
INIT_13 => X"41401E240665750440C9488280254530314080C2C601040420352148A00501B1",
INIT_14 => X"500811204D000700114204A70422016149916011008CAA8858850B00C32591C0",
INIT_15 => X"FFC06E60AC0496022300233104663040808E991765205000070121D41D18D098",
INIT_16 => X"40100401004010040100401004010040102090010008000001C0E010020007DF",
INIT_17 => X"0100401004010040100401004010040100401004010040100401004010040100",
INIT_18 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_19 => X"FFEF9FEEFF7FFDF7FF3E3DFDF7E0000000000000000000000000401004010040",
INIT_1A => X"BEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBFFDFDFFFCF3CF3F",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFEFF7FBFDFEFF7FBFDFEFBEF",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000FFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0001000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E954AA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0004",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA0004154BAFFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"52E974BA0804000AAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0004174BAFF",
INIT_2B => X"FFFFFFFFFFFFFFFFEF552E954AA000400000007FFFFFFFFFFFFFFFFFFFFFFEF5",
INIT_2C => X"A082E95400007FFFFFFFFFFFFFFFFFFFFDFEF5D2E974BA002E97400007FFFFFF",
INIT_2D => X"FFFFFBFDFEF5D2A954AA002E974BA087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFBFDFFF5D2E954BA007FC00BA5D7FFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA000002000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080005000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"A974AA0000104AAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974BA0000174AAFFFF",
INIT_32 => X"FFFFFFFFFFFFDFEF552E954BA080A000AAE3FFFFFFFFFFFFFFFFFFFFFFFEF552",
INIT_33 => X"02A95400087FFFFFFFFFFFFFFFFFFBFDFEF5D2E974AA000A07000007FFFFFFFF",
INIT_34 => X"F7FBFDFFF5D2A954AA082A924281C7FFFFFFFFFFFFFFFFFFBFDFEF5D2A974BA0",
INIT_35 => X"A557FFFFFFFFFFFFFFFF7FBFDFFF552E974BA0020924BA1C7FFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000E3FFFFFFFFFFFFFFEFF7FBFFFFF552E974AA0071C50B",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0000020000000000000000000000000000",
INIT_38 => X"74BA0000174BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954AA080017410FFFFFF",
INIT_39 => X"FFFFFFFFFFDFEF552E954AA0004000AAF7FFFFFFFFFFFFFFFFFFFFFFFEF552A9",
INIT_3A => X"E95410087FFFFFFFFFFFFFFFF7FBFDFEF5D2A954BA082E800AAA2FFFFFFFFFFF",
INIT_3B => X"FBFFFFF552E954BA002E97410087FFFFFFFFFFFFFEFF7FBFDFFF5D2A974AA002",
INIT_3C => X"57FFFFFFFFFFFDFEFF7FBFFFEF552E974AA082A820AA557FFFFFFFFFFFFFEFF7",
INIT_3D => X"5D2E954AA0051554BA5D7FFFFFFFFFBFDFEFF7FFFFFEF5D2A974BA0000020AA5",
INIT_3E => X"0000000000000000000000000000000000000AAFFFFFFFFFFBFDFEFFFFFFDFEF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_4,               -- Port A enable input
WEA      => wbe_a_hi_1024_4(2),               -- Port A write enable input
DIA(0)   => data_write_a(21),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_4(21),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_4,               -- Port B enable input
WEB      => wbe_b_hi_1024_4(2),               -- Port B write enable input
DIB(0)   => data_write_b(21),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_4(21),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_22_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"5290F4CDE914905A14A43D33F488243E17122300F55FEB189B343A1140548380",
INIT_01 => X"A54007B259F6A975386262000C344BA9573C6FF57B18A5FB0ABFCD3C2C5F4F0C",
INIT_02 => X"021DFF8C38B3C009D203551040030071869D0040180AA2DC53DB89BEA8204001",
INIT_03 => X"2603475A969D0475A969D0460EAA401005111011BD506954EDB40F5EF41434C0",
INIT_04 => X"922D9002100ED69E443D988B0D5400103E48003D0800011E803B06B5B9125A15",
INIT_05 => X"281B5A0C06000408F4DF9422010D8802022F2124A8022492580040440002021C",
INIT_06 => X"F780C4C052881ADA0E05440205DA50930FA182010004700083E220800440B588",
INIT_07 => X"049D028B93FB561833D8094A02F5EA92FD7247E10305C40040D136E6A023F7FC",
INIT_08 => X"00028241680A0E002A9400803A884B5B5206B7C2E53CA25144009007A64EBD64",
INIT_09 => X"41008810240240C6694008010392354010000560141801002028A83D2A08E06D",
INIT_0A => X"34000000848BCA6902A29C54539C020E11810098D4067EFF9FF284D483E2AB41",
INIT_0B => X"500001840000C80B410014088040F4A944B1AA313C0022AA0011C0DC00028001",
INIT_0C => X"80B14004D158C8CA24A1C2A870AA1C2A870AA1C2A870AA1C2A872550E1543800",
INIT_0D => X"80A14050A01509E050854498B5281A1C34E506A2C6898B52A154DAC6B6000850",
INIT_0E => X"0B03001A483A4146603050080410089180008800143D83888281A2034A850142",
INIT_0F => X"A4160600349075238473F1210006133835E92273612B3482C090068A0E84AC56",
INIT_10 => X"30060181BA1B13959DC08DA902458870201970B29602562B0581200D141D0959",
INIT_11 => X"E042021C040D0152C8058B3840F044708E7E1C20A0106EA166C13AFC14AA3804",
INIT_12 => X"080E004B0C17C1439A9838301DC1A8438EA32C009DC1A8255300650458A1D588",
INIT_13 => X"018010E186F110A908E3A8CB0026C9A610A908E6A60F0807626610E160589C4C",
INIT_14 => X"2A701667334005800B1605F043858125E0D04110408D2485CA034681E43A1E40",
INIT_15 => X"00646002304244A91102C93A2D608D2A258DF8034188200C050171A41108F084",
INIT_16 => X"110441104411044110441104411044110466C440446CA06951D4EA8010009804",
INIT_17 => X"0040100401004411044110441104411044110441104411044110441104411044",
INIT_18 => X"0401004010040100401004010040100401004010040100401004010040100401",
INIT_19 => X"F7DFBFDEFE8FF1F7DEBDDF7DF7D05122890000000003FFFFFFFF900401004010",
INIT_1A => X"9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7BFFDFD7DDDF7DF7D",
INIT_1B => X"F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE79E7",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000003F9FCFE7F3F9FCFE7F3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA000400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0800",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000002000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2A954BA000015400FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080402010FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2A954BA0004154BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A0004174BAFFFFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0800154AAFFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF552A974AA0000174BAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974A",
INIT_2E => X"000007FFFFFFFFFFFFFFFFFFFFFFEF552E974BA0804000AAA2FFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080400010000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E954AA080005000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000402010FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2A954BA000417410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"804154BAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974BA0000174AAFFFFFFFFFFF",
INIT_34 => X"FFFFFFFEF552A974AA0000104AAE3FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0",
INIT_35 => X"AA2FFFFFFFFFFFFFFFFFFFFFFFEF552E954BA000E124BAE3FFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000007FFFFFFFFFFFFFFFFFFFFDFEF552E954BA080A000A",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804000100000000000000000000000000",
INIT_38 => X"54AA000400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2A954AA080017410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"0174BAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A954BA000415400FFFFFFFFFFFFF",
INIT_3B => X"FFFDFEF552E974AA0804174AAF7FFFFFFFFFFFFFFFFFFFFFFFEF552A974BA000",
INIT_3C => X"2FFFFFFFFFFFFFFFFFFFFFDFEF552E954AA0004000AAA2FFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2A954BA082E800AAAAFFFFFFFFFFFFFFFFFFFBFDFEF5D2E954BA002A820BAA",
INIT_3E => X"0000000000000000000000000000000000000087FFFFFFFFFFFFFFFF7FBFDFEF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_4,               -- Port A enable input
WEA      => wbe_a_hi_1024_4(2),               -- Port A write enable input
DIA(0)   => data_write_a(22),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_4(22),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_4,               -- Port B enable input
WEB      => wbe_b_hi_1024_4(2),               -- Port B write enable input
DIB(0)   => data_write_b(22),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_4(22),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_23_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"EF20906D902424807BC8241BC81801B97D38AD3C0800103362A6741C80A12A02",
INIT_01 => X"001FFF8409F089003B4422000D80C80106804A7951C5B9D1C828043EA28838F9",
INIT_02 => X"E01CEE21649C82C40800000F9FFEFF8E72CA7F5FC2E22809925A0D3611C877F8",
INIT_03 => X"24000400402670400402670D48222DC1764446838624000080007460C40001BF",
INIT_04 => X"68403FFC020560E0443E21037C01FFFC0002EE00628BF0E02FAD781014085014",
INIT_05 => X"0112000202FBFFF00920017FF0F0628BFF8488890979800002F702002BB807A0",
INIT_06 => X"EF85788B681FC000000001FFF0010000000001F7CBC385F87C0BFFFF20040001",
INIT_07 => X"F6E200000000C1440E3AE408009120071070FA07A1CB23FFA403F0C4D23BF7C0",
INIT_08 => X"0BF87CA400804000003FF7FFD8880A034AC09662305AB10555421006891A1089",
INIT_09 => X"BE1F5FEA10092C0896A243FFC0008087FFBEF2000000001DFFC612C0C0400100",
INIT_0A => X"41FF0C2060501000600000000001BFFA800808189A657EF81DD0C00079CC8001",
INIT_0B => X"018C24110A860006C620C0312241C482B20400CC52492710CC80060020A81BFE",
INIT_0C => X"0C08866907048320C20C10030400C10030400C10030400C10030400608018210",
INIT_0D => X"040002000041500300100040000500C000801000C02400000952800001FFBF04",
INIT_0E => X"FC850015385380380CDB86106502C5043FFD5FFF00A04BC010A7724B10000800",
INIT_0F => X"89F90A002A70A710A51C01C05904014861433602A1CAF13F2110055614C72FC0",
INIT_10 => X"E02D02001C1E14981B43253EE50C8220180F1082E06397E07E42200AAC298E57",
INIT_11 => X"8421802400A90022B0070FAE18019214A380344920080B21A58B02AC60BACDF0",
INIT_12 => X"0A2A000C480B0704B54028101AC49C84BB4100009AC49C80857A82D20CE8CB22",
INIT_13 => X"01E00C8103416445C12ED0400027C5292445C12D500B0005A62D344CB241D095",
INIT_14 => X"132C907425604680038706A35132C94BDD011010404428886AC91B11311C8280",
INIT_15 => X"FF000470BE0692020328CA0028042054A92771C50FC070110001C1680809591D",
INIT_16 => X"00802008020080200802008020080200800800200200000000000008004807DF",
INIT_17 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_18 => X"8020080200802008020080200802008020080200802008020080200802008020",
INIT_19 => X"0000000000000000000000000000000000000000000000000000008020080200",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080002010FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974AA000400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000400010FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974AA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080000010FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E954AA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954A",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA000015400FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080002010FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974AA000400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000402010FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E954AA080005000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA080407000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA00041741",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080000010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000402010FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2A954AA080002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954AA080017410FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"552A954BA000415400F7FFFFFFFFFFFFFFFFFFFFFFFFF552A954BA080015410F",
INIT_3E => X"0000000000000000000000000000000000000F7FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_4,               -- Port A enable input
WEA      => wbe_a_hi_1024_4(2),               -- Port A write enable input
DIA(0)   => data_write_a(23),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_4(23),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_4,               -- Port B enable input
WEB      => wbe_b_hi_1024_4(2),               -- Port B write enable input
DIB(0)   => data_write_b(23),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_4(23),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_24_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100600007FFF000080108004000800020000840041000080808",
INIT_02 => X"FC5CA803400EB8209000000F9FFEFF8E7240FF1FC22409EA04018E50074017F0",
INIT_03 => X"11100400000000400000000D00002CC07400000090C080019001010A000001BF",
INIT_04 => X"68003FFC00040000000000008001FFFC0002EE00000370E007A100000000E468",
INIT_05 => X"0000000000F8BFF00920004DF0F00001DF8000000079800000F3000029980780",
INIT_06 => X"6E461803081FC000000001FFF0000000000001F7C3C380F87C019FFF00000000",
INIT_07 => X"600C2400013649609C8000980040814210254000A00B21FF2003F2A80D500000",
INIT_08 => X"0BF80000000000000003F7FFD88D2B4A02C0940062EC2804001610020408178B",
INIT_09 => X"8E1F5FE010092C0892A041FFC0000001FFBEF0000000001DFFC002C000000000",
INIT_0A => X"41FF0C0000000000600000000001BFFA0000005501AA00000CE2000009400000",
INIT_0B => X"018C0411020600048620C030020502000200000400490510CC00040020201BF4",
INIT_0C => X"0808064106040300C00C10030400C10030400C10030400C10030400608018210",
INIT_0D => X"0000000000004003000000000000001200580000000000000000000001FFBE00",
INIT_0E => X"0086C022005381380FDB96516140C6043FFD5BFF000041000000004110000000",
INIT_0F => X"80010D804400A7240C840C201D0210840043B4804012500021E0088014C04940",
INIT_10 => X"4109038041021C980200D06410C1924030008142E06024A00043C01100298092",
INIT_11 => X"587CC200002100C14428090A1D02348190814C09C010104025AA40041A0D8005",
INIT_12 => X"022E0030300B0E46177004208000D8C61D7004300000D884817B00011306B2D9",
INIT_13 => X"01E003060344710009875C018100013831000985DC000C20003C310006143B70",
INIT_14 => X"4001850EDC004780144806A64400186CBF8961104000C3807884000846EB9500",
INIT_15 => X"FF0006E08C063C0220002201490418082010A57263E0100008000290161E711C",
INIT_16 => X"00000000000000000000000000000000000000000000000000000000000007DF",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"F2D0AEEAF6E7CC1132CDB4441990000000000000000000000000000000000000",
INIT_1A => X"BEFBE79E79E79E79E79EFBEFBEFBEFBEFBEF9EF9EF9EF9EFA69861219575D75F",
INIT_1B => X"783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1EFBEF",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000783C1E0F0783C1E0F0",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0201000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A000400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA000400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000400000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402010000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"00002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080002010FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000400010FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA00040000",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020100000000000000000000000000",
INIT_38 => X"74BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"000010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA000002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974AA000402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000002010F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_4,               -- Port A enable input
WEA      => wbe_a_hi_1024_4(3),               -- Port A write enable input
DIA(0)   => data_write_a(24),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_4(24),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_4,               -- Port B enable input
WEB      => wbe_b_hi_1024_4(3),               -- Port B write enable input
DIB(0)   => data_write_b(24),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_4(24),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_25_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100200002000000080100004000000020000800041000080808",
INIT_02 => X"FC400086000000800000000F9FFEFF8E738FFF1FC204010000000111568DD7F8",
INIT_03 => X"00000400000000400000000D00002CC4740000008000000080000000000001BF",
INIT_04 => X"68003FFF64A564AC000000000001FFFE0082EF00010370E007A1000000004000",
INIT_05 => X"0A00040148F8BFF80920804DF0F00101DFC040000079C92484F30499299837C1",
INIT_06 => X"66041803081FC0E0801101FFFD000E41002299F7E3C380F87C019FFF81200096",
INIT_07 => X"000000080480AE00000080000000000000000000A00B21FF2003E00000000000",
INIT_08 => X"1BF80000400A02000003F7FFFA0008000200A0400008A0000014100200081000",
INIT_09 => X"8E1F5FFA53EFBCACB2E369FFE0010001FFBEF80C40630C7DFFEEBAF000800202",
INIT_0A => X"41FF0C0600000000600000000001BFFE00301000000000000CC020000140000C",
INIT_0B => X"01DCCC31222730A49620C030020100000200000400490D10EC00040220201BF4",
INIT_0C => X"0808064106240300C00C10030400C10030400C10030400C10030400608018210",
INIT_0D => X"0883044582114013412080000000000000000000000000000012800001FFBE00",
INIT_0E => X"00040020000180380FC386106140C6043FFD5BFF00A04B80608003CB120C1106",
INIT_0F => X"0000080040000200040400000100000000009480000240000100080000400900",
INIT_10 => X"0001000000000808000000240000020000000100006004800002001000008012",
INIT_11 => X"0001001808220000002004001900000080800008000000000022400000088000",
INIT_12 => X"0010000000000E00110000000000408009000000000040808063004000008200",
INIT_13 => X"6000000000046100000240000000001021000004400000000010210000001010",
INIT_14 => X"4000000404000800000000060400000088000001800000001084000000088000",
INIT_15 => X"FF800C608C041002000002000006100000002100000000180600000000100018",
INIT_16 => X"4110441104411044110441104411044510629041040D180400000010028047DF",
INIT_17 => X"1104411044110441104411044110441104411044110441104411044110441104",
INIT_18 => X"1044110441104411044110441104411044110441104411044110441104411044",
INIT_19 => X"FBA2894A196A8C5A2932EC15DA080800002FFFFFFFFFFFFFFFFFC11044110441",
INIT_1A => X"2492492492492492492410410410410410410492410492412000531215A69A6B",
INIT_1B => X"158AC562B158AC562B158AC562B158AC562B1588C46231188C46231188C49249",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000B158AC562B158AC562B",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080000010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000010FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08000000",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_4,               -- Port A enable input
WEA      => wbe_a_hi_1024_4(3),               -- Port A write enable input
DIA(0)   => data_write_a(25),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_4(25),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_4,               -- Port B enable input
WEB      => wbe_b_hi_1024_4(3),               -- Port B write enable input
DIB(0)   => data_write_b(25),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_4(25),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_26_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"E9264EAB20190CA3BA4997AA9002AE9C001006B0778015CFA17E0811039879C7",
INIT_01 => X"2FFFF9BB1F773C7F9BB07DFFFDD863FC5FFF3FEFFBBF9FFB22FFFBC7B9F30686",
INIT_02 => X"E06CCC62052E708180F6FFBFFFFCFFFFF9C7FF7FC24332E642090000074037F6",
INIT_03 => X"428003739CD9863739CD9869FE2B7DEAF300029E4E300DFE69A6E644E6FF473F",
INIT_04 => X"7C2FEFFFF5BA124F003DD31EAFFFFFEE9FF7EE6F4C0770FFD7DC7CA53997B2B1",
INIT_05 => X"DFFB5421C1F8BBFAFDBFFACDF0FFCC05DDDBFF3690F9EDB7F5F7AFF639BD7DE3",
INIT_06 => X"EFD044ABC817C3E3A74667FDFFB6FF5727CC3BFEF7C3FAF87FF59F7FFBFEF69F",
INIT_07 => X"00003002132462052E708180EF060C18E5BEFB051225CDFF7002C4EEDE77F6E0",
INIT_08 => X"3FFF7D5000EC75088ED3FF7FC8790E46426CE06CB1F8E041051831FA3068D77E",
INIT_09 => X"C05FD7FF9BEFBDCEFBEE59FEF44F6603EFBEFAFCC2E35E7FDFD147CCF3F583FA",
INIT_0A => X"67FF1C7FBFADEB31E35768E8ED6BFDF3EB3EBF9DDBCE7FDC1DF8A760F3EACC02",
INIT_0B => X"5BDDCC3B336F7C548667D47B7737AF3FD62601EDC25B3533DCEB07F262213FFC",
INIT_0C => X"5F9A06E19F4D93A0EA0F78C35E30D78C35E30D78C35E30D78C35E986BC61AE31",
INIT_0D => X"5FD7AFEFDFFAF59B6FF28FE1D80D73D840607307DCFE1D80EF69A004DFFFF7FF",
INIT_0E => X"0004001F8041897B2FFFC6D86D70CE04FFFFF3FF1F5F5475BD7F72E4D75EBFAF",
INIT_0F => X"F60008003F008237B0040A00010003E020023E0201F45EC0010007E01047D17B",
INIT_10 => X"00010001DC0004C81003DE050A700200001DC0006863E8BD8002000FC0208FA2",
INIT_11 => X"2200E400002801E1A00004C21C0206F60081800800007B00010F02007EC09A0E",
INIT_12 => X"0880007E000807C7C1A612001E0015C7C19C22001E0015C59DFE82011A311AA0",
INIT_13 => X"00001BC00101F60409F0670840070809760409F06984800780097604067D0010",
INIT_14 => X"81019F40042100001F800203D81019EC085614000085C80023D81009CF008A74",
INIT_15 => X"FF802FFDFFAFD082003B032FB987E04021D481D4000819060801E0D00001231D",
INIT_16 => X"EBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEFFBFBFBFBBFCFBB0FFDFEFFEF2DFFFFFB",
INIT_17 => X"BFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAF",
INIT_18 => X"FAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFE",
INIT_19 => X"475B15BCF491E166CC8553F86EDB5C88646FFFFFFFFFFFFFFFFFEBFAFEBFAFEB",
INIT_1A => X"861861861861861861861861861861861861869A69A61861AFBD54D5F871C71D",
INIT_1B => X"984C26130984C26130984C26130984C26130984C26130984C26130984C261861",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000984C26130984C26130",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040201",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_4,               -- Port A enable input
WEA      => wbe_a_hi_1024_4(3),               -- Port A write enable input
DIA(0)   => data_write_a(26),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_4(26),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_4,               -- Port B enable input
WEB      => wbe_b_hi_1024_4(3),               -- Port B write enable input
DIB(0)   => data_write_b(26),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_4(26),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_27_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"00080A40000A41248002029000050A088000008242A0004404480002000A1155",
INIT_01 => X"2FFFF1C11F781C129C107DFFFE0860941E81258CA2B71C2220EC1B86E1A00002",
INIT_02 => X"E1000000810000014400FF6FFFF0FFFFF8007F1FC21110005080200000221FF0",
INIT_03 => X"4080026318C18226318C1821302232EAE00002BE001115FE48620040840A863F",
INIT_04 => X"643D4FFC2530000F003D821C0BFFFF8E9EF79E6D440748FED70060842105B0B0",
INIT_05 => X"D6F39020D1F8A3FAFDBFBACDC8FDC405D1DB7F1490E5EDB7D5CBADB2385D79C3",
INIT_06 => X"6FE000A38007C3032646EFF1F0B6FF46A78C39F8E723F2E47FE59C7F9ADA2612",
INIT_07 => X"00002820000000810000014401060C180190310540118DFF1000C0849673F6C0",
INIT_08 => X"3FF779100062B12A8EC3F47FC80208808210880C00082050000110023068D030",
INIT_09 => X"005F07E09BFFBD07FBAC09F8E42922038F7DF8BEC2E39C5F1FD047CEF1B582D8",
INIT_0A => X"63FF5D5F9FADE911E81C09818109E1F16B16B71092CE7ED81CF403601228C402",
INIT_0B => X"1BFDCC39732F3554866AD57C37BEAF1C152201A4C05B7531D56B05B06A213FF8",
INIT_0C => X"5BCA06F18FC59380F00E34430D10C34430D10C34430D10C34430F0861A2186B5",
INIT_0D => X"5B56ADAB5FAAE58B2F628EA0C80FA3F04040510768EA0C80CC61A0044DFFC6EB",
INIT_0E => X"0004001D800188792CE79715710AE4047FFD23FF315D54358D593474955AB6AD",
INIT_0F => X"520008003B000297B0040200010003E020001F0201E44A400100076000579129",
INIT_10 => X"00010001DC00004A10035E0408300200001DC000086BC8948002000EC000AF22",
INIT_11 => X"02002400002801E1A00000C01E0202F60080800800007B00000782006EC0820A",
INIT_12 => X"0080007E000006A7C10602001E0001A7C10C02001E0001C18DE282010A311AA0",
INIT_13 => X"00001BC00000FE0401F04300400708007E0401F04180800780007E04047D0010",
INIT_14 => X"81011F40040100001F800002F81011EC080604000085C80001F810094F008034",
INIT_15 => X"FF800C6DDDAFD082001B03249887E04001D481D4000009020801E0D00001021F",
INIT_16 => X"AB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6BF1EBDABD8E270BF84A25C6ACB777E3",
INIT_17 => X"B6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6AD",
INIT_18 => X"6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADA",
INIT_19 => X"490E2168100481CA860402104A471688747FFFFFFFFFFFFFFFFFAB6ADAB6ADAB",
INIT_1A => X"000000000000000000000000000000000008200000000000200072F210000001",
INIT_1B => X"05028140A05028140A05028140A05028140A0500804020100804020100800000",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000A05028140A05028140A",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040201",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_4,               -- Port A enable input
WEA      => wbe_a_hi_1024_4(3),               -- Port A write enable input
DIA(0)   => data_write_a(27),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_4(27),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_4,               -- Port B enable input
WEB      => wbe_b_hi_1024_4(3),               -- Port B write enable input
DIB(0)   => data_write_b(27),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_4(27),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_28_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"02200AA400180030808802A900002A08001280A08A801044104A1000001818C3",
INIT_01 => X"0AA00011460214428114180000882214413D0A71592A01D92213D28005210202",
INIT_02 => X"0451110A012100884000AA30200000000C100040104112101100008888200000",
INIT_03 => X"448000318C52A20318C52A20148810200111100C211004AA00034204200A2200",
INIT_04 => X"04004001001A90110000121402AA0000003C00000500000040080421080D0080",
INIT_05 => X"4060000C8001000000002E000000050000001610300000010000802202040012",
INIT_06 => X"1000002080001111001222000425A1040026A008000000000000000009328280",
INIT_07 => X"2491008A00491201210088400122448908A20402000408001000040820000000",
INIT_08 => X"20058310402A160026500000028040101004200C840082115554000112244814",
INIT_09 => X"4140000800000060000720000102028000000490160801020002200011100010",
INIT_0A => X"020000081B34211082B694D4D294000020020381040000000200032040004400",
INIT_0B => X"4800210C19808400500010009110091500020B408810000100200020408B0000",
INIT_0C => X"01028000080118020023604858121604858121604858121604858090B0242C00",
INIT_0D => X"010000800920040804020A6058003108402043058C460580653020005A004039",
INIT_0E => X"00000002800008014004104104420A00C000200005000010040A0020CC000200",
INIT_0F => X"520000000500000010000200000000000000280000040A40000000A000001029",
INIT_10 => X"00000000000000C0000002000830000000000000480008148000000140000020",
INIT_11 => X"020024000000000000000440000000020000800000000000000C00000040020A",
INIT_12 => X"00800000000001804006020000000500400C0200000005400A90000000100000",
INIT_13 => X"0000000000018200001003004000000142000010018080000001420000200000",
INIT_14 => X"8000080000010000000000018800008000060400000000000310000008000034",
INIT_15 => X"000002040080000000110006B081400000400000000009020000000000002200",
INIT_16 => X"802008020080200802008020080200802101210810C39A66A90A85420413A820",
INIT_17 => X"0200802008020080200802008020080200802008020080200802008020080200",
INIT_18 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_19 => X"DE21102C110A00246972BD89A40A0C22E1000000000000000000002008020080",
INIT_1A => X"2082082082082082082082082082082082082082082082080D35050758C30C31",
INIT_1B => X"0582C160B0582C160B0582C160B0582C160B0580C06030180C06030180C08208",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000B0582C160B0582C160B",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_4,               -- Port A enable input
WEA      => wbe_a_hi_1024_4(3),               -- Port A write enable input
DIA(0)   => data_write_a(28),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_4(28),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_4,               -- Port B enable input
WEB      => wbe_b_hi_1024_4(3),               -- Port B write enable input
DIB(0)   => data_write_b(28),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_4(28),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_29_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"79964E4BA01DACAB9E659792D00AAE160002829C7FDFEFCEE97C2815039D70C3",
INIT_01 => X"0ABFF9AB0775343F9AB01DF80D5821FC0FFF3FEFD1AF9FF1207FFBC7B9720586",
INIT_02 => X"002CCC60050E700080F6AAA7BFFC007189C7FF2FC00330E602800000074037F6",
INIT_03 => X"468003210868A63210868A68DA017D207200021C4E200CAA6186A40042FF4300",
INIT_04 => X"7C2FE002F0900001003C5316A6ABFFE21F36E02F0D03701F47D41800109FB281",
INIT_05 => X"4979440580F9B808F49F6A4DF00F8D01DC4B97369078249370F482E62BA41462",
INIT_06 => X"B250442BC81001E1870223FC0BF7F11507C423FE33C078F803F19F00E936721D",
INIT_07 => X"00011080012460050E700080EF020408EC8CFA01122149FF700200665A35D260",
INIT_08 => X"2BFD055040A452000443FF00007906464068406C31F84000000831FA1028575A",
INIT_09 => X"805FD017102690AA694551FE30444681E0820AD40201423FC00122C493500172",
INIT_0A => X"0600002AFFBE2330815568A8AD6ABC02A02A0B0CCB463B4C0748A720B1EA4C00",
INIT_0B => X"0850400A11414C005005000B51158936D20601A98A10200308A002E240010BFC",
INIT_0C => X"05928020194918A22A2268C81A32068C81A32068C81A32068C81A99034640C00",
INIT_0D => X"058102C48970541944B20FA1580561D040406305587A158046282000DBFFF13D",
INIT_0E => X"000000028040890327DCD28928324400DFFFF0001F1F0050342D42A086040B02",
INIT_0F => X"F60000000500802010000A000000000000022A0000141EC0000000A01000507B",
INIT_10 => X"00000000000004C0000082010A700000000000006800283D80000001402000A0",
INIT_11 => X"2200E4000000000000000442040004020001800000000000010D000010401A0E",
INIT_12 => X"08800000000801C040A6120000001540409C2200000015441DAC800010100000",
INIT_13 => X"0000000001019600081027084000000956000810298480000009560002200000",
INIT_14 => X"800088000021000000000201D800088000561400000000002358000088000A74",
INIT_15 => X"00802594A282C0000033010FB181E00020400000000819060000000000002305",
INIT_16 => X"C0B02C0B02C0B02C0B02C0B02C0B02C4B12B312912831A27FCFE7FFB175B6FF8",
INIT_17 => X"0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02",
INIT_18 => X"B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C",
INIT_19 => X"BBCF9F96EE7FFDF7FE783FFDFFEA0C00602FFFFFFFFFFFFFFFFFC0B02C0B02C0",
INIT_1A => X"EFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEEBAEBAEBAEBAEBBFFDF9FBEFFFFFFE",
INIT_1B => X"BFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFBEFB",
INIT_1C => X"FFFFFFFFFFFFFFF800000000000000000000000000000FBFDFEFF7FBFDFEFF7F",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_4,               -- Port A enable input
WEA      => wbe_a_hi_1024_4(3),               -- Port A write enable input
DIA(0)   => data_write_a(29),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_4(29),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_4,               -- Port B enable input
WEB      => wbe_b_hi_1024_4(3),               -- Port B write enable input
DIB(0)   => data_write_b(29),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_4(29),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_30_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"F7FFBFFEFF9FE1F7FFBFFFFDFFD0000000000000000000000000000000000000",
INIT_1A => X"9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7AFBD75F5FDF7DF7F",
INIT_1B => X"F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE79E7",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000003F9FCFE7F3F9FCFE7F3",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_4,               -- Port A enable input
WEA      => wbe_a_hi_1024_4(3),               -- Port A write enable input
DIA(0)   => data_write_a(30),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_4(30),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_4,               -- Port B enable input
WEB      => wbe_b_hi_1024_4(3),               -- Port B write enable input
DIB(0)   => data_write_b(30),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_4(30),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_31_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"129000008004A00804A40000400800020000000C005FEA005800200400050100",
INIT_01 => X"255FF18019700810180065FFFC0040801E80258CA2951C2200EC0906A0804140",
INIT_02 => X"E0000000000000011000550FDFF0FFFFF0007F1FC200000044000000000817F0",
INIT_03 => X"0000024210A30024210A3001002220C06044469200040154482000408400043F",
INIT_04 => X"602D0FFC2420000E003D80080955FF8E1ECA8E2D400340FE870060842100B030",
INIT_05 => X"0213100040F8A3F8FDBF944DC0FDC001D1CB6904A061EDB6D4C30490281831C1",
INIT_06 => X"6FC000830007C202060445F1F0D25E4207A099F0E303F0E07FE19C7F80402412",
INIT_07 => X"0000200000000000000001100004081001103107000185FF0000C0849673F6C0",
INIT_08 => X"1BF27A00000000000883F47FC800080002008000000820440000100220489020",
INIT_09 => X"011F07E013EFBC06FBA009F8E00120038F3CF82C44630C5D1FC002CCE0808248",
INIT_0A => X"61FF0C06C48BC801600000000001A1F00110101092CE7ED81CF0004012288000",
INIT_0B => X"11DCCC31222730048620C4382204A608142002A440492530C401049020221BF8",
INIT_0C => X"0888066187448380E00C10030400C10030400C10030400C10030600608018210",
INIT_0D => X"080204010200418301208480800D02D00040100240A808008840800405FF8640",
INIT_0E => X"0004001D000180780CE386106100C4043FFD03FF101D40008001304018081004",
INIT_0F => X"000008003A000217A0040000010003E02000160201E040000100074000478100",
INIT_10 => X"00010001DC00000810035C0400000200001DC0000063C0800002000E80008F02",
INIT_11 => X"00000000002801E1A00000801C0202F40080000800007B00000302006E808000",
INIT_12 => X"0000007E00000607810000001E000087810000001E000081846282010A211AA0",
INIT_13 => X"00001BC00000740401E0400000070800340401E04000000780003404045D0010",
INIT_14 => X"01011740040000001F8000025010116C080000000085C80000C8100947008000",
INIT_15 => X"FF800C609C06D082000A03200806A040019481D4000000000801E0D00001001D",
INIT_16 => X"010040100401004010040100401004010060C040040C200950402090128057C3",
INIT_17 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_18 => X"0040100401004010040100401004010040100401004010040100401004010040",
INIT_19 => X"00000000000000000000000000001000802FFFFFFFFFFFFFFFFF810040100401",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_25 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFF",
INIT_27 => X"0200000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_2B => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_2C => X"A080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_2D => X"FFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974B",
INIT_2E => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFF",
INIT_2F => X"FFFF5D2E974BA080402000000000000000000000000000000000000000000000",
INIT_30 => X"FFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFF",
INIT_31 => X"E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFF",
INIT_32 => X"FFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2",
INIT_33 => X"80402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFF",
INIT_34 => X"FFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0",
INIT_35 => X"0FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFF",
INIT_36 => X"00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200",
INIT_37 => X"FFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000000",
INIT_38 => X"74BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFF",
INIT_39 => X"FFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E9",
INIT_3A => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFF",
INIT_3B => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_3D => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_3E => X"0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_1024_4,               -- Port A enable input
WEA      => wbe_a_hi_1024_4(3),               -- Port A write enable input
DIA(0)   => data_write_a(31),        -- Port A data input
DOA(0)   => data_read_a_hi_1024_4(31),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_1024_4,               -- Port B enable input
WEB      => wbe_b_hi_1024_4(3),               -- Port B write enable input
DIB(0)   => data_write_b(31),        -- Port B data input
DOB(0)   => data_read_b_hi_1024_4(31),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


end;