library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_misc.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library UNISIM;
use UNISIM.vcomponents.all;

entity ram_master is
	port(clk             : in  std_logic;
        address_a       : in  std_logic_vector(31 downto 2);
        enable_a        : in  std_logic;
        wbe_a           : in  std_logic_vector(3 downto 0);
        data_write_a    : in  std_logic_vector(31 downto 0);
        data_read_a     : out std_logic_vector(31 downto 0);

        address_b       : in  std_logic_vector(31 downto 2);
        enable_b        : in  std_logic;
        wbe_b           : in  std_logic_vector(3 downto 0);
        data_write_b    : in  std_logic_vector(31 downto 0);
        data_read_b     : out std_logic_vector(31 downto 0));
end; --entity ram     

architecture ram_master of ram_master is
signal enable_a_lo       : std_logic;
signal wbe_a_lo          : std_logic_vector(3 downto 0);
signal data_write_a_lo   : std_logic_vector(31 downto 0);
signal data_read_a_lo    : std_logic_vector(31 downto 0);
signal enable_b_lo       : std_logic;
signal wbe_b_lo          : std_logic_vector(3 downto 0);
signal data_read_b_lo    : std_logic_vector(31 downto 0);
signal enable_a_hi       : std_logic;
signal wbe_a_hi          : std_logic_vector(3 downto 0);
signal data_read_a_hi   : std_logic_vector(31 downto 0);
signal enable_b_hi       : std_logic;
signal wbe_b_hi          : std_logic_vector(3 downto 0);
signal data_read_b_hi    : std_logic_vector(31 downto 0);
signal address_a_reg     : std_logic_vector(31 downto 2);
signal address_b_reg     : std_logic_vector(31 downto 2);
signal enable_a_lo_256       : std_logic;
signal wbe_a_lo_256          : std_logic_vector(3 downto 0);
signal data_write_a_lo_256   : std_logic_vector(31 downto 0);
signal data_read_a_lo_256    : std_logic_vector(31 downto 0);
signal enable_b_lo_256       : std_logic;
signal wbe_b_lo_256          : std_logic_vector(3 downto 0);
signal data_read_b_lo_256    : std_logic_vector(31 downto 0);
signal enable_a_hi_256       : std_logic;
signal wbe_a_hi_256          : std_logic_vector(3 downto 0);
signal data_read_a_hi_256   : std_logic_vector(31 downto 0);
signal enable_b_hi_256       : std_logic;
signal wbe_b_hi_256          : std_logic_vector(3 downto 0);
signal data_read_b_hi_256    : std_logic_vector(31 downto 0);
signal enable_a_lo_512       : std_logic;
signal wbe_a_lo_512          : std_logic_vector(3 downto 0);
signal data_write_a_lo_512   : std_logic_vector(31 downto 0);
signal data_read_a_lo_512    : std_logic_vector(31 downto 0);
signal enable_b_lo_512       : std_logic;
signal wbe_b_lo_512          : std_logic_vector(3 downto 0);
signal data_read_b_lo_512    : std_logic_vector(31 downto 0);
signal enable_a_hi_512       : std_logic;
signal wbe_a_hi_512          : std_logic_vector(3 downto 0);
signal data_read_a_hi_512   : std_logic_vector(31 downto 0);
signal enable_b_hi_512       : std_logic;
signal wbe_b_hi_512          : std_logic_vector(3 downto 0);
signal data_read_b_hi_512    : std_logic_vector(31 downto 0);
signal enable_a_lo_512_2       : std_logic;
signal wbe_a_lo_512_2          : std_logic_vector(3 downto 0);
signal data_write_a_lo_512_2   : std_logic_vector(31 downto 0);
signal data_read_a_lo_512_2    : std_logic_vector(31 downto 0);
signal enable_b_lo_512_2       : std_logic;
signal wbe_b_lo_512_2          : std_logic_vector(3 downto 0);
signal data_read_b_lo_512_2    : std_logic_vector(31 downto 0);
signal enable_a_hi_512_2       : std_logic;
signal wbe_a_hi_512_2          : std_logic_vector(3 downto 0);
signal data_read_a_hi_512_2   : std_logic_vector(31 downto 0);
signal enable_b_hi_512_2       : std_logic;
signal wbe_b_hi_512_2          : std_logic_vector(3 downto 0);
signal data_read_b_hi_512_2    : std_logic_vector(31 downto 0);
begin
process(clk)
begin
if rising_edge(clk) then
	address_a_reg <= address_a;
	address_b_reg <= address_b;
	end if;
end process;
data_read_a <= data_read_a_lo when (address_a_reg < x"0001000"&"00") else
data_read_a_hi when ((address_a_reg >= x"0001000"&"00") and (address_a_reg < x"0002000"&"00")) else 
data_read_a_lo_256 when ((address_a_reg >= x"0002000"&"00") and (address_a_reg < x"0003000"&"00")) else 
data_read_a_hi_256 when ((address_a_reg >= x"0003000"&"00") and (address_a_reg < x"0004000"&"00")) else 
data_read_a_lo_512 when ((address_a_reg >= x"0004000"&"00") and (address_a_reg < x"0005000"&"00")) else 
data_read_a_hi_512 when ((address_a_reg >= x"0005000"&"00") and (address_a_reg < x"0006000"&"00")) else 
data_read_a_lo_512_2 when ((address_a_reg >= x"0006000"&"00") and (address_a_reg < x"0007000"&"00")) else 
data_read_a_hi_512_2 when ((address_a_reg >= x"0007000"&"00") and (address_a_reg < x"0008000"&"00")); 
data_read_b <= data_read_b_lo when (address_b_reg < x"0001000"&"00") else
data_read_b_hi when ((address_b_reg >= x"0001000"&"00") and (address_b_reg < x"0002000"&"00")) else
data_read_b_lo_256 when ((address_b_reg >= x"0002000"&"00") and (address_a_reg < x"0003000"&"00")) else 
data_read_b_hi_256 when ((address_b_reg >= x"0003000"&"00") and (address_b_reg< x"0004000"&"00")) else 
data_read_b_lo_512 when ((address_b_reg >= x"0004000"&"00") and (address_b_reg< x"0005000"&"00")) else 
data_read_b_hi_512 when ((address_b_reg >= x"0005000"&"00") and (address_b_reg< x"0006000"&"00")) else 
data_read_b_lo_512_2 when ((address_b_reg >= x"0006000"&"00") and (address_b_reg< x"0007000"&"00")) else 
data_read_b_hi_512_2 when ((address_b_reg >= x"0007000"&"00") and (address_b_reg< x"0008000"&"00")); 
enable_a_lo <= enable_a when (address_a < x"0001000"&"00") else '0';
enable_b_lo <= enable_b when (address_b < x"0001000"&"00") else '0';
enable_a_hi <= enable_a when ((address_a >= x"0001000"&"00") and (address_a < x"0002000"&"00")) else '0';
enable_b_hi <= enable_b when ((address_b >= x"0001000"&"00") and (address_b < x"0002000"&"00")) else '0';
enable_a_lo_256 <= enable_a when ((address_a >= x"0002000"&"00") and (address_a < x"0003000"&"00")) else '0';
enable_b_lo_256 <= enable_b when ((address_b >= x"0002000"&"00") and (address_b < x"0003000"&"00")) else '0';
enable_a_hi_256 <= enable_a when ((address_a >= x"0003000"&"00") and (address_a < x"0004000"&"00")) else '0';
enable_b_hi_256 <= enable_b when ((address_b >= x"0003000"&"00") and (address_b < x"0004000"&"00")) else '0';
enable_a_lo_512 <= enable_a when ((address_a >= x"0004000"&"00") and (address_a < x"0005000"&"00")) else '0';
enable_b_lo_512 <= enable_b when ((address_b >= x"0004000"&"00") and (address_b < x"0005000"&"00")) else '0';
enable_a_hi_512 <= enable_a when ((address_a >= x"0005000"&"00") and (address_a < x"0006000"&"00")) else '0';
enable_b_hi_512 <= enable_b when ((address_b >= x"0005000"&"00") and (address_b < x"0006000"&"00")) else '0';
enable_a_lo_512_2 <= enable_a when ((address_a >= x"0006000"&"00") and (address_a < x"0007000"&"00")) else '0';
enable_b_lo_512_2 <= enable_b when ((address_b >= x"0006000"&"00") and (address_b < x"0007000"&"00")) else '0';
enable_a_hi_512_2 <= enable_a when ((address_a >= x"0007000"&"00") and (address_a < x"0008000"&"00")) else '0';
enable_b_hi_512_2 <= enable_b when ((address_b >= x"0007000"&"00") and (address_b < x"0008000"&"00")) else '0';
wbe_a_lo <= wbe_a when  enable_a_lo='1' else x"0";
wbe_a_hi <= wbe_a when  enable_a_hi='1' else x"0";
wbe_b_lo <= wbe_b when  enable_b_lo='1' else x"0";
wbe_b_hi <= wbe_b when  enable_b_hi='1' else x"0";
wbe_a_lo_256 <= wbe_a when  enable_a_lo_256='1' else x"0";
wbe_a_hi_256 <= wbe_a when  enable_a_hi_256='1' else x"0";
wbe_b_lo_256 <= wbe_b when  enable_b_lo_256='1' else x"0";
wbe_b_hi_256 <= wbe_b when  enable_b_hi_256='1' else x"0";
wbe_a_lo_512 <= wbe_a when  enable_a_lo_512='1' else x"0";
wbe_a_hi_512 <= wbe_a when  enable_a_hi_512='1' else x"0";
wbe_b_lo_512 <= wbe_b when  enable_b_lo_512='1' else x"0";
wbe_b_hi_512 <= wbe_b when  enable_b_hi_512='1' else x"0";
wbe_a_lo_512_2 <= wbe_a when  enable_a_lo_512_2='1' else x"0";
wbe_a_hi_512_2 <= wbe_a when  enable_a_hi_512_2='1' else x"0";
wbe_b_lo_512_2 <= wbe_b when  enable_b_lo_512_2='1' else x"0";
wbe_b_hi_512_2 <= wbe_b when  enable_b_hi_512_2='1' else x"0";



ram_bit_0_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"ED39BA795990D275FB4A6E96ACC4731DEA4598B0AFB54867F6EE4618C3749803",
INIT_01 => X"58A0047C8607844847CA180001E4A2404042106208408208C2002069161734B3",
INIT_02 => X"8B1EC9562121F8051500147A0E5629A302CF28400615F5787B09FBF999BB1EFD",
INIT_03 => X"404EFC0A2AD6100F01A88E851CE47803C280110521898F6996088862C7B22221",
INIT_04 => X"C0D001C0100AEC83C008E7880D01A64661800002C21A52C590D2012194804844",
INIT_05 => X"650002C3F08754001B51981E007910070F01C1E003980015A204C22F32328BAF",
INIT_06 => X"BCDA4677CAEE7CF5BB870E1DDB9889C5FBFC440129A0604442180238203F70C1",
INIT_07 => X"7AAE0088B02000C2EC3A0E829836E0AF3325372E2AA8FDF3C18306758B24197A",
INIT_08 => X"D7E40002F7AE005FFB4730010411400A61080000F7F4C464B58294901606D5A5",
INIT_09 => X"C4801C40469B0CA9881A28C141118000C5A85A60444210123820B43B40804274",
INIT_0A => X"400800219010107ED453C041B13216656074EA560F0092A24856B05312226900",
INIT_0B => X"27122C3E04E03383E2781EA781E2781EA781E2781EA781E2781C33C0613C0E29",
INIT_0C => X"74EB1F50D0758A9650E520610A6A57A5529E2B439499CF96B086000000B09870",
INIT_0D => X"04F07E024108F4E28638EC57250004480155C1375A97A9121F8BA749D3A4E9D2",
INIT_0E => X"04F07E42177EFDF8570184071575970F8FC07D5BFF078004F07E007D5BFF0780",
INIT_0F => X"8F85ECB1FE047F5FB7B30E0700461E5AF8007D5BFF078004F07E007D5BFF0780",
INIT_10 => X"C0184D07C1DF15C7E3E2177EFDF8C3C03009C3CDD47C7F403FB3FDF89701C011",
INIT_11 => X"4F80FE659C6104C6D7103F9D1D064189B5924418D65FE45DEE55BBEDE34CF900",
INIT_12 => X"6395F64207F3A3A1483136B881FCCB38C2098DACA01FFF603F80001F80FDC81F",
INIT_13 => X"FED151E01015C3BB507D3F811FBEC32B81840714F8D91F4FC513F37C8AE07002",
INIT_14 => X"61692F293185D8D724E15D3FCC6B7C236FE0691A9500125C1F83F8CC1F4FC507",
INIT_15 => X"E93A4E93A4E93A4E93A4E93A4F942F90E9628540052090650525A0000066A00B",
INIT_16 => X"93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4",
INIT_17 => X"3A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E",
INIT_18 => X"09B56C74DAB15D1CF13501AA495000000000000000003A4E93A4E93A4E93A4E9",
INIT_19 => X"2082082082082082082082082082082082082082082084E41DC71C7155F3898E",
INIT_1A => X"3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F8208208208208",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE5294A5294A52800003E1F0F87C3E1F0F87C3E1F0F87C",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000030FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"A975EFFFAABDE00FFAEBDFFF5D2EAAAAAF7AEBDEBA0000000000000000000000",
INIT_22 => X"8000155087FC0155F7D168B55007BFDF45085168ABA002E82145085155545F7A",
INIT_23 => X"FFFD7545AA8028A00A2802AABAFF8028BEF5D7FFFE10005542145557FD5545FF",
INIT_24 => X"F7AEAAAAAA2FFFDF4500043FE105D2E954BAF7FFC0010080017555555568AAAF",
INIT_25 => X"A5D5168A00A2D142155005142010FFAE820AAFF842AABAA2AE95545FFD168ABA",
INIT_26 => X"FF5D2A821550000000BA007FD55FF5D7FC0145007FD7400550415410002E974B",
INIT_27 => X"F455D5142000082E82145FFD17DFEFFFD168BFFF780000BA007FE8AAAFF803FF",
INIT_28 => X"0000000000000000000000000000000000000000AAFBEAA00007BFDFFF082EBD",
INIT_29 => X"AABEA495FC716F002A975FFE3AA95E00EBAEBDFD75D2AA8A80EA8E2FE3F00000",
INIT_2A => X"56A16D557BC257D415E0216FA3F1E8FC0145B68B551475FAF6D1C556F0AA1C24",
INIT_2B => X"7FD24AFE3D02DAAAE12BD5545A2803AA0000542A0070071C50BAFEF1FAE0016D",
INIT_2C => X"A8B50F55A2F150005A3A438BD04AFAB8F550A8010E004924874825D7FEAA8548",
INIT_2D => X"A2A5504001C74BA42A1571E8028E3DB7816D0120155EA568E870BAEB8A05A2AE",
INIT_2E => X"2FFAFD2A82485FD2415A105C21451ED42A002545E055FFBE81D0BE8EA8A3AA05",
INIT_2F => X"100AA1D0F6F480B6A555A2A57A002A3D5FDB6A5C7E3DFFFE90B45B47ABA497A8",
INIT_30 => X"A0AFE80A8B0A000000000000000000000000000000000000000000000B55EAAA",
INIT_31 => X"ABEF5D557FEBA55022A3F70C6B405F4D2AE975EFAAAAB5E1AF3AABFF45592E88",
INIT_32 => X"411A8DED57CE1055555E5F58EFFC01FE2CACB65F520EBE9EF67D7BEA1FD5D556",
INIT_33 => X"A4AD0079C75D6070CC5CBB0280C029ABAA3EBC114728007521170821CE0FDE69",
INIT_34 => X"2A95E02A2AAB5EB0F280800EFAEE9F5D18F3142341D5DEEBEF55080034E0A592",
INIT_35 => X"B69C30E02116220415A9540AA854140A0A2047F353AAF6C77F7F20D968BF5781",
INIT_36 => X"ABEBE1B4D792A4AD1183454180DD3FDCAAAB7C91565455C141E41887D58AC448",
INIT_37 => X"F0000001FF01EABC4B8014174FF7DA80F52FEDE6BE93172D7D625B556EEAB157",
INIT_38 => X"FF0000001FF0000001FF0000001FF0000001FF0000001FF0000001FF0000001F",
INIT_39 => X"0000000000000000000000000001FF0000001FF0000001FF0000001FF0000001",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000100000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(0),        -- Port A data input
DOA(0)   => data_read_a_lo(0),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(0),        -- Port B data input
DOB(0)   => data_read_b_lo(0),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_1_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"212C001411984004084D000508C53810A03D1450E839B003342114428A000803",
INIT_01 => X"08000011400A100A81160000008C005400400002000000000000028001340000",
INIT_02 => X"C084484000002014400205851002007030450E0000A606C8C44CB4C6666C00E0",
INIT_03 => X"33DF380008164004000002000C80400002031943000101091608463061120118",
INIT_04 => X"4140008000000002000064000400004201000000000210458010070080100433",
INIT_05 => X"8500101040200000010009100000000508000100000000002010600100208D04",
INIT_06 => X"B5EDFDE24618AD433060C182BA860044204C000008A004100008000820280020",
INIT_07 => X"581E02100020000A81244890AA20263030517F122AA801F0983060AC564BF808",
INIT_08 => X"00820800C7A00045B103200000140A02234808000584000004808400020011A4",
INIT_09 => X"0000104000020082800808111008400000200204100000100820800144000414",
INIT_0A => X"12804062945211441E13C051156E800008402802060C94000040901102800000",
INIT_0B => X"24002006406401918C191AC191A4191A4191AC191AC191A4191A00C8560C8D29",
INIT_0C => X"0408010040050880383820080F105F05800302E0E08842422006000000041032",
INIT_0D => X"05000600000090C1841808172580000000008008020084082080204010200810",
INIT_0E => X"0500066210000178470184000000878402C000001E07800500062000001E0780",
INIT_0F => X"00003C404600000011A30E0700000009382000001E07800500062000001E0780",
INIT_10 => X"C0180000012010C20022100000F0C3C03000000055200340000000F88701C000",
INIT_11 => X"05800241186100004D100098190240001290002050068000001010486140F900",
INIT_12 => X"0000164A001303204800026880048230C2000094A0000F601F8000000001C908",
INIT_13 => X"12D051E01000000154200580003C030381840000004B08014401025480E07000",
INIT_14 => X"40082300218450C2800010094000482142E0601895001000000041C408014400",
INIT_15 => X"0802008020080200802008020080008208600500A82A15008000000000468000",
INIT_16 => X"8020080200802008020080200802008020080200802008020080200802008020",
INIT_17 => X"0200802008020080200802008020080200802008020080200802008020080200",
INIT_18 => X"BABEFC54A0810C7452B5420A1000000000000000000002008020080200802008",
INIT_19 => X"AAAAAAAAAAAAAAAAAAAAAAAAAAA28A28A28A28A2A8218D2C0C92492581328A46",
INIT_1A => X"2E974BA5D2E974BA5D2E974BA5D2E975BADD6EB75BADD6EB75BAAAAAAAAAAAAA",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFF6318C6318C63000002E974BA5D2E974BA5D2E974BA5D",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"00000000000000000000000C0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"002155557FFFFFF007FC21EFA2FFD74AAAAD5555550000000000000000000000",
INIT_22 => X"7FD75FFAAAA800AAF7AA974BAFFFBE8B45F7AEBDF455D2EAABEFF7FFE8BFF5D0",
INIT_23 => X"0557DF45AAD1400BAA2AE801550051555EFF7AA95400552AAAABAFFD1574105D",
INIT_24 => X"FFFBEAB55F780020AAAA80020AA082EAAB5500517DF555D2EAAA105500001550",
INIT_25 => X"AF7AE820AA0851574BAA2D1574AA5D7BFDEBAFFD540155557FD5400F78028BFF",
INIT_26 => X"FFFFD56AAAAFFFFD7555AAD168B45AAAEAAABAFF842ABEF5D517DF55552A974A",
INIT_27 => X"4BAF7AE80010082A97410557FEABFFAAFBE8BEFAAD1575EF557FFFE10557FFFF",
INIT_28 => X"00000000000000000000000000000000000000005D7FFDF4500043FE105D2E95",
INIT_29 => X"A8BC2EBDFEAF7F1F840017D4975D2FEF147FC51C7A2FBD5490BFD1C056A00000",
INIT_2A => X"AA8AAAE3D145410F7F1D55D71C002DABAEBAA974BAF7FFEFB45FFAABDF55492A",
INIT_2B => X"0E2AE85028B40155145F7AF6DBED5450AA1C2080BEF495FC71D54124924385FA",
INIT_2C => X"571D2E28E38E0216FA2D1E8E80140F45082B4002D082082AB8B6DBEDB7DF7F54",
INIT_2D => X"A97F7AF6D417E92482BF84020BA495557E3FF78E021FF1471FDEAAFFD56F16D5",
INIT_2E => X"7002FD74951D71EDFFABFD16FAAAE92BD5545A2DA3FB7DAAD4AAAAF487BC70BF",
INIT_2F => X"550A8010E00492487482FFFE82A85EBAE2FFC55554ADBD7A2FFC7BEFF6FFD7FC",
INIT_30 => X"400FBF9424F7000000000000000000000000000000000000000000000547AB8F",
INIT_31 => X"DF55F7AABFF55082CA8B4DF6C1E8F5E5400021EF005162BEF047FD5545AAFBF7",
INIT_32 => X"404547184164AA5D2EBEEB0A2D555410D3555714F8338AAAA1D0AE974AAF7FFF",
INIT_33 => X"AEABFFDF79DCBF755962010BDCBBC21455D7FEABEF75550ACBB7582225FF5843",
INIT_34 => X"D57D412F7D55F5E50C7F401BAAE8403CF5A3FFEAAEB083BC1000FF8409000512",
INIT_35 => X"2AA9FEAFDF7F431A9F7FFE81FF013A8001AFF801F8BA0C57740BDAA0688E5405",
INIT_36 => X"A2FBF7FED2C7F955445079E280A00C56145EF5D16BABAA3EBC3157ABD5FFE55F",
INIT_37 => X"0000000000596EBEF55080034E0A592A4AD00FB863550229BCABEB7DA403FFFD",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000100000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(1),        -- Port A data input
DOA(0)   => data_read_a_lo(1),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(1),        -- Port B data input
DOB(0)   => data_read_b_lo(1),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_2_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10E006600180111284380310006289800480032283E000A34301002001A0817",
INIT_01 => X"A14AC00A1079284D04A044A54E504368404000720885800802000006ECD10200",
INIT_02 => X"92250052A0348C310102048800A8507000040C8550200000480E0080001321E0",
INIT_03 => X"020204E4593C0824400C2220483042809292430400440180000890A4C9400242",
INIT_04 => X"486854B141002252142241502460480031B94420634850069A42241009610A04",
INIT_05 => X"800504244080892105AA6010A44882144840910A21220A8C820025E4A0000B00",
INIT_06 => X"A000442802280000340810209C444804206000AC800088096A0EA8C022208012",
INIT_07 => X"309820A848E0AA09826489A5CC49002001020112028201F8A20488260000108A",
INIT_08 => X"2400582881E0C1419D12041455509341A539C42A0D8208099002801700D10103",
INIT_09 => X"110D525861263100009200151409130A3C80C8C8096A06B8C12088400A9C2080",
INIT_0A => X"0451394CD0391A441583C04B580040089581001342801044877200D002A00DE0",
INIT_0B => X"144423040240450114901149013C9011C9013C9011C90134901144801A4808A5",
INIT_0C => X"D8A5345206D2C10082080A90C00000188150100C202A4640000E2B4081969420",
INIT_0D => X"050080400A0391A51240C480000AA902AA009028C83220008086952B4285A54A",
INIT_0E => X"05008021C00000000040000000020288000500000008000500802A0000000800",
INIT_0F => X"0002300000428000000040000000000D002A0000000800050080250000000800",
INIT_10 => X"0000000001204004000508000000100000000002054000130000000000800000",
INIT_11 => X"000C00000000000068144000000000001A000106200010021002000000000080",
INIT_12 => X"0002004A880000000000034098000000000000D024A000000000000001000900",
INIT_13 => X"00000000000000041400000A8000000000000000010A00000284000000000000",
INIT_14 => X"012100000002000280000000011080C000000000000000000000430000000260",
INIT_15 => X"A769DA769DA769DA368DA36CDA3A9A13A14801404134DA84A024024155000399",
INIT_16 => X"168DA769DA769DA769DA368DA368DA368DA769DA769DA769DA368DA368DA368D",
INIT_17 => X"68DA168DA169DA569DA569DA568DA168DA168DA169DA569DA569DA568DA168DA",
INIT_18 => X"138D70C030B51C50C7D000A2012F81F81F83F03F03F069DA569DA569DA568DA1",
INIT_19 => X"1041041041041041041041041041041041041041024860208165965975960040",
INIT_1A => X"25128944A25128944A25128944A25128944A25128944A2512894104104104104",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFF8421084210840703F25128944A25128944A25128944A",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"00000000000000000000000F0FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"415555087BFFF55A2AA800BAFFAE9540008002AA000000000000000000000000",
INIT_22 => X"7FE8B555551421455D0002145552EBFEBA007FC21EFA2FFD75EFAA8415410AA8",
INIT_23 => X"FFFE8B45552EBDF45FFAEAABFFF7FFE8B55F784155EFA2AEBDEAAA2FBEAABA5D",
INIT_24 => X"5D2AAAAAA5D2E820BAA2FBEAB5555557DF55A2AEBDF555D2E954BAA2AA974BAF",
INIT_25 => X"A5D04021EF557FC21FFAA8428BFFAAAA954AAAAAAAAAAAFFD1574105D7FFFF55",
INIT_26 => X"EFF7800215500557DF55AA80001FFAA80001550055575EFFF84021555D043DEA",
INIT_27 => X"B5500517DF555D042AA10A284154005D0015410085568A00FF80175FFA2D17DF",
INIT_28 => X"00000000000000000000000000000000000000005D00020AAAA80020AA082EAA",
INIT_29 => X"D55D2BE800042AFE8E1557D0075D2F45BEAA800AAFFAA9543A080038A2A00000",
INIT_2A => X"0BDEAAA2FBF8AAA557BE8B6D5D5FFABEF49040017D5D20B8EAA007FC51C7A2FB",
INIT_2B => X"0E174BFA02A974BAF7F5EFB455D2ABDF55492AA8BC7EBDFEAFEFFD00105FFBC2",
INIT_2C => X"3D155E105571D55D71C002DABA5524820BAB6FFEFB6D555578F7DB6A0BDF7D48",
INIT_2D => X"092A071555D5E3AE821D00001FF0871C016DBED1FDE90E3A497492B6AAADAAAE",
INIT_2E => X"0E3DA3DFD5E3DFFFBD5A38A021551C5F7AF6DBE8F401D7B6A0001470155C51D0",
INIT_2F => X"82B4002D082082AB8B6D1C5B7DF7FF78E075C5BE8555400550A38428007FED00",
INIT_30 => X"4AA00042AAA2000000000000000000000000000000000000000000000410F450",
INIT_31 => X"AAAA007FD5555AAFBD7545FBB8020A3F7AE975EF005560B55F7AA800AAF7AA95",
INIT_32 => X"E8F5EFF84165EFF7802BAB0A2FFEAABA557BEABEF057D68F5F5A00021EF55042",
INIT_33 => X"52ABFFFF841FFE75CA882108202E974AAF7D57DF55D7AABFF5428ACA8F45A6C1",
INIT_34 => X"84174A8FFAEBFEB0A2D55541051555694F002CA8AA80800020AAF7FBFFFEF045",
INIT_35 => X"7AAA155F595542455512A975455D3AA8A005500151FF0C57401E5F3D1E00A1A8",
INIT_36 => X"5D2A8A0B882FFFFE10AAAAAB755A66B6AF56A2AA801455D7FE8BFFF680800FFF",
INIT_37 => X"00000000000C3BC1000FF8409000512AEABFF5D79FCAF774AE005BE789555400",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000200000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(2),        -- Port A data input
DOA(0)   => data_read_a_lo(2),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(2),        -- Port B data input
DOB(0)   => data_read_b_lo(2),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_3_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"210C44A20020248B08431120001604B8156023104C4077133420400A02380202",
INIT_01 => X"015A2A424080216D3C2462C99E104B49404040028804A0080A000C16A0D90A0C",
INIT_02 => X"C0A4065000F0A95011000D1501005270B4045AB330860281CC08008222170060",
INIT_03 => X"AD22014098340394A4021320080841C40B411B4298042180002846B06900811A",
INIT_04 => X"244B32A86D20014A0D20403194904900071A24110F0BF400F85F92420E0C946E",
INIT_05 => X"80331030442898B4812840D0500008C528280B063006A64CA30004E5A4E40304",
INIT_06 => X"90016CA00E380042302040A0BC47160424428198C0038C89904E640023600816",
INIT_07 => X"1288020843A66620816049908AA0061011CA0142000009F0A810292E7402F088",
INIT_08 => X"20003C9984A0AC411102014D34EC2200214D5099048823019603A01A49410103",
INIT_09 => X"001CD74C4826220010A8891451284B661CA24A4C899046740121824004100080",
INIT_0A => X"44C9516DC0135C45159BE45F112B48804DC10203021290400772C0F402820D4C",
INIT_0B => X"B400624402404501A49018490184901A4901A4901849018C901A648056480C2D",
INIT_0C => X"D7A9B54000D7C10820680D08C420180381211081A022160000266723E1909021",
INIT_0D => X"400080200E199A4A2CA2994C0399981666409800CA52E4890806BD6B56BDAB52",
INIT_0E => X"40008008E00000000000000000024008000C8000000000400080028000000000",
INIT_0F => X"000A000000588000000000000000200400088000000000400080078000000000",
INIT_10 => X"0000001000004004000D800000000000000000022040000B4000000000000000",
INIT_11 => X"001A0000000000082006C000000000020804087220000122000A000000000000",
INIT_12 => X"00020800B8000000000041002E00000000001040466000000000000001020080",
INIT_13 => X"00000000000000048200004A600000000000000003008000320C000000000000",
INIT_14 => X"432900000222200871028000210400C4000000000000000000080200800030E0",
INIT_15 => X"AF6A5AF6A5AF6A5AF6A5AF6E5AFADA91AB68000101B4D20C08EC461733804A19",
INIT_16 => X"B6B5AF6A5AF6A5AF6A5AF6A5AF6A5AF6A5AB6B5AB6B5AB6B5AB6B5AB6B5AB6B5",
INIT_17 => X"6BDAB6B5A96ADAF6A5AD6ADAF6A5AD6ADAF6A5AD6BDAB6B5A96BDAB6B5A96BDA",
INIT_18 => X"C78C706428A14C586290008A044D54AAB556AA9556AAEBDAB6B5A96BDAB6B5A9",
INIT_19 => X"92492492492492492492492492410410410410412821600001249249015303C0",
INIT_1A => X"351A8D46A351A8D46A351A8D46A351A9D4EA753A9D4EA753A9D4924924924924",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000001543B351A8D46A351A8D46A351A8D46A",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"43DF55FFAA955EFA2D168B55557BEAA000055420000000000000000000000000",
INIT_22 => X"7BE8BFFA2D155410AA8415555087BFFF55A2AA800BAFFAE9554508002AA00AA8",
INIT_23 => X"52ABFEBA007FC21EF007FD75FFAA841541008002AB55AAAA955EF005568A0008",
INIT_24 => X"005168B455D042AB45F7FFD741000042AA10AAAABFF5508003FF555D00021455",
INIT_25 => X"0A2D1575FFF7AA975555D2E80145F78415545082EBDEAAA2FBEAABA5D7FC0155",
INIT_26 => X"55552A954BAFFFFE8B55552EBDE00F7AEAABFFF7FBEAB55F7AABDEBA5D7FC201",
INIT_27 => X"F55A2AEBDF555D2E954BA002EAAABA002A821EF5555554AA087BC01FFFFAAAAB",
INIT_28 => X"0000000000000000000000000000000000000000082E820BAA2FBEAB5555557D",
INIT_29 => X"95578080038A2AA28E3AF55E3A0BA5D7AADB6FB7D5D7FEAA3808554203A00000",
INIT_2A => X"0925D7085F6AA10087FEABD7AAD57AEBAB68E1557D1475FAF45BEAA800AAFFAA",
INIT_2B => X"04AAFFA41040017D5D20B8EAA007FC51C7A2FBD55D7BE80004AA1E8E2AB55B6A",
INIT_2C => X"2FBE80AA557BE8B6D5D5FFABEF49002FB55FFF5D0438140E2FA38B6AEBFF6D1D",
INIT_2D => X"AB8ABAE925D21C7010EADB525D7FFAE975C75D0A901FFFF801557D1C20B8EAAA",
INIT_2E => X"20875C21D5EB8AA8FFF012A954BAFFF5EFB455D20BDE00EBAAA8BC7EBDFEAFEF",
INIT_2F => X"BAB6FFEFB6D555578F7DB6A0BDF7DEB8E125FF002EADA921420871D74971D248",
INIT_30 => X"ABA0051400A20000000000000000000000000000000000000000000001C24820",
INIT_31 => X"8B55F7AA800BAF7AA955EF00042AAA2A2AEAAB55A28408145AAFFFFFFF5D7FEA",
INIT_32 => X"020A35D2ABEF55F7800015F087FEAA00007FEAB55FAD568AA2AFAE975EF55516",
INIT_33 => X"ABFEAAF7AE9DFF759A82AEF70800021EF55042AAAA007FD55558A7BD7145FBB8",
INIT_34 => X"84175EF55002AAB0A2FFEAABA557BEA3EF057968F575D003FF55F7D5420BA5D2",
INIT_35 => X"A8429F45A7D5EAF5FFBAEAAA10554155400AAFFD5145FBAC9755F05040255FFD",
INIT_36 => X"550415557085540000005156155FE90A8F5C082E974AAF7D57DF45552A3FF10A",
INIT_37 => X"00000000005500020AAF7FBFFFEF04552ABFFFF843FFE77C80825BC052ABFE10",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000100000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(3),        -- Port A data input
DOA(0)   => data_read_a_lo(3),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(3),        -- Port B data input
DOB(0)   => data_read_b_lo(3),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_4_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"A108400020612C80284210081034849800A000303100048B3432C82904204002",
INIT_01 => X"21066802000820491C00650E1E004360403008418984014902030906A8D10200",
INIT_02 => X"120404E00E4C0600000206100008402005040C00F104008040080080001310E0",
INIT_03 => X"DCA201514D1C0D706C5CF010083A0708BA0841945004010000080084C1000002",
INIT_04 => X"5C4CF21C48B133483C80417570D000083A62488074C1350EA60D785C0A6B0619",
INIT_05 => X"000F0400028083B381A60001E5546EB5C0E2B81E4166DE000139200004E50940",
INIT_06 => X"80004408020800023000102098000204A040038600018019004B800123208806",
INIT_07 => X"120C20204665E1008024188488800000001A01520000A1F08044892400001088",
INIT_08 => X"0801007AC0A1EB413102063CF3E0B3028D29F407059B0B000205A801C2200102",
INIT_09 => X"106052400922D00406BE1002C6150F41200280001900439001FD8A0004142000",
INIT_0A => X"047F2201D899BA503583504B58AB80804540001202805544314041B48A888EC5",
INIT_0B => X"1441E3443043410C5010C3010C1010C3010C1010C1010C3010C14086980861A5",
INIT_0C => X"020000A02600000805400502C0A0004A00625015000A12000026E1E180011220",
INIT_0D => X"400000000E43930C20C20188120782861E4004A800600401A030001008080400",
INIT_0E => X"40000021A8800000000000000000400800170024000000400000310024000000",
INIT_0F => X"0008000000AA80200800000000002000003400240000004000003B0024000000",
INIT_10 => X"00000010000000040004A080000000000000000020400006C008020000000000",
INIT_11 => X"002C008200000008001B4020200000020000090760000200110A040010000000",
INIT_12 => X"00000803E004040000004000E801040000001000086000000000000000020040",
INIT_13 => X"0000000000000000810000164001008000000000020040002240008020000000",
INIT_14 => X"04001040026026004000000002940040000410000000000000080000400000B8",
INIT_15 => X"040080201004008060000001806AC000004890015124D880100886D8F0014420",
INIT_16 => X"4010000180600000018020100400802010000080601000008020000401802000",
INIT_17 => X"0100000004008020180600000000000180600802010000000401802018020000",
INIT_18 => X"3807E05000140634504048820064B261934D964C326980004010000080600806",
INIT_19 => X"AAAAAAAAAAAAAAAAAAAAAAAAAAA28A28A28A28A2934C8D0CCD145144C0A28A06",
INIT_1A => X"068341A0D068341A0D068341A0D068351A8D46A351A8D46A351AAAAAAAAAAAAA",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000000173F068341A0D068341A0D068341A0D",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"57FE10FFFBEAA10007FD7410FFAA97555082A800AA0000000000000000000000",
INIT_22 => X"7FEAA00007BE8AAAAA843DF55FFAA955EFA2D168B55557BEAB45005542000005",
INIT_23 => X"87BFFF55A2AA800BAFFAE9555508002AA000055574105D2A800AA00043FEBA5D",
INIT_24 => X"A2D17DE1000517FE10AAAAA8AAA002E97545557BC00AAA2FFEAAAAAA84155550",
INIT_25 => X"0A2D157400AAAE974AAAAAA974BA08002AB55A2AA955EF005568A00087BE8BFF",
INIT_26 => X"BA080002145552ABFEAA007FC21EF007FD75FFAA8417410A2D140000F7FBC201",
INIT_27 => X"A10AAAABFF5508003FF55F7D568A00552EA8BEFA2AABDEAA087BEAAAAA2FBD54",
INIT_28 => X"000000000000000000000000000000000000000055042AB45F7FFD741000042A",
INIT_29 => X"EAB7808554203A145178E00FFFBE8A101475D5400F7A49057D0824850B800000",
INIT_2A => X"E8008200043FE925571EFA380871C7028A28E3AF55F7A0925D7AADB6FB7D5D7F",
INIT_2B => X"F5FDA38BE8E1557D1475FAF45BEAA800AAFFAA9557D080038AAA145157428492",
INIT_2C => X"85F6AA10087FEABD7AAD57AEBA08517DE00AAAEA8A9200249056D4175C5092AA",
INIT_2D => X"FEDB42028EBFBC2028BED152438AAA092492AAA4954281C0E2FB55B6A0925D70",
INIT_2E => X"A0875EDA80BEF1C743840040017D5520B8EAA007FC51C7007BD55D7BE80004AA",
INIT_2F => X"55FFF5D0438140E2FA38B6AEBFF6DBE84AAEBAF7DF6AA00412EAABFFAA803DEB",
INIT_30 => X"1EF0800154B200000000000000000000000000000000000000000000041002FB",
INIT_31 => X"0145AAFFFFFEF5D7FEABFF0051400A25D5568A00FFFFEAA105D5155410FF8402",
INIT_32 => X"2AAA25555410BA082E8201000043FE005D517DEBA0851574B2AAAEAAB55F7840",
INIT_33 => X"4001FF005575408AA557FEB2FFAE975EF555168B55F7AA800BAF7AA955EF0004",
INIT_34 => X"2ABFF55F7800015F087FEAA00007FEAB55FAD568AA200557DE00AAAAAAA00080",
INIT_35 => X"87BD6145FAAC000A2A6FBC00BAAAFBC00BAF7D1550AAAA8002010F2AC154B25F",
INIT_36 => X"082EA8BFFAA843FEBA08517DE00F3F9574B30800021EF55042AAAA007FD55550",
INIT_37 => X"000000000008003FF55F7D5420BA5D2ABFEAAF7AEBDFF779A82AA43F7FBE8A00",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000200000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(4),        -- Port A data input
DOA(0)   => data_read_a_lo(4),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(4),        -- Port B data input
DOB(0)   => data_read_b_lo(4),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_5_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50DF4A0791B3FCB694379283C81FD996A091832102004A337A20E07C0C1E006",
INIT_01 => X"294014468000A04D5C6A60000C34C24841280A00084000C8C212892EEAD53235",
INIT_02 => X"50AE41540CA1D9100002171C1F0A5171134E2A200D8633F8CD09DBFBBB970E7C",
INIT_03 => X"214E3C521D16021B64430CC51C45B8154689094241898749920842946B90010A",
INIT_04 => X"A2F20F7D7A314CB5C208E28A1BF0224A448920028A185340D0C20B2690000C22",
INIT_05 => X"7520B430B20B984809A8886E230C6106371146E1829941C58310402C600381CF",
INIT_06 => X"9CC96CD7C63A7495B9A356ACBC4601C57FD44F8549A46490261C4B39203F7080",
INIT_07 => X"12A88800B029E0C0A12C4B92AA36A2111167357C220095F3C8952A2E5D26F078",
INIT_08 => X"F3F00503B4AE105B534711820C0C0A1043080300F7E0E728B1829C2FEA0A95A1",
INIT_09 => X"C5184F084136848C9298A8560688F480C58858449026145B3830F40944906234",
INIT_0A => X"50EB4124D2B3902BF5C9700C1199DCA84DF46A974F92C7E28F1630D38088A438",
INIT_0B => X"B3144E5636E3178C86B8CC6B8CA6B8CE6B8C86B8CE6B8CA6B8CC15C6435C670C",
INIT_0C => X"79E51E70E070AA8132252008360A7E91504104C8948047D6B0AE1FE440B28A71",
INIT_0D => X"05F0FE40014090400400080329FF8089FF49611F589765923E139F09C78CE7C6",
INIT_0E => X"05F0FE64037FFD7857418407157797878F005F0DFF0F8005F0FE205F0DFF0F80",
INIT_0F => X"8F87FCB1F8053FDEB9B34E0700461E5FF8205F29FF0F8005F0FE205F29FF0F80",
INIT_10 => X"C0184D07C1FF55C3E3E0037FFCF8D3C03009C3CFD53C7E001FF2FAF89781C011",
INIT_11 => X"4E0CDF47186104C6FF177BD939024189BF900401165D645CEEF5BBCDF148F980",
INIT_12 => X"6397F64AEF7F2320483137F8A9BF8A30C2098DFCA06FFFE01F80001F81FDC94F",
INIT_13 => X"FFD051E01015C3BF553D3E0E5FFE838381840714F9DB4F4FA213F774A0E07002",
INIT_14 => X"8B652E2B3120C81284641D3E8DBF7D636FE070189500125C1F83FBCC4F4F80EF",
INIT_15 => X"E7394E339CE138CE5394E33D4E1E0E30E1208C251134921C12A44103F064014B",
INIT_16 => X"7384E3394E338CE538CE1394E3384E738CE139CE1394E7384E339CE139CE5384",
INIT_17 => X"38CE139CE1384E7384E7394E3384E738CE539CE139CE538CE5384E3394E7384E",
INIT_18 => X"7F7B9DB7FF3A1B6DB7ED438A9C3124B2DA6924965B4D384E7384E339CE138CE5",
INIT_19 => X"FBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEF9F7CFDFDDCF3CF3DF5E5BB4E",
INIT_1A => X"7BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEFBEFBEFBEFBE",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE000000000000118D27BBDDEEF77BBDDEEF77BBDDEEF7",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"E955450055421FFFFFBC0010AAD5574BA557FFDFFF0000000000000000000000",
INIT_22 => X"D5575EF55517FF5500557FE10FFFBEAA10007FD7410FFAA97410082A800AAAAA",
INIT_23 => X"FAA955EFA2D168B55557BEAB55005542000007FD74000055574BA5D7FD7555A2",
INIT_24 => X"007BC00AAAAAEBDF45A28428B45FFD168BFF00002AABA5D2ABFFFFAA843DF55F",
INIT_25 => X"AFF80174BAAAD1555EF5555555550055574105D2A800AA00043FEBA5D7FEAA00",
INIT_26 => X"FFAA8415555087BFFF55A2AA800BAFFAE95555080028A00A2FFFDE00F7D57FEB",
INIT_27 => X"545557BC00AAA2FFEAAAA082A97545F7D5420BA5D2E821FFA2D5554BA557BD75",
INIT_28 => X"000000000000000000000000000000000000000000517FE10AAAAA8AAA002E97",
INIT_29 => X"9043D0824850B8A2AE9756D145B401FFFFFFC7010BEDF524AA5571FDFEF00000",
INIT_2A => X"1524BA5571D757DB6D5525EF555178F6D145178E00EBFBE8A101475D5400F7A4",
INIT_2B => X"24BFFFFA28E3AF55F7A0925D7AADB6FB7D5D7FEAB7D0855420BA1471D7438085",
INIT_2C => X"0043FE925571EFA380871C7028B6AEBDF45B68A28B6DEBDF6DBEF1C0A28AAA55",
INIT_2D => X"A2FBF8E10EBD578EAAFF8415482BED1555EF55555057D145152428492E800820",
INIT_2E => X"FB6DF574A85575C55EFBE8E1557D1475FAF45BEAA800AAFFAA9557D080038AAA",
INIT_2F => X"00AAAEA8A9200249056D4175C50920875FDA381C209256DFFDF420BA552A821F",
INIT_30 => X"0BA55557DFF700000000000000000000000000000000000000000000008517DE",
INIT_31 => X"AA105D5155410FF84020AA0800154B2AAAA975FF5D7BC21EFF7FBD7400F7FBC0",
INIT_32 => X"400A25551554BA0051400BA5551575EFF7D1401FF5D5568BE7555568A00AAFFE",
INIT_33 => X"FFDFFF552EA8AAA55043DFF7AAAEAAB55F78400145AAFFFFFEF5D7FEABFF0051",
INIT_34 => X"55400BA082E8201000043FE005D517DEBA0851574B2FFAABFF45FFAAAABFFAAF",
INIT_35 => X"7AA955EF00002AAA2A2FBE8A00A2D16AAAAFF8002410FFD5575EF5555421E755",
INIT_36 => X"FFFFC00BA552A821EFFFFFD74BA5D51575F7FFAE975EF555168B55F7AA800BAF",
INIT_37 => X"000000000000557DE00AAAAAAA000804001FF0055554088A557FEB25D00021FF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000C00000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(5),        -- Port A data input
DOA(0)   => data_read_a_lo(5),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(5),        -- Port B data input
DOB(0)   => data_read_b_lo(5),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_6_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10800B0061A01002840002C03002818000402322520070B313301C4389B2082",
INIT_01 => X"274008482009404C18A160000C52424841000000090800090210000008510200",
INIT_02 => X"102430600C800110000006100009D070012408000000000648080000001210E0",
INIT_03 => X"000200501D1D02140C420200480140040608010040400104681A0084490C4802",
INIT_04 => X"404402820021000A00824002141000980500000808001114C000080624600600",
INIT_05 => X"120024204209981001A806500304610528000500000080000000300000012940",
INIT_06 => X"2000440832280002300010209C4400142061207A024008900008000220600220",
INIT_07 => X"130C8A220FF41F00902008808800182001020150000001F0800408264000100A",
INIT_08 => X"001BF002C4A01041B1120101000010128568837F04842B080020890008080342",
INIT_09 => X"011847140126805432A62A1596C8B5DF10000008900000100220C00084000008",
INIT_0A => X"44EB4104D09392053589F11C59898888454010830212C54081000410A0088C00",
INIT_0B => X"B0044245B25B456C0096C0096C4096C4096C2096C2096C6096C444B6004B600C",
INIT_0C => X"09040020280010000B3002820110101D0012402CC00802410C26800860070621",
INIT_0D => X"0500819D0000900208201040C4007920004884080000448C281018100C000200",
INIT_0E => X"05008182100000000000000000022AE800C00004000000050081A00004000000",
INIT_0F => X"0002330006000000080000000000000D07A00020000000050081A00020000000",
INIT_10 => X"0000000001204A340002100000000000000000020F4001400000020000000000",
INIT_11 => X"019300020000000068D08000200000001A692121000280000000000010000000",
INIT_12 => X"000201FA100400000000034696010000000000D3478000000000000001003F00",
INIT_13 => X"00000000000000043C0001C0A000008000000000012E000054AC000020000000",
INIT_14 => X"0200000040A410C2810800016000809400001000000000000000433300007600",
INIT_15 => X"060180400000008060180404002AC0200208940041309210B28048180F028000",
INIT_16 => X"2008000100601802000000100601800000000180600800000020180600000000",
INIT_17 => X"0180600000008040100200800000060100000802010040180200002018040100",
INIT_18 => X"7F8FF0F4FA955F7CF7F40A80907638C31C71C718638E00006018040080200004",
INIT_19 => X"38E38E38E38E38E38E38E38E38E38E38E38E38E39B6CEDECDDF7DF7DF5F78BCE",
INIT_1A => X"3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE38E38E38E38E",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFF000000000000196A03F9FCFE7F3F9FCFE7F3F9FCFE7F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"00000000000000000000000C0FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"BFDF45F7AA974AAAAAA97555F784174BAF7D5555FF0000000000000000000000",
INIT_22 => X"FBD7410AA8428AAAAAAE955450055421FFFFFBC0010AAD5574BA557FFDFFF087",
INIT_23 => X"FFBEAA10007FD7410FFAA97400082A800AA08515555508043FE00F7AA97555A2",
INIT_24 => X"55517FF55A2AA97400552AAAB45082E80155F7D1575EFFFAA9555500557FE10F",
INIT_25 => X"FF7AAA8A10082EAAB45A2FFC2000007FD74000055574BA5D7FD7555A2D5575EF",
INIT_26 => X"FFAA843DF55FFAA955EFA2D168B55557BEAB5500554200000003DE10FFD5401F",
INIT_27 => X"BFF00002AABA5D2ABFFFF087BD5545007BFDE10AA803FE105D516AABAFF843FF",
INIT_28 => X"0000000000000000000000000000000000000000AAAEBDF45A28428B45FFD168",
INIT_29 => X"524AA5571FDFEF1C7BFFF55FFA095482B6A49256DEB84104BAFFD1525FF00000",
INIT_2A => X"03DE28F7A49057DAAF5D2428A2842AAAAA2AE9756D145B401FFFFFFC7010BEDF",
INIT_2B => X"A49756D145178E00EBFBE8A101475D5400F7A4904380824850381C5B5057D1C0",
INIT_2C => X"571D757DB6D5525EF555178F6DAAA495428412AAFB451C2A8017DE3DF525FFFF",
INIT_2D => X"1C0E3FE00E3DB471EFE3AAAAA00082EA8B6DA2F1C50381471D74380851524BA5",
INIT_2E => X"049516AAB8FF8428FEFA28E3AF55F7A0925D7AADB6FB7D5D7FEAB7D0855420BA",
INIT_2F => X"45B68A28B6DEBDF6DBEF1C0A28AAA5524BFFFF1C7BD057D1C71FFE10A28038E1",
INIT_30 => X"0AAFFD1401E7000000000000000000000000000000000000000000000B6AEBDF",
INIT_31 => X"21EFF7FBD7400F7FBC00BA55557DFF7557BFDF55F78017400F780001FFAA8400",
INIT_32 => X"154B2557FC01EF55043FEAAFF80021EFA2D1420BAAA8428AA2AAAA975FF5D7BC",
INIT_33 => X"A821EFAAFBC01FFF780155F7555568A00AAFFEAA105D5155410FF84020AA0800",
INIT_34 => X"51554BA0051400BA5551575EFF7D1401FF5D5568BE7AA80174AA082ABDF555D2",
INIT_35 => X"D7FEABFF0051400A25D2EBFE10AAFFD55EFA2AEA8A10082EA8BEFAAD5554B255",
INIT_36 => X"55557DE00AA842AA0000516AABAFF8428BE7AAAEAAB55F78400145AAFFFFFEF5",
INIT_37 => X"0000000000FFAABFF45FFAAAABFFAAFFFDFFF552EA8AAA55043DFF7557BC01EF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000900000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(6),        -- Port A data input
DOA(0)   => data_read_a_lo(6),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(6),        -- Port B data input
DOB(0)   => data_read_b_lo(6),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_7_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10844B00482258A2842112C02450418800002300500030B313300C418992002",
INIT_01 => X"234008422008604D1C20E0000E11426840000000080000080200090000110204",
INIT_02 => X"1025207000B08910000206101188D03080144880010400044808000000122160",
INIT_03 => X"000200401914821004420000CA01000C0600010000605114291A008449484802",
INIT_04 => X"40440200002100080006500210101019040000000B085024D842080244000000",
INIT_05 => X"1A8024200009981001A8224001040104200204000000800CC2092CE4A0004900",
INIT_06 => X"A000440822280002340010209C040014A061200052500810000C490323208E28",
INIT_07 => X"128802020028000890240980A809102001020140000009F0800408264000100A",
INIT_08 => X"001A0602C4A01051B13281010408881203480200448423199046821008082351",
INIT_09 => X"336784144126811054809C1040140A001C8648481000045903318B80A400310A",
INIT_0A => X"000800009010100014114110312388984502148282A08415B032095048008100",
INIT_0B => X"20CDC1C483484D201192011920119201192051920519205192074C9018C90188",
INIT_0C => X"D8A5B44001D2C12901228F82F005310D293054048A2212004466000DA1908528",
INIT_0D => X"800F8108A0D09802082010408580008000000008C85264010816851B428DA146",
INIT_0E => X"800F81321000020000261900E28A204040E000A0000007800F814000A0000007",
INIT_0F => X"7072024807000020400000581C01C1A406400084000007800F81400084000007",
INIT_10 => X"060180E83800E820101210000200000CC3003C32080201C0000C000000160700",
INIT_11 => X"81DD00804086423120B74020023090644840A34000828800000004000420020B",
INIT_12 => X"1C6A0186E8000446120C8905BA0004810C84624237E00010001878007F0030C0",
INIT_13 => X"00080208E4083C44230201AEE0010040261900E30520C0806EAC0082000984C0",
INIT_14 => X"0121011088A600C032128201519480D40005802448160403E0700622C0806EE8",
INIT_15 => X"A1685A1685A168DA368DA36CDA30DA13A108810111349A943AA4401000928A19",
INIT_16 => X"368DA768DA1685A1685A5685A368DA368DA7685A1685A1685A768DA368DA368D",
INIT_17 => X"685A1685A169DA368DA1685A1695A368DA3685A1685A168DA368DA1685A1685A",
INIT_18 => X"00000000000000000000400A8448410400020820800069DA1685A168DA369DA3",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000003667B000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"0155EFAAAEA8ABAAAFBFDE0055556AA005D04155550000000000000000000000",
INIT_22 => X"556AA00FFAE95555087BFDF45F7AA974AAAAAA97555F784174BAF7D5555FFF78",
INIT_23 => X"055421FFFFFBC0010AAD5574BA557FFDFFF5555555EFAAFFFDFEFAAAAAAB455D",
INIT_24 => X"AA8428AAA557BFDFFF55003DFFFF7FBEAA00002EAAAAA082EA8A00AAAE955450",
INIT_25 => X"0552EBDE00007BEAAAAA2D14000008515555508043FE00F7AA97555A2FBD7410",
INIT_26 => X"FF00557FE10FFFBEAA10007FD7410FFAA97400082A800AAF7AE975FFA2800001",
INIT_27 => X"155F7D1575EFFFAA955555D51574AAAAFFD5545087FEAB455D516AB55557BD55",
INIT_28 => X"0000000000000000000000000000000000000000A2AA97400552AAAB45082E80",
INIT_29 => X"104BAFFD1525FFFF8E175C7A2AAAAA82A2F1FAE105D556AA10410E1755500000",
INIT_2A => X"1FFFD7AAAAAFB7D495F6AA10E3AE905551C7BFFF55FFA095482B6A49256DEB84",
INIT_2B => X"2EAAA00A2AE9756D145B401FFFFFFC7010BEDF524AA5571FDFEF415B575D7AAF",
INIT_2C => X"7A49057DAAF5D2428A2842AAAA497BFAFFF49003AFEFEBFBEAA001C2EA8A821C",
INIT_2D => X"F7A4905C7A28A070384120BDE100075EAA82BEDB470101C5B5057D1C003DE28F",
INIT_2E => X"D555F6AB57417BC05D7145178E00EBFBE8A101475D5400F7A490438082485038",
INIT_2F => X"28412AAFB451C2A8017DE3DF525FFFFA49756D495150492BEF1D2555087BE8B7",
INIT_30 => X"A10002E9754D000000000000000000000000000000000000000000000AAA4954",
INIT_31 => X"7400F780001FFAA84000AAFFD1401E7FFAA97555A2AEA8A10AAD568A00555168",
INIT_32 => X"7DFF7007BD5555AAD57DF55AAAEBDFEF007BE8A10AAAE8215D557BFDF55F7801",
INIT_33 => X"FEAA105D2EAAA005D2AAAA18AAAA975FF5D7BC21EFF7FBD7400F7FBC00BA5555",
INIT_34 => X"7FC01EF55043FEAAFF80021EFA2D1420BAAA8428AA2007FE8BFF080028BFFAAF",
INIT_35 => X"F84020AA0800154B2FF8402145A2AA954AA00043DE0000516AA10F7FBD740855",
INIT_36 => X"FFD140145007FE8BEF557BEAB55087FC215D555568A00AAFFEAA105D5155410F",
INIT_37 => X"0000000000AA80174AA082ABDF555D2A821EFAAFBC01FFF780155F7005140000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000000FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(7),        -- Port A data input
DOA(0)   => data_read_a_lo(7),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(7),        -- Port B data input
DOB(0)   => data_read_b_lo(7),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_8_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00000648E2840112C00000418000002700500030B3132000400812086",
INIT_01 => X"214009C21838284D042100000212026840000000180800080200080040510204",
INIT_02 => X"1021004000900110000006100088503000240800014400004808000000122160",
INIT_03 => X"0002004019110214044A82000121400C86000000000000860188008448400002",
INIT_04 => X"000402800031200A0000090214100889A5000000490090104800000224000400",
INIT_05 => X"10C025204289981000A820500344010428008500010080080909304040202004",
INIT_06 => X"8000440003280000340010208C04003420600000C6180810000C490703200010",
INIT_07 => X"130002000028000890240980A809012001020050000009F08004082640000082",
INIT_08 => X"20100402C4201041310041010008801201480200051023090024811008090A1A",
INIT_09 => X"0100001001248100308214528148A48008000008100004590711C04034000083",
INIT_0A => X"10804000801210140001C0103001088845010482004000008420041020008900",
INIT_0B => X"0004404002004400448000480004800048000480004800048000440022400200",
INIT_0C => X"880420000880204909004502D100A10C04205424010216010C26800805000004",
INIT_0D => X"8000801100509802082010400400018000488428800004082014000200010000",
INIT_0E => X"8000800A00000207A8BE7B00000200082040808000F07F80008000808000F07F",
INIT_0F => X"0002000402100000404CB1F8FC0000040000808000F07F80008000808000F07F",
INIT_10 => X"3E07800000004004080A000002072C3FCF0000020040804800040007687E3F00",
INIT_11 => X"10800018639EC00020100002C2F9B0000801016001008100000040120CB3067F",
INIT_12 => X"000200020000585EB6000100800030C73D8000402000001FC07FF80001000080",
INIT_13 => X"002EAE1FEC0000040200408000003C547E7B00000100801004000803551F8FC0",
INIT_14 => X"00000000440610C8000A808040000208901B86E568FE0C000000020080100400",
INIT_15 => X"0040100401004090240902449028D0230249850101349A98BAC0481000888810",
INIT_16 => X"0401004010040100401004010240902409024090240902409004010040100401",
INIT_17 => X"4010040100409024090240902409004010040100401004090240902409024090",
INIT_18 => X"543EBC57A10A1E75D6440A889050000000000000000040902409024010040100",
INIT_19 => X"79E79E79E79E79E79E79E79E79E79E79E79E79E7BF3CCD8DF5B2DB2CA4028A0A",
INIT_1A => X"4F87D3E1F4F87D3E1F4F87D3E1F4F87C3E1F0F87C3E1F0F87C3E79E79E79E79E",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000000D3E94F87D3E1F4F87D3E1F4F87D3E1F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"000000087BEAA10F7803DE00FFAEBFFFF0800155FF0000000000000000000000",
INIT_22 => X"7FC2145005155555F780155EFAAAEA8ABAAAFBFDE0055556AA005D0415555080",
INIT_23 => X"7AA974AAAAAA97555F784174BAF7D5555FF552AA8AAA557FC0010F780154105D",
INIT_24 => X"FFAE95555AAFFE8A00552EBFE00F7D17FF45F7FFFFF55AA80155FF087BFDF45F",
INIT_25 => X"5F7D140010552E821EFAAAABDF555555555EFAAFFFDFEFAAAAAAB455D556AA00",
INIT_26 => X"00AAAE955450055421FFFFFBC0010AAD5574BA557FFDFFF5504000AAAAAAA8B5",
INIT_27 => X"A00002EAAAAA082EA8A00002AA8A10F78402155AA8028A00A2D57FF45557BE8A",
INIT_28 => X"0000000000000000000000000000000000000000557BFDFFF55003DFFFF7FBEA",
INIT_29 => X"6AA10410E17555080E000280071E8A00EB8E3FE10F7AEBAFFF080A175D700000",
INIT_2A => X"1C2000FF8A17400557FC015514555757DFF8E175C7A2AAAAA82A2F1FAE105D55",
INIT_2B => X"8A105D71C7BFFF55FFA095482B6A49256DEB84104BAFFD1525FF492EA8AAA557",
INIT_2C => X"AAAAFB7D495F6AA10E3AE90555A2FBE8A38492ABDE10EBDF7AF6DE3FFF8F7DB6",
INIT_2D => X"550E00082B6A0AFB55F7D1420104124821D7AAA0BDF6D415B575D7AAF1FFFD7A",
INIT_2E => X"0B6D578F6D557FFDA00A2AE9756D145B401FFFFFFC7010BEDF524AA5571FDFEF",
INIT_2F => X"FF49003AFEFEBFBEAA001C2EA8A821C2EAAA001C2EA8A00F7800017DA2842FA0",
INIT_30 => X"BEF082E95545000000000000000000000000000000000000000000000497BFAF",
INIT_31 => X"8A10AAD568A00555168A10002E9754D082E820BA08556AA00AAAABFE00F7AEAA",
INIT_32 => X"401E7082EAAABA5D5140010F7AE974105D7BC21555D51575EFFFAA97555A2AEA",
INIT_33 => X"BEABFFAAFBEABFFF7AA80145557BFDF55F78017400F780001FFAA84000AAFFD1",
INIT_34 => X"7BD5555AAD57DF55AAAEBDFEF007BE8A10AAAE8215DA2FFE8ABA082ABFE00AAF",
INIT_35 => X"7FBC00BA55557DFF75D2E82010F7843DF45FFD540000000402145AA843FFFF00",
INIT_36 => X"F780021FFA2803DE10FFD16ABFF5D7BFDE10AAAA975FF5D7BC21EFF7FBD7400F",
INIT_37 => X"0000000000007FE8BFF080028BFFAAFFEAA105D2EAAA005D2AAAA185D2AAAA10",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000400000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(8),        -- Port A data input
DOA(0)   => data_read_a_lo(8),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(8),        -- Port B data input
DOB(0)   => data_read_b_lo(8),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_9_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000B0001800002840002C0000281800000030000000033022000000000002",
INIT_01 => X"8000098218302849180060000C004240413C0A61590001D90213C90008510200",
INIT_02 => X"000008700CB089100002061031200074810448800104008048080080001210E2",
INIT_03 => X"000200140C1822000A028010408100000628000140402080041A100040024840",
INIT_04 => X"41040000000400080002040200080800040000000B08D1055842080604600700",
INIT_05 => X"10002024000020102400010000026104200004000400800C8B0024E4E0010C40",
INIT_06 => X"8000440802280002700800008A840004A0610000C0000810000C590103600810",
INIT_07 => X"538600220028001890240980A80800200102025000000BF08200002440000883",
INIT_08 => X"00000402C220104131102101040810028528820005100003900E884000010007",
INIT_09 => X"00000005E000000600BCA284140200800C834948100004590111824404012080",
INIT_0A => X"04080000901012100A1141005922000245410002008880000032005080000800",
INIT_0B => X"2000020040044010440104401004010440100401044010040104400802008208",
INIT_0C => X"D1A1344420D2E100000808000000000481000000202002400006800825908402",
INIT_0D => X"0500000000109000000000000580008000080000C852240100068D0B4685A342",
INIT_0E => X"0500000A00000000000000000000028000408020000000050000208020000000",
INIT_0F => X"0000304002100020000000000000000900208004000000050000208004000000",
INIT_10 => X"0000000001200000000A00000000000000000000050000480008000000000000",
INIT_11 => X"009F0080000000004807C0200000000012000020000081000000040000000000",
INIT_12 => X"00000048F8000400000002403E0004000000009067E000000000000000000900",
INIT_13 => X"0000000000000000140000CEE001000000000000000A000036AC008000000000",
INIT_14 => X"03210000000400CA81000000619480D4000400000000000000004100000036E8",
INIT_15 => X"A368DA368DA3685A1685A1685A121A11A1419001512490040024001000008019",
INIT_16 => X"1685A1685A1685A1685A1685A368DA368DA368DA368DA368DA368DA368DA368D",
INIT_17 => X"685A1685A168DA368DA368DA368DA368DA368DA368DA3685A1685A1685A1685A",
INIT_18 => X"CCF48DE68A895C38E250080000000000000000000000685A1685A1685A1685A1",
INIT_19 => X"514514514514514514514514514D34D34D34D34D28E10040392482090157344C",
INIT_1A => X"4D268341A0D069349A0D069349A0D068341A0D068341A0D06834514514514514",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000001654D0D069349A0D068341A4D268341A",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"BE8B45002A974AAAA803DFFFAA843DF45FFFFEAABA0000000000000000000000",
INIT_22 => X"AEBDE00AAFBEAABA080000000087BEAA10F7803DE00FFAEBFFFF0800155FFAAF",
INIT_23 => X"AAEA8ABAAAFBFDE0055556AA005D0415555087BFDE00A2FBD7400F7FBFDFFFA2",
INIT_24 => X"005155555557BE8BEF007FFDEAAAAD1555EF0055401FFF7AEAAA10F780155EFA",
INIT_25 => X"0F7AA974AA082E80010A2AAAAA10552AA8AAA557FC0010F780154105D7FC2145",
INIT_26 => X"BA087BFDF45F7AA974AAAAAA97555F784174BAF7D5555FFF780154AA5D2AA8A1",
INIT_27 => X"F45F7FFFFF55AA80155FF080400145FFFBEAABAF7D17FEBAA2AEBDF45002EAAA",
INIT_28 => X"0000000000000000000000000000000000000000AAFFE8A00552EBFE00F7D17F",
INIT_29 => X"BAFFF080A175D7BEF1E8B6D002090482B68E38FC7BE8A3DF7DF7F5E8A9200000",
INIT_2A => X"BD0400FFF5FDFC7B6A0BDE38B6F5E8A92080E000280071E8A00EB8E3FE10F7AE",
INIT_2B => X"AAA8A38FF8E175C7A2AAAAA82A2F1FAE105D556AA10410E175550871FFE00A2F",
INIT_2C => X"F8A17400557FC015514555757D5D71E8BEF147BFAE82A2DB555C71C5B451D7FF",
INIT_2D => X"FF84174BA5D20AAA00E3AA904BA142A87010A2AEADA38492EA8AAA5571C2000F",
INIT_2E => X"AAAA0BFF7D0024ADA921C7BFFF55FFA095482B6A49256DEB84104BAFFD1525FF",
INIT_2F => X"38492ABDE10EBDF7AF6DE3FFF8F7DB68A105D7000400155FFFBEDA82FFD57DEB",
INIT_30 => X"FEFF7D16AA00000000000000000000000000000000000000000000000A2FBE8A",
INIT_31 => X"AA00AAAABFE00F7AEAABEF082E95545F7D568BEF080402000F7AAA8B55FFAABD",
INIT_32 => X"9754D00517DE00A2FFC2000F7D17FF55FF803FEAAFFD16AA00082E820BA08556",
INIT_33 => X"FD55555D7FD5555FFAAA8AAAFFAA97555A2AEA8A10AAD568A00555168A10002E",
INIT_34 => X"2EAAABA5D5140010F7AE974105D7BC21555D51575EF555568BEF5D7FE8A10AAF",
INIT_35 => X"A84000AAFFD1401E7FF80174AA5D0028A00AAAE800AA552A97400A2AEBDEAA08",
INIT_36 => X"F7FBFFE00FFD17FEAAA2803DFEF08043FE00557BFDF55F78017400F780001FFA",
INIT_37 => X"0000000000A2FFE8ABA082ABFE00AAFBEABFFAAFBEABFFF7AA80145080002145",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000800000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(9),        -- Port A data input
DOA(0)   => data_read_a_lo(9),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(9),        -- Port B data input
DOB(0)   => data_read_b_lo(9),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_10_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000B0001800002840002C0000281800020030000000033022000000180006",
INIT_01 => X"000008000000004C002000000010026840000000080000080200000000110200",
INIT_02 => X"0000004000800110000006100000003000040800010400004808000000120060",
INIT_03 => X"000200000810020000020000400100000600000000400000001A000040004800",
INIT_04 => X"0004000000000008000200020000000004000000080010004000000200000000",
INIT_05 => X"1000202000011010000000000000010520000400000080000000200000200004",
INIT_06 => X"80004408022800023000000088040004A061000040000810000C490103600000",
INIT_07 => X"120420020028000890240980A808002001020050000009F08000002440000082",
INIT_08 => X"00000402C0201051311001000000020201080200440400000000800000000000",
INIT_09 => X"0000105808000000000000000000008000008088100004590111800004000000",
INIT_0A => X"00804000801210440003C1411008800045000002000014000040009002800000",
INIT_0B => X"0400200000000000000004000040000000000000040000400000000000000221",
INIT_0C => X"0100802000000000000002802000000400100000000002000026000840011400",
INIT_0D => X"0500000000409002082010400400008000400008002044082000081004080204",
INIT_0E => X"0500000200000000000000000000028000400000000000050000200000000000",
INIT_0F => X"0000304002000000000000000000000900200000000000050000200000000000",
INIT_10 => X"0000000001200000000200000000000000000000050000400000000000000000",
INIT_11 => X"0082000000000000480080000000000012000101000080000000000000000000",
INIT_12 => X"0000004810000000000002400400000000000090400000000000000000000940",
INIT_13 => X"0000000000000000150000C00000000000000000000A40001400000000000000",
INIT_14 => X"02000000002400C2810000006000000000000000000000000000410040001400",
INIT_15 => X"020080200802008020080200800800220200840001309A08A848001000008000",
INIT_16 => X"0000000000000000000000000200802008020080200802008020080200802008",
INIT_17 => X"0080200802000000000000000000000000000000000000000000000000000000",
INIT_18 => X"940FE0D397124355520542821010000000000000000000802008020080200802",
INIT_19 => X"28A28A28A28A28A28A28A28A28A28A28A28A28A29554199854514514F546890A",
INIT_1A => X"32994CA6532995CAE572B94CA6532994CA6532994CA6532994CA28A28A28A28A",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000001867172B94CA6532994CA6572B95CAE5",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FC2155F7D155545AA80001EFAAFBEAB45557FFDE100000000000000000000000",
INIT_22 => X"FBE8BFFF78402155AAFBE8B45002A974AAAA803DFFFAA843DF45FFFFEAABA007",
INIT_23 => X"87BEAA10F7803DE00FFAEBFFFF0800155FF00042AB55FFD168B55AA8000010FF",
INIT_24 => X"AAFBEAABAA2FFD741055003DFEFF7AA801FFAAD16AABA002ABDE100800000000",
INIT_25 => X"FF7FBC0145F78028A00A2D142155087BFDE00A2FBD7400F7FBFDFFFA2AEBDE00",
INIT_26 => X"BAF780155EFAAAEA8ABAAAFBFDE0055556AA005D0415555007FD74105555555E",
INIT_27 => X"5EF0055401FFF7AEAAA105D042ABFF5D556AB55AAD168ABA002A975FFF7AEBDE",
INIT_28 => X"0000000000000000000000000000000000000000557BE8BEF007FFDEAAAAD155",
INIT_29 => X"3DF7DF7F5E8A92007BC217DEBDB55555AA8E071D7AAFBEFB455D71F8E0000000",
INIT_2A => X"B6DB55BE8E05000EBFFE8BC7E38E07145BEF1E8B6D002090482B68E38FC7BE8A",
INIT_2B => X"2EB8E00080E000280071E8A00EB8E3FE10F7AEBAFFF080A175D700042AB7DEBD",
INIT_2C => X"FF5FDFC7B6A0BDE38B6F5E8A92B6FBD5410490A3DFD7F7A4821D7A2D16FA8214",
INIT_2D => X"0071D54104951555D7EBF5C5155E3842AA00BED1421450871FFE00A2FBD0400F",
INIT_2E => X"20820955EFE3AEBDEAAFF8E175C7A2AAAAA82A2F1FAE105D556AA10410E17555",
INIT_2F => X"EF147BFAE82A2DB555C71C5B451D7FFAAA8A38410E2ABD749516FB55BED16FA8",
INIT_30 => X"F455D556AA000000000000000000000000000000000000000000000005D71E8B",
INIT_31 => X"2000F7AAA8B55FFAABDFEFF7D16AA00087FC01EFA2FFD7545AAAE97555A2FBFD",
INIT_32 => X"9554500042ABFFA2FFFFF45F7AE97400AAFFE8B45AAAA95545F7D568BEF08040",
INIT_33 => X"400155A2D57FE00552EA8A00082E820BA08556AA00AAAABFE00F7AEAABEF082E",
INIT_34 => X"517DE00A2FFC2000F7D17FF55FF803FEAAFFD16AA00FFFBD5400082EBFF45F78",
INIT_35 => X"55168A10002E9754D085155410085557555AAD557555A2802AA10FFD54214500",
INIT_36 => X"08557DF55F7D17FE000804155FFAAAABDEAAFFAA97555A2AEA8A10AAD568A005",
INIT_37 => X"0000000000555568BEF5D7FE8A10AAFFD55555D7FD5555FFAAA8AAA002AAAB45",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000008FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(10),        -- Port A data input
DOA(0)   => data_read_a_lo(10),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(10),        -- Port B data input
DOB(0)   => data_read_b_lo(10),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_11_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10180B05A0010402840602C2D001019000000300000000330A20080EC180002",
INIT_01 => X"AB400986B830284D1820E0000C3642484000000008000008820009080A512220",
INIT_02 => X"102A68440080011000000618062AD03502640800010410424908136019920868",
INIT_03 => X"004A0846191B22120642000442C110044600000101E9225CDC9A10844A9A4842",
INIT_04 => X"0094024000250808800216021138000B848000000800100040000102A0600200",
INIT_05 => X"7E4024242008A8102CA88A44010401042200444000888000000028000002A002",
INIT_06 => X"8088445712280000B18812288E0400253855200045C86810000C5B0503286A28",
INIT_07 => X"10008822A028004880200A80880208200122006C000015F0C20408264902C840",
INIT_08 => X"9390040280241041D1754100000018108728820024002B3A01A89540080824C8",
INIT_09 => X"A1001C41A1348498B080801010000080D00301081000045B0511D28D94012339",
INIT_0A => X"44080000901012428003414158230CBA4576708241C010908040341322008000",
INIT_0B => X"040464D280144050C72A0872A0C72A0872A0C72A0C72A0872A0C595043950421",
INIT_0C => X"0804001400000820110A42822204880CD81040442900021704E6000800001D54",
INIT_0D => X"80C62D0500409002082010404580018000404012004004192C10000000000000",
INIT_0E => X"80C62D5803161C526DB40506C120A806ABB0D808CC334A80A54B70D408CC32D2",
INIT_0F => X"2B5144D0DD903C54916D15458C0513005570D408CC334A80A54B70D808CC32D2",
INIT_10 => X"52148C4DB05621E363F813961C20EDA944016558C2347A080B10D8DD6422AA10",
INIT_11 => X"1880144D3345C65593800319C18BD1ECA1C9010112566F10AC4183C340DAE02D",
INIT_12 => X"5810503000633830DE3C2C9C00289A66AA8DE50E0800360614AC281430890600",
INIT_13 => X"0CD2A9CEA8199B6B082B55900314140365320485C4F00AD544407241C175C402",
INIT_14 => X"0000074044C4801832701A89D20A38093631425969020855A281844E00540404",
INIT_15 => X"0000000000000000000000000020C00200088101513492101280401000400200",
INIT_16 => X"2008020080200802008020080000000000000000000000000000000000000000",
INIT_17 => X"0080200802008020080200802008020080200802008020080200802008020080",
INIT_18 => X"804180C0B10A4210420140028400000000000000000000802008020080200802",
INIT_19 => X"000000000000000000000000000820820820820801C414947000000055062608",
INIT_1A => X"0000000004020000000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000001F87E000000000000010080000000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"ABDF5508557DF45002ABDFFFF7803DE10AA80000AA0000000000000000000000",
INIT_22 => X"FFE8A10A28000000007FC2155F7D155545AA80001EFAAFBEAB45557FFDE10082",
INIT_23 => X"02A974AAAA803DFFFAA843DF45FFFFEAABAA2AEBFF45FFAEBFEAA002A801FFF7",
INIT_24 => X"F78402155AAD155555A28428BFF002ABDE00A2AABFE10082ABFFEFAAFBE8B450",
INIT_25 => X"0002A80010A2842AAAA007BFFF4500042AB55FFD168B55AA8000010FFFBE8BFF",
INIT_26 => X"00080000000087BEAA10F7803DE00FFAEBFFFF0800155FF00557FF45557FC201",
INIT_27 => X"1FFAAD16AABA002ABDE10A2D168A10A284021FF5D00154BAF7FBE8BEFFFD5400",
INIT_28 => X"0000000000000000000000000000000000000000A2FFD741055003DFEFF7AA80",
INIT_29 => X"EFB455D71F8E00002EBDF6D005B78F7D142ABDFC7F78E3FE28B684070AA00000",
INIT_2A => X"0BDEAA1C2A801C7E3FFEFA10B68407038007BC217DEBDB55555AA8E071D7AAFB",
INIT_2B => X"20B8FEFBEF1E8B6D002090482B68E38FC7BE8A3DF7DF7F5E8A92BEAEBFF7DEBA",
INIT_2C => X"E8E05000EBFFE8BC7E38E07145B6D15756DA28A28BFF082ABAE10B6AAB8E2808",
INIT_2D => X"08517DF7D497BC5028142A87000A28A2AA92007FF8F7D00042AB7DEBDB6DB55B",
INIT_2E => X"2FFFFEFBC7E3DF42028080E000280071E8A00EB8E3FE10F7AEBAFFF080A175D7",
INIT_2F => X"10490A3DFD7F7A4821D7A2D16FA82142EB8E00B6DB6AA28A280001FF5D0A1048",
INIT_30 => X"EAAF784154BA000000000000000000000000000000000000000000000B6FBD54",
INIT_31 => X"7545AAAE97555A2FBFDF455D556AA00082EBFFEF007BE8BFF5D2ABDF55F7AABD",
INIT_32 => X"6AA00FFAEBFFEFAA803DEBA5D2E82155A2FBFDE00FF84154BA087FC01EFA2FFD",
INIT_33 => X"AAAA00FFAAA8AAA080028BFFF7D568BEF080402000F7AAA8B55FFAABDFEFF7D1",
INIT_34 => X"042ABFFA2FFFFF45F7AE97400AAFFE8B45AAAA95545F7D5555FFAAAAA8BFF002",
INIT_35 => X"7AEAABEF082E9554508557DFFF007BD54BA5D2E95400A2AEA8A00007FEABFF00",
INIT_36 => X"AA80001FF5D2E82000F7FFFFF45AAFFC20BA082E820BA08556AA00AAAABFE00F",
INIT_37 => X"0000000000FFFBD5400082EBFF45F78400155A2D57FE00552EA8A00FFFFE8AAA",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000800000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(11),        -- Port A data input
DOA(0)   => data_read_a_lo(11),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(11),        -- Port B data input
DOB(0)   => data_read_b_lo(11),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_12_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"A500C4B01BC0268A6940312C0DE045196A831A300500032B333287E4FC812006",
INIT_01 => X"AF400D869830E84D5823E0000C1742484000000008000008820009280A553235",
INIT_02 => X"502A7144008001100000171C022BD13412762A000586235ECC09C8423B960866",
INIT_03 => X"31863846191BA218064204000281200406A10843010022DEDF0852944A9C014A",
INIT_04 => X"0014030000250409000014821038080B840000400800102040000302F0600233",
INIT_05 => X"7FC034348008A8102CA88F48010601042400048000188000000938000002E088",
INIT_06 => X"9CC96CC6F63A5001F12B56A0AC8601F47AC06400D1F80C10020C493F03343A38",
INIT_07 => X"1020002030280098A12048908A16BA311177124C000003F08A94282E5C262861",
INIT_08 => X"827A0602902A10491165E10000049010C52882008600A73A01E8974008092CF8",
INIT_09 => X"47000001A1248008F000000000000080000F010C100204593F11A6CDF48023BF",
INIT_0A => X"040000208010120ACA01400058010CBA4D277C86CCE802B380003C1360008000",
INIT_0B => X"011C46D3C7BC1EF083AF0C3AF083AF083AF0C3AF083AF083AF0C1D7861D78400",
INIT_0C => X"08040014C9001AE91D17E50AD79FEFC87C2154745F82131FFCCE00080000095E",
INIT_0D => X"807BF7118180984004000803D40001880001001400C005031010000000000000",
INIT_0E => X"807BF76A109C944B5891BF06C5EEB14FCBF0D90076D61C807BF7D0D80876D49C",
INIT_0F => X"6DE38EB9FB10350C00A99F7CA80757365E50D80876D61C807BF7D0D90076D49C",
INIT_10 => X"841BCC69A0D8C6F7F0AA001C943A65756A0976EB5A7E7FC8951018186334F311",
INIT_11 => X"D5A014481991C6A737D80211912970CDCDD1864116D6C7080651CB4661F33615",
INIT_12 => X"349E929300423224AE19B9BEC0289033238D4E6EA805892946A9B011A7B152CF",
INIT_13 => X"6244CD7AC01CAAA56B3E6D9001068715D64006D2A961CF9B44512A2504532182",
INIT_14 => X"00000439FDC25C58067A9FAB46095A0B5289A0282D2E1444ACB12A17CF9B4414",
INIT_15 => X"0000000000000000000000040026C00000288401513492909280401000F70A00",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"088881360A95090CB05442029010000000000000000000000000000000000000",
INIT_19 => X"1041041041041041041041041049249249249249200100002D4514510051B946",
INIT_1A => X"592C964B2592C964B2592C964B2592C86432190C86432190C864104104104104",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000002007F592C964B2592C964B2592C964B2",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"43FE0008557DFFF0800020105D557FEAA00557DE100000000000000000000000",
INIT_22 => X"557DFFFF7AA80000082ABDF5508557DF45002ABDFFFF7803DE10AA80000AAAA8",
INIT_23 => X"7D155545AA80001EFAAFBEAB45557FFDE10AAD5420000051555FFA2AA8200000",
INIT_24 => X"A28000000A2D155410F7FFFFEBA08003FE00082AA8AAAAAFFC00BA007FC2155F",
INIT_25 => X"0A2AABFE1055516ABEF5D517DEAAA2AEBFF45FFAEBFEAA002A801FFF7FFE8A10",
INIT_26 => X"55AAFBE8B45002A974AAAA803DFFFAA843DF45FFFFEAABA000028A105D2ABFE1",
INIT_27 => X"E00A2AABFE10082ABFFEF085542000000417555002A820AA08557DFFFF7AA821",
INIT_28 => X"0000000000000000000000000000000000000000AAD155555A28428BFF002ABD",
INIT_29 => X"3FE28B684070AABE803AE38145B78FD7000005010495B7AE921C517DE1000000",
INIT_2A => X"B505FFB6A487000005F7AFD7F7A482038002EBDF6D005B78F7D142ABDFC7F78E",
INIT_2B => X"F5C2082007BC217DEBDB55555AA8E071D7AAFBEFB455D71F8E00BED547038145",
INIT_2C => X"C2A801C7E3FFEFA10B68407038B6D550428FFF1FDE821C003FE001C2EAAAAAB6",
INIT_2D => X"00002FA285D20BDE28A2A4B8E10555B68BEF5D517DEAABEAEBFF7DEBA0BDEAA1",
INIT_2E => X"2005F7DFD7F7A482155BEF1E8B6D002090482B68E38FC7BE8A3DF7DF7F5E8A92",
INIT_2F => X"6DA28A28BFF082ABAE10B6AAB8E280820B8FEF085F4703814001055514208208",
INIT_30 => X"A0055517DE00000000000000000000000000000000000000000000000B6D1575",
INIT_31 => X"8BFF5D2ABDF55F7AABDEAAF784154BAF7802AABA5D7FEAB45080015410007FEA",
INIT_32 => X"6AA00F7D1554BA5D7BC01FFFF8015410007FEAB45F780020BA082EBFFEF007BE",
INIT_33 => X"43FE10552EAAAAAFFD140000087FC01EFA2FFD7545AAAE97555A2FBFDF455D55",
INIT_34 => X"AEBFFEFAA803DEBA5D2E82155A2FBFDE00FF84154BAF7D1400BAFFD57FE005D0",
INIT_35 => X"FAABDFEFF7D16AA0008003FEBA55003DEBAA28428A105D7FEABEF55557DEBAFF",
INIT_36 => X"550402145550000010087FFFF45F78402145F7D568BEF080402000F7AAA8B55F",
INIT_37 => X"0000000000F7D5555FFAAAAA8BFF002AAAA00FFAAA8AAA080028BFF087BD54AA",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000000FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(12),        -- Port A data input
DOA(0)   => data_read_a_lo(12),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(12),        -- Port B data input
DOB(0)   => data_read_b_lo(12),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_13_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10110A0441812402840402822007818000E00700000000330A3000000008042",
INIT_01 => X"A1400984B830C848180260000C0042604001000008220008A200100802110200",
INIT_02 => X"10A00860009141100000C6180C285035000E0800010431004908135980120C60",
INIT_03 => X"004E20441910221B06420C85D5013804060000000040324C441A108468024842",
INIT_04 => X"0184034010250089C00EA8021938325B04800002091090014880080200000900",
INIT_05 => X"18002424B008881024A8004E01040104270004E0000080090500604840000481",
INIT_06 => X"80004414022A2490B00A142C8C840005794540015E006810001C4B01032C7E20",
INIT_07 => X"510200028028004880280A808816002101022468000011F082040A264006C000",
INIT_08 => X"D2B00402B220104B531001000008001041080200B660E30B200C8040080A9206",
INIT_09 => X"A1000809A93484D21000000000000080C90391881000145B0111A30404015000",
INIT_0A => X"000000008010102A82014100101118BA4510008241480290882400900000A000",
INIT_0B => X"0284484000000000400000000040000000000000040000000000000020000000",
INIT_0C => X"A944AA2000A02000212800020000000D80004084A0000390002E001843210400",
INIT_0D => X"859C1881A04090000000000021800180010341179065441356150A1285094284",
INIT_0E => X"859C188810C65A72A617520252781EA02520D589B9A260859C1840DD81B9A0E0",
INIT_0F => X"0E71F1052D942748C19484E39442D15961C0DD81B9A260859C1840D589B9A0E0",
INIT_10 => X"E60605C0C12CBD400B0810C65A61AA459D0047398500D5889D26907356533C00",
INIT_11 => X"8F60CA1562094650CA28398A42C051E0332181010109294C8E1160CB8C80A561",
INIT_12 => X"2645056D073148580A3C065141942AC4128CA199180C5232575138094450AD0A",
INIT_13 => X"84CA93A2FC008962142B17301A9A1A5196A80245208E0AC5C853C8028163B8C0",
INIT_14 => X"0240034000E4DC8A84000014982372011FC1E475F0F0084A3961F5A80AC5C816",
INIT_15 => X"4250942509425094250942509428D421420882020120981812C8403000088212",
INIT_16 => X"2509425094250942509425094250942509425094250942509425094250942509",
INIT_17 => X"5094250942509425094250942509425094250942509425094250942509425094",
INIT_18 => X"FF3F7DF7FF3E9F7DF7E24502A800000000000000000050942509425094250942",
INIT_19 => X"EBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBF7DFDFDDD555555F7EFBBEE",
INIT_1A => X"7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAEBAEBAEBAEBA",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000000007F7EBF5FAFD7EBF5FAFD7EBF5FAFD",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5554BA087FFFF55557BD54AAF7FBC01FFA2802ABEF0000000000000000000000",
INIT_22 => X"2E80155AA802AB45AA843FE0008557DFFF0800020105D557FEAA00557DE10AAD",
INIT_23 => X"8557DF45002ABDFFFF7803DE10AA80000AA087BD75EF087FFFFEF557BEAB4555",
INIT_24 => X"F7AA80000AAD1420AA087BD7555FFD168AAAFFAE820AA5D5557555082ABDF550",
INIT_25 => X"5FFD157555085140010F7AEAABFFAAD5420000051555FFA2AA8200000557DFFF",
INIT_26 => X"45007FC2155F7D155545AA80001EFAAFBEAB45557FFDE10AAAEA8BFFA2FBD754",
INIT_27 => X"E00082AA8AAAAAFFC00BA00002AAAAF7D5574BA557BE8A10A284154BAFFAAAAB",
INIT_28 => X"0000000000000000000000000000000000000000A2D155410F7FFFFEBA08003F",
INIT_29 => X"7AE921C517DE10A2DB50482147FFAF554971D0492E3F1C71C7BE8A2ABD700000",
INIT_2A => X"FFAFD7497BE8B5555208217DBE8A2AB45BE803AE38145B78FD7000005010495B",
INIT_2B => X"5F5056D002EBDF6D005B78F7D142ABDFC7F78E3FE28B684070AA1C71D25D7007",
INIT_2C => X"6A487000005F7AFD7F7A482038AADF47092147FD257DFFD568A82FFA4870BA55",
INIT_2D => X"A2A0ADBC7A2FFD257DE3DF52555085142000FFAAAFBFFBED547038145B505FFB",
INIT_2E => X"0B680124BAFFAAAFB45007BC217DEBDB55555AA8E071D7AAFBEFB455D71F8E00",
INIT_2F => X"28FFF1FDE821C003FE001C2EAAAAAB6F5C20821C002AA92FFDF574824171EAA1",
INIT_30 => X"545F7AEA8B55000000000000000000000000000000000000000000000B6D5504",
INIT_31 => X"AB45080015410007FEAA0055517DE00A2FFC00105D7BE8B55085142010AAD157",
INIT_32 => X"154BA5D5140145007BE8B55087BEAB555D04001EFF7AAA8B55F7802AABA5D7FE",
INIT_33 => X"16AA10FF80174AA557FC21EF082EBFFEF007BE8BFF5D2ABDF55F7AABDEAAF784",
INIT_34 => X"D1554BA5D7BC01FFFF8015410007FEAB45F780020BAA2FFD54105D7FC21EFFFD",
INIT_35 => X"2FBFDF455D556AA00A2803FF45AAFFC21EFAAFBC0155085540000FFAEBFFEFF7",
INIT_36 => X"F7FBD5410085568A10FF80020AAFFAABFF55087FC01EFA2FFD7545AAAE97555A",
INIT_37 => X"0000000000F7D1400BAFFD57FE005D043FE10552EAAAAAFFD1400005D042AA00",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000CFFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(13),        -- Port A data input
DOA(0)   => data_read_a_lo(13),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(13),        -- Port B data input
DOB(0)   => data_read_b_lo(13),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_14_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10020A000180000284008280000281800000030000000033022000000580002",
INIT_01 => X"A140098018300848184860000C20C24040000000084000084200000000110200",
INIT_02 => X"1020006000900110000006102028503400040800010400204908012018120E64",
INIT_03 => X"000200441910221006420000400100040600000000E9E401209A108448004842",
INIT_04 => X"0004020000250008000200021038000804000000090090004800080200000000",
INIT_05 => X"500024240008881024A800400104010420000400000080080100204040000000",
INIT_06 => X"8000440102282015B10A10288E0400042345400040006810000C5901033D7880",
INIT_07 => X"1100000200280048802008828812002001220064000005F1C2850A2649204070",
INIT_08 => X"00B00402802010411110010000080010010802000400230B000C804008080002",
INIT_09 => X"01000009A92480001000000000000080C8038188100004590111B68404010000",
INIT_0A => X"0000000080101000000141001001088A45000082400000008020009000008000",
INIT_0B => X"0004404000000000400004000000000000004000000000000004000000000000",
INIT_0C => X"8904A0200080200001080002000000088000400420000200002E000841010400",
INIT_0D => X"0500000C80409000000000000000018000000000806044010014081204090204",
INIT_0E => X"0500005813A0210D072E8D012001028402908004000587050000108004000707",
INIT_0F => X"9004300044900812386A280E5800088980108020000587050000108020000707",
INIT_10 => X"DE00482E19E30002007813A02096038AE200880405200308828062A68C0BC700",
INIT_11 => X"00000E5A08E6000048001292B83280001208A1011004011060049A1C59192055",
INIT_12 => X"492060480256530650000240001DB011CC00009000032C4C979E3806180C0900",
INIT_13 => X"5A3433EDE00154181400000007BCBD858F120120541A0000000033757465B2C0",
INIT_14 => X"02002C000024008A84001A0902000422E3E99681004802115652594000000001",
INIT_15 => X"0240902409024090240902409028D021020880000120901812C8401000000210",
INIT_16 => X"2409024090240902409024090240902409024090240902409024090240902409",
INIT_17 => X"4090240902409024090240902409024090240902409024090240902409024090",
INIT_18 => X"5C8FF0F7BE9D5F7DF65040028000000000000000000040902409024090240902",
INIT_19 => X"79E79E79E79E79E79E79E79E79E79E79E79E79E7BF7DDDDDFCF3CF3DF5579B4E",
INIT_1A => X"3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE79E79E79E79E",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000003FF803F9FCFE7F3F9FCFE7F3F9FCFE7F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"BE8B55A2AE80000F7D5555555D2AAAABAAAD1420BA0000000000000000000000",
INIT_22 => X"00155EF0804155EFAAD5554BA087FFFF55557BD54AAF7FBC01FFA2802ABEFA2F",
INIT_23 => X"8557DFFF0800020105D557FEAA00557DE10A2AA801FFA28402000AAAE9554555",
INIT_24 => X"AA802AB4500516AA00A2AE800BAFFFFC20BAF7AEA8B45080417400AA843FE000",
INIT_25 => X"0A2843FEBAFFFBD7410A2D168BFF087BD75EF087FFFFEF557BEAB45552E80155",
INIT_26 => X"AA082ABDF5508557DF45002ABDFFFF7803DE10AA80000AA005568ABAA2840201",
INIT_27 => X"AAAFFAE820AA5D5557555002E80155A280000005D7FFDF4555517DFEF00043FE",
INIT_28 => X"0000000000000000000000000000000000000000AAD1420AA087BD7555FFD168",
INIT_29 => X"C71C7BE8A2ABD7A2FFEDB55B6A080038E3DB50555412AA8ABAAADB4009200000",
INIT_2A => X"402038AAAA955554900105FF0800175D7A2DB50482147FFAF554971D0492E3F1",
INIT_2B => X"0A12410BE803AE38145B78FD7000005010495B7AE921C517DE10A2AE851FFB68",
INIT_2C => X"97BE8B5555208217DBE8A2AB451C556FA00A2A0800BAE3F1C0092EBAAADB6D08",
INIT_2D => X"00516DABAA28402038B6803DE82F7F5D5410A2D568BC71C71D25D7007FFAFD74",
INIT_2E => X"55D5F78FD7000E3FEAA002EBDF6D005B78F7D142ABDFC7F78E3FE28B684070AA",
INIT_2F => X"92147FD257DFFD568A82FFA4870BA555F5056D002A80155B680000105D7FF8F4",
INIT_30 => X"AAAAAFFC2000000000000000000000000000000000000000000000000AADF470",
INIT_31 => X"8B55085142010AAD157545F7AEA8B55A2FBFFF55FF84000AAAAFBC0145002AA8",
INIT_32 => X"7DE00A2AA955FFFF80020BAAAAA975450800001EF080417555A2FFC00105D7BE",
INIT_33 => X"140000A2AEBFFEF082A82010F7802AABA5D7FEAB45080015410007FEAA005551",
INIT_34 => X"5140145007BE8B55087BEAB555D04001EFF7AAA8B555D557FE00A280020BAAAD",
INIT_35 => X"7AABDEAAF784154BA08557FEAAA284000AAFF803DE00FFD557400AAD56AB455D",
INIT_36 => X"F780020105D7BEAB45557BE8B45082EBFEBA082EBFFEF007BE8BFF5D2ABDF55F",
INIT_37 => X"0000000000A2FFD54105D7FC21EFFFD16AA10FF80174AA557FC21EF082A80145",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000000FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(14),        -- Port A data input
DOA(0)   => data_read_a_lo(14),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(14),        -- Port B data input
DOB(0)   => data_read_b_lo(14),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_15_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000A000000000284000280000001800020030000000033022000000180002",
INIT_01 => X"A140098018300848180060000C00424040000000080000080200000000110200",
INIT_02 => X"102100400C8011100000061000A8503401044880010430004808000180122378",
INIT_03 => X"000200541D102210064200000045000546080000400020000008108448400042",
INIT_04 => X"8094020000254C880000028A1018000844000000880013504000002600000000",
INIT_05 => X"10002424000AA81024A82040010C61062001440002988000000024808001004B",
INIT_06 => X"80004400022A00003C8912248E0400042854400040006810000C4901032B1800",
INIT_07 => X"50200000B0280048A0280A828801002101020040000005F38204082640000000",
INIT_08 => X"01F00402802610411100110000000010010802000400230A0008884008080004",
INIT_09 => X"01000001A12481041000000000000080C0030108100004590111820404000000",
INIT_0A => X"0000000080101000004140001001088A45000082000000008000001080008000",
INIT_0B => X"0004404000000000400004000040000400000000000000000004000020000200",
INIT_0C => X"0804000020024100012808020000000981004004A0200310000C000800000000",
INIT_0D => X"0000001180009000000000002100018000000000004004010010000000000000",
INIT_0E => X"00000008000002000000000000000000000080A40000000000000080A4000000",
INIT_0F => X"00000000001000204800000000000000000080A40000000000000080A4000000",
INIT_10 => X"000000000000000000080000020000000000000000000008000C020000000000",
INIT_11 => X"000000824000000000000020220000000001800100020300000004003420480A",
INIT_12 => X"0000000000040440000000000001048000000000000000100800400000000000",
INIT_13 => X"000800000000000000000000000100C220050000000000000000008220884400",
INIT_14 => X"000000000000000830000000000000000016101C5C1400000000000000000000",
INIT_15 => X"0000000000000000000000000020C00000088000012090101280401000000200",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000040028000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"000010082A954BA00003DFEF085155400F78428BEF0000000000000000000000",
INIT_22 => X"8015400FF84001EFA2FBE8B55A2AE80000F7D5555555D2AAAABAAAD1420BAFF8",
INIT_23 => X"87FFFF55557BD54AAF7FBC01FFA2802ABEFF7AE95555A2FBE8BEFA2843DE00AA",
INIT_24 => X"0804155EFFFFBE8BFF0800174AA557BFDE10A2FBEAB45F7D56AABAAAD5554BA0",
INIT_25 => X"5FFD568BEF087FE8A1055003FE00A2AA801FFA28402000AAAE955455500155EF",
INIT_26 => X"45AA843FE0008557DFFF0800020105D557FEAA00557DE10F7D1574AAA2D16AB5",
INIT_27 => X"0BAF7AEA8B45080417400FFFFC2145080015400AA802AA00AAAE800BA5D00155",
INIT_28 => X"000000000000000000000000000000000000000000516AA00A2AE800BAFFFFC2",
INIT_29 => X"A8ABAAADB40092E38E070280024904AA1C0438FD7005150438F78A2DBFF00000",
INIT_2A => X"FE8BC7BE8E38E10A28017400E38A051FFA2FFEDB55B6A080038E3DB50555412A",
INIT_2B => X"D16AABAA2DB50482147FFAF554971D0492E3F1C71C7BE8A2ABD7E3AA9257DA2F",
INIT_2C => X"AAA955554900105FF0800175D7E3FFEFBD70000124AA557FFDE10A2FBEDB6DF7",
INIT_2D => X"FFDF50482A2DB6AB45FFD56DBD7087BEAA38410038E38A2AE851FFB68402038A",
INIT_2E => X"0AAA085082550A1057DBE803AE38145B78FD7000005010495B7AE921C517DE10",
INIT_2F => X"00A2A0800BAE3F1C0092EBAAADB6D080A12410FFF1C017D140410400BE8E28A1",
INIT_30 => X"0AAF7AEBDFEF0000000000000000000000000000000000000000000001C556FA",
INIT_31 => X"00AAAAFBC0145002AA8AAAAAFFC2000AAAA974AA0800020BA550028B55085540",
INIT_32 => X"A8B55AAAE821EFAAFBEAB55F7AAA8A00AA8417400AAAE975EFA2FBFFF55FF840",
INIT_33 => X"BFFE10A2FFFFFEFF7D568ABAA2FFC00105D7BE8B55085142010AAD157545F7AE",
INIT_34 => X"AA955FFFF80020BAAAAA975450800001EF080417555AAFFFDF450804020AA557",
INIT_35 => X"07FEAA0055517DE00FFFBC2000AAFBE8B55F7D17DF45007FE8AAA08002AAAAA2",
INIT_36 => X"5D0000010F7AAA8A10AA8017400552A801EFF7802AABA5D7FEAB450800154100",
INIT_37 => X"00000000005D557FE00A280020BAAAD140000A2AEBFFEF082A82010FFD5421EF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000C00000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(15),        -- Port A data input
DOA(0)   => data_read_a_lo(15),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(15),        -- Port B data input
DOB(0)   => data_read_b_lo(15),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_16_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"DA22C618B1000482B688B186588884862A400438255FC38381441205BA803003",
INIT_01 => X"264AC80028404C211203A952A90341080B173340412000E1005D628000820484",
INIT_02 => X"400034C206C405000001A48202084004003008255040826EE008B440200E2042",
INIT_03 => X"A459C1240181AB20AD27315B7F1983CA1C900040422A005762010010000C0400",
INIT_04 => X"296E542B6E3A825C15FB385321B4ADFE16AB45FD2C400002E205231201290A28",
INIT_05 => X"B9E5815006028179808C00A0D2152B90707A1E0BD423CAC0000D610000000710",
INIT_06 => X"81F104A1415C292164280081C6AB88742086ACACDE240000A80090CE82A803B9",
INIT_07 => X"400800000ACCAA280940580400A37B8896CA4D000A80C1102A00001C14028009",
INIT_08 => X"0015452880C8D90409A02D965965200100104F2B00822512000000231520A024",
INIT_09 => X"A5AA80018120E00066000000000012C9000A0000D0A80000BF8028E87C1B9927",
INIT_0A => X"00520228080108039501200848002912300208092B940192D1000000000000A8",
INIT_0B => X"03561180063DB4F6110001100011000110001100011000110001080008800080",
INIT_0C => X"080200854409418B02ED0000502A02972000040BB401100010012B4C90000100",
INIT_0D => X"6D061A1F8D60D80820500101244AA8A2AA242E80000009200120000000000000",
INIT_0E => X"6D066210E5001DB4A5B400C7D553847165A99000C6564CDD051DC99000C65555",
INIT_0F => X"21D0C48F254946148107354292673D1F72C99000C6564CDD0565C99000C65555",
INIT_10 => X"952D2058F33225787810F5001D6121A9559224D1FF97D0272F04D89441A56D8A",
INIT_11 => X"6C1C74485B81E31306C71D1093AB8A64811BADC00992180D58033B1172F2A025",
INIT_12 => X"7B86DED8E3A212748F0E0CA638E890B7A8546120C0AFF5B548AC431FB1C7DB07",
INIT_13 => X"EFCE9B26DECA1AD36A2E4F40DF6AAAF260AF88899E8B8B93D12A877178DD0032",
INIT_14 => X"A8009F8B108C80A1021B9A8BB8056662CA1951596800FC01A38D4D4B072B922F",
INIT_15 => X"00000000000000000000000000044000102A0001148442A1108103595580A840",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"4C690DA64C1C4F68A36040000000000000000000000000000000000000000000",
INIT_19 => X"D14D14D14D14D14D14D14D14D14514514514514529E5F87869E79E78558D1154",
INIT_1A => X"3D1E8F47A7D3E9F4FA7D3E9F4FA7D3E9F47A7D1E9F47A7D1E9F4D14D14D14D14",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE000000000000000007D3E9F4FA7D3E8F47A3D1E8F47A",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFEFF7D168B55AAD17FFFF552EBFE00007FC00AA0000000000000000000000",
INIT_22 => X"04000BA552A821FFFF8000010082A954BA00003DFEF085155400F78428BEF087",
INIT_23 => X"2AE80000F7D5555555D2AAAABAAAD1420BA5D2E975EFF7D568BFFFF80175EF00",
INIT_24 => X"FF84001EF0000020AA5D00154005D043FF45555540000082EAABFFA2FBE8B55A",
INIT_25 => X"0087FD74BAAAAEBFFEF557FC00AAF7AE95555A2FBE8BEFA2843DE00AA8015400",
INIT_26 => X"FFAAD5554BA087FFFF55557BD54AAF7FBC01FFA2802ABEF557BEABEF5D041541",
INIT_27 => X"E10A2FBEAB45F7D56AABA082A97545F7D16ABFFFFAABFEAAFF84001FF002A821",
INIT_28 => X"0000000000000000000000000000000000000000FFFBE8BFF0800174AA557BFD",
INIT_29 => X"50438F78A2DBFF0871F8FC7E3D56AB6DBEDB7FFEF552AB8E38087FC209200000",
INIT_2A => X"16ABFFE38E175EF1400000BA412E871FFE38E070280024904AA1C0438FD70051",
INIT_2B => X"2EAFBD7A2FFEDB55B6A080038E3DB50555412AA8ABAAADB400924920925EFF7D",
INIT_2C => X"E8E38E10A28017400E38A051FF0804050BA410A1240055003FF6D5551420101C",
INIT_2D => X"4975EDBC7550E12410087FD74AAB6AABFFC7557FC00BAE3AA9257DA2FFE8BC7B",
INIT_2E => X"AF780051C70824851D7A2DB50482147FFAF554971D0492E3F1C71C7BE8A2ABD7",
INIT_2F => X"D70000124AA557FFDE10A2FBEDB6DF7D16AABA08249756DF7D168BC7F7AABAEA",
INIT_30 => X"AAA007BC0000000000000000000000000000000000000000000000000E3FFEFB",
INIT_31 => X"20BA550028B550855400AAF7AEBDFEF08516AB55A2D16ABEFFFFBFDFFF552AAA",
INIT_32 => X"C20000000021EFF7D568BFFA2AA955FF5D04020AA002A955EFAAAA974AA08000",
INIT_33 => X"03DFEF5D51420005D2ABFF45A2FBFFF55FF84000AAAAFBC0145002AA8AAAAAFF",
INIT_34 => X"AE821EFAAFBEAB55F7AAA8A00AA8417400AAAE975EF0800174BA002E820105D0",
INIT_35 => X"AD157545F7AEA8B5500557DF45552A82000007BD74AAF7AEBDF455D7BC20BAAA",
INIT_36 => X"F7D568B55FFAAAAABAFF8415545000015555A2FFC00105D7BE8B55085142010A",
INIT_37 => X"0000000000AAFFFDF450804020AA557BFFE10A2FFFFFEFF7D568ABA0804155FF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000400000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(16),        -- Port A data input
DOA(0)   => data_read_a_lo(16),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(16),        -- Port B data input
DOB(0)   => data_read_b_lo(16),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_17_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"5284CE4FB7BD2C8994A13392DBD02E14006B82AC7E800D44D3DD2FD5F9B961C0",
INIT_01 => X"F9BA301F7E03FC6793F2199B39FC233C11D93AE6F3BB92B32091DBC339B24542",
INIT_02 => X"1D5FC0C08F040404446965C0607FB8A217C400C33A908078551BD04222186338",
INIT_03 => X"8504930A37F65820CB24111B7F08014A0AB84A52B6D2AFF97C1B5AC757F06D6B",
INIT_04 => X"250834336D1E81500FDB38302292ADFE103B6DBD204037F202042075E2B1D00A",
INIT_05 => X"8F039786062C6CE092F5FE005236781C402A0807B4070670083DC68206D7E6D0",
INIT_06 => X"0CD26803C3582408962C58B183F8AEF42045919B30E085DD2ED57D4EED08CA6A",
INIT_07 => X"700000B30380670B8142500448E3E01E94EF1340A28AC1AC8156044D1400AA00",
INIT_08 => X"009F3A1B0120A1C51DFFC40C30E5F0182D0950190C0810BE00E9A76E4C6FFBE4",
INIT_09 => X"8FCCC200A59BDD2FFE3F3EC7C7DEF207000F00059D2ED56D7EED2ED3C9A867DC",
INIT_0A => X"0617112E46F05D02DD814102F800633F1D0A7CC9AE7A08BFF0001D35682AC0CE",
INIT_0B => X"8A3F06ABD73DBCF4FBCF4FBCF4FBCF4FBCF4FBCF4FBCF4FBCF4FBE7A7DE7A780",
INIT_0C => X"001000974F08518F5AFFC94B533FADA7FDE97D6BFF329E1B50FF99F086000D9E",
INIT_0D => X"F50B018F95EA3DED1652EC0B27E67F419E2E1E8000C0036340B8000000000000",
INIT_0E => X"F50B01C8DF7F96197DB4AFC8C8886AF672A1537F759299F50B03C1537F759199",
INIT_0F => X"6068331C5103E7EF0FBEED6BB6A9412007C1537F759299F50B03C1537F759199",
INIT_10 => X"21F2CD7F252CDABB3CE8CF7F963AB9FD6AD434201AA68B837FFD1F7B7125B68C",
INIT_11 => X"BD055EB6D555CB2949C15BA7270FF256526BBFD55BBE71D79F73C7AC6DB9BF37",
INIT_12 => X"94080BF82B74E4E1FE4ACA4E0ABD6DAAAB965293036FF6B652A99A6026027FBE",
INIT_13 => X"EF5CBA7A43482800FEFAFD06B8CFCCAB7550D0C2022EAEBD438697AD2EBA9168",
INIT_14 => X"AC00A8BBFC8B501CF7A0FED9A548FA19752C4A4EADAE42FCBC38C3B7BEBF42CF",
INIT_15 => X"0000000000000000000000000026E100002F382DBD9ECFE117805F20CFDAAB00",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"09EDCC4052E917114F981800C000000000000000000000000000000000000000",
INIT_19 => X"EBA69AEBA69A69AEBA69AEBA69A69A69A69A69A68698686981D75D7443720030",
INIT_1A => X"46A351A8D068341A0D068341A0D068341A0D46A341A0D46A341A69AEBA69A69A",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000000000046A351A8D46A351A8D46A351A8D",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFEFF7FBEAB450804001EFAAD57FEAA0000000000000000000000",
INIT_22 => X"51401EF087FD74AA087FFFFEFF7D168B55AAD17FFFF552EBFE00007FC00AA087",
INIT_23 => X"82A954BA00003DFEF085155400F78428BEFAAD168A000004020AA5D7BE8B4500",
INIT_24 => X"552A821FF5D00020BA552A82000552A821555D7FEAB55FF80175EFFF80000100",
INIT_25 => X"FAAFBC01EF5D0015555557BFDEBA5D2E975EFF7D568BFFFF80175EF0004000BA",
INIT_26 => X"BAA2FBE8B55A2AE80000F7D5555555D2AAAABAAAD1420BAFFFFFDF45AAD17FFF",
INIT_27 => X"F45555540000082EAABFF00516AA10552E820BA007FEABEF005555555A2D1554",
INIT_28 => X"00000000000000000000000000000000000000000000020AA5D00154005D043F",
INIT_29 => X"B8E38087FC2092147FFFFFFFFFBFDFC7EBF5E8B550000071EFB6DF7AE9200000",
INIT_2A => X"A07082497FEFB6D1451471EF007BD04920871F8FC7E3D56AB6DBEDB7FFEF552A",
INIT_2B => X"8E175FFE38E070280024904AA1C0438FD7005150438F78A2DBFFBED16AA381C0",
INIT_2C => X"38E175EF1400000BA412E871FF550A00092492A850105D2A80155417BEFB6DEB",
INIT_2D => X"FFF5FFF6DAADF7FFD7B6F1C71EF55001756D5D7BFAEBA4920925EFF7D16ABFFE",
INIT_2E => X"700515556DA2DF50492A2FFEDB55B6A080038E3DB50555412AA8ABAAADB40092",
INIT_2F => X"BA410A1240055003FF6D5551420101C2EAFBD7145B6AA28492487082007FEDBD",
INIT_30 => X"5EFFFFBEAA000000000000000000000000000000000000000000000000804050",
INIT_31 => X"ABEFFFFBFDFFF552AAAAAA007BC0000557FFDFEFF7FBFFF55A2D16AB55000017",
INIT_32 => X"BDFEFF7D568AAA5D2A97410007BFFFFF5551555EF087FC200008516AB55A2D16",
INIT_33 => X"A82155087FFFFEFAAAA975EFAAAA974AA0800020BA550028B550855400AAF7AE",
INIT_34 => X"00021EFF7D568BFFA2AA955FF5D04020AA002A955EF5D2E80010002A954005D2",
INIT_35 => X"02AA8AAAAAFFC2000FFD57DFFFAAFFFDF55FFD1575FF5504175EF5D7FEAAAA00",
INIT_36 => X"000415410007BFFF450051555EFA2FBC0000A2FBFFF55FF84000AAAAFBC01450",
INIT_37 => X"00000000000800174BA002E820105D003DFEF5D51420005D2ABFF45557FE8AAA",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000CFFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(17),        -- Port A data input
DOA(0)   => data_read_a_lo(17),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(17),        -- Port B data input
DOB(0)   => data_read_b_lo(17),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_18_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"69844019080000A21A611406840014122A641074155FC28A2024001001801003",
INIT_01 => X"01067920034004180005E9E3C90360C0041C0181002001602025800008440084",
INIT_02 => X"40AC3CAA22D605200000856E2481902400344A20F802C22054001000021E2379",
INIT_03 => X"A54C23B34C81EB2076471000800981140C010101750D1007E58040102B0E0100",
INIT_04 => X"22660C1C0065003C04040013236E105016A028402D618803EB092B9201490B2A",
INIT_05 => X"B8E080000000005889AC41E04508A99070200E010001C1CA11803850C8000100",
INIT_06 => X"800A4CE301545001F40050216C09950004C2047BCF1C8090C02800C0120886B3",
INIT_07 => X"814A0080064C1F300020080182001A9E02C03400082002700000217294007101",
INIT_08 => X"000117088080990419002D86184A01018030430700802541420440022030041A",
INIT_09 => X"7030C30B885200D274004008080003C32A10A19090C02010E102294406168800",
INIT_0A => X"00602A01880980037109700C04C44C92A88DCC2211E44174112840880000060D",
INIT_0B => X"11C0D95C20C2030A003080030800308003080030800308003080018400184004",
INIT_0C => X"8304E02809832E6021002020404042000F00008400811824AD4007ECD9436261",
INIT_0D => X"0AFCE5D22A82B20000520100C801F8A07E103000A1285C84000418360C1B060D",
INIT_0E => X"0AFCFD8CB17E5B4F045557575E6EFBE3942C1040A41D660AFCE1CC1040A41E66",
INIT_0F => X"8E7FFBB385661C08D1455ABA91E6FF5FDFCC1040A41D660AFCF9CC1040A41E66",
INIT_10 => X"015F82C006C3AF31E64CB17E5A9655017F1FC73FAF1D61B1040294C58AD1FF5F",
INIT_11 => X"B95454005BAA36DCF8E519001BF80DEB3EE2020EA678189C6EC32881F7F75648",
INIT_12 => X"67D7EDFCA320037E81BD77D728A800B7546DBDFF12904747A351145FC53ABF8D",
INIT_13 => X"92B764225C57C97EBE76E1254F0C0D4514A84F5573FE9DBA4A38E247C522CC0E",
INIT_14 => X"BE84370001B6922070440556B15F7FABBC40151D7C747D8220673C3B9DB84B20",
INIT_15 => X"06C1B06C1B06C1B06C1B06C1B0491069068000004060300A005A01183F240014",
INIT_16 => X"6C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B",
INIT_17 => X"C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B0",
INIT_18 => X"B80EE173C2300F7DF16000000000000000000000000041B06C1B06C1B06C1B06",
INIT_19 => X"AAAAAA28A28A28AAAAAAA28A28A28A28A28A28A2910591505C104104B28BBECE",
INIT_1A => X"128944A25128944A25128944A25128944A2552A954AA5128944AAAA28A28A28A",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000128944A25128944A25128944A25",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFDFEF5D2A974BA082E954000000000000000000000000",
INIT_22 => X"0028B55002E82000087FFFFFFFFFFFFFEFF7FBEAB450804001EFAAD57FEAA087",
INIT_23 => X"7D168B55AAD17FFFF552EBFE00007FC00AA087FFFFFFFFFBFDF45AAD568B5508",
INIT_24 => X"087FD74AAAAFFFDF45A2D16AB55F7FFFFFFF00043DE10AA843DE00087FFFFEFF",
INIT_25 => X"A55042ABEF5D7FD75FFAAD540145AAD168A000004020AA5D7BE8B450051401EF",
INIT_26 => X"45FF8000010082A954BA00003DFEF085155400F78428BEFAA80000000804154B",
INIT_27 => X"1555D7FEAB55FF80175EF5D00020105D2A97400082E95555085168A10557FD75",
INIT_28 => X"00000000000000000000000000000000000000005D00020BA552A82000552A82",
INIT_29 => X"071EFB6DF7AE921C7FFFFFFFFFFFFFFFF7FBFDFFF5D2A954AA082A9242800000",
INIT_2A => X"1FAF55A2DF6DB7D1C002AB7D002A82028147FFFFFFFFFBFDFC7EBF5E8B550000",
INIT_2B => X"8E38E280871F8FC7E3D56AB6DBEDB7FFEF552AB8E38087FC2092087FFDFC7E3F",
INIT_2C => X"97FEFB6D1451471EF007BD0492B6F1F8F55AADF6DB7DE3F5FAFC708003DE28B6",
INIT_2D => X"A28407038140410492550A2ABC7497BD25FFAADF4516DBED16AA381C0A070824",
INIT_2E => X"D1C516FA28417BD5545E38E070280024904AA1C0438FD7005150438F78A2DBFF",
INIT_2F => X"92492A850105D2A80155417BEFB6DEB8E175FF5D0E05000492097428002E9557",
INIT_30 => X"4AA082A820AA000000000000000000000000000000000000000000000550A000",
INIT_31 => X"FF55A2D16AB550000175EFFFFBEAA00557FFFFFFFFFFFDFEFF7FBFFFEF552E97",
INIT_32 => X"C0000087BFDF45AAD568B55AAFBFDFEF55042ABEF002A800AA557FFDFEFF7FBF",
INIT_33 => X"16AB4500043DEAAFFAEAAAAA08516AB55A2D16ABEFFFFBFDFFF552AAAAAA007B",
INIT_34 => X"D568AAA5D2A97410007BFFFFF5551555EF087FC2000FFD56AB45A2FFFDFFFAAD",
INIT_35 => X"855400AAF7AEBDFEFA280154BA550400000552AA8B45087FC01EFA2FFD55EFF7",
INIT_36 => X"0804154BA082A975EF5D517DEAA007BD5545AAAA974AA0800020BA550028B550",
INIT_37 => X"00000000005D2E80010002A954005D2A82155087FFFFEFAAAA975EF5D2E97400",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000400000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(18),        -- Port A data input
DOA(0)   => data_read_a_lo(18),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(18),        -- Port B data input
DOB(0)   => data_read_b_lo(18),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_19_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"042200000000000041088001001AA00000000000000000000000500802000003",
INIT_01 => X"074018000024000000000404000000000A22000800000800004A200000000001",
INIT_02 => X"0000048002C405000000000006A84000000000200893C246A20000000020031A",
INIT_03 => X"082A58E411004B2000071000000981000C000000002045000200000000000000",
INIT_04 => X"200604000000001C0400001320000000162000002C4000026201201200090800",
INIT_05 => X"1020800000000058840200204000099070200E010001C0400000000000000000",
INIT_06 => X"0012048037805421402850001402498820022802400480405008901100A00102",
INIT_07 => X"00000000020C0130481204919200010C82000000000006002A548902A0020109",
INIT_08 => X"0001150800009900000005861840000000004301000B000000000001C1C00000",
INIT_09 => X"001F00002024B20002000000000002C300000000405000103010204000000000",
INIT_0A => X"00000000000000000000000000000040002000044000000000000000000002F0",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000420003B00000000000000000040012C80000000",
INIT_0D => X"45001A03C0825A0D20800000000018A006001000000000000000000000000000",
INIT_0E => X"450002131E01A1F6EA0A0020211146E069C2ACC01AE80045001D82ACC01AE800",
INIT_0F => X"1188340C3E1CFAD27CC2E004481020892282ACC01AE80045000582ACC01AE800",
INIT_10 => X"DEA03228D810007019931E01A1E5BA02802008C06F029D4C7B76639CEC0A0020",
INIT_11 => X"428AA3592000000206C2A4DAC00000008113C246A181C03FE4662A84575768DF",
INIT_12 => X"08201090549B5800000000261546B24000000000C53807E7CC06618018C51210",
INIT_13 => X"13F6A185A0A0168128411ACB800C0E108A0720288C011046B5986247C5452291",
INIT_14 => X"0000C220010808C10D9A92A74CD7CF4A080031B1515B212143D841431046B58A",
INIT_15 => X"00000000000000000000000000000000000000000000000000000118030004E0",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"3F0C7010C660C744192000000000000000000000000000000000000000000000",
INIT_19 => X"1861861861869A61861861861861861861861861A8208C4C1534D34C07208BBA",
INIT_1A => X"0984C26130984C26130984C26130984D26930984C26130984C261861861869A6",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE000000000000000000984C26130984C26130984C2613",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF552A974AA0004174BA0000000000000000000000",
INIT_22 => X"2E974BAA2FFFFE10087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974BA082E95400F7F",
INIT_23 => X"FFFFFFEFF7FBEAB450804001EFAAD57FEAAF7FFFFFFFFFFFFFFFFF7FBFDFFF55",
INIT_24 => X"002E82000F7FFFFFFFFFFFFDFEFA2D568B550004001EFAAAEA8ABA087FFFFFFF",
INIT_25 => X"5AAD16ABEF5D2ABFF55080402010087FFFFFFFFFBFDF45AAD568B55080028B55",
INIT_26 => X"BA087FFFFEFF7D168B55AAD17FFFF552EBFE00007FC00AAF7FFFFFFFF7FBE8B5",
INIT_27 => X"FFF00043DE10AA843DE00557FFDFEFA2D16AB55A2FFFDFEF5D2EBFE00AAFFFFE",
INIT_28 => X"0000000000000000000000000000000000000000AAFFFDF45A2D16AB55F7FFFF",
INIT_29 => X"954AA082A92428E3FFFFFFFFFFFFFFFFFFFFFFFEF552A974AA0000104AA00000",
INIT_2A => X"FFDFEFF7F5FAFC7492A974AAB6F5F8E101C7FFFFFFFFFFFFFFFF7FBFDFFF5D2A",
INIT_2B => X"A4A8AAA147FFFFFFFFFBFDFC7EBF5E8B550000071EFB6DF7AE92EBFFFFFFFFFF",
INIT_2C => X"2DF6DB7D1C002AB7D002A82028FFFFFFFEFF7F1F8FD7AAD16AB450000001FFBE",
INIT_2D => X"F7FBF8FC7E3F5EAB45B6DF6FBEF5D2AB8F7D000000010087FFDFC7E3F1FAF55A",
INIT_2E => X"7412ABFE28B6F5F8E820871F8FC7E3D56AB6DBEDB7FFEF552AB8E38087FC2092",
INIT_2F => X"55AADF6DB7DE3F5FAFC708003DE28B68E38E284971F8FC7AAD56DB6DBEF5F8FD",
INIT_30 => X"4AA0004000AA000000000000000000000000000000000000000000000B6F1F8F",
INIT_31 => X"DFEFF7FBFFFEF552E974AA082A820AAA2FFFFFFFFFFFFFFFFFFFFFDFEF552E95",
INIT_32 => X"EAA00A2FFFFFFFF7FBFDFFFFFD568B55002A954AAF7D568A00557FFFFFFFFFFF",
INIT_33 => X"56AB450004001EFFF842AAAA557FFDFEFF7FBFFF55A2D16AB550000175EFFFFB",
INIT_34 => X"7BFDF45AAD568B55AAFBFDFEF55042ABEF002A800AAF7FBFDFEFF7D56AB45AAD",
INIT_35 => X"52AAAAAA007BC0000FFFBE8B55AAD168B55F7FFFFFFF552AA8BEF08040200008",
INIT_36 => X"A2D57FFFFF7D568B45002ABDEAAFFD16AA0008516AB55A2D16ABEFFFFBFDFFF5",
INIT_37 => X"0000000000FFD56AB45A2FFFDFFFAAD16AB4500043DEAAFFAEAAAAA08556AB55",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000800000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(19),        -- Port A data input
DOA(0)   => data_read_a_lo(19),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(19),        -- Port B data input
DOB(0)   => data_read_b_lo(19),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_20_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000003",
INIT_01 => X"A65FF80000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000048002CC070000000000000000000000002FF86100200000000220002362",
INIT_03 => X"0000000000080F6000977060009B87A03C000000000000000000000000000000",
INIT_04 => X"3F2EFC040388137C3E20C477600142019E6000003CC0000A6601601A000B0000",
INIT_05 => X"102F91D10802ABFB80000021C8010FB0F0F43E1FE867DFC04400390210000220",
INIT_06 => X"90492261000080003400000010008000004203FE400580000000803000200006",
INIT_07 => X"401000004FFDFF28C4300C0010200100004000002AA001F00000000014000000",
INIT_08 => X"0801F5780259FB00000007BEFBC010002008FF7F00000000010018A81000041C",
INIT_09 => X"00000000020000000000000000000ADF00000020000000800000802830011023",
INIT_0A => X"0000000000000200020000000000000000000000000000000200200290000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"08120000B9090A700000200000004000000400000080002000407FED80000000",
INIT_0D => X"000079804000F00000000000C01FF8A7FE003000000004008100000000000000",
INIT_0E => X"0000798201000000100000000135386000401000010000000079801000010000",
INIT_0F => X"0185C300020004000010000000000252C7801000010000000079801000010000",
INIT_10 => X"00000010C1F30F300002010000080000000000CD8A0000400400000010000000",
INIT_11 => X"008040000000000292C0080000000000A5604000000284000818505200080000",
INIT_12 => X"0015E1B00100000000001496008000000000052B000048080000000000FC3600",
INIT_13 => X"80000000000002BA280000800830300000000000B8B400000401881010000000",
INIT_14 => X"00000000020020020001000040283024E6FB8604020080000383383B00000400",
INIT_15 => X"000000000000000000000004010201001003020200000000000127DBFF004000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"038200010089120104D204002000000000000000000000000000000000000000",
INIT_19 => X"B2CB2CB2CB2CB2CB2CB2CB2CB2C30C30C30C30C306982121A1E79E79A0700030",
INIT_1A => X"432190C86432190C86432190C86432190C86432190C86432190CB2CB2CB2CB2C",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000432190C86432190C86432190C86",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA0804020100000000000000000000000",
INIT_22 => X"2E954AA000400000F7FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0004174BAFFF",
INIT_23 => X"FFFFFFFFFFFFFDFEF5D2A974BA082E95400007FFFFFFFFFFFFFFFFFFFFFFEF55",
INIT_24 => X"A2FFFFE10FFFFFFFFFFFFFFFFFFFFFBFDFFF5D2E954BA007FC00BA087FFFFFFF",
INIT_25 => X"FF7FBFFF550800020BAAAD56AAAAF7FFFFFFFFFFFFFFFFF7FBFDFFF552E974BA",
INIT_26 => X"10087FFFFFFFFFFFFFEFF7FBEAB450804001EFAAD57FEAA007FFFFFFFFFFFFFE",
INIT_27 => X"B550004001EFAAAEA8ABA5D7FFFFFFFFFFFDFEFF7D56AB450000021EFA2D57DE",
INIT_28 => X"0000000000000000000000000000000000000000F7FFFFFFFFFFFFDFEFA2D568",
INIT_29 => X"974AA0000104AAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA08000500000000",
INIT_2A => X"FFFFFFFFFBFDFEF5D2E974AA000A07000E3FFFFFFFFFFFFFFFFFFFFFFFEF552A",
INIT_2B => X"71C50BA1C7FFFFFFFFFFFFFFFF7FBFDFFF5D2A954AA082A92428087FFFFFFFFF",
INIT_2C => X"7F5FAFC7492A974AAB6F5F8E10E3FFFFFFFFFFFFFFEFF7FBFFFFF552E974AA00",
INIT_2D => X"1C7FFFFFFFFFBFDFEFE3F5F8F450004050AABEDF6FABAEBFFFFFFFFFFFFDFEFF",
INIT_2E => X"50804021FFB6D57DE28147FFFFFFFFFBFDFC7EBF5E8B550000071EFB6DF7AE92",
INIT_2F => X"EFF7F1F8FD7AAD16AB450000001FFBEA4A8AAA497FFFFFFF7FBF8FC7EBD168B4",
INIT_30 => X"4AA080017410000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFDFEF552E954AA0004000AAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A95",
INIT_32 => X"820AA087FFFFFFFFFFFFFEFF7FBFDFFF5D2A974AA002E95410A2FFFFFFFFFFFF",
INIT_33 => X"FFDFEF5D2E954AA0051554BA557FFFFFFFFFFFDFEFF7FBFFFEF552E974AA082A",
INIT_34 => X"FFFFFFFF7FBFDFFFFFD568B55002A954AAF7D568A00AAFFFFFFFFFFBFDFEFFFF",
INIT_35 => X"000175EFFFFBEAA005D7FFFFEFF7FBFDFFFAAD16AB450804174AAFFFFFFEBAA2",
INIT_36 => X"F7FFEAB45A2D568B550804001EFF7D57DEBA557FFDFEFF7FBFFF55A2D16AB550",
INIT_37 => X"0000000000F7FBFDFEFF7D56AB45AAD56AB450004001EFFF842AAAA087BFDFEF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000000FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(20),        -- Port A data input
DOA(0)   => data_read_a_lo(20),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(20),        -- Port B data input
DOB(0)   => data_read_b_lo(20),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_21_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"4A302428B824900A128C090A5C1800261500213C005FE812D10420054085A202",
INIT_01 => X"081FFE3440B609703B0427F801A40B8115BC4F655300340288A40D30040E4DD8",
INIT_02 => X"04CA478082CC1740002019824E0203100640303FF8C0B31061096E21A1840814",
INIT_03 => X"8C329E9204020FE002577800405B87047D5042129D8D0248903200013290C800",
INIT_04 => X"3E7FFE02482553FC3C020277E128080A1E6000003CC0000A6601E03A8B0F0008",
INIT_05 => X"F43F8140000203FFC806C8A1C1048FF0F0E07E1F00F7FFC00024010000468310",
INIT_06 => X"08710C10015E083D01A24404786BE0014114C3FE4187A009A663A680100B3096",
INIT_07 => X"200800008FDFFF00290000100211019812E210488228000000900260026C6058",
INIT_08 => X"0EF1F5FA0041FF080AC707FEFBC110008420F7FF388B70A20389346FE8000580",
INIT_09 => X"917FC30010107688862A28C54518DBFF00020004C0A6044901112A0908AA0A30",
INIT_0A => X"006309044081A001B188300E20806520398C6021569249C4B3007127080806FF",
INIT_0B => X"904595123203040D9228D9228D9228D9228D9228D9228D9228D99146C9146C84",
INIT_0C => X"88042090068008003120000806001402504110C48002403601887FEF80022A51",
INIT_0D => X"26C0AC404E43032CA0C205880A7FFAB7FE01409400400C0594A4002200110008",
INIT_0E => X"26C0AC086A170250454004C6012280129B034A080C0B0016A0D20346080C0A80",
INIT_0F => X"0B064092D85938C0112144050224120C500346080C0B0016A0D2034A080C0A80",
INIT_10 => X"40702E058355458967E86A170220D1800093414B0414782E4B5000D81480809A",
INIT_11 => X"081B1545104135443306C35901024F88A88049062A747512B76783C5D040E080",
INIT_12 => X"40160040D86B202049B22198362A8A208279854400A036801480031401900800",
INIT_13 => X"0DD001C002D38334000914028354008301008C0CF1480245108C7640A0604032",
INIT_14 => X"AC0496022300233104662848808E191526205018030060540284FA0C0044022C",
INIT_15 => X"004010040100401004010040102090010008000001C0E010020007DFFFC06E60",
INIT_16 => X"0401004010040100401004010040100401004010040100401004010040100401",
INIT_17 => X"4010040100401004010040100401004010040100401004010040100401004010",
INIT_18 => X"FF7FFDF7FF3E3DFDF7E000000000000000000000000040100401004010040100",
INIT_19 => X"FBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBFFDFDFFFCF3CF3FFFEF9FEE",
INIT_1A => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFEFF7FBFDFEFF7FBFDFEFBEFBEFBEFBE",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0004000100000000000000000000000",
INIT_22 => X"2A954BA0004154BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080402010FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF552A974AA0004174BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"000400000007FFFFFFFFFFFFFFFFFFFFFFEF552E974BA0804000AAF7FFFFFFFF",
INIT_25 => X"FFFFFFDFEF5D2E974BA002E97400007FFFFFFFFFFFFFFFFFFFFFFEF552E954AA",
INIT_26 => X"BA087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974BA082E95400007FFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2E954BA007FC00BA5D7FFFFFFFFFFFFFFFFFFBFDFEF5D2A954AA002E974",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFBFD",
INIT_29 => X"954AA080005000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA00000200000000",
INIT_2A => X"FFFFFFFFFFFFFFF552A974BA0000174AAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0A000AAE3FFFFFFFFFFFFFFFFFFFFFFFEF552A974AA0000104AAF7FFFFFFFFFF",
INIT_2C => X"FFBFDFEF5D2E974AA000A07000007FFFFFFFFFFFFFFFFFFFFDFEF552E954BA08",
INIT_2D => X"1C7FFFFFFFFFFFFFFFFFFBFDFEF5D2A974BA002A95400087FFFFFFFFFFFFFFFF",
INIT_2E => X"F552E974BA0020924BA1C7FFFFFFFFFFFFFFFF7FBFDFFF5D2A954AA082A92428",
INIT_2F => X"FFFFFFFFFEFF7FBFFFFF552E974AA0071C50BA557FFFFFFFFFFFFFFFF7FBFDFF",
INIT_30 => X"4BA000002000000000000000000000000000000000000000000000000E3FFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2A954AA080017410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"000AAF7FFFFFFFFFFFFFFFFFFFFFFFEF552A974BA0000174BAFFFFFFFFFFFFFF",
INIT_33 => X"BFDFEF5D2A954BA082E800AAA2FFFFFFFFFFFFFFFFFFFFFDFEF552E954AA0004",
INIT_34 => X"7FFFFFFFFFFFFFEFF7FBFDFFF5D2A974AA002E95410087FFFFFFFFFFFFFFFF7F",
INIT_35 => X"52E974AA082A820AA557FFFFFFFFFFFFFEFF7FBFFFFF552E954BA002E9741008",
INIT_36 => X"FFFBFDFEFF7FFFFFEF5D2A974BA0000020AA557FFFFFFFFFFFDFEFF7FBFFFEF5",
INIT_37 => X"0000000000AAFFFFFFFFFFBFDFEFFFFFFDFEF5D2E954AA0051554BA5D7FFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(21),        -- Port A data input
DOA(0)   => data_read_a_lo(21),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(21),        -- Port B data input
DOB(0)   => data_read_b_lo(21),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_22_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"5290F4CDE914905A14A43D33F488243E17122300F55FEB189B343A1140548380",
INIT_01 => X"A94007B259F6A975386262000C344BA9573C6FF57B18A5FB0ABFCD3C2C5F4F0C",
INIT_02 => X"D56B4302AC01005111011BD506AA5205274056900596A539584E2E6DFE4B2418",
INIT_03 => X"6B03F2F6151A2081F24001E8400008F401CB10C6594423C8923AD6B55AD0EB5A",
INIT_04 => X"8001023D37E50880436200808BC8492A0089249600101100008087248B64426E",
INIT_05 => X"A51035B41C0A88046CAEE8C23C08E040011C0020F8882001102D620A06D68301",
INIT_06 => X"B93FF975CF7889D085E997A2144E8FC2060B880081A26DCD4047EFF9EF018980",
INIT_07 => X"283800AA500200E8024AD03546A3262FB5AA5542A882040C7A64CBD64065F028",
INIT_08 => X"141008801018040E48D500400015805060040080A2A0F4A82381B4000A0905A0",
INIT_09 => X"4D0000002126F30C902A29C54539C020E11810098D4067EFF9FF284D483E2AB4",
INIT_0A => X"1400006100003202D040050220103D2A512C6A8C4F0008AA800470370000A000",
INIT_0B => X"013456520CA09281C2A81C2A81C2A81C2A81C2A81C2A81C2A81C9540E1540E00",
INIT_0C => X"A1402A13C0A10A893165281A1C2A7283516344C594A85536B1AD800214202C50",
INIT_0D => X"3C70FC20515808A0100820112300011000287B071105034406950A0285014280",
INIT_0E => X"3C70FC48E11CFC48400184CE0D6783139B0959A41606003C70FA0958AC160480",
INIT_0F => X"0D87E8B3B811B52048B10E0402AE1606D80958AC1606003C70FA0959A4160480",
INIT_10 => X"80F84E0185594581E088E11CFC38414020DD42CF909D7E0A551C02180300C0DD",
INIT_11 => X"441154C258012D86F3044A3133004A99BD8455300654458A1D588C4061403000",
INIT_12 => X"A096A240894626600953379822A984B0025B0DEC0345C9200680027181B44887",
INIT_13 => X"E2404160035482BE521C2C04A90783C18000D610B9D8070B12B1A2A62040202A",
INIT_14 => X"304244A91102C93A2D608D2A258DF8034284200C050070E40C80620C870B02C4",
INIT_15 => X"4411044110441104411044110466C440446CA06951D4EA801000980400646002",
INIT_16 => X"0100441104411044110441104411044110441104411044110441104411044110",
INIT_17 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_18 => X"FE8FF1F7DEBDDF7DF7D05122890000000003FFFFFFFF90040100401004010040",
INIT_19 => X"79E79E79E79E79E79E79E79E79E79E79E79E79E7BFFDFD7DDDF7DF7DF7DFBFDE",
INIT_1A => X"3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE79E79E79E79E",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE000000000000000003F9FCFE7F3F9FCFE7F3F9FCFE7F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0800000000000000000000000000000",
INIT_22 => X"2E974AA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000400010FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E954AA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"0004154BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA000015400FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF552A974AA0800154AAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA",
INIT_26 => X"BAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0004174BAFFFFFFFFFFFFFFFFF",
INIT_27 => X"FEF552E974BA0804000AAA2FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0000174",
INIT_28 => X"0000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040001000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E954AA000402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0417410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080005000FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF552A974BA0000174AAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA00",
INIT_2D => X"E3FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0804154BAF7FFFFFFFFFFFFFFFFF",
INIT_2E => X"F552E954BA000E124BAE3FFFFFFFFFFFFFFFFFFFFFFFEF552A974AA0000104AA",
INIT_2F => X"FFFFFFFFFFFFFFFFDFEF552E954BA080A000AAA2FFFFFFFFFFFFFFFFFFFFFFFE",
INIT_30 => X"4BA080400010000000000000000000000000000000000000000000000007FFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"17410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000400010FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF552A954BA000415400FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954AA0800",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFEF552A974BA0000174BAF7FFFFFFFFFFFFFFFFFFF",
INIT_35 => X"52E954AA0004000AAA2FFFFFFFFFFFFFFFFFFFFFDFEF552E974AA0804174AAF7",
INIT_36 => X"FFFFFFFFFFFFBFDFEF5D2E954BA002A820BAA2FFFFFFFFFFFFFFFFFFFFFDFEF5",
INIT_37 => X"0000000000087FFFFFFFFFFFFFFFF7FBFDFEF5D2A954BA082E800AAAAFFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000000FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(22),        -- Port A data input
DOA(0)   => data_read_a_lo(22),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(22),        -- Port B data input
DOB(0)   => data_read_b_lo(22),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_23_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"EF20906D902424807BC8241BC81801B97D38AD3C0800103362A6741C80A12A02",
INIT_01 => X"001FFF8409F089003B4422000D80C80106804A7951C5B9D1C828043EA28838F9",
INIT_02 => X"028406A002DC176444683862400003111001303FFC00F240D50146013B300500",
INIT_03 => X"001B243004080FE000177003145F87017D584B10D804034800200200A1008008",
INIT_04 => X"BEFFFC0248005FFC3C18A2FFE12222425E600000BDC0800AEE01E81A100F0A00",
INIT_05 => X"D03F8000000003FF810640A1C0008FF2F0E17E1F02FFFFC80100004044800080",
INIT_06 => X"800264B4854650040123428C204BF40F439647FF4807E189A477EF81DF0AF116",
INIT_07 => X"01000000FFDFFFE800401005C0A0008F86C60840AAAA100C68D1810C9F4A0020",
INIT_08 => X"1BE1F5F80003FF0002021FFEFBC80000000077FF184B03010004002FE1F29002",
INIT_09 => X"907FC308181204800600000000001BFFA800808189A657EF81DD0C00079CC800",
INIT_0A => X"0063090442A18001B188300C48907120AC810033149249C433200180082A06FF",
INIT_0B => X"9A41C1443243050C1010C1010C1010C1010C1010C1010C1010C1008608086084",
INIT_0C => X"000082A00600200080000500C000400800601200000254A000007FEFC1030221",
INIT_0D => X"0A9080400E0BF30C20CA858E087FFABFFE01409780214EE49620001000080004",
INIT_0E => X"0A908044294700701641005218521210150E5789F90A000A90800E5F81F90880",
INIT_0F => X"0E0220036864A7DCA190440301E2105C000E5F81F90A000A90800E5789F90880",
INIT_10 => X"C1400500C6CE5400032429470068924010164302048156305D66F8701681000E",
INIT_11 => X"2E0CCB0500013440600339C800004D8018000857A82920CE8CB220C81400A180",
INIT_12 => X"220344406739000009B0030019960A00026880C0422C52B01700044901488822",
INIT_13 => X"85C811A010428104128996465ADA020180804A040108A2658217C4008060300C",
INIT_14 => X"BE0692020328CA0028042054A92771C50FC070109000C1C819078280A265920E",
INIT_15 => X"020080200802008020080200800800200200000000000008004807DFFF000470",
INIT_16 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_17 => X"0080200802008020080200802008020080200802008020080200802008020080",
INIT_18 => X"0000000000000000000000000000000000000000000000802008020080200802",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000",
INIT_22 => X"2E974BA080002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E974BA000400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000400000FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF5D2E954AA080000010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA",
INIT_26 => X"10FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080402010FFFFFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2A954BA000015400FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA0804000",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E974BA080002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF5D2E954AA000402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA00",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080002010FFFFFFFFFFFFFFFFFFF",
INIT_2E => X"F5D2A954BA080407000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080005000",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF5D2A954BA000417410FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA080402000000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"02000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000010FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF5D2E974AA000402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0000",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000400010FFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"D2A954AA080017410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954AA080002000FF",
INIT_36 => X"FFFFFFFFFFFFFFFFFF552A954BA080015410FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_37 => X"0000000000F7FFFFFFFFFFFFFFFFFFFFFFFFF552A954BA000415400F7FFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000000FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(23),        -- Port A data input
DOA(0)   => data_read_a_lo(23),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(23),        -- Port B data input
DOB(0)   => data_read_b_lo(23),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_24_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100600007FFF000080108004000800020000840041000080808",
INIT_02 => X"0000068002CC07400000090C080002000000103FF811F150231000520ABE4404",
INIT_03 => X"8428180000080FE000177000001B87003D4000000E8B84010020000000008000",
INIT_04 => X"3E2FFC024800137C3C000077E00000001E6000003CC0000A6601E01A000F0200",
INIT_05 => X"103F8000000003FF80000021C0000FF0F0E03E1F0067FFC00000000000000000",
INIT_06 => X"00132412079001AD00810005E8000001401643FE4007E5501AA00000DC8C3006",
INIT_07 => X"000000000FDFFF62695A5685C094831D966000008002100C2040A178B600C240",
INIT_08 => X"08E1F5F80001FF00000007FEFBC00000000077FF000B00000000002FE0000000",
INIT_09 => X"107FC300000000000600000000001BFFA0000005501AA00000CE200000940000",
INIT_0A => X"00630104408180012188300C00814080008000010012414433000100080806FD",
INIT_0B => X"904181003003000C1000C1000C1000C1000C1000C1000C1000C1000608006084",
INIT_0C => X"00000080060000000000000012002C00000000000000000000007FEF80020201",
INIT_0D => X"440082404E0B332CA2C20188087FFAB7FE000082000000008220000000000000",
INIT_0E => X"4400824903210308074084210002460402009280010D80440084009280010F00",
INIT_0F => X"800A2400401A0C82183248060010280C20009280010D80440084009280010F00",
INIT_10 => X"C0A078160000404A0469032102981380202080026420020D06C002A08481C020",
INIT_11 => X"00164F400860000824059AD01802000208104817B00011306B2D9B0DD5082080",
INIT_12 => X"41021800B35A0300400041202C9E8010C0001040C5836CC01780018601030088",
INIT_13 => X"DB1011E000A140058220004AEFFC8101810021084301880030A8B77400603011",
INIT_14 => X"8C063C0220002201490418082010A57263E010000201033016085A40880030A1",
INIT_15 => X"000000000000000000000000000000000000000000000000000007DFFF0006E0",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"F6E7CC1132CDB444199000000000000000000000000000000000000000000000",
INIT_19 => X"79E79E79E79EFBEFBEFBEFBEFBEF9EF9EF9EF9EFA69861219575D75FF2D0AEEA",
INIT_1A => X"0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1EFBEFBEFBE79E",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE000000000000000000783C1E0F0783C1E0F0783C1E0F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020100000000000000000000000",
INIT_22 => X"2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"080002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_26 => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000400010FFFFFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2E974AA000400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0004000",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040201000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF5D2E974BA080002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFF",
INIT_2E => X"F5D2E974AA000400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF5D2E974AA000400000FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA080402010000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"00010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000010FFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002010FF",
INIT_36 => X"FFFFFFFFFFFFFFFFFF5D2E974AA000002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_37 => X"0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000402010FFFFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(24),        -- Port A data input
DOA(0)   => data_read_a_lo(24),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(24),        -- Port B data input
DOB(0)   => data_read_b_lo(24),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_25_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100200002000000080100004000000020000800041000080808",
INIT_02 => X"0000068002CC474000000800000002000000103FFCE302008000000880844A04",
INIT_03 => X"00000101C0200FF004177800081B87003D400000080000000020000000008000",
INIT_04 => X"3E2FFE024820137C3C004077F01000001E7249213CC1264A660DF05A000F9000",
INIT_05 => X"103F81C1002203FF80000021C1140FF8F0E03E1F0067FFE04800258280010052",
INIT_06 => X"80480AE20000000100000001C8608001401643FE4007C00000000000CC083006",
INIT_07 => X"280800000FDFFFEA4050140540B00100840000080002A00C2040810000000010",
INIT_08 => X"C8E1F5FA21C9FF80040007FEFBE031018C31F7FFBAEBC0020008086FE0000100",
INIT_09 => X"107FC301800000000600000000001BFFE00301000000000000CC020000140000",
INIT_0A => X"0077330C4889CC292588300C0080400000800001001243443B000100880806FD",
INIT_0B => X"904189003003000C1000C1000C1000C1000C1000C1000C1000C1000608006084",
INIT_0C => X"8B04228026824100000000000000000000000000000004A000007FEF80020201",
INIT_0D => X"400000400E03C30C20C2818C087FFAB7FE01409700C10007962418220C110608",
INIT_0E => X"4000000001010000004000000000400400001200000800400000001200000800",
INIT_0F => X"0008000000000480000040000000200000001200000800400000001200000800",
INIT_10 => X"0000001001000002000001010000100000000000202000000440000000800000",
INIT_11 => X"0000410000000008000008400000000200000806300400000820000020004880",
INIT_12 => X"0000080001080000000040000082000000001000000040800800000000020008",
INIT_13 => X"8100000000000000802000000840000200040000020008000000840000804000",
INIT_14 => X"8C04100200000200000610000000210000000018140000000008000008000000",
INIT_15 => X"04411044110441104411044510629041040D180400000010028047DFFF800C60",
INIT_16 => X"4411044110441104411044110441104411044110441104411044110441104411",
INIT_17 => X"4110441104411044110441104411044110441104411044110441104411044110",
INIT_18 => X"196A8C5A2932EC15DA080800002FFFFFFFFFFFFFFFFFC1104411044110441104",
INIT_19 => X"92492492492410410410410410410492410492412000531215A69A6BFBA2894A",
INIT_1A => X"B158AC562B158AC562B158AC562B1588C46231188C46231188C4924924924924",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000B158AC562B158AC562B158AC562",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000",
INIT_22 => X"2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF5D2E974BA080400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_26 => X"10FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0800000",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400000FFFFFFFFFFFFFFFFFFF",
INIT_2E => X"F5D2E974BA080000010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA080402000000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"02000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400000FF",
INIT_36 => X"FFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_37 => X"0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000000FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(25),        -- Port A data input
DOA(0)   => data_read_a_lo(25),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(25),        -- Port B data input
DOB(0)   => data_read_b_lo(25),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_26_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"E9264EAB20190CA3BA4997AA9002AE9C001006B0778015CFA17E0811039879C7",
INIT_01 => X"F1FFF9BB1F773C7F9BB07DFFFDD863FC5FFF3FEFFBBF9FFB22FFFBC7B9F30686",
INIT_02 => X"9B3184F8AFDEAF300029E4E300FC78A6258548EFFA71C00172082400003A2161",
INIT_03 => X"0213C3FDFFFC7F74FFBF737A603B87FEBE1A5294F65628A0001B9CE6CC606E73",
INIT_04 => X"7E2EFEBF6FFEB37C3FF3017776FFCDA43E7B6DFD7DEBFD8E6F5F78DF0BFBD644",
INIT_05 => X"902F87C74E8CCFFBB6FF70E1FE61FFBDF0FEBE1FFD67DFFEFFBDA7F7FED50870",
INIT_06 => X"213246200BCC8920360C1831CD7DF60A244B9BFEE00589DDBCEFEDC1DFA08957",
INIT_07 => X"B1D4223B4FFDFF21CC721C85DCE1458E8782484020A2C1FCA3468D77E0000300",
INIT_08 => X"2C05FD7BC471FBD13D980FBEFBEBF30B8D79FF7F451F33CFD60FE8FFFDF54003",
INIT_09 => X"19FFC71FEFED7B251E35768E8ED6BFDF3EB3EBF9DDBCE7FDC1DF8A760F3EACC0",
INIT_0A => X"56F7730ECCDBDF152199F51EDDCDEBCFF589807B7096CD4CF73AC1FC98884FFF",
INIT_0B => X"B867D3683A03A40F78C0D78C0D78C0D78C0D78C0D78C0D78C0D7A606BC606B8C",
INIT_0C => X"DFBFF5EB36DFE51FC3A80D73D840303983EE7F0EA03BDA680137FFFDFFD7E681",
INIT_0D => X"3F0080425E6BFF8DB0DAE19C09FFFFE7FE3EBEA8EB7AFEE5C9AEBD7F5EBFAF5F",
INIT_0E => X"3F00800DEC010280004000F808020290100FA2F60008003F00800FA2F6000800",
INIT_0F => X"00023002007BC0A14E00400003B8000D000FA2F60008003F00800FA2F6000800",
INIT_10 => X"01E0320007204008040DEC010300100000F600020581003F604D0700008000EE",
INIT_11 => X"201F21A2C40039006807C46426040E101A0259DFE82011A311AA042016040080",
INIT_12 => X"80020048F88C84C101C203403E434588007200D047F00090200007E0010009B0",
INIT_13 => X"0109000003E2000416C0804FE04140E80000F808010AB02033AC048A2A00003D",
INIT_14 => X"FFAFD082003B032FB987E04021D481D4000419060201E1A000044300B02033E8",
INIT_15 => X"AFEBFAFEBFAFEBFAFEBFAFEFFBFBFBFBBFCFBB0FFDFEFFEF2DFFFFFBFF802FFD",
INIT_16 => X"FEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBF",
INIT_17 => X"EBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFA",
INIT_18 => X"F491E166CC8553F86EDB5C88646FFFFFFFFFFFFFFFFFEBFAFEBFAFEBFAFEBFAF",
INIT_19 => X"1861861861861861861861861861869A69A61861AFBD54D5F871C71D475B15BC",
INIT_1A => X"0984C26130984C26130984C26130984C26130984C26130984C26186186186186",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE000000000000000000984C26130984C26130984C2613",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000",
INIT_22 => X"2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_26 => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFF",
INIT_2E => X"F5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA080402000000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"02010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_36 => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_37 => X"0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(26),        -- Port A data input
DOA(0)   => data_read_a_lo(26),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(26),        -- Port B data input
DOB(0)   => data_read_b_lo(26),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_27_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"00080A40000A41248002029000050A088000008242A0004404480002000A1155",
INIT_01 => X"F1FFF1C11F781C129C107DFFFE0860941E81258CA2B71C2220EC1B86E1A00002",
INIT_02 => X"183080988B2EAE00002BE001117C78C6848140CFFA0000800042008000011081",
INIT_03 => X"000003FDF3E47C74F7BCF36A203A47F6B8184210B6160820001318C60C204C63",
INIT_04 => X"7E28FEBF6FEEB3723F71017476DFC524397B6DF572EB6C8E175E70D90F539600",
INIT_05 => X"000F86064C8DDFE3B6FF50D1FC61DE39C8FCB91FF9671FE6B68984B5BCE40834",
INIT_06 => X"0000000800000042020C18300520620A80231BFE200181092CE7ED80DFC00147",
INIT_07 => X"8AC4AA3B0FD1FF201044110560884000840200520002080C23468D0300000282",
INIT_08 => X"2005F0784411E390A4880E3DF7E2FB0B8E717C7F411F3BC6D60B60FFDDE44001",
INIT_09 => X"18FFD757E7ED7A211E81C09818109E1F16B16B71092CE7ED81CF403601228C40",
INIT_0A => X"46FF730E5CCBCD55219AB55F0DEFABC7054880693016DD4C755AC16C1A884FFE",
INIT_0B => X"BC63F1683803C00E3440C3440C3440C3440C3440C3440C3440C3C2061A2061AD",
INIT_0C => X"56BF55CB165EC51D41880FA3F040202883B475062033186801137FF1BAD6F281",
INIT_0D => X"3B0000421E2B0F2E2AE215C808FFFA47FE62BAA86B1AB268E92AB56D5AB6AD5B",
INIT_0E => X"3B000025EC010080004000F808000098100F22520008003B00002F2252000800",
INIT_0F => X"00001042006BC0810600400003B80001002F22520008003B00002F2252000800",
INIT_10 => X"01E032000620000C0405EC010100100000F6000001C1003760410500008000EE",
INIT_11 => X"201D2120840039000817444404040E10020218DE282010A311AA002002040080",
INIT_12 => X"8000000AE888808101C20040BA4241080072001027F00080200007E0000001F0",
INIT_13 => X"0101000003E2000007C0800FE04040280000F8080002F02023AC04080A00003D",
INIT_14 => X"DDAFD082001B03249887E04001D481D4000009020201E1A000040100F02023E8",
INIT_15 => X"ADAB6ADAB6ADAB6ADAB6ADAB6BF1EBDABD8E270BF84A25C6ACB777E3FF800C6D",
INIT_16 => X"DAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6",
INIT_17 => X"AB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6A",
INIT_18 => X"100481CA860402104A471688747FFFFFFFFFFFFFFFFFAB6ADAB6ADAB6ADAB6AD",
INIT_19 => X"0000000000000000000000000008200000000000200072F210000001490E2168",
INIT_1A => X"A05028140A05028140A05028140A050080402010080402010080000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000A05028140A05028140A05028140",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000",
INIT_22 => X"2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_26 => X"10FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFF",
INIT_2E => X"F5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA080402000000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"02000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FF",
INIT_36 => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_37 => X"0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000000FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(27),        -- Port A data input
DOA(0)   => data_read_a_lo(27),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(27),        -- Port B data input
DOB(0)   => data_read_b_lo(27),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_28_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"02200AA400180030808802A900002A08001280A08A801044104A1000001818C3",
INIT_01 => X"50A00011460214428114180000882214413D0A71592A01D92213D28005210202",
INIT_02 => X"8A54800A210200111100C2110054289220810440030404010844000444410001",
INIT_03 => X"4200040822D4500001E0000028000002000211842010092000018C6295200631",
INIT_04 => X"00400000000B8000000140000005840C00000040002008808100048100100044",
INIT_05 => X"0000222200244400135110000135100000000000000000024CA0A01018000320",
INIT_06 => X"A004912008208040024489121144080400081000200008104000000020000041",
INIT_07 => X"A85800994000000A0200802004204420210001022AA8A0001122448142491008",
INIT_08 => X"0414000201800004080A000000124058200408000880004440004080160C4100",
INIT_09 => X"0080000206CB0821082B694D4D29400002002038104000000020003204000440",
INIT_0A => X"12000843066021001400040024440245400082D022040000400800081022C000",
INIT_0B => X"0002002C004001036050160501605016050160501605016050160280B0280B00",
INIT_0C => X"0012400810080414C0A800310840102182C62302A0194C08001680100E4040A0",
INIT_0D => X"05000002003004208208841401800040000A0000200814004198000400020001",
INIT_0E => X"0500000004000080000000000000028000002052000000050000002052000000",
INIT_0F => X"0000300000004001060000000000000900002052000000050000002052000000",
INIT_10 => X"0000000001200000000004000100000000000000050000002001050000000000",
INIT_11 => X"00002020840000004800040404040000120200A9000000010000002002040000",
INIT_12 => X"0000004800808081000002400040410800000090001000002000000000000910",
INIT_13 => X"0001000000000000144000010000402800000000000A1000010000080A000000",
INIT_14 => X"0080000000110006B08140000040000000000902000000000000410010000100",
INIT_15 => X"0080200802008020080200802101210810C39A66A90A85420413A82000000204",
INIT_16 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_17 => X"8020080200802008020080200802008020080200802008020080200802008020",
INIT_18 => X"110A00246972BD89A40A0C22E100000000000000000000200802008020080200",
INIT_19 => X"82082082082082082082082082082082082082080D35050758C30C31DE21102C",
INIT_1A => X"B0582C160B0582C160B0582C160B0580C06030180C06030180C0820820820820",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000B0582C160B0582C160B0582C160",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000",
INIT_22 => X"2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_26 => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFF",
INIT_2E => X"F5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA080402000000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"02000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_36 => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_37 => X"0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000000FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(28),        -- Port A data input
DOA(0)   => data_read_a_lo(28),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(28),        -- Port B data input
DOB(0)   => data_read_b_lo(28),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_29_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"79964E4BA01DACAB9E659792D00AAE160002829C7FDFEFCEE97C2815039D70C3",
INIT_01 => X"50BFF9AB0775343F9AB01DF80D5821FC0FFF3FEFD1AF9FF1207FFBC7B9720586",
INIT_02 => X"0D15846807D207200021C4E200D428A2018408600271C000720A0000003A2161",
INIT_03 => X"0002C009EEFC5F10F9B70178681B80FA3E000100765029A00019084345606421",
INIT_04 => X"3E6E023D27DA937C03E3407712E5CDA41E0924DC3D20B98AE905189F0BF8C000",
INIT_05 => X"902003C30E0447F877F930203E213F8CF01E3E00FC67C03A4D9C87525E510160",
INIT_06 => X"0012460003CC002036040811D919F402244293FEE00400CCB46BA4C164A08857",
INIT_07 => X"914800110FFC0001CC320C81D841418E82800100000041FCA1428575A0001108",
INIT_08 => X"0805FD0180E1F8C1111A0782082B50080508FF00048B124D4005C8AFF4154102",
INIT_09 => X"0180000ABFEF89250815568A8AD6ABC02A02A0B0CCB463B4C0748A720B1EA4C0",
INIT_0A => X"021410028450530014014002D445624DB481806A62840800C22800B8900042FF",
INIT_0B => X"0806522C0A40A50268D0068D0068D0068D0068D0068D0068D006A68034680300",
INIT_0C => X"8912E0A83289641F42A80561D040203182AC3D0AA0118A080036FFFC4F4164A0",
INIT_0D => X"050080424069F5A51250648801BFFFE0003E3E00A0685A85410C0816040B0205",
INIT_0E => X"050080080400028000000000000202900000A0F600000005008000A0F6000000",
INIT_0F => X"00023000001040214E0000000000000D0000A0F600000005008000A0F6000000",
INIT_10 => X"000000000120400800080400030000000000000205800008200D070000000000",
INIT_11 => X"000220A2C400000068008424260400001A0241DAC80001010000042016040000",
INIT_12 => X"00020048108484C10000034004414588000000D04010001020000000010009B0",
INIT_13 => X"000900000000000416C00041000140E800000000010AB0001100008A2A000000",
INIT_14 => X"A282C0000033010FB181E00020400000000419060000000000004300B0001100",
INIT_15 => X"02C0B02C0B02C0B02C0B02C4B12B312912831A27FCFE7FFB175B6FF800802594",
INIT_16 => X"2C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B",
INIT_17 => X"C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B0",
INIT_18 => X"EE7FFDF7FE783FFDFFEA0C00602FFFFFFFFFFFFFFFFFC0B02C0B02C0B02C0B02",
INIT_19 => X"BEFBEFBEFBEFBEFBEFBEFBEFBEEBAEBAEBAEBAEBBFFDF9FBEFFFFFFEBBCF9F96",
INIT_1A => X"FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFBEFBEFBEFBEF",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000FBFDFEFF7FBFDFEFF7FBFDFEFF7",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000",
INIT_22 => X"2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_26 => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFF",
INIT_2E => X"F5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA080402000000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"02000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_36 => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_37 => X"0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(29),        -- Port A data input
DOA(0)   => data_read_a_lo(29),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(29),        -- Port B data input
DOB(0)   => data_read_b_lo(29),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_30_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"FF9FE1F7FFBFFFFDFFD000000000000000000000000000000000000000000000",
INIT_19 => X"79E79E79E79E79E79E79E79E79E79E79E79E79E7AFBD75F5FDF7DF7FF7FFBFFE",
INIT_1A => X"3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE79E79E79E79E",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE000000000000000003F9FCFE7F3F9FCFE7F3F9FCFE7F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000",
INIT_22 => X"2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_26 => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFF",
INIT_2E => X"F5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA080402000000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"02000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_36 => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_37 => X"0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(30),        -- Port A data input
DOA(0)   => data_read_a_lo(30),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(30),        -- Port B data input
DOB(0)   => data_read_b_lo(30),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_31_8 : RAMB16_S1_S1
generic map (
INIT_00 => X"129000008004A00804A40000400800020000000C005FEA005800200400050100",
INIT_01 => X"A15FF18019700810180065FFFC0040801E80258CA2951C2200EC0906A0804140",
INIT_02 => X"146000808A0C060444692000402850040400408FF80000000010000000004000",
INIT_03 => X"000003F5D1202C70F654716A001A07F438184210960600000012108518004842",
INIT_04 => X"3E28FE3F6FE513703F70007472DA4128187B6DB530C1240A060C70580B439200",
INIT_05 => X"000F84040C088BE3E4AE40C1FD04CE38C0FC381FF8671FE01009048084C40010",
INIT_06 => X"0000000000000008000810200420620E00030BFE000181092CE7ED80DF800106",
INIT_07 => X"000000220FD1FF200040100540800000840200408002000C2244890200000200",
INIT_08 => X"0011F0780011E38004800E3CF3E0B1118C31747F000B33820209206FC9E80000",
INIT_09 => X"187FC301B124F2001600000000001A1F00110101092CE7ED81CF000401228800",
INIT_0A => X"0477330C4889CC012188310E08812982050800A91012494C31004124080886FE",
INIT_0B => X"9861D1403803800C1000C1000C1000C1000C1000C1000C1000C1800608006084",
INIT_0C => X"020400830602410901000D02D0002008012054040022102001017FE190022201",
INIT_0D => X"3A0000401E030B0C20C20188087FFA07FE203A80010002608030102008100408",
INIT_0E => X"3A000005E8010000004000F808000010100F02000008003A00000F0200000800",
INIT_0F => X"00000002006B80800000400003B80000000F02000008003A00000F0200000800",
INIT_10 => X"01E03200060000080405E8010000100000F600000081003740400000008000EE",
INIT_11 => X"201D0100000039000007404000000E1000001846282010A211AA000000000080",
INIT_12 => X"80000000E808000001C200003A0200000072000007E00080000007E0000000A0",
INIT_13 => X"0100000003E200000280800EE04000000000F8080000A02022AC04000000003D",
INIT_14 => X"9C06D082000A03200806A040019481D4000000000201E1A000040000A02022E8",
INIT_15 => X"0401004010040100401004010060C040040C200950402090128057C3FF800C60",
INIT_16 => X"4010040100401004010040100401004010040100401004010040100401004010",
INIT_17 => X"0100401004010040100401004010040100401004010040100401004010040100",
INIT_18 => X"000000000000000000001000802FFFFFFFFFFFFFFFFF81004010040100401004",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000",
INIT_22 => X"2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_26 => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFF",
INIT_2E => X"F5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA080402000000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"02000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_36 => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_37 => X"0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(31),        -- Port A data input
DOA(0)   => data_read_a_lo(31),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(31),        -- Port B data input
DOB(0)   => data_read_b_lo(31),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_0_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"ED39BA795990D275FB4A6E96ACC4731DEA4598B0AFB54867F6EE4618C3749803",
INIT_01 => X"58A0047C8607844847CA180001E4A2404042106208408208C2002069161734B3",
INIT_02 => X"8B1EC9562121F8051500147A0E5629A302CF28400615F5787B09FBF999BB1EFD",
INIT_03 => X"404EFC0A2AD6100F01A88E851CE47803C280110521898F6996088862C7B22221",
INIT_04 => X"C0D001C0100AEC83C008E7880D01A64661800002C21A52C590D2012194804844",
INIT_05 => X"650002C3F08754001B51981E007910070F01C1E003980015A204C22F32328BAF",
INIT_06 => X"BCDA4677CAEE7CF5BB870E1DDB9889C5FBFC440129A0604442180238203F70C1",
INIT_07 => X"7AAE0088B02000C2EC3A0E829836E0AF3325372E2AA8FDF3C18306758B24197A",
INIT_08 => X"D7E40002F7AE005FFB4730010411400A61080000F7F4C464B58294901606D5A5",
INIT_09 => X"C4801C40469B0CA9881A28C141118000C5A85A60444210123820B43B40804274",
INIT_0A => X"400800219010107ED453C041B13216656074EA560F0092A24856B05312226900",
INIT_0B => X"27122C3E04E03383E2781EA781E2781EA781E2781EA781E2781C33C0613C0E29",
INIT_0C => X"74EB1F50D0758A9650E520610A6A57A5529E2B439499CF96B086000000B09870",
INIT_0D => X"04F07E024108F4E28638EC57250004480155C1375A97A9121F8BA749D3A4E9D2",
INIT_0E => X"04F07E42177EFDF8570184071575970F8FC07D5BFF078004F07E007D5BFF0780",
INIT_0F => X"8F85ECB1FE047F5FB7B30E0700461E5AF8007D5BFF078004F07E007D5BFF0780",
INIT_10 => X"C0184D07C1DF15C7E3E2177EFDF8C3C03009C3CDD47C7F403FB3FDF89701C011",
INIT_11 => X"4F80FE659C6104C6D7103F9D1D064189B5924418D65FE45DEE55BBEDE34CF900",
INIT_12 => X"6395F64207F3A3A1483136B881FCCB38C2098DACA01FFF603F80001F80FDC81F",
INIT_13 => X"FED151E01015C3BB507D3F811FBEC32B81840714F8D91F4FC513F37C8AE07002",
INIT_14 => X"61692F293185D8D724E15D3FCC6B7C236FE0691A9500125C1F83F8CC1F4FC507",
INIT_15 => X"E93A4E93A4E93A4E93A4E93A4F942F90E9628540052090650525A0000066A00B",
INIT_16 => X"93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4",
INIT_17 => X"3A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E",
INIT_18 => X"09B56C74DAB15D1CF13501AA495000000000000000003A4E93A4E93A4E93A4E9",
INIT_19 => X"2082082082082082082082082082082082082082082084E41DC71C7155F3898E",
INIT_1A => X"3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F8208208208208",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE5294A5294A52800003E1F0F87C3E1F0F87C3E1F0F87C",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000030FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"A975EFFFAABDE00FFAEBDFFF5D2EAAAAAF7AEBDEBA0000000000000000000000",
INIT_22 => X"8000155087FC0155F7D168B55007BFDF45085168ABA002E82145085155545F7A",
INIT_23 => X"FFFD7545AA8028A00A2802AABAFF8028BEF5D7FFFE10005542145557FD5545FF",
INIT_24 => X"F7AEAAAAAA2FFFDF4500043FE105D2E954BAF7FFC0010080017555555568AAAF",
INIT_25 => X"A5D5168A00A2D142155005142010FFAE820AAFF842AABAA2AE95545FFD168ABA",
INIT_26 => X"FF5D2A821550000000BA007FD55FF5D7FC0145007FD7400550415410002E974B",
INIT_27 => X"F455D5142000082E82145FFD17DFEFFFD168BFFF780000BA007FE8AAAFF803FF",
INIT_28 => X"0000000000000000000000000000000000000000AAFBEAA00007BFDFFF082EBD",
INIT_29 => X"AABEA495FC716F002A975FFE3AA95E00EBAEBDFD75D2AA8A80EA8E2FE3F00000",
INIT_2A => X"56A16D557BC257D415E0216FA3F1E8FC0145B68B551475FAF6D1C556F0AA1C24",
INIT_2B => X"7FD24AFE3D02DAAAE12BD5545A2803AA0000542A0070071C50BAFEF1FAE0016D",
INIT_2C => X"A8B50F55A2F150005A3A438BD04AFAB8F550A8010E004924874825D7FEAA8548",
INIT_2D => X"A2A5504001C74BA42A1571E8028E3DB7816D0120155EA568E870BAEB8A05A2AE",
INIT_2E => X"2FFAFD2A82485FD2415A105C21451ED42A002545E055FFBE81D0BE8EA8A3AA05",
INIT_2F => X"100AA1D0F6F480B6A555A2A57A002A3D5FDB6A5C7E3DFFFE90B45B47ABA497A8",
INIT_30 => X"A0AFE80A8B0A000000000000000000000000000000000000000000000B55EAAA",
INIT_31 => X"ABEF5D557FEBA55022A3F70C6B405F4D2AE975EFAAAAB5E1AF3AABFF45592E88",
INIT_32 => X"411A8DED57CE1055555E5F58EFFC01FE2CACB65F520EBE9EF67D7BEA1FD5D556",
INIT_33 => X"A4AD0079C75D6070CC5CBB0280C029ABAA3EBC114728007521170821CE0FDE69",
INIT_34 => X"2A95E02A2AAB5EB0F280800EFAEE9F5D18F3142341D5DEEBEF55080034E0A592",
INIT_35 => X"B69C30E02116220415A9540AA854140A0A2047F353AAF6C77F7F20D968BF5781",
INIT_36 => X"ABEBE1B4D792A4AD1183454180DD3FDCAAAB7C91565455C141E41887D58AC448",
INIT_37 => X"F0000001FF01EABC4B8014174FF7DA80F52FEDE6BE93172D7D625B556EEAB157",
INIT_38 => X"FF0000001FF0000001FF0000001FF0000001FF0000001FF0000001FF0000001F",
INIT_39 => X"0000000000000000000000000001FF0000001FF0000001FF0000001FF0000001",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000100000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(0),        -- Port A data input
DOA(0)   => data_read_a_hi(0),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(0),        -- Port B data input
DOB(0)   => data_read_b_hi(0),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_1_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"212C001411984004084D000508C53810A03D1450E839B003342114428A000803",
INIT_01 => X"08000011400A100A81160000008C005400400002000000000000028001340000",
INIT_02 => X"C084484000002014400205851002007030450E0000A606C8C44CB4C6666C00E0",
INIT_03 => X"33DF380008164004000002000C80400002031943000101091608463061120118",
INIT_04 => X"4140008000000002000064000400004201000000000210458010070080100433",
INIT_05 => X"8500101040200000010009100000000508000100000000002010600100208D04",
INIT_06 => X"B5EDFDE24618AD433060C182BA860044204C000008A004100008000820280020",
INIT_07 => X"581E02100020000A81244890AA20263030517F122AA801F0983060AC564BF808",
INIT_08 => X"00820800C7A00045B103200000140A02234808000584000004808400020011A4",
INIT_09 => X"0000104000020082800808111008400000200204100000100820800144000414",
INIT_0A => X"12804062945211441E13C051156E800008402802060C94000040901102800000",
INIT_0B => X"24002006406401918C191AC191A4191A4191AC191AC191A4191A00C8560C8D29",
INIT_0C => X"0408010040050880383820080F105F05800302E0E08842422006000000041032",
INIT_0D => X"05000600000090C1841808172580000000008008020084082080204010200810",
INIT_0E => X"0500066210000178470184000000878402C000001E07800500062000001E0780",
INIT_0F => X"00003C404600000011A30E0700000009382000001E07800500062000001E0780",
INIT_10 => X"C0180000012010C20022100000F0C3C03000000055200340000000F88701C000",
INIT_11 => X"05800241186100004D100098190240001290002050068000001010486140F900",
INIT_12 => X"0000164A001303204800026880048230C2000094A0000F601F8000000001C908",
INIT_13 => X"12D051E01000000154200580003C030381840000004B08014401025480E07000",
INIT_14 => X"40082300218450C2800010094000482142E0601895001000000041C408014400",
INIT_15 => X"0802008020080200802008020080008208600500A82A15008000000000468000",
INIT_16 => X"8020080200802008020080200802008020080200802008020080200802008020",
INIT_17 => X"0200802008020080200802008020080200802008020080200802008020080200",
INIT_18 => X"BABEFC54A0810C7452B5420A1000000000000000000002008020080200802008",
INIT_19 => X"AAAAAAAAAAAAAAAAAAAAAAAAAAA28A28A28A28A2A8218D2C0C92492581328A46",
INIT_1A => X"2E974BA5D2E974BA5D2E974BA5D2E975BADD6EB75BADD6EB75BAAAAAAAAAAAAA",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFF6318C6318C63000002E974BA5D2E974BA5D2E974BA5D",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"00000000000000000000000C0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"002155557FFFFFF007FC21EFA2FFD74AAAAD5555550000000000000000000000",
INIT_22 => X"7FD75FFAAAA800AAF7AA974BAFFFBE8B45F7AEBDF455D2EAABEFF7FFE8BFF5D0",
INIT_23 => X"0557DF45AAD1400BAA2AE801550051555EFF7AA95400552AAAABAFFD1574105D",
INIT_24 => X"FFFBEAB55F780020AAAA80020AA082EAAB5500517DF555D2EAAA105500001550",
INIT_25 => X"AF7AE820AA0851574BAA2D1574AA5D7BFDEBAFFD540155557FD5400F78028BFF",
INIT_26 => X"FFFFD56AAAAFFFFD7555AAD168B45AAAEAAABAFF842ABEF5D517DF55552A974A",
INIT_27 => X"4BAF7AE80010082A97410557FEABFFAAFBE8BEFAAD1575EF557FFFE10557FFFF",
INIT_28 => X"00000000000000000000000000000000000000005D7FFDF4500043FE105D2E95",
INIT_29 => X"A8BC2EBDFEAF7F1F840017D4975D2FEF147FC51C7A2FBD5490BFD1C056A00000",
INIT_2A => X"AA8AAAE3D145410F7F1D55D71C002DABAEBAA974BAF7FFEFB45FFAABDF55492A",
INIT_2B => X"0E2AE85028B40155145F7AF6DBED5450AA1C2080BEF495FC71D54124924385FA",
INIT_2C => X"571D2E28E38E0216FA2D1E8E80140F45082B4002D082082AB8B6DBEDB7DF7F54",
INIT_2D => X"A97F7AF6D417E92482BF84020BA495557E3FF78E021FF1471FDEAAFFD56F16D5",
INIT_2E => X"7002FD74951D71EDFFABFD16FAAAE92BD5545A2DA3FB7DAAD4AAAAF487BC70BF",
INIT_2F => X"550A8010E00492487482FFFE82A85EBAE2FFC55554ADBD7A2FFC7BEFF6FFD7FC",
INIT_30 => X"400FBF9424F7000000000000000000000000000000000000000000000547AB8F",
INIT_31 => X"DF55F7AABFF55082CA8B4DF6C1E8F5E5400021EF005162BEF047FD5545AAFBF7",
INIT_32 => X"404547184164AA5D2EBEEB0A2D555410D3555714F8338AAAA1D0AE974AAF7FFF",
INIT_33 => X"AEABFFDF79DCBF755962010BDCBBC21455D7FEABEF75550ACBB7582225FF5843",
INIT_34 => X"D57D412F7D55F5E50C7F401BAAE8403CF5A3FFEAAEB083BC1000FF8409000512",
INIT_35 => X"2AA9FEAFDF7F431A9F7FFE81FF013A8001AFF801F8BA0C57740BDAA0688E5405",
INIT_36 => X"A2FBF7FED2C7F955445079E280A00C56145EF5D16BABAA3EBC3157ABD5FFE55F",
INIT_37 => X"0000000000596EBEF55080034E0A592A4AD00FB863550229BCABEB7DA403FFFD",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000100000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(1),        -- Port A data input
DOA(0)   => data_read_a_hi(1),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(1),        -- Port B data input
DOB(0)   => data_read_b_hi(1),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_2_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10E006600180111284380310006289800480032283E000A34301002001A0817",
INIT_01 => X"A14AC00A1079284D04A044A54E504368404000720885800802000006ECD10200",
INIT_02 => X"92250052A0348C310102048800A8507000040C8550200000480E0080001321E0",
INIT_03 => X"020204E4593C0824400C2220483042809292430400440180000890A4C9400242",
INIT_04 => X"486854B141002252142241502460480031B94420634850069A42241009610A04",
INIT_05 => X"800504244080892105AA6010A44882144840910A21220A8C820025E4A0000B00",
INIT_06 => X"A000442802280000340810209C444804206000AC800088096A0EA8C022208012",
INIT_07 => X"309820A848E0AA09826489A5CC49002001020112028201F8A20488260000108A",
INIT_08 => X"2400582881E0C1419D12041455509341A539C42A0D8208099002801700D10103",
INIT_09 => X"110D525861263100009200151409130A3C80C8C8096A06B8C12088400A9C2080",
INIT_0A => X"0451394CD0391A441583C04B580040089581001342801044877200D002A00DE0",
INIT_0B => X"144423040240450114901149013C9011C9013C9011C90134901144801A4808A5",
INIT_0C => X"D8A5345206D2C10082080A90C00000188150100C202A4640000E2B4081969420",
INIT_0D => X"050080400A0391A51240C480000AA902AA009028C83220008086952B4285A54A",
INIT_0E => X"05008021C00000000040000000020288000500000008000500802A0000000800",
INIT_0F => X"0002300000428000000040000000000D002A0000000800050080250000000800",
INIT_10 => X"0000000001204004000508000000100000000002054000130000000000800000",
INIT_11 => X"000C00000000000068144000000000001A000106200010021002000000000080",
INIT_12 => X"0002004A880000000000034098000000000000D024A000000000000001000900",
INIT_13 => X"00000000000000041400000A8000000000000000010A00000284000000000000",
INIT_14 => X"012100000002000280000000011080C000000000000000000000430000000260",
INIT_15 => X"A769DA769DA769DA368DA36CDA3A9A13A14801404134DA84A024024155000399",
INIT_16 => X"168DA769DA769DA769DA368DA368DA368DA769DA769DA769DA368DA368DA368D",
INIT_17 => X"68DA168DA169DA569DA569DA568DA168DA168DA169DA569DA569DA568DA168DA",
INIT_18 => X"138D70C030B51C50C7D000A2012F81F81F83F03F03F069DA569DA569DA568DA1",
INIT_19 => X"1041041041041041041041041041041041041041024860208165965975960040",
INIT_1A => X"25128944A25128944A25128944A25128944A25128944A2512894104104104104",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFF8421084210840703F25128944A25128944A25128944A",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"00000000000000000000000F0FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"415555087BFFF55A2AA800BAFFAE9540008002AA000000000000000000000000",
INIT_22 => X"7FE8B555551421455D0002145552EBFEBA007FC21EFA2FFD75EFAA8415410AA8",
INIT_23 => X"FFFE8B45552EBDF45FFAEAABFFF7FFE8B55F784155EFA2AEBDEAAA2FBEAABA5D",
INIT_24 => X"5D2AAAAAA5D2E820BAA2FBEAB5555557DF55A2AEBDF555D2E954BAA2AA974BAF",
INIT_25 => X"A5D04021EF557FC21FFAA8428BFFAAAA954AAAAAAAAAAAFFD1574105D7FFFF55",
INIT_26 => X"EFF7800215500557DF55AA80001FFAA80001550055575EFFF84021555D043DEA",
INIT_27 => X"B5500517DF555D042AA10A284154005D0015410085568A00FF80175FFA2D17DF",
INIT_28 => X"00000000000000000000000000000000000000005D00020AAAA80020AA082EAA",
INIT_29 => X"D55D2BE800042AFE8E1557D0075D2F45BEAA800AAFFAA9543A080038A2A00000",
INIT_2A => X"0BDEAAA2FBF8AAA557BE8B6D5D5FFABEF49040017D5D20B8EAA007FC51C7A2FB",
INIT_2B => X"0E174BFA02A974BAF7F5EFB455D2ABDF55492AA8BC7EBDFEAFEFFD00105FFBC2",
INIT_2C => X"3D155E105571D55D71C002DABA5524820BAB6FFEFB6D555578F7DB6A0BDF7D48",
INIT_2D => X"092A071555D5E3AE821D00001FF0871C016DBED1FDE90E3A497492B6AAADAAAE",
INIT_2E => X"0E3DA3DFD5E3DFFFBD5A38A021551C5F7AF6DBE8F401D7B6A0001470155C51D0",
INIT_2F => X"82B4002D082082AB8B6D1C5B7DF7FF78E075C5BE8555400550A38428007FED00",
INIT_30 => X"4AA00042AAA2000000000000000000000000000000000000000000000410F450",
INIT_31 => X"AAAA007FD5555AAFBD7545FBB8020A3F7AE975EF005560B55F7AA800AAF7AA95",
INIT_32 => X"E8F5EFF84165EFF7802BAB0A2FFEAABA557BEABEF057D68F5F5A00021EF55042",
INIT_33 => X"52ABFFFF841FFE75CA882108202E974AAF7D57DF55D7AABFF5428ACA8F45A6C1",
INIT_34 => X"84174A8FFAEBFEB0A2D55541051555694F002CA8AA80800020AAF7FBFFFEF045",
INIT_35 => X"7AAA155F595542455512A975455D3AA8A005500151FF0C57401E5F3D1E00A1A8",
INIT_36 => X"5D2A8A0B882FFFFE10AAAAAB755A66B6AF56A2AA801455D7FE8BFFF680800FFF",
INIT_37 => X"00000000000C3BC1000FF8409000512AEABFF5D79FCAF774AE005BE789555400",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000200000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(2),        -- Port A data input
DOA(0)   => data_read_a_hi(2),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(2),        -- Port B data input
DOB(0)   => data_read_b_hi(2),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_3_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"210C44A20020248B08431120001604B8156023104C4077133420400A02380202",
INIT_01 => X"015A2A424080216D3C2462C99E104B49404040028804A0080A000C16A0D90A0C",
INIT_02 => X"C0A4065000F0A95011000D1501005270B4045AB330860281CC08008222170060",
INIT_03 => X"AD22014098340394A4021320080841C40B411B4298042180002846B06900811A",
INIT_04 => X"244B32A86D20014A0D20403194904900071A24110F0BF400F85F92420E0C946E",
INIT_05 => X"80331030442898B4812840D0500008C528280B063006A64CA30004E5A4E40304",
INIT_06 => X"90016CA00E380042302040A0BC47160424428198C0038C89904E640023600816",
INIT_07 => X"1288020843A66620816049908AA0061011CA0142000009F0A810292E7402F088",
INIT_08 => X"20003C9984A0AC411102014D34EC2200214D5099048823019603A01A49410103",
INIT_09 => X"001CD74C4826220010A8891451284B661CA24A4C899046740121824004100080",
INIT_0A => X"44C9516DC0135C45159BE45F112B48804DC10203021290400772C0F402820D4C",
INIT_0B => X"B400624402404501A49018490184901A4901A4901849018C901A648056480C2D",
INIT_0C => X"D7A9B54000D7C10820680D08C420180381211081A022160000266723E1909021",
INIT_0D => X"400080200E199A4A2CA2994C0399981666409800CA52E4890806BD6B56BDAB52",
INIT_0E => X"40008008E00000000000000000024008000C8000000000400080028000000000",
INIT_0F => X"000A000000588000000000000000200400088000000000400080078000000000",
INIT_10 => X"0000001000004004000D800000000000000000022040000B4000000000000000",
INIT_11 => X"001A0000000000082006C000000000020804087220000122000A000000000000",
INIT_12 => X"00020800B8000000000041002E00000000001040466000000000000001020080",
INIT_13 => X"00000000000000048200004A600000000000000003008000320C000000000000",
INIT_14 => X"432900000222200871028000210400C4000000000000000000080200800030E0",
INIT_15 => X"AF6A5AF6A5AF6A5AF6A5AF6E5AFADA91AB68000101B4D20C08EC461733804A19",
INIT_16 => X"B6B5AF6A5AF6A5AF6A5AF6A5AF6A5AF6A5AB6B5AB6B5AB6B5AB6B5AB6B5AB6B5",
INIT_17 => X"6BDAB6B5A96ADAF6A5AD6ADAF6A5AD6ADAF6A5AD6BDAB6B5A96BDAB6B5A96BDA",
INIT_18 => X"C78C706428A14C586290008A044D54AAB556AA9556AAEBDAB6B5A96BDAB6B5A9",
INIT_19 => X"92492492492492492492492492410410410410412821600001249249015303C0",
INIT_1A => X"351A8D46A351A8D46A351A8D46A351A9D4EA753A9D4EA753A9D4924924924924",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000001543B351A8D46A351A8D46A351A8D46A",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"43DF55FFAA955EFA2D168B55557BEAA000055420000000000000000000000000",
INIT_22 => X"7BE8BFFA2D155410AA8415555087BFFF55A2AA800BAFFAE9554508002AA00AA8",
INIT_23 => X"52ABFEBA007FC21EF007FD75FFAA841541008002AB55AAAA955EF005568A0008",
INIT_24 => X"005168B455D042AB45F7FFD741000042AA10AAAABFF5508003FF555D00021455",
INIT_25 => X"0A2D1575FFF7AA975555D2E80145F78415545082EBDEAAA2FBEAABA5D7FC0155",
INIT_26 => X"55552A954BAFFFFE8B55552EBDE00F7AEAABFFF7FBEAB55F7AABDEBA5D7FC201",
INIT_27 => X"F55A2AEBDF555D2E954BA002EAAABA002A821EF5555554AA087BC01FFFFAAAAB",
INIT_28 => X"0000000000000000000000000000000000000000082E820BAA2FBEAB5555557D",
INIT_29 => X"95578080038A2AA28E3AF55E3A0BA5D7AADB6FB7D5D7FEAA3808554203A00000",
INIT_2A => X"0925D7085F6AA10087FEABD7AAD57AEBAB68E1557D1475FAF45BEAA800AAFFAA",
INIT_2B => X"04AAFFA41040017D5D20B8EAA007FC51C7A2FBD55D7BE80004AA1E8E2AB55B6A",
INIT_2C => X"2FBE80AA557BE8B6D5D5FFABEF49002FB55FFF5D0438140E2FA38B6AEBFF6D1D",
INIT_2D => X"AB8ABAE925D21C7010EADB525D7FFAE975C75D0A901FFFF801557D1C20B8EAAA",
INIT_2E => X"20875C21D5EB8AA8FFF012A954BAFFF5EFB455D20BDE00EBAAA8BC7EBDFEAFEF",
INIT_2F => X"BAB6FFEFB6D555578F7DB6A0BDF7DEB8E125FF002EADA921420871D74971D248",
INIT_30 => X"ABA0051400A20000000000000000000000000000000000000000000001C24820",
INIT_31 => X"8B55F7AA800BAF7AA955EF00042AAA2A2AEAAB55A28408145AAFFFFFFF5D7FEA",
INIT_32 => X"020A35D2ABEF55F7800015F087FEAA00007FEAB55FAD568AA2AFAE975EF55516",
INIT_33 => X"ABFEAAF7AE9DFF759A82AEF70800021EF55042AAAA007FD55558A7BD7145FBB8",
INIT_34 => X"84175EF55002AAB0A2FFEAABA557BEA3EF057968F575D003FF55F7D5420BA5D2",
INIT_35 => X"A8429F45A7D5EAF5FFBAEAAA10554155400AAFFD5145FBAC9755F05040255FFD",
INIT_36 => X"550415557085540000005156155FE90A8F5C082E974AAF7D57DF45552A3FF10A",
INIT_37 => X"00000000005500020AAF7FBFFFEF04552ABFFFF843FFE77C80825BC052ABFE10",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000100000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(3),        -- Port A data input
DOA(0)   => data_read_a_hi(3),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(3),        -- Port B data input
DOB(0)   => data_read_b_hi(3),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_4_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"A108400020612C80284210081034849800A000303100048B3432C82904204002",
INIT_01 => X"21066802000820491C00650E1E004360403008418984014902030906A8D10200",
INIT_02 => X"120404E00E4C0600000206100008402005040C00F104008040080080001310E0",
INIT_03 => X"DCA201514D1C0D706C5CF010083A0708BA0841945004010000080084C1000002",
INIT_04 => X"5C4CF21C48B133483C80417570D000083A62488074C1350EA60D785C0A6B0619",
INIT_05 => X"000F0400028083B381A60001E5546EB5C0E2B81E4166DE000139200004E50940",
INIT_06 => X"80004408020800023000102098000204A040038600018019004B800123208806",
INIT_07 => X"120C20204665E1008024188488800000001A01520000A1F08044892400001088",
INIT_08 => X"0801007AC0A1EB413102063CF3E0B3028D29F407059B0B000205A801C2200102",
INIT_09 => X"106052400922D00406BE1002C6150F41200280001900439001FD8A0004142000",
INIT_0A => X"047F2201D899BA503583504B58AB80804540001202805544314041B48A888EC5",
INIT_0B => X"1441E3443043410C5010C3010C1010C3010C1010C1010C3010C14086980861A5",
INIT_0C => X"020000A02600000805400502C0A0004A00625015000A12000026E1E180011220",
INIT_0D => X"400000000E43930C20C20188120782861E4004A800600401A030001008080400",
INIT_0E => X"40000021A8800000000000000000400800170024000000400000310024000000",
INIT_0F => X"0008000000AA80200800000000002000003400240000004000003B0024000000",
INIT_10 => X"00000010000000040004A080000000000000000020400006C008020000000000",
INIT_11 => X"002C008200000008001B4020200000020000090760000200110A040010000000",
INIT_12 => X"00000803E004040000004000E801040000001000086000000000000000020040",
INIT_13 => X"0000000000000000810000164001008000000000020040002240008020000000",
INIT_14 => X"04001040026026004000000002940040000410000000000000080000400000B8",
INIT_15 => X"040080201004008060000001806AC000004890015124D880100886D8F0014420",
INIT_16 => X"4010000180600000018020100400802010000080601000008020000401802000",
INIT_17 => X"0100000004008020180600000000000180600802010000000401802018020000",
INIT_18 => X"3807E05000140634504048820064B261934D964C326980004010000080600806",
INIT_19 => X"AAAAAAAAAAAAAAAAAAAAAAAAAAA28A28A28A28A2934C8D0CCD145144C0A28A06",
INIT_1A => X"068341A0D068341A0D068341A0D068351A8D46A351A8D46A351AAAAAAAAAAAAA",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000000173F068341A0D068341A0D068341A0D",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"57FE10FFFBEAA10007FD7410FFAA97555082A800AA0000000000000000000000",
INIT_22 => X"7FEAA00007BE8AAAAA843DF55FFAA955EFA2D168B55557BEAB45005542000005",
INIT_23 => X"87BFFF55A2AA800BAFFAE9555508002AA000055574105D2A800AA00043FEBA5D",
INIT_24 => X"A2D17DE1000517FE10AAAAA8AAA002E97545557BC00AAA2FFEAAAAAA84155550",
INIT_25 => X"0A2D157400AAAE974AAAAAA974BA08002AB55A2AA955EF005568A00087BE8BFF",
INIT_26 => X"BA080002145552ABFEAA007FC21EF007FD75FFAA8417410A2D140000F7FBC201",
INIT_27 => X"A10AAAABFF5508003FF55F7D568A00552EA8BEFA2AABDEAA087BEAAAAA2FBD54",
INIT_28 => X"000000000000000000000000000000000000000055042AB45F7FFD741000042A",
INIT_29 => X"EAB7808554203A145178E00FFFBE8A101475D5400F7A49057D0824850B800000",
INIT_2A => X"E8008200043FE925571EFA380871C7028A28E3AF55F7A0925D7AADB6FB7D5D7F",
INIT_2B => X"F5FDA38BE8E1557D1475FAF45BEAA800AAFFAA9557D080038AAA145157428492",
INIT_2C => X"85F6AA10087FEABD7AAD57AEBA08517DE00AAAEA8A9200249056D4175C5092AA",
INIT_2D => X"FEDB42028EBFBC2028BED152438AAA092492AAA4954281C0E2FB55B6A0925D70",
INIT_2E => X"A0875EDA80BEF1C743840040017D5520B8EAA007FC51C7007BD55D7BE80004AA",
INIT_2F => X"55FFF5D0438140E2FA38B6AEBFF6DBE84AAEBAF7DF6AA00412EAABFFAA803DEB",
INIT_30 => X"1EF0800154B200000000000000000000000000000000000000000000041002FB",
INIT_31 => X"0145AAFFFFFEF5D7FEABFF0051400A25D5568A00FFFFEAA105D5155410FF8402",
INIT_32 => X"2AAA25555410BA082E8201000043FE005D517DEBA0851574B2AAAEAAB55F7840",
INIT_33 => X"4001FF005575408AA557FEB2FFAE975EF555168B55F7AA800BAF7AA955EF0004",
INIT_34 => X"2ABFF55F7800015F087FEAA00007FEAB55FAD568AA200557DE00AAAAAAA00080",
INIT_35 => X"87BD6145FAAC000A2A6FBC00BAAAFBC00BAF7D1550AAAA8002010F2AC154B25F",
INIT_36 => X"082EA8BFFAA843FEBA08517DE00F3F9574B30800021EF55042AAAA007FD55550",
INIT_37 => X"000000000008003FF55F7D5420BA5D2ABFEAAF7AEBDFF779A82AA43F7FBE8A00",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000200000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(4),        -- Port A data input
DOA(0)   => data_read_a_hi(4),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(4),        -- Port B data input
DOB(0)   => data_read_b_hi(4),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_5_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50DF4A0791B3FCB694379283C81FD996A091832102004A337A20E07C0C1E006",
INIT_01 => X"294014468000A04D5C6A60000C34C24841280A00084000C8C212892EEAD53235",
INIT_02 => X"50AE41540CA1D9100002171C1F0A5171134E2A200D8633F8CD09DBFBBB970E7C",
INIT_03 => X"214E3C521D16021B64430CC51C45B8154689094241898749920842946B90010A",
INIT_04 => X"A2F20F7D7A314CB5C208E28A1BF0224A448920028A185340D0C20B2690000C22",
INIT_05 => X"7520B430B20B984809A8886E230C6106371146E1829941C58310402C600381CF",
INIT_06 => X"9CC96CD7C63A7495B9A356ACBC4601C57FD44F8549A46490261C4B39203F7080",
INIT_07 => X"12A88800B029E0C0A12C4B92AA36A2111167357C220095F3C8952A2E5D26F078",
INIT_08 => X"F3F00503B4AE105B534711820C0C0A1043080300F7E0E728B1829C2FEA0A95A1",
INIT_09 => X"C5184F084136848C9298A8560688F480C58858449026145B3830F40944906234",
INIT_0A => X"50EB4124D2B3902BF5C9700C1199DCA84DF46A974F92C7E28F1630D38088A438",
INIT_0B => X"B3144E5636E3178C86B8CC6B8CA6B8CE6B8C86B8CE6B8CA6B8CC15C6435C670C",
INIT_0C => X"79E51E70E070AA8132252008360A7E91504104C8948047D6B0AE1FE440B28A71",
INIT_0D => X"05F0FE40014090400400080329FF8089FF49611F589765923E139F09C78CE7C6",
INIT_0E => X"05F0FE64037FFD7857418407157797878F005F0DFF0F8005F0FE205F0DFF0F80",
INIT_0F => X"8F87FCB1F8053FDEB9B34E0700461E5FF8205F29FF0F8005F0FE205F29FF0F80",
INIT_10 => X"C0184D07C1FF55C3E3E0037FFCF8D3C03009C3CFD53C7E001FF2FAF89781C011",
INIT_11 => X"4E0CDF47186104C6FF177BD939024189BF900401165D645CEEF5BBCDF148F980",
INIT_12 => X"6397F64AEF7F2320483137F8A9BF8A30C2098DFCA06FFFE01F80001F81FDC94F",
INIT_13 => X"FFD051E01015C3BF553D3E0E5FFE838381840714F9DB4F4FA213F774A0E07002",
INIT_14 => X"8B652E2B3120C81284641D3E8DBF7D636FE070189500125C1F83FBCC4F4F80EF",
INIT_15 => X"E7394E339CE138CE5394E33D4E1E0E30E1208C251134921C12A44103F064014B",
INIT_16 => X"7384E3394E338CE538CE1394E3384E738CE139CE1394E7384E339CE139CE5384",
INIT_17 => X"38CE139CE1384E7384E7394E3384E738CE539CE139CE538CE5384E3394E7384E",
INIT_18 => X"7F7B9DB7FF3A1B6DB7ED438A9C3124B2DA6924965B4D384E7384E339CE138CE5",
INIT_19 => X"FBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEF9F7CFDFDDCF3CF3DF5E5BB4E",
INIT_1A => X"7BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEFBEFBEFBEFBE",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE000000000000118D27BBDDEEF77BBDDEEF77BBDDEEF7",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"E955450055421FFFFFBC0010AAD5574BA557FFDFFF0000000000000000000000",
INIT_22 => X"D5575EF55517FF5500557FE10FFFBEAA10007FD7410FFAA97410082A800AAAAA",
INIT_23 => X"FAA955EFA2D168B55557BEAB55005542000007FD74000055574BA5D7FD7555A2",
INIT_24 => X"007BC00AAAAAEBDF45A28428B45FFD168BFF00002AABA5D2ABFFFFAA843DF55F",
INIT_25 => X"AFF80174BAAAD1555EF5555555550055574105D2A800AA00043FEBA5D7FEAA00",
INIT_26 => X"FFAA8415555087BFFF55A2AA800BAFFAE95555080028A00A2FFFDE00F7D57FEB",
INIT_27 => X"545557BC00AAA2FFEAAAA082A97545F7D5420BA5D2E821FFA2D5554BA557BD75",
INIT_28 => X"000000000000000000000000000000000000000000517FE10AAAAA8AAA002E97",
INIT_29 => X"9043D0824850B8A2AE9756D145B401FFFFFFC7010BEDF524AA5571FDFEF00000",
INIT_2A => X"1524BA5571D757DB6D5525EF555178F6D145178E00EBFBE8A101475D5400F7A4",
INIT_2B => X"24BFFFFA28E3AF55F7A0925D7AADB6FB7D5D7FEAB7D0855420BA1471D7438085",
INIT_2C => X"0043FE925571EFA380871C7028B6AEBDF45B68A28B6DEBDF6DBEF1C0A28AAA55",
INIT_2D => X"A2FBF8E10EBD578EAAFF8415482BED1555EF55555057D145152428492E800820",
INIT_2E => X"FB6DF574A85575C55EFBE8E1557D1475FAF45BEAA800AAFFAA9557D080038AAA",
INIT_2F => X"00AAAEA8A9200249056D4175C50920875FDA381C209256DFFDF420BA552A821F",
INIT_30 => X"0BA55557DFF700000000000000000000000000000000000000000000008517DE",
INIT_31 => X"AA105D5155410FF84020AA0800154B2AAAA975FF5D7BC21EFF7FBD7400F7FBC0",
INIT_32 => X"400A25551554BA0051400BA5551575EFF7D1401FF5D5568BE7555568A00AAFFE",
INIT_33 => X"FFDFFF552EA8AAA55043DFF7AAAEAAB55F78400145AAFFFFFEF5D7FEABFF0051",
INIT_34 => X"55400BA082E8201000043FE005D517DEBA0851574B2FFAABFF45FFAAAABFFAAF",
INIT_35 => X"7AA955EF00002AAA2A2FBE8A00A2D16AAAAFF8002410FFD5575EF5555421E755",
INIT_36 => X"FFFFC00BA552A821EFFFFFD74BA5D51575F7FFAE975EF555168B55F7AA800BAF",
INIT_37 => X"000000000000557DE00AAAAAAA000804001FF0055554088A557FEB25D00021FF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000C00000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(5),        -- Port A data input
DOA(0)   => data_read_a_hi(5),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(5),        -- Port B data input
DOB(0)   => data_read_b_hi(5),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_6_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10800B0061A01002840002C03002818000402322520070B313301C4389B2082",
INIT_01 => X"274008482009404C18A160000C52424841000000090800090210000008510200",
INIT_02 => X"102430600C800110000006100009D070012408000000000648080000001210E0",
INIT_03 => X"000200501D1D02140C420200480140040608010040400104681A0084490C4802",
INIT_04 => X"404402820021000A00824002141000980500000808001114C000080624600600",
INIT_05 => X"120024204209981001A806500304610528000500000080000000300000012940",
INIT_06 => X"2000440832280002300010209C4400142061207A024008900008000220600220",
INIT_07 => X"130C8A220FF41F00902008808800182001020150000001F0800408264000100A",
INIT_08 => X"001BF002C4A01041B1120101000010128568837F04842B080020890008080342",
INIT_09 => X"011847140126805432A62A1596C8B5DF10000008900000100220C00084000008",
INIT_0A => X"44EB4104D09392053589F11C59898888454010830212C54081000410A0088C00",
INIT_0B => X"B0044245B25B456C0096C0096C4096C4096C2096C2096C6096C444B6004B600C",
INIT_0C => X"09040020280010000B3002820110101D0012402CC00802410C26800860070621",
INIT_0D => X"0500819D0000900208201040C4007920004884080000448C281018100C000200",
INIT_0E => X"05008182100000000000000000022AE800C00004000000050081A00004000000",
INIT_0F => X"0002330006000000080000000000000D07A00020000000050081A00020000000",
INIT_10 => X"0000000001204A340002100000000000000000020F4001400000020000000000",
INIT_11 => X"019300020000000068D08000200000001A692121000280000000000010000000",
INIT_12 => X"000201FA100400000000034696010000000000D3478000000000000001003F00",
INIT_13 => X"00000000000000043C0001C0A000008000000000012E000054AC000020000000",
INIT_14 => X"0200000040A410C2810800016000809400001000000000000000433300007600",
INIT_15 => X"060180400000008060180404002AC0200208940041309210B28048180F028000",
INIT_16 => X"2008000100601802000000100601800000000180600800000020180600000000",
INIT_17 => X"0180600000008040100200800000060100000802010040180200002018040100",
INIT_18 => X"7F8FF0F4FA955F7CF7F40A80907638C31C71C718638E00006018040080200004",
INIT_19 => X"38E38E38E38E38E38E38E38E38E38E38E38E38E39B6CEDECDDF7DF7DF5F78BCE",
INIT_1A => X"3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE38E38E38E38E",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFF000000000000196A03F9FCFE7F3F9FCFE7F3F9FCFE7F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"00000000000000000000000C0FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"BFDF45F7AA974AAAAAA97555F784174BAF7D5555FF0000000000000000000000",
INIT_22 => X"FBD7410AA8428AAAAAAE955450055421FFFFFBC0010AAD5574BA557FFDFFF087",
INIT_23 => X"FFBEAA10007FD7410FFAA97400082A800AA08515555508043FE00F7AA97555A2",
INIT_24 => X"55517FF55A2AA97400552AAAB45082E80155F7D1575EFFFAA9555500557FE10F",
INIT_25 => X"FF7AAA8A10082EAAB45A2FFC2000007FD74000055574BA5D7FD7555A2D5575EF",
INIT_26 => X"FFAA843DF55FFAA955EFA2D168B55557BEAB5500554200000003DE10FFD5401F",
INIT_27 => X"BFF00002AABA5D2ABFFFF087BD5545007BFDE10AA803FE105D516AABAFF843FF",
INIT_28 => X"0000000000000000000000000000000000000000AAAEBDF45A28428B45FFD168",
INIT_29 => X"524AA5571FDFEF1C7BFFF55FFA095482B6A49256DEB84104BAFFD1525FF00000",
INIT_2A => X"03DE28F7A49057DAAF5D2428A2842AAAAA2AE9756D145B401FFFFFFC7010BEDF",
INIT_2B => X"A49756D145178E00EBFBE8A101475D5400F7A4904380824850381C5B5057D1C0",
INIT_2C => X"571D757DB6D5525EF555178F6DAAA495428412AAFB451C2A8017DE3DF525FFFF",
INIT_2D => X"1C0E3FE00E3DB471EFE3AAAAA00082EA8B6DA2F1C50381471D74380851524BA5",
INIT_2E => X"049516AAB8FF8428FEFA28E3AF55F7A0925D7AADB6FB7D5D7FEAB7D0855420BA",
INIT_2F => X"45B68A28B6DEBDF6DBEF1C0A28AAA5524BFFFF1C7BD057D1C71FFE10A28038E1",
INIT_30 => X"0AAFFD1401E7000000000000000000000000000000000000000000000B6AEBDF",
INIT_31 => X"21EFF7FBD7400F7FBC00BA55557DFF7557BFDF55F78017400F780001FFAA8400",
INIT_32 => X"154B2557FC01EF55043FEAAFF80021EFA2D1420BAAA8428AA2AAAA975FF5D7BC",
INIT_33 => X"A821EFAAFBC01FFF780155F7555568A00AAFFEAA105D5155410FF84020AA0800",
INIT_34 => X"51554BA0051400BA5551575EFF7D1401FF5D5568BE7AA80174AA082ABDF555D2",
INIT_35 => X"D7FEABFF0051400A25D2EBFE10AAFFD55EFA2AEA8A10082EA8BEFAAD5554B255",
INIT_36 => X"55557DE00AA842AA0000516AABAFF8428BE7AAAEAAB55F78400145AAFFFFFEF5",
INIT_37 => X"0000000000FFAABFF45FFAAAABFFAAFFFDFFF552EA8AAA55043DFF7557BC01EF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000900000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(6),        -- Port A data input
DOA(0)   => data_read_a_hi(6),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(6),        -- Port B data input
DOB(0)   => data_read_b_hi(6),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_7_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10844B00482258A2842112C02450418800002300500030B313300C418992002",
INIT_01 => X"234008422008604D1C20E0000E11426840000000080000080200090000110204",
INIT_02 => X"1025207000B08910000206101188D03080144880010400044808000000122160",
INIT_03 => X"000200401914821004420000CA01000C0600010000605114291A008449484802",
INIT_04 => X"40440200002100080006500210101019040000000B085024D842080244000000",
INIT_05 => X"1A8024200009981001A8224001040104200204000000800CC2092CE4A0004900",
INIT_06 => X"A000440822280002340010209C040014A061200052500810000C490323208E28",
INIT_07 => X"128802020028000890240980A809102001020140000009F0800408264000100A",
INIT_08 => X"001A0602C4A01051B13281010408881203480200448423199046821008082351",
INIT_09 => X"336784144126811054809C1040140A001C8648481000045903318B80A400310A",
INIT_0A => X"000800009010100014114110312388984502148282A08415B032095048008100",
INIT_0B => X"20CDC1C483484D201192011920119201192051920519205192074C9018C90188",
INIT_0C => X"D8A5B44001D2C12901228F82F005310D293054048A2212004466000DA1908528",
INIT_0D => X"800F8108A0D09802082010408580008000000008C85264010816851B428DA146",
INIT_0E => X"800F81321000020000261900E28A204040E000A0000007800F814000A0000007",
INIT_0F => X"7072024807000020400000581C01C1A406400084000007800F81400084000007",
INIT_10 => X"060180E83800E820101210000200000CC3003C32080201C0000C000000160700",
INIT_11 => X"81DD00804086423120B74020023090644840A34000828800000004000420020B",
INIT_12 => X"1C6A0186E8000446120C8905BA0004810C84624237E00010001878007F0030C0",
INIT_13 => X"00080208E4083C44230201AEE0010040261900E30520C0806EAC0082000984C0",
INIT_14 => X"0121011088A600C032128201519480D40005802448160403E0700622C0806EE8",
INIT_15 => X"A1685A1685A168DA368DA36CDA30DA13A108810111349A943AA4401000928A19",
INIT_16 => X"368DA768DA1685A1685A5685A368DA368DA7685A1685A1685A768DA368DA368D",
INIT_17 => X"685A1685A169DA368DA1685A1695A368DA3685A1685A168DA368DA1685A1685A",
INIT_18 => X"00000000000000000000400A8448410400020820800069DA1685A168DA369DA3",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000003667B000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"0155EFAAAEA8ABAAAFBFDE0055556AA005D04155550000000000000000000000",
INIT_22 => X"556AA00FFAE95555087BFDF45F7AA974AAAAAA97555F784174BAF7D5555FFF78",
INIT_23 => X"055421FFFFFBC0010AAD5574BA557FFDFFF5555555EFAAFFFDFEFAAAAAAB455D",
INIT_24 => X"AA8428AAA557BFDFFF55003DFFFF7FBEAA00002EAAAAA082EA8A00AAAE955450",
INIT_25 => X"0552EBDE00007BEAAAAA2D14000008515555508043FE00F7AA97555A2FBD7410",
INIT_26 => X"FF00557FE10FFFBEAA10007FD7410FFAA97400082A800AAF7AE975FFA2800001",
INIT_27 => X"155F7D1575EFFFAA955555D51574AAAAFFD5545087FEAB455D516AB55557BD55",
INIT_28 => X"0000000000000000000000000000000000000000A2AA97400552AAAB45082E80",
INIT_29 => X"104BAFFD1525FFFF8E175C7A2AAAAA82A2F1FAE105D556AA10410E1755500000",
INIT_2A => X"1FFFD7AAAAAFB7D495F6AA10E3AE905551C7BFFF55FFA095482B6A49256DEB84",
INIT_2B => X"2EAAA00A2AE9756D145B401FFFFFFC7010BEDF524AA5571FDFEF415B575D7AAF",
INIT_2C => X"7A49057DAAF5D2428A2842AAAA497BFAFFF49003AFEFEBFBEAA001C2EA8A821C",
INIT_2D => X"F7A4905C7A28A070384120BDE100075EAA82BEDB470101C5B5057D1C003DE28F",
INIT_2E => X"D555F6AB57417BC05D7145178E00EBFBE8A101475D5400F7A490438082485038",
INIT_2F => X"28412AAFB451C2A8017DE3DF525FFFFA49756D495150492BEF1D2555087BE8B7",
INIT_30 => X"A10002E9754D000000000000000000000000000000000000000000000AAA4954",
INIT_31 => X"7400F780001FFAA84000AAFFD1401E7FFAA97555A2AEA8A10AAD568A00555168",
INIT_32 => X"7DFF7007BD5555AAD57DF55AAAEBDFEF007BE8A10AAAE8215D557BFDF55F7801",
INIT_33 => X"FEAA105D2EAAA005D2AAAA18AAAA975FF5D7BC21EFF7FBD7400F7FBC00BA5555",
INIT_34 => X"7FC01EF55043FEAAFF80021EFA2D1420BAAA8428AA2007FE8BFF080028BFFAAF",
INIT_35 => X"F84020AA0800154B2FF8402145A2AA954AA00043DE0000516AA10F7FBD740855",
INIT_36 => X"FFD140145007FE8BEF557BEAB55087FC215D555568A00AAFFEAA105D5155410F",
INIT_37 => X"0000000000AA80174AA082ABDF555D2A821EFAAFBC01FFF780155F7005140000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000000FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(7),        -- Port A data input
DOA(0)   => data_read_a_hi(7),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(7),        -- Port B data input
DOB(0)   => data_read_b_hi(7),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_8_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00000648E2840112C00000418000002700500030B3132000400812086",
INIT_01 => X"214009C21838284D042100000212026840000000180800080200080040510204",
INIT_02 => X"1021004000900110000006100088503000240800014400004808000000122160",
INIT_03 => X"0002004019110214044A82000121400C86000000000000860188008448400002",
INIT_04 => X"000402800031200A0000090214100889A5000000490090104800000224000400",
INIT_05 => X"10C025204289981000A820500344010428008500010080080909304040202004",
INIT_06 => X"8000440003280000340010208C04003420600000C6180810000C490703200010",
INIT_07 => X"130002000028000890240980A809012001020050000009F08004082640000082",
INIT_08 => X"20100402C4201041310041010008801201480200051023090024811008090A1A",
INIT_09 => X"0100001001248100308214528148A48008000008100004590711C04034000083",
INIT_0A => X"10804000801210140001C0103001088845010482004000008420041020008900",
INIT_0B => X"0004404002004400448000480004800048000480004800048000440022400200",
INIT_0C => X"880420000880204909004502D100A10C04205424010216010C26800805000004",
INIT_0D => X"8000801100509802082010400400018000488428800004082014000200010000",
INIT_0E => X"8000800A00000207A8BE7B00000200082040808000F07F80008000808000F07F",
INIT_0F => X"0002000402100000404CB1F8FC0000040000808000F07F80008000808000F07F",
INIT_10 => X"3E07800000004004080A000002072C3FCF0000020040804800040007687E3F00",
INIT_11 => X"10800018639EC00020100002C2F9B0000801016001008100000040120CB3067F",
INIT_12 => X"000200020000585EB6000100800030C73D8000402000001FC07FF80001000080",
INIT_13 => X"002EAE1FEC0000040200408000003C547E7B00000100801004000803551F8FC0",
INIT_14 => X"00000000440610C8000A808040000208901B86E568FE0C000000020080100400",
INIT_15 => X"0040100401004090240902449028D0230249850101349A98BAC0481000888810",
INIT_16 => X"0401004010040100401004010240902409024090240902409004010040100401",
INIT_17 => X"4010040100409024090240902409004010040100401004090240902409024090",
INIT_18 => X"543EBC57A10A1E75D6440A889050000000000000000040902409024010040100",
INIT_19 => X"79E79E79E79E79E79E79E79E79E79E79E79E79E7BF3CCD8DF5B2DB2CA4028A0A",
INIT_1A => X"4F87D3E1F4F87D3E1F4F87D3E1F4F87C3E1F0F87C3E1F0F87C3E79E79E79E79E",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000000D3E94F87D3E1F4F87D3E1F4F87D3E1F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"000000087BEAA10F7803DE00FFAEBFFFF0800155FF0000000000000000000000",
INIT_22 => X"7FC2145005155555F780155EFAAAEA8ABAAAFBFDE0055556AA005D0415555080",
INIT_23 => X"7AA974AAAAAA97555F784174BAF7D5555FF552AA8AAA557FC0010F780154105D",
INIT_24 => X"FFAE95555AAFFE8A00552EBFE00F7D17FF45F7FFFFF55AA80155FF087BFDF45F",
INIT_25 => X"5F7D140010552E821EFAAAABDF555555555EFAAFFFDFEFAAAAAAB455D556AA00",
INIT_26 => X"00AAAE955450055421FFFFFBC0010AAD5574BA557FFDFFF5504000AAAAAAA8B5",
INIT_27 => X"A00002EAAAAA082EA8A00002AA8A10F78402155AA8028A00A2D57FF45557BE8A",
INIT_28 => X"0000000000000000000000000000000000000000557BFDFFF55003DFFFF7FBEA",
INIT_29 => X"6AA10410E17555080E000280071E8A00EB8E3FE10F7AEBAFFF080A175D700000",
INIT_2A => X"1C2000FF8A17400557FC015514555757DFF8E175C7A2AAAAA82A2F1FAE105D55",
INIT_2B => X"8A105D71C7BFFF55FFA095482B6A49256DEB84104BAFFD1525FF492EA8AAA557",
INIT_2C => X"AAAAFB7D495F6AA10E3AE90555A2FBE8A38492ABDE10EBDF7AF6DE3FFF8F7DB6",
INIT_2D => X"550E00082B6A0AFB55F7D1420104124821D7AAA0BDF6D415B575D7AAF1FFFD7A",
INIT_2E => X"0B6D578F6D557FFDA00A2AE9756D145B401FFFFFFC7010BEDF524AA5571FDFEF",
INIT_2F => X"FF49003AFEFEBFBEAA001C2EA8A821C2EAAA001C2EA8A00F7800017DA2842FA0",
INIT_30 => X"BEF082E95545000000000000000000000000000000000000000000000497BFAF",
INIT_31 => X"8A10AAD568A00555168A10002E9754D082E820BA08556AA00AAAABFE00F7AEAA",
INIT_32 => X"401E7082EAAABA5D5140010F7AE974105D7BC21555D51575EFFFAA97555A2AEA",
INIT_33 => X"BEABFFAAFBEABFFF7AA80145557BFDF55F78017400F780001FFAA84000AAFFD1",
INIT_34 => X"7BD5555AAD57DF55AAAEBDFEF007BE8A10AAAE8215DA2FFE8ABA082ABFE00AAF",
INIT_35 => X"7FBC00BA55557DFF75D2E82010F7843DF45FFD540000000402145AA843FFFF00",
INIT_36 => X"F780021FFA2803DE10FFD16ABFF5D7BFDE10AAAA975FF5D7BC21EFF7FBD7400F",
INIT_37 => X"0000000000007FE8BFF080028BFFAAFFEAA105D2EAAA005D2AAAA185D2AAAA10",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000400000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(8),        -- Port A data input
DOA(0)   => data_read_a_hi(8),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(8),        -- Port B data input
DOB(0)   => data_read_b_hi(8),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_9_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000B0001800002840002C0000281800000030000000033022000000000002",
INIT_01 => X"8000098218302849180060000C004240413C0A61590001D90213C90008510200",
INIT_02 => X"000008700CB089100002061031200074810448800104008048080080001210E2",
INIT_03 => X"000200140C1822000A028010408100000628000140402080041A100040024840",
INIT_04 => X"41040000000400080002040200080800040000000B08D1055842080604600700",
INIT_05 => X"10002024000020102400010000026104200004000400800C8B0024E4E0010C40",
INIT_06 => X"8000440802280002700800008A840004A0610000C0000810000C590103600810",
INIT_07 => X"538600220028001890240980A80800200102025000000BF08200002440000883",
INIT_08 => X"00000402C220104131102101040810028528820005100003900E884000010007",
INIT_09 => X"00000005E000000600BCA284140200800C834948100004590111824404012080",
INIT_0A => X"04080000901012100A1141005922000245410002008880000032005080000800",
INIT_0B => X"2000020040044010440104401004010440100401044010040104400802008208",
INIT_0C => X"D1A1344420D2E100000808000000000481000000202002400006800825908402",
INIT_0D => X"0500000000109000000000000580008000080000C852240100068D0B4685A342",
INIT_0E => X"0500000A00000000000000000000028000408020000000050000208020000000",
INIT_0F => X"0000304002100020000000000000000900208004000000050000208004000000",
INIT_10 => X"0000000001200000000A00000000000000000000050000480008000000000000",
INIT_11 => X"009F0080000000004807C0200000000012000020000081000000040000000000",
INIT_12 => X"00000048F8000400000002403E0004000000009067E000000000000000000900",
INIT_13 => X"0000000000000000140000CEE001000000000000000A000036AC008000000000",
INIT_14 => X"03210000000400CA81000000619480D4000400000000000000004100000036E8",
INIT_15 => X"A368DA368DA3685A1685A1685A121A11A1419001512490040024001000008019",
INIT_16 => X"1685A1685A1685A1685A1685A368DA368DA368DA368DA368DA368DA368DA368D",
INIT_17 => X"685A1685A168DA368DA368DA368DA368DA368DA368DA3685A1685A1685A1685A",
INIT_18 => X"CCF48DE68A895C38E250080000000000000000000000685A1685A1685A1685A1",
INIT_19 => X"514514514514514514514514514D34D34D34D34D28E10040392482090157344C",
INIT_1A => X"4D268341A0D069349A0D069349A0D068341A0D068341A0D06834514514514514",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000001654D0D069349A0D068341A4D268341A",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"BE8B45002A974AAAA803DFFFAA843DF45FFFFEAABA0000000000000000000000",
INIT_22 => X"AEBDE00AAFBEAABA080000000087BEAA10F7803DE00FFAEBFFFF0800155FFAAF",
INIT_23 => X"AAEA8ABAAAFBFDE0055556AA005D0415555087BFDE00A2FBD7400F7FBFDFFFA2",
INIT_24 => X"005155555557BE8BEF007FFDEAAAAD1555EF0055401FFF7AEAAA10F780155EFA",
INIT_25 => X"0F7AA974AA082E80010A2AAAAA10552AA8AAA557FC0010F780154105D7FC2145",
INIT_26 => X"BA087BFDF45F7AA974AAAAAA97555F784174BAF7D5555FFF780154AA5D2AA8A1",
INIT_27 => X"F45F7FFFFF55AA80155FF080400145FFFBEAABAF7D17FEBAA2AEBDF45002EAAA",
INIT_28 => X"0000000000000000000000000000000000000000AAFFE8A00552EBFE00F7D17F",
INIT_29 => X"BAFFF080A175D7BEF1E8B6D002090482B68E38FC7BE8A3DF7DF7F5E8A9200000",
INIT_2A => X"BD0400FFF5FDFC7B6A0BDE38B6F5E8A92080E000280071E8A00EB8E3FE10F7AE",
INIT_2B => X"AAA8A38FF8E175C7A2AAAAA82A2F1FAE105D556AA10410E175550871FFE00A2F",
INIT_2C => X"F8A17400557FC015514555757D5D71E8BEF147BFAE82A2DB555C71C5B451D7FF",
INIT_2D => X"FF84174BA5D20AAA00E3AA904BA142A87010A2AEADA38492EA8AAA5571C2000F",
INIT_2E => X"AAAA0BFF7D0024ADA921C7BFFF55FFA095482B6A49256DEB84104BAFFD1525FF",
INIT_2F => X"38492ABDE10EBDF7AF6DE3FFF8F7DB68A105D7000400155FFFBEDA82FFD57DEB",
INIT_30 => X"FEFF7D16AA00000000000000000000000000000000000000000000000A2FBE8A",
INIT_31 => X"AA00AAAABFE00F7AEAABEF082E95545F7D568BEF080402000F7AAA8B55FFAABD",
INIT_32 => X"9754D00517DE00A2FFC2000F7D17FF55FF803FEAAFFD16AA00082E820BA08556",
INIT_33 => X"FD55555D7FD5555FFAAA8AAAFFAA97555A2AEA8A10AAD568A00555168A10002E",
INIT_34 => X"2EAAABA5D5140010F7AE974105D7BC21555D51575EF555568BEF5D7FE8A10AAF",
INIT_35 => X"A84000AAFFD1401E7FF80174AA5D0028A00AAAE800AA552A97400A2AEBDEAA08",
INIT_36 => X"F7FBFFE00FFD17FEAAA2803DFEF08043FE00557BFDF55F78017400F780001FFA",
INIT_37 => X"0000000000A2FFE8ABA082ABFE00AAFBEABFFAAFBEABFFF7AA80145080002145",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000800000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(9),        -- Port A data input
DOA(0)   => data_read_a_hi(9),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(9),        -- Port B data input
DOB(0)   => data_read_b_hi(9),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_10_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000B0001800002840002C0000281800020030000000033022000000180006",
INIT_01 => X"000008000000004C002000000010026840000000080000080200000000110200",
INIT_02 => X"0000004000800110000006100000003000040800010400004808000000120060",
INIT_03 => X"000200000810020000020000400100000600000000400000001A000040004800",
INIT_04 => X"0004000000000008000200020000000004000000080010004000000200000000",
INIT_05 => X"1000202000011010000000000000010520000400000080000000200000200004",
INIT_06 => X"80004408022800023000000088040004A061000040000810000C490103600000",
INIT_07 => X"120420020028000890240980A808002001020050000009F08000002440000082",
INIT_08 => X"00000402C0201051311001000000020201080200440400000000800000000000",
INIT_09 => X"0000105808000000000000000000008000008088100004590111800004000000",
INIT_0A => X"00804000801210440003C1411008800045000002000014000040009002800000",
INIT_0B => X"0400200000000000000004000040000000000000040000400000000000000221",
INIT_0C => X"0100802000000000000002802000000400100000000002000026000840011400",
INIT_0D => X"0500000000409002082010400400008000400008002044082000081004080204",
INIT_0E => X"0500000200000000000000000000028000400000000000050000200000000000",
INIT_0F => X"0000304002000000000000000000000900200000000000050000200000000000",
INIT_10 => X"0000000001200000000200000000000000000000050000400000000000000000",
INIT_11 => X"0082000000000000480080000000000012000101000080000000000000000000",
INIT_12 => X"0000004810000000000002400400000000000090400000000000000000000940",
INIT_13 => X"0000000000000000150000C00000000000000000000A40001400000000000000",
INIT_14 => X"02000000002400C2810000006000000000000000000000000000410040001400",
INIT_15 => X"020080200802008020080200800800220200840001309A08A848001000008000",
INIT_16 => X"0000000000000000000000000200802008020080200802008020080200802008",
INIT_17 => X"0080200802000000000000000000000000000000000000000000000000000000",
INIT_18 => X"940FE0D397124355520542821010000000000000000000802008020080200802",
INIT_19 => X"28A28A28A28A28A28A28A28A28A28A28A28A28A29554199854514514F546890A",
INIT_1A => X"32994CA6532995CAE572B94CA6532994CA6532994CA6532994CA28A28A28A28A",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000001867172B94CA6532994CA6572B95CAE5",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FC2155F7D155545AA80001EFAAFBEAB45557FFDE100000000000000000000000",
INIT_22 => X"FBE8BFFF78402155AAFBE8B45002A974AAAA803DFFFAA843DF45FFFFEAABA007",
INIT_23 => X"87BEAA10F7803DE00FFAEBFFFF0800155FF00042AB55FFD168B55AA8000010FF",
INIT_24 => X"AAFBEAABAA2FFD741055003DFEFF7AA801FFAAD16AABA002ABDE100800000000",
INIT_25 => X"FF7FBC0145F78028A00A2D142155087BFDE00A2FBD7400F7FBFDFFFA2AEBDE00",
INIT_26 => X"BAF780155EFAAAEA8ABAAAFBFDE0055556AA005D0415555007FD74105555555E",
INIT_27 => X"5EF0055401FFF7AEAAA105D042ABFF5D556AB55AAD168ABA002A975FFF7AEBDE",
INIT_28 => X"0000000000000000000000000000000000000000557BE8BEF007FFDEAAAAD155",
INIT_29 => X"3DF7DF7F5E8A92007BC217DEBDB55555AA8E071D7AAFBEFB455D71F8E0000000",
INIT_2A => X"B6DB55BE8E05000EBFFE8BC7E38E07145BEF1E8B6D002090482B68E38FC7BE8A",
INIT_2B => X"2EB8E00080E000280071E8A00EB8E3FE10F7AEBAFFF080A175D700042AB7DEBD",
INIT_2C => X"FF5FDFC7B6A0BDE38B6F5E8A92B6FBD5410490A3DFD7F7A4821D7A2D16FA8214",
INIT_2D => X"0071D54104951555D7EBF5C5155E3842AA00BED1421450871FFE00A2FBD0400F",
INIT_2E => X"20820955EFE3AEBDEAAFF8E175C7A2AAAAA82A2F1FAE105D556AA10410E17555",
INIT_2F => X"EF147BFAE82A2DB555C71C5B451D7FFAAA8A38410E2ABD749516FB55BED16FA8",
INIT_30 => X"F455D556AA000000000000000000000000000000000000000000000005D71E8B",
INIT_31 => X"2000F7AAA8B55FFAABDFEFF7D16AA00087FC01EFA2FFD7545AAAE97555A2FBFD",
INIT_32 => X"9554500042ABFFA2FFFFF45F7AE97400AAFFE8B45AAAA95545F7D568BEF08040",
INIT_33 => X"400155A2D57FE00552EA8A00082E820BA08556AA00AAAABFE00F7AEAABEF082E",
INIT_34 => X"517DE00A2FFC2000F7D17FF55FF803FEAAFFD16AA00FFFBD5400082EBFF45F78",
INIT_35 => X"55168A10002E9754D085155410085557555AAD557555A2802AA10FFD54214500",
INIT_36 => X"08557DF55F7D17FE000804155FFAAAABDEAAFFAA97555A2AEA8A10AAD568A005",
INIT_37 => X"0000000000555568BEF5D7FE8A10AAFFD55555D7FD5555FFAAA8AAA002AAAB45",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000008FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(10),        -- Port A data input
DOA(0)   => data_read_a_hi(10),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(10),        -- Port B data input
DOB(0)   => data_read_b_hi(10),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_11_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10180B05A0010402840602C2D001019000000300000000330A20080EC180002",
INIT_01 => X"AB400986B830284D1820E0000C3642484000000008000008820009080A512220",
INIT_02 => X"102A68440080011000000618062AD03502640800010410424908136019920868",
INIT_03 => X"004A0846191B22120642000442C110044600000101E9225CDC9A10844A9A4842",
INIT_04 => X"0094024000250808800216021138000B848000000800100040000102A0600200",
INIT_05 => X"7E4024242008A8102CA88A44010401042200444000888000000028000002A002",
INIT_06 => X"8088445712280000B18812288E0400253855200045C86810000C5B0503286A28",
INIT_07 => X"10008822A028004880200A80880208200122006C000015F0C20408264902C840",
INIT_08 => X"9390040280241041D1754100000018108728820024002B3A01A89540080824C8",
INIT_09 => X"A1001C41A1348498B080801010000080D00301081000045B0511D28D94012339",
INIT_0A => X"44080000901012428003414158230CBA4576708241C010908040341322008000",
INIT_0B => X"040464D280144050C72A0872A0C72A0872A0C72A0C72A0872A0C595043950421",
INIT_0C => X"0804001400000820110A42822204880CD81040442900021704E6000800001D54",
INIT_0D => X"80C62D0500409002082010404580018000404012004004192C10000000000000",
INIT_0E => X"80C62D5803161C526DB40506C120A806ABB0D808CC334A80A54B70D408CC32D2",
INIT_0F => X"2B5144D0DD903C54916D15458C0513005570D408CC334A80A54B70D808CC32D2",
INIT_10 => X"52148C4DB05621E363F813961C20EDA944016558C2347A080B10D8DD6422AA10",
INIT_11 => X"1880144D3345C65593800319C18BD1ECA1C9010112566F10AC4183C340DAE02D",
INIT_12 => X"5810503000633830DE3C2C9C00289A66AA8DE50E0800360614AC281430890600",
INIT_13 => X"0CD2A9CEA8199B6B082B55900314140365320485C4F00AD544407241C175C402",
INIT_14 => X"0000074044C4801832701A89D20A38093631425969020855A281844E00540404",
INIT_15 => X"0000000000000000000000000020C00200088101513492101280401000400200",
INIT_16 => X"2008020080200802008020080000000000000000000000000000000000000000",
INIT_17 => X"0080200802008020080200802008020080200802008020080200802008020080",
INIT_18 => X"804180C0B10A4210420140028400000000000000000000802008020080200802",
INIT_19 => X"000000000000000000000000000820820820820801C414947000000055062608",
INIT_1A => X"0000000004020000000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000001F87E000000000000010080000000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"ABDF5508557DF45002ABDFFFF7803DE10AA80000AA0000000000000000000000",
INIT_22 => X"FFE8A10A28000000007FC2155F7D155545AA80001EFAAFBEAB45557FFDE10082",
INIT_23 => X"02A974AAAA803DFFFAA843DF45FFFFEAABAA2AEBFF45FFAEBFEAA002A801FFF7",
INIT_24 => X"F78402155AAD155555A28428BFF002ABDE00A2AABFE10082ABFFEFAAFBE8B450",
INIT_25 => X"0002A80010A2842AAAA007BFFF4500042AB55FFD168B55AA8000010FFFBE8BFF",
INIT_26 => X"00080000000087BEAA10F7803DE00FFAEBFFFF0800155FF00557FF45557FC201",
INIT_27 => X"1FFAAD16AABA002ABDE10A2D168A10A284021FF5D00154BAF7FBE8BEFFFD5400",
INIT_28 => X"0000000000000000000000000000000000000000A2FFD741055003DFEFF7AA80",
INIT_29 => X"EFB455D71F8E00002EBDF6D005B78F7D142ABDFC7F78E3FE28B684070AA00000",
INIT_2A => X"0BDEAA1C2A801C7E3FFEFA10B68407038007BC217DEBDB55555AA8E071D7AAFB",
INIT_2B => X"20B8FEFBEF1E8B6D002090482B68E38FC7BE8A3DF7DF7F5E8A92BEAEBFF7DEBA",
INIT_2C => X"E8E05000EBFFE8BC7E38E07145B6D15756DA28A28BFF082ABAE10B6AAB8E2808",
INIT_2D => X"08517DF7D497BC5028142A87000A28A2AA92007FF8F7D00042AB7DEBDB6DB55B",
INIT_2E => X"2FFFFEFBC7E3DF42028080E000280071E8A00EB8E3FE10F7AEBAFFF080A175D7",
INIT_2F => X"10490A3DFD7F7A4821D7A2D16FA82142EB8E00B6DB6AA28A280001FF5D0A1048",
INIT_30 => X"EAAF784154BA000000000000000000000000000000000000000000000B6FBD54",
INIT_31 => X"7545AAAE97555A2FBFDF455D556AA00082EBFFEF007BE8BFF5D2ABDF55F7AABD",
INIT_32 => X"6AA00FFAEBFFEFAA803DEBA5D2E82155A2FBFDE00FF84154BA087FC01EFA2FFD",
INIT_33 => X"AAAA00FFAAA8AAA080028BFFF7D568BEF080402000F7AAA8B55FFAABDFEFF7D1",
INIT_34 => X"042ABFFA2FFFFF45F7AE97400AAFFE8B45AAAA95545F7D5555FFAAAAA8BFF002",
INIT_35 => X"7AEAABEF082E9554508557DFFF007BD54BA5D2E95400A2AEA8A00007FEABFF00",
INIT_36 => X"AA80001FF5D2E82000F7FFFFF45AAFFC20BA082E820BA08556AA00AAAABFE00F",
INIT_37 => X"0000000000FFFBD5400082EBFF45F78400155A2D57FE00552EA8A00FFFFE8AAA",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000800000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(11),        -- Port A data input
DOA(0)   => data_read_a_hi(11),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(11),        -- Port B data input
DOB(0)   => data_read_b_hi(11),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_12_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"A500C4B01BC0268A6940312C0DE045196A831A300500032B333287E4FC812006",
INIT_01 => X"AF400D869830E84D5823E0000C1742484000000008000008820009280A553235",
INIT_02 => X"502A7144008001100000171C022BD13412762A000586235ECC09C8423B960866",
INIT_03 => X"31863846191BA218064204000281200406A10843010022DEDF0852944A9C014A",
INIT_04 => X"0014030000250409000014821038080B840000400800102040000302F0600233",
INIT_05 => X"7FC034348008A8102CA88F48010601042400048000188000000938000002E088",
INIT_06 => X"9CC96CC6F63A5001F12B56A0AC8601F47AC06400D1F80C10020C493F03343A38",
INIT_07 => X"1020002030280098A12048908A16BA311177124C000003F08A94282E5C262861",
INIT_08 => X"827A0602902A10491165E10000049010C52882008600A73A01E8974008092CF8",
INIT_09 => X"47000001A1248008F000000000000080000F010C100204593F11A6CDF48023BF",
INIT_0A => X"040000208010120ACA01400058010CBA4D277C86CCE802B380003C1360008000",
INIT_0B => X"011C46D3C7BC1EF083AF0C3AF083AF083AF0C3AF083AF083AF0C1D7861D78400",
INIT_0C => X"08040014C9001AE91D17E50AD79FEFC87C2154745F82131FFCCE00080000095E",
INIT_0D => X"807BF7118180984004000803D40001880001001400C005031010000000000000",
INIT_0E => X"807BF76A109C944B5891BF06C5EEB14FCBF0D90076D61C807BF7D0D80876D49C",
INIT_0F => X"6DE38EB9FB10350C00A99F7CA80757365E50D80876D61C807BF7D0D90076D49C",
INIT_10 => X"841BCC69A0D8C6F7F0AA001C943A65756A0976EB5A7E7FC8951018186334F311",
INIT_11 => X"D5A014481991C6A737D80211912970CDCDD1864116D6C7080651CB4661F33615",
INIT_12 => X"349E929300423224AE19B9BEC0289033238D4E6EA805892946A9B011A7B152CF",
INIT_13 => X"6244CD7AC01CAAA56B3E6D9001068715D64006D2A961CF9B44512A2504532182",
INIT_14 => X"00000439FDC25C58067A9FAB46095A0B5289A0282D2E1444ACB12A17CF9B4414",
INIT_15 => X"0000000000000000000000040026C00000288401513492909280401000F70A00",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"088881360A95090CB05442029010000000000000000000000000000000000000",
INIT_19 => X"1041041041041041041041041049249249249249200100002D4514510051B946",
INIT_1A => X"592C964B2592C964B2592C964B2592C86432190C86432190C864104104104104",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000002007F592C964B2592C964B2592C964B2",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"43FE0008557DFFF0800020105D557FEAA00557DE100000000000000000000000",
INIT_22 => X"557DFFFF7AA80000082ABDF5508557DF45002ABDFFFF7803DE10AA80000AAAA8",
INIT_23 => X"7D155545AA80001EFAAFBEAB45557FFDE10AAD5420000051555FFA2AA8200000",
INIT_24 => X"A28000000A2D155410F7FFFFEBA08003FE00082AA8AAAAAFFC00BA007FC2155F",
INIT_25 => X"0A2AABFE1055516ABEF5D517DEAAA2AEBFF45FFAEBFEAA002A801FFF7FFE8A10",
INIT_26 => X"55AAFBE8B45002A974AAAA803DFFFAA843DF45FFFFEAABA000028A105D2ABFE1",
INIT_27 => X"E00A2AABFE10082ABFFEF085542000000417555002A820AA08557DFFFF7AA821",
INIT_28 => X"0000000000000000000000000000000000000000AAD155555A28428BFF002ABD",
INIT_29 => X"3FE28B684070AABE803AE38145B78FD7000005010495B7AE921C517DE1000000",
INIT_2A => X"B505FFB6A487000005F7AFD7F7A482038002EBDF6D005B78F7D142ABDFC7F78E",
INIT_2B => X"F5C2082007BC217DEBDB55555AA8E071D7AAFBEFB455D71F8E00BED547038145",
INIT_2C => X"C2A801C7E3FFEFA10B68407038B6D550428FFF1FDE821C003FE001C2EAAAAAB6",
INIT_2D => X"00002FA285D20BDE28A2A4B8E10555B68BEF5D517DEAABEAEBFF7DEBA0BDEAA1",
INIT_2E => X"2005F7DFD7F7A482155BEF1E8B6D002090482B68E38FC7BE8A3DF7DF7F5E8A92",
INIT_2F => X"6DA28A28BFF082ABAE10B6AAB8E280820B8FEF085F4703814001055514208208",
INIT_30 => X"A0055517DE00000000000000000000000000000000000000000000000B6D1575",
INIT_31 => X"8BFF5D2ABDF55F7AABDEAAF784154BAF7802AABA5D7FEAB45080015410007FEA",
INIT_32 => X"6AA00F7D1554BA5D7BC01FFFF8015410007FEAB45F780020BA082EBFFEF007BE",
INIT_33 => X"43FE10552EAAAAAFFD140000087FC01EFA2FFD7545AAAE97555A2FBFDF455D55",
INIT_34 => X"AEBFFEFAA803DEBA5D2E82155A2FBFDE00FF84154BAF7D1400BAFFD57FE005D0",
INIT_35 => X"FAABDFEFF7D16AA0008003FEBA55003DEBAA28428A105D7FEABEF55557DEBAFF",
INIT_36 => X"550402145550000010087FFFF45F78402145F7D568BEF080402000F7AAA8B55F",
INIT_37 => X"0000000000F7D5555FFAAAAA8BFF002AAAA00FFAAA8AAA080028BFF087BD54AA",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000000FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(12),        -- Port A data input
DOA(0)   => data_read_a_hi(12),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(12),        -- Port B data input
DOB(0)   => data_read_b_hi(12),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_13_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10110A0441812402840402822007818000E00700000000330A3000000008042",
INIT_01 => X"A1400984B830C848180260000C0042604001000008220008A200100802110200",
INIT_02 => X"10A00860009141100000C6180C285035000E0800010431004908135980120C60",
INIT_03 => X"004E20441910221B06420C85D5013804060000000040324C441A108468024842",
INIT_04 => X"0184034010250089C00EA8021938325B04800002091090014880080200000900",
INIT_05 => X"18002424B008881024A8004E01040104270004E0000080090500604840000481",
INIT_06 => X"80004414022A2490B00A142C8C840005794540015E006810001C4B01032C7E20",
INIT_07 => X"510200028028004880280A808816002101022468000011F082040A264006C000",
INIT_08 => X"D2B00402B220104B531001000008001041080200B660E30B200C8040080A9206",
INIT_09 => X"A1000809A93484D21000000000000080C90391881000145B0111A30404015000",
INIT_0A => X"000000008010102A82014100101118BA4510008241480290882400900000A000",
INIT_0B => X"0284484000000000400000000040000000000000040000000000000020000000",
INIT_0C => X"A944AA2000A02000212800020000000D80004084A0000390002E001843210400",
INIT_0D => X"859C1881A04090000000000021800180010341179065441356150A1285094284",
INIT_0E => X"859C188810C65A72A617520252781EA02520D589B9A260859C1840DD81B9A0E0",
INIT_0F => X"0E71F1052D942748C19484E39442D15961C0DD81B9A260859C1840D589B9A0E0",
INIT_10 => X"E60605C0C12CBD400B0810C65A61AA459D0047398500D5889D26907356533C00",
INIT_11 => X"8F60CA1562094650CA28398A42C051E0332181010109294C8E1160CB8C80A561",
INIT_12 => X"2645056D073148580A3C065141942AC4128CA199180C5232575138094450AD0A",
INIT_13 => X"84CA93A2FC008962142B17301A9A1A5196A80245208E0AC5C853C8028163B8C0",
INIT_14 => X"0240034000E4DC8A84000014982372011FC1E475F0F0084A3961F5A80AC5C816",
INIT_15 => X"4250942509425094250942509428D421420882020120981812C8403000088212",
INIT_16 => X"2509425094250942509425094250942509425094250942509425094250942509",
INIT_17 => X"5094250942509425094250942509425094250942509425094250942509425094",
INIT_18 => X"FF3F7DF7FF3E9F7DF7E24502A800000000000000000050942509425094250942",
INIT_19 => X"EBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBF7DFDFDDD555555F7EFBBEE",
INIT_1A => X"7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAEBAEBAEBAEBA",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000000007F7EBF5FAFD7EBF5FAFD7EBF5FAFD",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5554BA087FFFF55557BD54AAF7FBC01FFA2802ABEF0000000000000000000000",
INIT_22 => X"2E80155AA802AB45AA843FE0008557DFFF0800020105D557FEAA00557DE10AAD",
INIT_23 => X"8557DF45002ABDFFFF7803DE10AA80000AA087BD75EF087FFFFEF557BEAB4555",
INIT_24 => X"F7AA80000AAD1420AA087BD7555FFD168AAAFFAE820AA5D5557555082ABDF550",
INIT_25 => X"5FFD157555085140010F7AEAABFFAAD5420000051555FFA2AA8200000557DFFF",
INIT_26 => X"45007FC2155F7D155545AA80001EFAAFBEAB45557FFDE10AAAEA8BFFA2FBD754",
INIT_27 => X"E00082AA8AAAAAFFC00BA00002AAAAF7D5574BA557BE8A10A284154BAFFAAAAB",
INIT_28 => X"0000000000000000000000000000000000000000A2D155410F7FFFFEBA08003F",
INIT_29 => X"7AE921C517DE10A2DB50482147FFAF554971D0492E3F1C71C7BE8A2ABD700000",
INIT_2A => X"FFAFD7497BE8B5555208217DBE8A2AB45BE803AE38145B78FD7000005010495B",
INIT_2B => X"5F5056D002EBDF6D005B78F7D142ABDFC7F78E3FE28B684070AA1C71D25D7007",
INIT_2C => X"6A487000005F7AFD7F7A482038AADF47092147FD257DFFD568A82FFA4870BA55",
INIT_2D => X"A2A0ADBC7A2FFD257DE3DF52555085142000FFAAAFBFFBED547038145B505FFB",
INIT_2E => X"0B680124BAFFAAAFB45007BC217DEBDB55555AA8E071D7AAFBEFB455D71F8E00",
INIT_2F => X"28FFF1FDE821C003FE001C2EAAAAAB6F5C20821C002AA92FFDF574824171EAA1",
INIT_30 => X"545F7AEA8B55000000000000000000000000000000000000000000000B6D5504",
INIT_31 => X"AB45080015410007FEAA0055517DE00A2FFC00105D7BE8B55085142010AAD157",
INIT_32 => X"154BA5D5140145007BE8B55087BEAB555D04001EFF7AAA8B55F7802AABA5D7FE",
INIT_33 => X"16AA10FF80174AA557FC21EF082EBFFEF007BE8BFF5D2ABDF55F7AABDEAAF784",
INIT_34 => X"D1554BA5D7BC01FFFF8015410007FEAB45F780020BAA2FFD54105D7FC21EFFFD",
INIT_35 => X"2FBFDF455D556AA00A2803FF45AAFFC21EFAAFBC0155085540000FFAEBFFEFF7",
INIT_36 => X"F7FBD5410085568A10FF80020AAFFAABFF55087FC01EFA2FFD7545AAAE97555A",
INIT_37 => X"0000000000F7D1400BAFFD57FE005D043FE10552EAAAAAFFD1400005D042AA00",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000CFFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(13),        -- Port A data input
DOA(0)   => data_read_a_hi(13),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(13),        -- Port B data input
DOB(0)   => data_read_b_hi(13),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_14_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10020A000180000284008280000281800000030000000033022000000580002",
INIT_01 => X"A140098018300848184860000C20C24040000000084000084200000000110200",
INIT_02 => X"1020006000900110000006102028503400040800010400204908012018120E64",
INIT_03 => X"000200441910221006420000400100040600000000E9E401209A108448004842",
INIT_04 => X"0004020000250008000200021038000804000000090090004800080200000000",
INIT_05 => X"500024240008881024A800400104010420000400000080080100204040000000",
INIT_06 => X"8000440102282015B10A10288E0400042345400040006810000C5901033D7880",
INIT_07 => X"1100000200280048802008828812002001220064000005F1C2850A2649204070",
INIT_08 => X"00B00402802010411110010000080010010802000400230B000C804008080002",
INIT_09 => X"01000009A92480001000000000000080C8038188100004590111B68404010000",
INIT_0A => X"0000000080101000000141001001088A45000082400000008020009000008000",
INIT_0B => X"0004404000000000400004000000000000004000000000000004000000000000",
INIT_0C => X"8904A0200080200001080002000000088000400420000200002E000841010400",
INIT_0D => X"0500000C80409000000000000000018000000000806044010014081204090204",
INIT_0E => X"0500005813A0210D072E8D012001028402908004000587050000108004000707",
INIT_0F => X"9004300044900812386A280E5800088980108020000587050000108020000707",
INIT_10 => X"DE00482E19E30002007813A02096038AE200880405200308828062A68C0BC700",
INIT_11 => X"00000E5A08E6000048001292B83280001208A1011004011060049A1C59192055",
INIT_12 => X"492060480256530650000240001DB011CC00009000032C4C979E3806180C0900",
INIT_13 => X"5A3433EDE00154181400000007BCBD858F120120541A0000000033757465B2C0",
INIT_14 => X"02002C000024008A84001A0902000422E3E99681004802115652594000000001",
INIT_15 => X"0240902409024090240902409028D021020880000120901812C8401000000210",
INIT_16 => X"2409024090240902409024090240902409024090240902409024090240902409",
INIT_17 => X"4090240902409024090240902409024090240902409024090240902409024090",
INIT_18 => X"5C8FF0F7BE9D5F7DF65040028000000000000000000040902409024090240902",
INIT_19 => X"79E79E79E79E79E79E79E79E79E79E79E79E79E7BF7DDDDDFCF3CF3DF5579B4E",
INIT_1A => X"3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE79E79E79E79E",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000003FF803F9FCFE7F3F9FCFE7F3F9FCFE7F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"BE8B55A2AE80000F7D5555555D2AAAABAAAD1420BA0000000000000000000000",
INIT_22 => X"00155EF0804155EFAAD5554BA087FFFF55557BD54AAF7FBC01FFA2802ABEFA2F",
INIT_23 => X"8557DFFF0800020105D557FEAA00557DE10A2AA801FFA28402000AAAE9554555",
INIT_24 => X"AA802AB4500516AA00A2AE800BAFFFFC20BAF7AEA8B45080417400AA843FE000",
INIT_25 => X"0A2843FEBAFFFBD7410A2D168BFF087BD75EF087FFFFEF557BEAB45552E80155",
INIT_26 => X"AA082ABDF5508557DF45002ABDFFFF7803DE10AA80000AA005568ABAA2840201",
INIT_27 => X"AAAFFAE820AA5D5557555002E80155A280000005D7FFDF4555517DFEF00043FE",
INIT_28 => X"0000000000000000000000000000000000000000AAD1420AA087BD7555FFD168",
INIT_29 => X"C71C7BE8A2ABD7A2FFEDB55B6A080038E3DB50555412AA8ABAAADB4009200000",
INIT_2A => X"402038AAAA955554900105FF0800175D7A2DB50482147FFAF554971D0492E3F1",
INIT_2B => X"0A12410BE803AE38145B78FD7000005010495B7AE921C517DE10A2AE851FFB68",
INIT_2C => X"97BE8B5555208217DBE8A2AB451C556FA00A2A0800BAE3F1C0092EBAAADB6D08",
INIT_2D => X"00516DABAA28402038B6803DE82F7F5D5410A2D568BC71C71D25D7007FFAFD74",
INIT_2E => X"55D5F78FD7000E3FEAA002EBDF6D005B78F7D142ABDFC7F78E3FE28B684070AA",
INIT_2F => X"92147FD257DFFD568A82FFA4870BA555F5056D002A80155B680000105D7FF8F4",
INIT_30 => X"AAAAAFFC2000000000000000000000000000000000000000000000000AADF470",
INIT_31 => X"8B55085142010AAD157545F7AEA8B55A2FBFFF55FF84000AAAAFBC0145002AA8",
INIT_32 => X"7DE00A2AA955FFFF80020BAAAAA975450800001EF080417555A2FFC00105D7BE",
INIT_33 => X"140000A2AEBFFEF082A82010F7802AABA5D7FEAB45080015410007FEAA005551",
INIT_34 => X"5140145007BE8B55087BEAB555D04001EFF7AAA8B555D557FE00A280020BAAAD",
INIT_35 => X"7AABDEAAF784154BA08557FEAAA284000AAFF803DE00FFD557400AAD56AB455D",
INIT_36 => X"F780020105D7BEAB45557BE8B45082EBFEBA082EBFFEF007BE8BFF5D2ABDF55F",
INIT_37 => X"0000000000A2FFD54105D7FC21EFFFD16AA10FF80174AA557FC21EF082A80145",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000000FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(14),        -- Port A data input
DOA(0)   => data_read_a_hi(14),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(14),        -- Port B data input
DOB(0)   => data_read_b_hi(14),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_15_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000A000000000284000280000001800020030000000033022000000180002",
INIT_01 => X"A140098018300848180060000C00424040000000080000080200000000110200",
INIT_02 => X"102100400C8011100000061000A8503401044880010430004808000180122378",
INIT_03 => X"000200541D102210064200000045000546080000400020000008108448400042",
INIT_04 => X"8094020000254C880000028A1018000844000000880013504000002600000000",
INIT_05 => X"10002424000AA81024A82040010C61062001440002988000000024808001004B",
INIT_06 => X"80004400022A00003C8912248E0400042854400040006810000C4901032B1800",
INIT_07 => X"50200000B0280048A0280A828801002101020040000005F38204082640000000",
INIT_08 => X"01F00402802610411100110000000010010802000400230A0008884008080004",
INIT_09 => X"01000001A12481041000000000000080C0030108100004590111820404000000",
INIT_0A => X"0000000080101000004140001001088A45000082000000008000001080008000",
INIT_0B => X"0004404000000000400004000040000400000000000000000004000020000200",
INIT_0C => X"0804000020024100012808020000000981004004A0200310000C000800000000",
INIT_0D => X"0000001180009000000000002100018000000000004004010010000000000000",
INIT_0E => X"00000008000002000000000000000000000080A40000000000000080A4000000",
INIT_0F => X"00000000001000204800000000000000000080A40000000000000080A4000000",
INIT_10 => X"000000000000000000080000020000000000000000000008000C020000000000",
INIT_11 => X"000000824000000000000020220000000001800100020300000004003420480A",
INIT_12 => X"0000000000040440000000000001048000000000000000100800400000000000",
INIT_13 => X"000800000000000000000000000100C220050000000000000000008220884400",
INIT_14 => X"000000000000000830000000000000000016101C5C1400000000000000000000",
INIT_15 => X"0000000000000000000000000020C00000088000012090101280401000000200",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000040028000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"000010082A954BA00003DFEF085155400F78428BEF0000000000000000000000",
INIT_22 => X"8015400FF84001EFA2FBE8B55A2AE80000F7D5555555D2AAAABAAAD1420BAFF8",
INIT_23 => X"87FFFF55557BD54AAF7FBC01FFA2802ABEFF7AE95555A2FBE8BEFA2843DE00AA",
INIT_24 => X"0804155EFFFFBE8BFF0800174AA557BFDE10A2FBEAB45F7D56AABAAAD5554BA0",
INIT_25 => X"5FFD568BEF087FE8A1055003FE00A2AA801FFA28402000AAAE955455500155EF",
INIT_26 => X"45AA843FE0008557DFFF0800020105D557FEAA00557DE10F7D1574AAA2D16AB5",
INIT_27 => X"0BAF7AEA8B45080417400FFFFC2145080015400AA802AA00AAAE800BA5D00155",
INIT_28 => X"000000000000000000000000000000000000000000516AA00A2AE800BAFFFFC2",
INIT_29 => X"A8ABAAADB40092E38E070280024904AA1C0438FD7005150438F78A2DBFF00000",
INIT_2A => X"FE8BC7BE8E38E10A28017400E38A051FFA2FFEDB55B6A080038E3DB50555412A",
INIT_2B => X"D16AABAA2DB50482147FFAF554971D0492E3F1C71C7BE8A2ABD7E3AA9257DA2F",
INIT_2C => X"AAA955554900105FF0800175D7E3FFEFBD70000124AA557FFDE10A2FBEDB6DF7",
INIT_2D => X"FFDF50482A2DB6AB45FFD56DBD7087BEAA38410038E38A2AE851FFB68402038A",
INIT_2E => X"0AAA085082550A1057DBE803AE38145B78FD7000005010495B7AE921C517DE10",
INIT_2F => X"00A2A0800BAE3F1C0092EBAAADB6D080A12410FFF1C017D140410400BE8E28A1",
INIT_30 => X"0AAF7AEBDFEF0000000000000000000000000000000000000000000001C556FA",
INIT_31 => X"00AAAAFBC0145002AA8AAAAAFFC2000AAAA974AA0800020BA550028B55085540",
INIT_32 => X"A8B55AAAE821EFAAFBEAB55F7AAA8A00AA8417400AAAE975EFA2FBFFF55FF840",
INIT_33 => X"BFFE10A2FFFFFEFF7D568ABAA2FFC00105D7BE8B55085142010AAD157545F7AE",
INIT_34 => X"AA955FFFF80020BAAAAA975450800001EF080417555AAFFFDF450804020AA557",
INIT_35 => X"07FEAA0055517DE00FFFBC2000AAFBE8B55F7D17DF45007FE8AAA08002AAAAA2",
INIT_36 => X"5D0000010F7AAA8A10AA8017400552A801EFF7802AABA5D7FEAB450800154100",
INIT_37 => X"00000000005D557FE00A280020BAAAD140000A2AEBFFEF082A82010FFD5421EF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000C00000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(15),        -- Port A data input
DOA(0)   => data_read_a_hi(15),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(15),        -- Port B data input
DOB(0)   => data_read_b_hi(15),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_16_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"DA22C618B1000482B688B186588884862A400438255FC38381441205BA803003",
INIT_01 => X"264AC80028404C211203A952A90341080B173340412000E1005D628000820484",
INIT_02 => X"400034C206C405000001A48202084004003008255040826EE008B440200E2042",
INIT_03 => X"A459C1240181AB20AD27315B7F1983CA1C900040422A005762010010000C0400",
INIT_04 => X"296E542B6E3A825C15FB385321B4ADFE16AB45FD2C400002E205231201290A28",
INIT_05 => X"B9E5815006028179808C00A0D2152B90707A1E0BD423CAC0000D610000000710",
INIT_06 => X"81F104A1415C292164280081C6AB88742086ACACDE240000A80090CE82A803B9",
INIT_07 => X"400800000ACCAA280940580400A37B8896CA4D000A80C1102A00001C14028009",
INIT_08 => X"0015452880C8D90409A02D965965200100104F2B00822512000000231520A024",
INIT_09 => X"A5AA80018120E00066000000000012C9000A0000D0A80000BF8028E87C1B9927",
INIT_0A => X"00520228080108039501200848002912300208092B940192D1000000000000A8",
INIT_0B => X"03561180063DB4F6110001100011000110001100011000110001080008800080",
INIT_0C => X"080200854409418B02ED0000502A02972000040BB401100010012B4C90000100",
INIT_0D => X"6D061A1F8D60D80820500101244AA8A2AA242E80000009200120000000000000",
INIT_0E => X"6D066210E5001DB4A5B400C7D553847165A99000C6564CDD051DC99000C65555",
INIT_0F => X"21D0C48F254946148107354292673D1F72C99000C6564CDD0565C99000C65555",
INIT_10 => X"952D2058F33225787810F5001D6121A9559224D1FF97D0272F04D89441A56D8A",
INIT_11 => X"6C1C74485B81E31306C71D1093AB8A64811BADC00992180D58033B1172F2A025",
INIT_12 => X"7B86DED8E3A212748F0E0CA638E890B7A8546120C0AFF5B548AC431FB1C7DB07",
INIT_13 => X"EFCE9B26DECA1AD36A2E4F40DF6AAAF260AF88899E8B8B93D12A877178DD0032",
INIT_14 => X"A8009F8B108C80A1021B9A8BB8056662CA1951596800FC01A38D4D4B072B922F",
INIT_15 => X"00000000000000000000000000044000102A0001148442A1108103595580A840",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"4C690DA64C1C4F68A36040000000000000000000000000000000000000000000",
INIT_19 => X"D14D14D14D14D14D14D14D14D14514514514514529E5F87869E79E78558D1154",
INIT_1A => X"3D1E8F47A7D3E9F4FA7D3E9F4FA7D3E9F47A7D1E9F47A7D1E9F4D14D14D14D14",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE000000000000000007D3E9F4FA7D3E8F47A3D1E8F47A",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFEFF7D168B55AAD17FFFF552EBFE00007FC00AA0000000000000000000000",
INIT_22 => X"04000BA552A821FFFF8000010082A954BA00003DFEF085155400F78428BEF087",
INIT_23 => X"2AE80000F7D5555555D2AAAABAAAD1420BA5D2E975EFF7D568BFFFF80175EF00",
INIT_24 => X"FF84001EF0000020AA5D00154005D043FF45555540000082EAABFFA2FBE8B55A",
INIT_25 => X"0087FD74BAAAAEBFFEF557FC00AAF7AE95555A2FBE8BEFA2843DE00AA8015400",
INIT_26 => X"FFAAD5554BA087FFFF55557BD54AAF7FBC01FFA2802ABEF557BEABEF5D041541",
INIT_27 => X"E10A2FBEAB45F7D56AABA082A97545F7D16ABFFFFAABFEAAFF84001FF002A821",
INIT_28 => X"0000000000000000000000000000000000000000FFFBE8BFF0800174AA557BFD",
INIT_29 => X"50438F78A2DBFF0871F8FC7E3D56AB6DBEDB7FFEF552AB8E38087FC209200000",
INIT_2A => X"16ABFFE38E175EF1400000BA412E871FFE38E070280024904AA1C0438FD70051",
INIT_2B => X"2EAFBD7A2FFEDB55B6A080038E3DB50555412AA8ABAAADB400924920925EFF7D",
INIT_2C => X"E8E38E10A28017400E38A051FF0804050BA410A1240055003FF6D5551420101C",
INIT_2D => X"4975EDBC7550E12410087FD74AAB6AABFFC7557FC00BAE3AA9257DA2FFE8BC7B",
INIT_2E => X"AF780051C70824851D7A2DB50482147FFAF554971D0492E3F1C71C7BE8A2ABD7",
INIT_2F => X"D70000124AA557FFDE10A2FBEDB6DF7D16AABA08249756DF7D168BC7F7AABAEA",
INIT_30 => X"AAA007BC0000000000000000000000000000000000000000000000000E3FFEFB",
INIT_31 => X"20BA550028B550855400AAF7AEBDFEF08516AB55A2D16ABEFFFFBFDFFF552AAA",
INIT_32 => X"C20000000021EFF7D568BFFA2AA955FF5D04020AA002A955EFAAAA974AA08000",
INIT_33 => X"03DFEF5D51420005D2ABFF45A2FBFFF55FF84000AAAAFBC0145002AA8AAAAAFF",
INIT_34 => X"AE821EFAAFBEAB55F7AAA8A00AA8417400AAAE975EF0800174BA002E820105D0",
INIT_35 => X"AD157545F7AEA8B5500557DF45552A82000007BD74AAF7AEBDF455D7BC20BAAA",
INIT_36 => X"F7D568B55FFAAAAABAFF8415545000015555A2FFC00105D7BE8B55085142010A",
INIT_37 => X"0000000000AAFFFDF450804020AA557BFFE10A2FFFFFEFF7D568ABA0804155FF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000400000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(16),        -- Port A data input
DOA(0)   => data_read_a_hi(16),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(16),        -- Port B data input
DOB(0)   => data_read_b_hi(16),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_17_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"5284CE4FB7BD2C8994A13392DBD02E14006B82AC7E800D44D3DD2FD5F9B961C0",
INIT_01 => X"F9BA301F7E03FC6793F2199B39FC233C11D93AE6F3BB92B32091DBC339B24542",
INIT_02 => X"1D5FC0C08F040404446965C0607FB8A217C400C33A908078551BD04222186338",
INIT_03 => X"8504930A37F65820CB24111B7F08014A0AB84A52B6D2AFF97C1B5AC757F06D6B",
INIT_04 => X"250834336D1E81500FDB38302292ADFE103B6DBD204037F202042075E2B1D00A",
INIT_05 => X"8F039786062C6CE092F5FE005236781C402A0807B4070670083DC68206D7E6D0",
INIT_06 => X"0CD26803C3582408962C58B183F8AEF42045919B30E085DD2ED57D4EED08CA6A",
INIT_07 => X"700000B30380670B8142500448E3E01E94EF1340A28AC1AC8156044D1400AA00",
INIT_08 => X"009F3A1B0120A1C51DFFC40C30E5F0182D0950190C0810BE00E9A76E4C6FFBE4",
INIT_09 => X"8FCCC200A59BDD2FFE3F3EC7C7DEF207000F00059D2ED56D7EED2ED3C9A867DC",
INIT_0A => X"0617112E46F05D02DD814102F800633F1D0A7CC9AE7A08BFF0001D35682AC0CE",
INIT_0B => X"8A3F06ABD73DBCF4FBCF4FBCF4FBCF4FBCF4FBCF4FBCF4FBCF4FBE7A7DE7A780",
INIT_0C => X"001000974F08518F5AFFC94B533FADA7FDE97D6BFF329E1B50FF99F086000D9E",
INIT_0D => X"F50B018F95EA3DED1652EC0B27E67F419E2E1E8000C0036340B8000000000000",
INIT_0E => X"F50B01C8DF7F96197DB4AFC8C8886AF672A1537F759299F50B03C1537F759199",
INIT_0F => X"6068331C5103E7EF0FBEED6BB6A9412007C1537F759299F50B03C1537F759199",
INIT_10 => X"21F2CD7F252CDABB3CE8CF7F963AB9FD6AD434201AA68B837FFD1F7B7125B68C",
INIT_11 => X"BD055EB6D555CB2949C15BA7270FF256526BBFD55BBE71D79F73C7AC6DB9BF37",
INIT_12 => X"94080BF82B74E4E1FE4ACA4E0ABD6DAAAB965293036FF6B652A99A6026027FBE",
INIT_13 => X"EF5CBA7A43482800FEFAFD06B8CFCCAB7550D0C2022EAEBD438697AD2EBA9168",
INIT_14 => X"AC00A8BBFC8B501CF7A0FED9A548FA19752C4A4EADAE42FCBC38C3B7BEBF42CF",
INIT_15 => X"0000000000000000000000000026E100002F382DBD9ECFE117805F20CFDAAB00",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"09EDCC4052E917114F981800C000000000000000000000000000000000000000",
INIT_19 => X"EBA69AEBA69A69AEBA69AEBA69A69A69A69A69A68698686981D75D7443720030",
INIT_1A => X"46A351A8D068341A0D068341A0D068341A0D46A341A0D46A341A69AEBA69A69A",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000000000046A351A8D46A351A8D46A351A8D",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFEFF7FBEAB450804001EFAAD57FEAA0000000000000000000000",
INIT_22 => X"51401EF087FD74AA087FFFFEFF7D168B55AAD17FFFF552EBFE00007FC00AA087",
INIT_23 => X"82A954BA00003DFEF085155400F78428BEFAAD168A000004020AA5D7BE8B4500",
INIT_24 => X"552A821FF5D00020BA552A82000552A821555D7FEAB55FF80175EFFF80000100",
INIT_25 => X"FAAFBC01EF5D0015555557BFDEBA5D2E975EFF7D568BFFFF80175EF0004000BA",
INIT_26 => X"BAA2FBE8B55A2AE80000F7D5555555D2AAAABAAAD1420BAFFFFFDF45AAD17FFF",
INIT_27 => X"F45555540000082EAABFF00516AA10552E820BA007FEABEF005555555A2D1554",
INIT_28 => X"00000000000000000000000000000000000000000000020AA5D00154005D043F",
INIT_29 => X"B8E38087FC2092147FFFFFFFFFBFDFC7EBF5E8B550000071EFB6DF7AE9200000",
INIT_2A => X"A07082497FEFB6D1451471EF007BD04920871F8FC7E3D56AB6DBEDB7FFEF552A",
INIT_2B => X"8E175FFE38E070280024904AA1C0438FD7005150438F78A2DBFFBED16AA381C0",
INIT_2C => X"38E175EF1400000BA412E871FF550A00092492A850105D2A80155417BEFB6DEB",
INIT_2D => X"FFF5FFF6DAADF7FFD7B6F1C71EF55001756D5D7BFAEBA4920925EFF7D16ABFFE",
INIT_2E => X"700515556DA2DF50492A2FFEDB55B6A080038E3DB50555412AA8ABAAADB40092",
INIT_2F => X"BA410A1240055003FF6D5551420101C2EAFBD7145B6AA28492487082007FEDBD",
INIT_30 => X"5EFFFFBEAA000000000000000000000000000000000000000000000000804050",
INIT_31 => X"ABEFFFFBFDFFF552AAAAAA007BC0000557FFDFEFF7FBFFF55A2D16AB55000017",
INIT_32 => X"BDFEFF7D568AAA5D2A97410007BFFFFF5551555EF087FC200008516AB55A2D16",
INIT_33 => X"A82155087FFFFEFAAAA975EFAAAA974AA0800020BA550028B550855400AAF7AE",
INIT_34 => X"00021EFF7D568BFFA2AA955FF5D04020AA002A955EF5D2E80010002A954005D2",
INIT_35 => X"02AA8AAAAAFFC2000FFD57DFFFAAFFFDF55FFD1575FF5504175EF5D7FEAAAA00",
INIT_36 => X"000415410007BFFF450051555EFA2FBC0000A2FBFFF55FF84000AAAAFBC01450",
INIT_37 => X"00000000000800174BA002E820105D003DFEF5D51420005D2ABFF45557FE8AAA",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000CFFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(17),        -- Port A data input
DOA(0)   => data_read_a_hi(17),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(17),        -- Port B data input
DOB(0)   => data_read_b_hi(17),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_18_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"69844019080000A21A611406840014122A641074155FC28A2024001001801003",
INIT_01 => X"01067920034004180005E9E3C90360C0041C0181002001602025800008440084",
INIT_02 => X"40AC3CAA22D605200000856E2481902400344A20F802C22054001000021E2379",
INIT_03 => X"A54C23B34C81EB2076471000800981140C010101750D1007E58040102B0E0100",
INIT_04 => X"22660C1C0065003C04040013236E105016A028402D618803EB092B9201490B2A",
INIT_05 => X"B8E080000000005889AC41E04508A99070200E010001C1CA11803850C8000100",
INIT_06 => X"800A4CE301545001F40050216C09950004C2047BCF1C8090C02800C0120886B3",
INIT_07 => X"814A0080064C1F300020080182001A9E02C03400082002700000217294007101",
INIT_08 => X"000117088080990419002D86184A01018030430700802541420440022030041A",
INIT_09 => X"7030C30B885200D274004008080003C32A10A19090C02010E102294406168800",
INIT_0A => X"00602A01880980037109700C04C44C92A88DCC2211E44174112840880000060D",
INIT_0B => X"11C0D95C20C2030A003080030800308003080030800308003080018400184004",
INIT_0C => X"8304E02809832E6021002020404042000F00008400811824AD4007ECD9436261",
INIT_0D => X"0AFCE5D22A82B20000520100C801F8A07E103000A1285C84000418360C1B060D",
INIT_0E => X"0AFCFD8CB17E5B4F045557575E6EFBE3942C1040A41D660AFCE1CC1040A41E66",
INIT_0F => X"8E7FFBB385661C08D1455ABA91E6FF5FDFCC1040A41D660AFCF9CC1040A41E66",
INIT_10 => X"015F82C006C3AF31E64CB17E5A9655017F1FC73FAF1D61B1040294C58AD1FF5F",
INIT_11 => X"B95454005BAA36DCF8E519001BF80DEB3EE2020EA678189C6EC32881F7F75648",
INIT_12 => X"67D7EDFCA320037E81BD77D728A800B7546DBDFF12904747A351145FC53ABF8D",
INIT_13 => X"92B764225C57C97EBE76E1254F0C0D4514A84F5573FE9DBA4A38E247C522CC0E",
INIT_14 => X"BE84370001B6922070440556B15F7FABBC40151D7C747D8220673C3B9DB84B20",
INIT_15 => X"06C1B06C1B06C1B06C1B06C1B0491069068000004060300A005A01183F240014",
INIT_16 => X"6C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B",
INIT_17 => X"C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B0",
INIT_18 => X"B80EE173C2300F7DF16000000000000000000000000041B06C1B06C1B06C1B06",
INIT_19 => X"AAAAAA28A28A28AAAAAAA28A28A28A28A28A28A2910591505C104104B28BBECE",
INIT_1A => X"128944A25128944A25128944A25128944A2552A954AA5128944AAAA28A28A28A",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000128944A25128944A25128944A25",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFDFEF5D2A974BA082E954000000000000000000000000",
INIT_22 => X"0028B55002E82000087FFFFFFFFFFFFFEFF7FBEAB450804001EFAAD57FEAA087",
INIT_23 => X"7D168B55AAD17FFFF552EBFE00007FC00AA087FFFFFFFFFBFDF45AAD568B5508",
INIT_24 => X"087FD74AAAAFFFDF45A2D16AB55F7FFFFFFF00043DE10AA843DE00087FFFFEFF",
INIT_25 => X"A55042ABEF5D7FD75FFAAD540145AAD168A000004020AA5D7BE8B450051401EF",
INIT_26 => X"45FF8000010082A954BA00003DFEF085155400F78428BEFAA80000000804154B",
INIT_27 => X"1555D7FEAB55FF80175EF5D00020105D2A97400082E95555085168A10557FD75",
INIT_28 => X"00000000000000000000000000000000000000005D00020BA552A82000552A82",
INIT_29 => X"071EFB6DF7AE921C7FFFFFFFFFFFFFFFF7FBFDFFF5D2A954AA082A9242800000",
INIT_2A => X"1FAF55A2DF6DB7D1C002AB7D002A82028147FFFFFFFFFBFDFC7EBF5E8B550000",
INIT_2B => X"8E38E280871F8FC7E3D56AB6DBEDB7FFEF552AB8E38087FC2092087FFDFC7E3F",
INIT_2C => X"97FEFB6D1451471EF007BD0492B6F1F8F55AADF6DB7DE3F5FAFC708003DE28B6",
INIT_2D => X"A28407038140410492550A2ABC7497BD25FFAADF4516DBED16AA381C0A070824",
INIT_2E => X"D1C516FA28417BD5545E38E070280024904AA1C0438FD7005150438F78A2DBFF",
INIT_2F => X"92492A850105D2A80155417BEFB6DEB8E175FF5D0E05000492097428002E9557",
INIT_30 => X"4AA082A820AA000000000000000000000000000000000000000000000550A000",
INIT_31 => X"FF55A2D16AB550000175EFFFFBEAA00557FFFFFFFFFFFDFEFF7FBFFFEF552E97",
INIT_32 => X"C0000087BFDF45AAD568B55AAFBFDFEF55042ABEF002A800AA557FFDFEFF7FBF",
INIT_33 => X"16AB4500043DEAAFFAEAAAAA08516AB55A2D16ABEFFFFBFDFFF552AAAAAA007B",
INIT_34 => X"D568AAA5D2A97410007BFFFFF5551555EF087FC2000FFD56AB45A2FFFDFFFAAD",
INIT_35 => X"855400AAF7AEBDFEFA280154BA550400000552AA8B45087FC01EFA2FFD55EFF7",
INIT_36 => X"0804154BA082A975EF5D517DEAA007BD5545AAAA974AA0800020BA550028B550",
INIT_37 => X"00000000005D2E80010002A954005D2A82155087FFFFEFAAAA975EF5D2E97400",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000400000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(18),        -- Port A data input
DOA(0)   => data_read_a_hi(18),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(18),        -- Port B data input
DOB(0)   => data_read_b_hi(18),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_19_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"042200000000000041088001001AA00000000000000000000000500802000003",
INIT_01 => X"074018000024000000000404000000000A22000800000800004A200000000001",
INIT_02 => X"0000048002C405000000000006A84000000000200893C246A20000000020031A",
INIT_03 => X"082A58E411004B2000071000000981000C000000002045000200000000000000",
INIT_04 => X"200604000000001C0400001320000000162000002C4000026201201200090800",
INIT_05 => X"1020800000000058840200204000099070200E010001C0400000000000000000",
INIT_06 => X"0012048037805421402850001402498820022802400480405008901100A00102",
INIT_07 => X"00000000020C0130481204919200010C82000000000006002A548902A0020109",
INIT_08 => X"0001150800009900000005861840000000004301000B000000000001C1C00000",
INIT_09 => X"001F00002024B20002000000000002C300000000405000103010204000000000",
INIT_0A => X"00000000000000000000000000000040002000044000000000000000000002F0",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000420003B00000000000000000040012C80000000",
INIT_0D => X"45001A03C0825A0D20800000000018A006001000000000000000000000000000",
INIT_0E => X"450002131E01A1F6EA0A0020211146E069C2ACC01AE80045001D82ACC01AE800",
INIT_0F => X"1188340C3E1CFAD27CC2E004481020892282ACC01AE80045000582ACC01AE800",
INIT_10 => X"DEA03228D810007019931E01A1E5BA02802008C06F029D4C7B76639CEC0A0020",
INIT_11 => X"428AA3592000000206C2A4DAC00000008113C246A181C03FE4662A84575768DF",
INIT_12 => X"08201090549B5800000000261546B24000000000C53807E7CC06618018C51210",
INIT_13 => X"13F6A185A0A0168128411ACB800C0E108A0720288C011046B5986247C5452291",
INIT_14 => X"0000C220010808C10D9A92A74CD7CF4A080031B1515B212143D841431046B58A",
INIT_15 => X"00000000000000000000000000000000000000000000000000000118030004E0",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"3F0C7010C660C744192000000000000000000000000000000000000000000000",
INIT_19 => X"1861861861869A61861861861861861861861861A8208C4C1534D34C07208BBA",
INIT_1A => X"0984C26130984C26130984C26130984D26930984C26130984C261861861869A6",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE000000000000000000984C26130984C26130984C2613",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF552A974AA0004174BA0000000000000000000000",
INIT_22 => X"2E974BAA2FFFFE10087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974BA082E95400F7F",
INIT_23 => X"FFFFFFEFF7FBEAB450804001EFAAD57FEAAF7FFFFFFFFFFFFFFFFF7FBFDFFF55",
INIT_24 => X"002E82000F7FFFFFFFFFFFFDFEFA2D568B550004001EFAAAEA8ABA087FFFFFFF",
INIT_25 => X"5AAD16ABEF5D2ABFF55080402010087FFFFFFFFFBFDF45AAD568B55080028B55",
INIT_26 => X"BA087FFFFEFF7D168B55AAD17FFFF552EBFE00007FC00AAF7FFFFFFFF7FBE8B5",
INIT_27 => X"FFF00043DE10AA843DE00557FFDFEFA2D16AB55A2FFFDFEF5D2EBFE00AAFFFFE",
INIT_28 => X"0000000000000000000000000000000000000000AAFFFDF45A2D16AB55F7FFFF",
INIT_29 => X"954AA082A92428E3FFFFFFFFFFFFFFFFFFFFFFFEF552A974AA0000104AA00000",
INIT_2A => X"FFDFEFF7F5FAFC7492A974AAB6F5F8E101C7FFFFFFFFFFFFFFFF7FBFDFFF5D2A",
INIT_2B => X"A4A8AAA147FFFFFFFFFBFDFC7EBF5E8B550000071EFB6DF7AE92EBFFFFFFFFFF",
INIT_2C => X"2DF6DB7D1C002AB7D002A82028FFFFFFFEFF7F1F8FD7AAD16AB450000001FFBE",
INIT_2D => X"F7FBF8FC7E3F5EAB45B6DF6FBEF5D2AB8F7D000000010087FFDFC7E3F1FAF55A",
INIT_2E => X"7412ABFE28B6F5F8E820871F8FC7E3D56AB6DBEDB7FFEF552AB8E38087FC2092",
INIT_2F => X"55AADF6DB7DE3F5FAFC708003DE28B68E38E284971F8FC7AAD56DB6DBEF5F8FD",
INIT_30 => X"4AA0004000AA000000000000000000000000000000000000000000000B6F1F8F",
INIT_31 => X"DFEFF7FBFFFEF552E974AA082A820AAA2FFFFFFFFFFFFFFFFFFFFFDFEF552E95",
INIT_32 => X"EAA00A2FFFFFFFF7FBFDFFFFFD568B55002A954AAF7D568A00557FFFFFFFFFFF",
INIT_33 => X"56AB450004001EFFF842AAAA557FFDFEFF7FBFFF55A2D16AB550000175EFFFFB",
INIT_34 => X"7BFDF45AAD568B55AAFBFDFEF55042ABEF002A800AAF7FBFDFEFF7D56AB45AAD",
INIT_35 => X"52AAAAAA007BC0000FFFBE8B55AAD168B55F7FFFFFFF552AA8BEF08040200008",
INIT_36 => X"A2D57FFFFF7D568B45002ABDEAAFFD16AA0008516AB55A2D16ABEFFFFBFDFFF5",
INIT_37 => X"0000000000FFD56AB45A2FFFDFFFAAD16AB4500043DEAAFFAEAAAAA08556AB55",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000800000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(19),        -- Port A data input
DOA(0)   => data_read_a_hi(19),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(19),        -- Port B data input
DOB(0)   => data_read_b_hi(19),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_20_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000003",
INIT_01 => X"A65FF80000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000048002CC070000000000000000000000002FF86100200000000220002362",
INIT_03 => X"0000000000080F6000977060009B87A03C000000000000000000000000000000",
INIT_04 => X"3F2EFC040388137C3E20C477600142019E6000003CC0000A6601601A000B0000",
INIT_05 => X"102F91D10802ABFB80000021C8010FB0F0F43E1FE867DFC04400390210000220",
INIT_06 => X"90492261000080003400000010008000004203FE400580000000803000200006",
INIT_07 => X"401000004FFDFF28C4300C0010200100004000002AA001F00000000014000000",
INIT_08 => X"0801F5780259FB00000007BEFBC010002008FF7F00000000010018A81000041C",
INIT_09 => X"00000000020000000000000000000ADF00000020000000800000802830011023",
INIT_0A => X"0000000000000200020000000000000000000000000000000200200290000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"08120000B9090A700000200000004000000400000080002000407FED80000000",
INIT_0D => X"000079804000F00000000000C01FF8A7FE003000000004008100000000000000",
INIT_0E => X"0000798201000000100000000135386000401000010000000079801000010000",
INIT_0F => X"0185C300020004000010000000000252C7801000010000000079801000010000",
INIT_10 => X"00000010C1F30F300002010000080000000000CD8A0000400400000010000000",
INIT_11 => X"008040000000000292C0080000000000A5604000000284000818505200080000",
INIT_12 => X"0015E1B00100000000001496008000000000052B000048080000000000FC3600",
INIT_13 => X"80000000000002BA280000800830300000000000B8B400000401881010000000",
INIT_14 => X"00000000020020020001000040283024E6FB8604020080000383383B00000400",
INIT_15 => X"000000000000000000000004010201001003020200000000000127DBFF004000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"038200010089120104D204002000000000000000000000000000000000000000",
INIT_19 => X"B2CB2CB2CB2CB2CB2CB2CB2CB2C30C30C30C30C306982121A1E79E79A0700030",
INIT_1A => X"432190C86432190C86432190C86432190C86432190C86432190CB2CB2CB2CB2C",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000432190C86432190C86432190C86",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA0804020100000000000000000000000",
INIT_22 => X"2E954AA000400000F7FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0004174BAFFF",
INIT_23 => X"FFFFFFFFFFFFFDFEF5D2A974BA082E95400007FFFFFFFFFFFFFFFFFFFFFFEF55",
INIT_24 => X"A2FFFFE10FFFFFFFFFFFFFFFFFFFFFBFDFFF5D2E954BA007FC00BA087FFFFFFF",
INIT_25 => X"FF7FBFFF550800020BAAAD56AAAAF7FFFFFFFFFFFFFFFFF7FBFDFFF552E974BA",
INIT_26 => X"10087FFFFFFFFFFFFFEFF7FBEAB450804001EFAAD57FEAA007FFFFFFFFFFFFFE",
INIT_27 => X"B550004001EFAAAEA8ABA5D7FFFFFFFFFFFDFEFF7D56AB450000021EFA2D57DE",
INIT_28 => X"0000000000000000000000000000000000000000F7FFFFFFFFFFFFDFEFA2D568",
INIT_29 => X"974AA0000104AAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA08000500000000",
INIT_2A => X"FFFFFFFFFBFDFEF5D2E974AA000A07000E3FFFFFFFFFFFFFFFFFFFFFFFEF552A",
INIT_2B => X"71C50BA1C7FFFFFFFFFFFFFFFF7FBFDFFF5D2A954AA082A92428087FFFFFFFFF",
INIT_2C => X"7F5FAFC7492A974AAB6F5F8E10E3FFFFFFFFFFFFFFEFF7FBFFFFF552E974AA00",
INIT_2D => X"1C7FFFFFFFFFBFDFEFE3F5F8F450004050AABEDF6FABAEBFFFFFFFFFFFFDFEFF",
INIT_2E => X"50804021FFB6D57DE28147FFFFFFFFFBFDFC7EBF5E8B550000071EFB6DF7AE92",
INIT_2F => X"EFF7F1F8FD7AAD16AB450000001FFBEA4A8AAA497FFFFFFF7FBF8FC7EBD168B4",
INIT_30 => X"4AA080017410000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFDFEF552E954AA0004000AAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A95",
INIT_32 => X"820AA087FFFFFFFFFFFFFEFF7FBFDFFF5D2A974AA002E95410A2FFFFFFFFFFFF",
INIT_33 => X"FFDFEF5D2E954AA0051554BA557FFFFFFFFFFFDFEFF7FBFFFEF552E974AA082A",
INIT_34 => X"FFFFFFFF7FBFDFFFFFD568B55002A954AAF7D568A00AAFFFFFFFFFFBFDFEFFFF",
INIT_35 => X"000175EFFFFBEAA005D7FFFFEFF7FBFDFFFAAD16AB450804174AAFFFFFFEBAA2",
INIT_36 => X"F7FFEAB45A2D568B550804001EFF7D57DEBA557FFDFEFF7FBFFF55A2D16AB550",
INIT_37 => X"0000000000F7FBFDFEFF7D56AB45AAD56AB450004001EFFF842AAAA087BFDFEF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000000FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(20),        -- Port A data input
DOA(0)   => data_read_a_hi(20),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(20),        -- Port B data input
DOB(0)   => data_read_b_hi(20),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_21_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"4A302428B824900A128C090A5C1800261500213C005FE812D10420054085A202",
INIT_01 => X"081FFE3440B609703B0427F801A40B8115BC4F655300340288A40D30040E4DD8",
INIT_02 => X"04CA478082CC1740002019824E0203100640303FF8C0B31061096E21A1840814",
INIT_03 => X"8C329E9204020FE002577800405B87047D5042129D8D0248903200013290C800",
INIT_04 => X"3E7FFE02482553FC3C020277E128080A1E6000003CC0000A6601E03A8B0F0008",
INIT_05 => X"F43F8140000203FFC806C8A1C1048FF0F0E07E1F00F7FFC00024010000468310",
INIT_06 => X"08710C10015E083D01A24404786BE0014114C3FE4187A009A663A680100B3096",
INIT_07 => X"200800008FDFFF00290000100211019812E210488228000000900260026C6058",
INIT_08 => X"0EF1F5FA0041FF080AC707FEFBC110008420F7FF388B70A20389346FE8000580",
INIT_09 => X"917FC30010107688862A28C54518DBFF00020004C0A6044901112A0908AA0A30",
INIT_0A => X"006309044081A001B188300E20806520398C6021569249C4B3007127080806FF",
INIT_0B => X"904595123203040D9228D9228D9228D9228D9228D9228D9228D99146C9146C84",
INIT_0C => X"88042090068008003120000806001402504110C48002403601887FEF80022A51",
INIT_0D => X"26C0AC404E43032CA0C205880A7FFAB7FE01409400400C0594A4002200110008",
INIT_0E => X"26C0AC086A170250454004C6012280129B034A080C0B0016A0D20346080C0A80",
INIT_0F => X"0B064092D85938C0112144050224120C500346080C0B0016A0D2034A080C0A80",
INIT_10 => X"40702E058355458967E86A170220D1800093414B0414782E4B5000D81480809A",
INIT_11 => X"081B1545104135443306C35901024F88A88049062A747512B76783C5D040E080",
INIT_12 => X"40160040D86B202049B22198362A8A208279854400A036801480031401900800",
INIT_13 => X"0DD001C002D38334000914028354008301008C0CF1480245108C7640A0604032",
INIT_14 => X"AC0496022300233104662848808E191526205018030060540284FA0C0044022C",
INIT_15 => X"004010040100401004010040102090010008000001C0E010020007DFFFC06E60",
INIT_16 => X"0401004010040100401004010040100401004010040100401004010040100401",
INIT_17 => X"4010040100401004010040100401004010040100401004010040100401004010",
INIT_18 => X"FF7FFDF7FF3E3DFDF7E000000000000000000000000040100401004010040100",
INIT_19 => X"FBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBFFDFDFFFCF3CF3FFFEF9FEE",
INIT_1A => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFEFF7FBFDFEFF7FBFDFEFBEFBEFBEFBE",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0004000100000000000000000000000",
INIT_22 => X"2A954BA0004154BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080402010FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF552A974AA0004174BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"000400000007FFFFFFFFFFFFFFFFFFFFFFEF552E974BA0804000AAF7FFFFFFFF",
INIT_25 => X"FFFFFFDFEF5D2E974BA002E97400007FFFFFFFFFFFFFFFFFFFFFFEF552E954AA",
INIT_26 => X"BA087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974BA082E95400007FFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2E954BA007FC00BA5D7FFFFFFFFFFFFFFFFFFBFDFEF5D2A954AA002E974",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFBFD",
INIT_29 => X"954AA080005000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA00000200000000",
INIT_2A => X"FFFFFFFFFFFFFFF552A974BA0000174AAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0A000AAE3FFFFFFFFFFFFFFFFFFFFFFFEF552A974AA0000104AAF7FFFFFFFFFF",
INIT_2C => X"FFBFDFEF5D2E974AA000A07000007FFFFFFFFFFFFFFFFFFFFDFEF552E954BA08",
INIT_2D => X"1C7FFFFFFFFFFFFFFFFFFBFDFEF5D2A974BA002A95400087FFFFFFFFFFFFFFFF",
INIT_2E => X"F552E974BA0020924BA1C7FFFFFFFFFFFFFFFF7FBFDFFF5D2A954AA082A92428",
INIT_2F => X"FFFFFFFFFEFF7FBFFFFF552E974AA0071C50BA557FFFFFFFFFFFFFFFF7FBFDFF",
INIT_30 => X"4BA000002000000000000000000000000000000000000000000000000E3FFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2A954AA080017410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"000AAF7FFFFFFFFFFFFFFFFFFFFFFFEF552A974BA0000174BAFFFFFFFFFFFFFF",
INIT_33 => X"BFDFEF5D2A954BA082E800AAA2FFFFFFFFFFFFFFFFFFFFFDFEF552E954AA0004",
INIT_34 => X"7FFFFFFFFFFFFFEFF7FBFDFFF5D2A974AA002E95410087FFFFFFFFFFFFFFFF7F",
INIT_35 => X"52E974AA082A820AA557FFFFFFFFFFFFFEFF7FBFFFFF552E954BA002E9741008",
INIT_36 => X"FFFBFDFEFF7FFFFFEF5D2A974BA0000020AA557FFFFFFFFFFFDFEFF7FBFFFEF5",
INIT_37 => X"0000000000AAFFFFFFFFFFBFDFEFFFFFFDFEF5D2E954AA0051554BA5D7FFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(21),        -- Port A data input
DOA(0)   => data_read_a_hi(21),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(21),        -- Port B data input
DOB(0)   => data_read_b_hi(21),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_22_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"5290F4CDE914905A14A43D33F488243E17122300F55FEB189B343A1140548380",
INIT_01 => X"A94007B259F6A975386262000C344BA9573C6FF57B18A5FB0ABFCD3C2C5F4F0C",
INIT_02 => X"D56B4302AC01005111011BD506AA5205274056900596A539584E2E6DFE4B2418",
INIT_03 => X"6B03F2F6151A2081F24001E8400008F401CB10C6594423C8923AD6B55AD0EB5A",
INIT_04 => X"8001023D37E50880436200808BC8492A0089249600101100008087248B64426E",
INIT_05 => X"A51035B41C0A88046CAEE8C23C08E040011C0020F8882001102D620A06D68301",
INIT_06 => X"B93FF975CF7889D085E997A2144E8FC2060B880081A26DCD4047EFF9EF018980",
INIT_07 => X"283800AA500200E8024AD03546A3262FB5AA5542A882040C7A64CBD64065F028",
INIT_08 => X"141008801018040E48D500400015805060040080A2A0F4A82381B4000A0905A0",
INIT_09 => X"4D0000002126F30C902A29C54539C020E11810098D4067EFF9FF284D483E2AB4",
INIT_0A => X"1400006100003202D040050220103D2A512C6A8C4F0008AA800470370000A000",
INIT_0B => X"013456520CA09281C2A81C2A81C2A81C2A81C2A81C2A81C2A81C9540E1540E00",
INIT_0C => X"A1402A13C0A10A893165281A1C2A7283516344C594A85536B1AD800214202C50",
INIT_0D => X"3C70FC20515808A0100820112300011000287B071105034406950A0285014280",
INIT_0E => X"3C70FC48E11CFC48400184CE0D6783139B0959A41606003C70FA0958AC160480",
INIT_0F => X"0D87E8B3B811B52048B10E0402AE1606D80958AC1606003C70FA0959A4160480",
INIT_10 => X"80F84E0185594581E088E11CFC38414020DD42CF909D7E0A551C02180300C0DD",
INIT_11 => X"441154C258012D86F3044A3133004A99BD8455300654458A1D588C4061403000",
INIT_12 => X"A096A240894626600953379822A984B0025B0DEC0345C9200680027181B44887",
INIT_13 => X"E2404160035482BE521C2C04A90783C18000D610B9D8070B12B1A2A62040202A",
INIT_14 => X"304244A91102C93A2D608D2A258DF8034284200C050070E40C80620C870B02C4",
INIT_15 => X"4411044110441104411044110466C440446CA06951D4EA801000980400646002",
INIT_16 => X"0100441104411044110441104411044110441104411044110441104411044110",
INIT_17 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_18 => X"FE8FF1F7DEBDDF7DF7D05122890000000003FFFFFFFF90040100401004010040",
INIT_19 => X"79E79E79E79E79E79E79E79E79E79E79E79E79E7BFFDFD7DDDF7DF7DF7DFBFDE",
INIT_1A => X"3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE79E79E79E79E",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE000000000000000003F9FCFE7F3F9FCFE7F3F9FCFE7F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0800000000000000000000000000000",
INIT_22 => X"2E974AA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000400010FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E954AA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"0004154BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA000015400FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF552A974AA0800154AAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA",
INIT_26 => X"BAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0004174BAFFFFFFFFFFFFFFFFF",
INIT_27 => X"FEF552E974BA0804000AAA2FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0000174",
INIT_28 => X"0000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040001000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E954AA000402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0417410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080005000FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF552A974BA0000174AAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA00",
INIT_2D => X"E3FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0804154BAF7FFFFFFFFFFFFFFFFF",
INIT_2E => X"F552E954BA000E124BAE3FFFFFFFFFFFFFFFFFFFFFFFEF552A974AA0000104AA",
INIT_2F => X"FFFFFFFFFFFFFFFFDFEF552E954BA080A000AAA2FFFFFFFFFFFFFFFFFFFFFFFE",
INIT_30 => X"4BA080400010000000000000000000000000000000000000000000000007FFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"17410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000400010FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF552A954BA000415400FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954AA0800",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFEF552A974BA0000174BAF7FFFFFFFFFFFFFFFFFFF",
INIT_35 => X"52E954AA0004000AAA2FFFFFFFFFFFFFFFFFFFFFDFEF552E974AA0804174AAF7",
INIT_36 => X"FFFFFFFFFFFFBFDFEF5D2E954BA002A820BAA2FFFFFFFFFFFFFFFFFFFFFDFEF5",
INIT_37 => X"0000000000087FFFFFFFFFFFFFFFF7FBFDFEF5D2A954BA082E800AAAAFFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000000FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(22),        -- Port A data input
DOA(0)   => data_read_a_hi(22),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(22),        -- Port B data input
DOB(0)   => data_read_b_hi(22),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_23_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"EF20906D902424807BC8241BC81801B97D38AD3C0800103362A6741C80A12A02",
INIT_01 => X"001FFF8409F089003B4422000D80C80106804A7951C5B9D1C828043EA28838F9",
INIT_02 => X"028406A002DC176444683862400003111001303FFC00F240D50146013B300500",
INIT_03 => X"001B243004080FE000177003145F87017D584B10D804034800200200A1008008",
INIT_04 => X"BEFFFC0248005FFC3C18A2FFE12222425E600000BDC0800AEE01E81A100F0A00",
INIT_05 => X"D03F8000000003FF810640A1C0008FF2F0E17E1F02FFFFC80100004044800080",
INIT_06 => X"800264B4854650040123428C204BF40F439647FF4807E189A477EF81DF0AF116",
INIT_07 => X"01000000FFDFFFE800401005C0A0008F86C60840AAAA100C68D1810C9F4A0020",
INIT_08 => X"1BE1F5F80003FF0002021FFEFBC80000000077FF184B03010004002FE1F29002",
INIT_09 => X"907FC308181204800600000000001BFFA800808189A657EF81DD0C00079CC800",
INIT_0A => X"0063090442A18001B188300C48907120AC810033149249C433200180082A06FF",
INIT_0B => X"9A41C1443243050C1010C1010C1010C1010C1010C1010C1010C1008608086084",
INIT_0C => X"000082A00600200080000500C000400800601200000254A000007FEFC1030221",
INIT_0D => X"0A9080400E0BF30C20CA858E087FFABFFE01409780214EE49620001000080004",
INIT_0E => X"0A908044294700701641005218521210150E5789F90A000A90800E5F81F90880",
INIT_0F => X"0E0220036864A7DCA190440301E2105C000E5F81F90A000A90800E5789F90880",
INIT_10 => X"C1400500C6CE5400032429470068924010164302048156305D66F8701681000E",
INIT_11 => X"2E0CCB0500013440600339C800004D8018000857A82920CE8CB220C81400A180",
INIT_12 => X"220344406739000009B0030019960A00026880C0422C52B01700044901488822",
INIT_13 => X"85C811A010428104128996465ADA020180804A040108A2658217C4008060300C",
INIT_14 => X"BE0692020328CA0028042054A92771C50FC070109000C1C819078280A265920E",
INIT_15 => X"020080200802008020080200800800200200000000000008004807DFFF000470",
INIT_16 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_17 => X"0080200802008020080200802008020080200802008020080200802008020080",
INIT_18 => X"0000000000000000000000000000000000000000000000802008020080200802",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000",
INIT_22 => X"2E974BA080002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E974BA000400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000400000FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF5D2E954AA080000010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA",
INIT_26 => X"10FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080402010FFFFFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2A954BA000015400FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA0804000",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E974BA080002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF5D2E954AA000402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA00",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080002010FFFFFFFFFFFFFFFFFFF",
INIT_2E => X"F5D2A954BA080407000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080005000",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF5D2A954BA000417410FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA080402000000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"02000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000010FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF5D2E974AA000402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0000",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000400010FFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"D2A954AA080017410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954AA080002000FF",
INIT_36 => X"FFFFFFFFFFFFFFFFFF552A954BA080015410FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_37 => X"0000000000F7FFFFFFFFFFFFFFFFFFFFFFFFF552A954BA000415400F7FFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000000FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(23),        -- Port A data input
DOA(0)   => data_read_a_hi(23),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(23),        -- Port B data input
DOB(0)   => data_read_b_hi(23),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_24_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100600007FFF000080108004000800020000840041000080808",
INIT_02 => X"0000068002CC07400000090C080002000000103FF811F150231000520ABE4404",
INIT_03 => X"8428180000080FE000177000001B87003D4000000E8B84010020000000008000",
INIT_04 => X"3E2FFC024800137C3C000077E00000001E6000003CC0000A6601E01A000F0200",
INIT_05 => X"103F8000000003FF80000021C0000FF0F0E03E1F0067FFC00000000000000000",
INIT_06 => X"00132412079001AD00810005E8000001401643FE4007E5501AA00000DC8C3006",
INIT_07 => X"000000000FDFFF62695A5685C094831D966000008002100C2040A178B600C240",
INIT_08 => X"08E1F5F80001FF00000007FEFBC00000000077FF000B00000000002FE0000000",
INIT_09 => X"107FC300000000000600000000001BFFA0000005501AA00000CE200000940000",
INIT_0A => X"00630104408180012188300C00814080008000010012414433000100080806FD",
INIT_0B => X"904181003003000C1000C1000C1000C1000C1000C1000C1000C1000608006084",
INIT_0C => X"00000080060000000000000012002C00000000000000000000007FEF80020201",
INIT_0D => X"440082404E0B332CA2C20188087FFAB7FE000082000000008220000000000000",
INIT_0E => X"4400824903210308074084210002460402009280010D80440084009280010F00",
INIT_0F => X"800A2400401A0C82183248060010280C20009280010D80440084009280010F00",
INIT_10 => X"C0A078160000404A0469032102981380202080026420020D06C002A08481C020",
INIT_11 => X"00164F400860000824059AD01802000208104817B00011306B2D9B0DD5082080",
INIT_12 => X"41021800B35A0300400041202C9E8010C0001040C5836CC01780018601030088",
INIT_13 => X"DB1011E000A140058220004AEFFC8101810021084301880030A8B77400603011",
INIT_14 => X"8C063C0220002201490418082010A57263E010000201033016085A40880030A1",
INIT_15 => X"000000000000000000000000000000000000000000000000000007DFFF0006E0",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"F6E7CC1132CDB444199000000000000000000000000000000000000000000000",
INIT_19 => X"79E79E79E79EFBEFBEFBEFBEFBEF9EF9EF9EF9EFA69861219575D75FF2D0AEEA",
INIT_1A => X"0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1EFBEFBEFBE79E",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE000000000000000000783C1E0F0783C1E0F0783C1E0F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020100000000000000000000000",
INIT_22 => X"2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"080002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_26 => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000400010FFFFFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2E974AA000400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0004000",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040201000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF5D2E974BA080002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFF",
INIT_2E => X"F5D2E974AA000400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF5D2E974AA000400000FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA080402010000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"00010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000010FFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002010FF",
INIT_36 => X"FFFFFFFFFFFFFFFFFF5D2E974AA000002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_37 => X"0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000402010FFFFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(24),        -- Port A data input
DOA(0)   => data_read_a_hi(24),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(24),        -- Port B data input
DOB(0)   => data_read_b_hi(24),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_25_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100200002000000080100004000000020000800041000080808",
INIT_02 => X"0000068002CC474000000800000002000000103FFCE302008000000880844A04",
INIT_03 => X"00000101C0200FF004177800081B87003D400000080000000020000000008000",
INIT_04 => X"3E2FFE024820137C3C004077F01000001E7249213CC1264A660DF05A000F9000",
INIT_05 => X"103F81C1002203FF80000021C1140FF8F0E03E1F0067FFE04800258280010052",
INIT_06 => X"80480AE20000000100000001C8608001401643FE4007C00000000000CC083006",
INIT_07 => X"280800000FDFFFEA4050140540B00100840000080002A00C2040810000000010",
INIT_08 => X"C8E1F5FA21C9FF80040007FEFBE031018C31F7FFBAEBC0020008086FE0000100",
INIT_09 => X"107FC301800000000600000000001BFFE00301000000000000CC020000140000",
INIT_0A => X"0077330C4889CC292588300C0080400000800001001243443B000100880806FD",
INIT_0B => X"904189003003000C1000C1000C1000C1000C1000C1000C1000C1000608006084",
INIT_0C => X"8B04228026824100000000000000000000000000000004A000007FEF80020201",
INIT_0D => X"400000400E03C30C20C2818C087FFAB7FE01409700C10007962418220C110608",
INIT_0E => X"4000000001010000004000000000400400001200000800400000001200000800",
INIT_0F => X"0008000000000480000040000000200000001200000800400000001200000800",
INIT_10 => X"0000001001000002000001010000100000000000202000000440000000800000",
INIT_11 => X"0000410000000008000008400000000200000806300400000820000020004880",
INIT_12 => X"0000080001080000000040000082000000001000000040800800000000020008",
INIT_13 => X"8100000000000000802000000840000200040000020008000000840000804000",
INIT_14 => X"8C04100200000200000610000000210000000018140000000008000008000000",
INIT_15 => X"04411044110441104411044510629041040D180400000010028047DFFF800C60",
INIT_16 => X"4411044110441104411044110441104411044110441104411044110441104411",
INIT_17 => X"4110441104411044110441104411044110441104411044110441104411044110",
INIT_18 => X"196A8C5A2932EC15DA080800002FFFFFFFFFFFFFFFFFC1104411044110441104",
INIT_19 => X"92492492492410410410410410410492410492412000531215A69A6BFBA2894A",
INIT_1A => X"B158AC562B158AC562B158AC562B1588C46231188C46231188C4924924924924",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000B158AC562B158AC562B158AC562",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000",
INIT_22 => X"2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF5D2E974BA080400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_26 => X"10FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0800000",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400000FFFFFFFFFFFFFFFFFFF",
INIT_2E => X"F5D2E974BA080000010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA080402000000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"02000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400000FF",
INIT_36 => X"FFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_37 => X"0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000000FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(25),        -- Port A data input
DOA(0)   => data_read_a_hi(25),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(25),        -- Port B data input
DOB(0)   => data_read_b_hi(25),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_26_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"E9264EAB20190CA3BA4997AA9002AE9C001006B0778015CFA17E0811039879C7",
INIT_01 => X"F1FFF9BB1F773C7F9BB07DFFFDD863FC5FFF3FEFFBBF9FFB22FFFBC7B9F30686",
INIT_02 => X"9B3184F8AFDEAF300029E4E300FC78A6258548EFFA71C00172082400003A2161",
INIT_03 => X"0213C3FDFFFC7F74FFBF737A603B87FEBE1A5294F65628A0001B9CE6CC606E73",
INIT_04 => X"7E2EFEBF6FFEB37C3FF3017776FFCDA43E7B6DFD7DEBFD8E6F5F78DF0BFBD644",
INIT_05 => X"902F87C74E8CCFFBB6FF70E1FE61FFBDF0FEBE1FFD67DFFEFFBDA7F7FED50870",
INIT_06 => X"213246200BCC8920360C1831CD7DF60A244B9BFEE00589DDBCEFEDC1DFA08957",
INIT_07 => X"B1D4223B4FFDFF21CC721C85DCE1458E8782484020A2C1FCA3468D77E0000300",
INIT_08 => X"2C05FD7BC471FBD13D980FBEFBEBF30B8D79FF7F451F33CFD60FE8FFFDF54003",
INIT_09 => X"19FFC71FEFED7B251E35768E8ED6BFDF3EB3EBF9DDBCE7FDC1DF8A760F3EACC0",
INIT_0A => X"56F7730ECCDBDF152199F51EDDCDEBCFF589807B7096CD4CF73AC1FC98884FFF",
INIT_0B => X"B867D3683A03A40F78C0D78C0D78C0D78C0D78C0D78C0D78C0D7A606BC606B8C",
INIT_0C => X"DFBFF5EB36DFE51FC3A80D73D840303983EE7F0EA03BDA680137FFFDFFD7E681",
INIT_0D => X"3F0080425E6BFF8DB0DAE19C09FFFFE7FE3EBEA8EB7AFEE5C9AEBD7F5EBFAF5F",
INIT_0E => X"3F00800DEC010280004000F808020290100FA2F60008003F00800FA2F6000800",
INIT_0F => X"00023002007BC0A14E00400003B8000D000FA2F60008003F00800FA2F6000800",
INIT_10 => X"01E0320007204008040DEC010300100000F600020581003F604D0700008000EE",
INIT_11 => X"201F21A2C40039006807C46426040E101A0259DFE82011A311AA042016040080",
INIT_12 => X"80020048F88C84C101C203403E434588007200D047F00090200007E0010009B0",
INIT_13 => X"0109000003E2000416C0804FE04140E80000F808010AB02033AC048A2A00003D",
INIT_14 => X"FFAFD082003B032FB987E04021D481D4000419060201E1A000044300B02033E8",
INIT_15 => X"AFEBFAFEBFAFEBFAFEBFAFEFFBFBFBFBBFCFBB0FFDFEFFEF2DFFFFFBFF802FFD",
INIT_16 => X"FEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBF",
INIT_17 => X"EBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFA",
INIT_18 => X"F491E166CC8553F86EDB5C88646FFFFFFFFFFFFFFFFFEBFAFEBFAFEBFAFEBFAF",
INIT_19 => X"1861861861861861861861861861869A69A61861AFBD54D5F871C71D475B15BC",
INIT_1A => X"0984C26130984C26130984C26130984C26130984C26130984C26186186186186",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE000000000000000000984C26130984C26130984C2613",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000",
INIT_22 => X"2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_26 => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFF",
INIT_2E => X"F5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA080402000000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"02010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_36 => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_37 => X"0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(26),        -- Port A data input
DOA(0)   => data_read_a_hi(26),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(26),        -- Port B data input
DOB(0)   => data_read_b_hi(26),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_27_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"00080A40000A41248002029000050A088000008242A0004404480002000A1155",
INIT_01 => X"F1FFF1C11F781C129C107DFFFE0860941E81258CA2B71C2220EC1B86E1A00002",
INIT_02 => X"183080988B2EAE00002BE001117C78C6848140CFFA0000800042008000011081",
INIT_03 => X"000003FDF3E47C74F7BCF36A203A47F6B8184210B6160820001318C60C204C63",
INIT_04 => X"7E28FEBF6FEEB3723F71017476DFC524397B6DF572EB6C8E175E70D90F539600",
INIT_05 => X"000F86064C8DDFE3B6FF50D1FC61DE39C8FCB91FF9671FE6B68984B5BCE40834",
INIT_06 => X"0000000800000042020C18300520620A80231BFE200181092CE7ED80DFC00147",
INIT_07 => X"8AC4AA3B0FD1FF201044110560884000840200520002080C23468D0300000282",
INIT_08 => X"2005F0784411E390A4880E3DF7E2FB0B8E717C7F411F3BC6D60B60FFDDE44001",
INIT_09 => X"18FFD757E7ED7A211E81C09818109E1F16B16B71092CE7ED81CF403601228C40",
INIT_0A => X"46FF730E5CCBCD55219AB55F0DEFABC7054880693016DD4C755AC16C1A884FFE",
INIT_0B => X"BC63F1683803C00E3440C3440C3440C3440C3440C3440C3440C3C2061A2061AD",
INIT_0C => X"56BF55CB165EC51D41880FA3F040202883B475062033186801137FF1BAD6F281",
INIT_0D => X"3B0000421E2B0F2E2AE215C808FFFA47FE62BAA86B1AB268E92AB56D5AB6AD5B",
INIT_0E => X"3B000025EC010080004000F808000098100F22520008003B00002F2252000800",
INIT_0F => X"00001042006BC0810600400003B80001002F22520008003B00002F2252000800",
INIT_10 => X"01E032000620000C0405EC010100100000F6000001C1003760410500008000EE",
INIT_11 => X"201D2120840039000817444404040E10020218DE282010A311AA002002040080",
INIT_12 => X"8000000AE888808101C20040BA4241080072001027F00080200007E0000001F0",
INIT_13 => X"0101000003E2000007C0800FE04040280000F8080002F02023AC04080A00003D",
INIT_14 => X"DDAFD082001B03249887E04001D481D4000009020201E1A000040100F02023E8",
INIT_15 => X"ADAB6ADAB6ADAB6ADAB6ADAB6BF1EBDABD8E270BF84A25C6ACB777E3FF800C6D",
INIT_16 => X"DAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6",
INIT_17 => X"AB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6A",
INIT_18 => X"100481CA860402104A471688747FFFFFFFFFFFFFFFFFAB6ADAB6ADAB6ADAB6AD",
INIT_19 => X"0000000000000000000000000008200000000000200072F210000001490E2168",
INIT_1A => X"A05028140A05028140A05028140A050080402010080402010080000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000A05028140A05028140A05028140",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000",
INIT_22 => X"2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_26 => X"10FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFF",
INIT_2E => X"F5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA080402000000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"02000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FF",
INIT_36 => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_37 => X"0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000000FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(27),        -- Port A data input
DOA(0)   => data_read_a_hi(27),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(27),        -- Port B data input
DOB(0)   => data_read_b_hi(27),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_28_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"02200AA400180030808802A900002A08001280A08A801044104A1000001818C3",
INIT_01 => X"50A00011460214428114180000882214413D0A71592A01D92213D28005210202",
INIT_02 => X"8A54800A210200111100C2110054289220810440030404010844000444410001",
INIT_03 => X"4200040822D4500001E0000028000002000211842010092000018C6295200631",
INIT_04 => X"00400000000B8000000140000005840C00000040002008808100048100100044",
INIT_05 => X"0000222200244400135110000135100000000000000000024CA0A01018000320",
INIT_06 => X"A004912008208040024489121144080400081000200008104000000020000041",
INIT_07 => X"A85800994000000A0200802004204420210001022AA8A0001122448142491008",
INIT_08 => X"0414000201800004080A000000124058200408000880004440004080160C4100",
INIT_09 => X"0080000206CB0821082B694D4D29400002002038104000000020003204000440",
INIT_0A => X"12000843066021001400040024440245400082D022040000400800081022C000",
INIT_0B => X"0002002C004001036050160501605016050160501605016050160280B0280B00",
INIT_0C => X"0012400810080414C0A800310840102182C62302A0194C08001680100E4040A0",
INIT_0D => X"05000002003004208208841401800040000A0000200814004198000400020001",
INIT_0E => X"0500000004000080000000000000028000002052000000050000002052000000",
INIT_0F => X"0000300000004001060000000000000900002052000000050000002052000000",
INIT_10 => X"0000000001200000000004000100000000000000050000002001050000000000",
INIT_11 => X"00002020840000004800040404040000120200A9000000010000002002040000",
INIT_12 => X"0000004800808081000002400040410800000090001000002000000000000910",
INIT_13 => X"0001000000000000144000010000402800000000000A1000010000080A000000",
INIT_14 => X"0080000000110006B08140000040000000000902000000000000410010000100",
INIT_15 => X"0080200802008020080200802101210810C39A66A90A85420413A82000000204",
INIT_16 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_17 => X"8020080200802008020080200802008020080200802008020080200802008020",
INIT_18 => X"110A00246972BD89A40A0C22E100000000000000000000200802008020080200",
INIT_19 => X"82082082082082082082082082082082082082080D35050758C30C31DE21102C",
INIT_1A => X"B0582C160B0582C160B0582C160B0580C06030180C06030180C0820820820820",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000B0582C160B0582C160B0582C160",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000",
INIT_22 => X"2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_26 => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFF",
INIT_2E => X"F5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA080402000000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"02000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_36 => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_37 => X"0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000000FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(28),        -- Port A data input
DOA(0)   => data_read_a_hi(28),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(28),        -- Port B data input
DOB(0)   => data_read_b_hi(28),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_29_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"79964E4BA01DACAB9E659792D00AAE160002829C7FDFEFCEE97C2815039D70C3",
INIT_01 => X"50BFF9AB0775343F9AB01DF80D5821FC0FFF3FEFD1AF9FF1207FFBC7B9720586",
INIT_02 => X"0D15846807D207200021C4E200D428A2018408600271C000720A0000003A2161",
INIT_03 => X"0002C009EEFC5F10F9B70178681B80FA3E000100765029A00019084345606421",
INIT_04 => X"3E6E023D27DA937C03E3407712E5CDA41E0924DC3D20B98AE905189F0BF8C000",
INIT_05 => X"902003C30E0447F877F930203E213F8CF01E3E00FC67C03A4D9C87525E510160",
INIT_06 => X"0012460003CC002036040811D919F402244293FEE00400CCB46BA4C164A08857",
INIT_07 => X"914800110FFC0001CC320C81D841418E82800100000041FCA1428575A0001108",
INIT_08 => X"0805FD0180E1F8C1111A0782082B50080508FF00048B124D4005C8AFF4154102",
INIT_09 => X"0180000ABFEF89250815568A8AD6ABC02A02A0B0CCB463B4C0748A720B1EA4C0",
INIT_0A => X"021410028450530014014002D445624DB481806A62840800C22800B8900042FF",
INIT_0B => X"0806522C0A40A50268D0068D0068D0068D0068D0068D0068D006A68034680300",
INIT_0C => X"8912E0A83289641F42A80561D040203182AC3D0AA0118A080036FFFC4F4164A0",
INIT_0D => X"050080424069F5A51250648801BFFFE0003E3E00A0685A85410C0816040B0205",
INIT_0E => X"050080080400028000000000000202900000A0F600000005008000A0F6000000",
INIT_0F => X"00023000001040214E0000000000000D0000A0F600000005008000A0F6000000",
INIT_10 => X"000000000120400800080400030000000000000205800008200D070000000000",
INIT_11 => X"000220A2C400000068008424260400001A0241DAC80001010000042016040000",
INIT_12 => X"00020048108484C10000034004414588000000D04010001020000000010009B0",
INIT_13 => X"000900000000000416C00041000140E800000000010AB0001100008A2A000000",
INIT_14 => X"A282C0000033010FB181E00020400000000419060000000000004300B0001100",
INIT_15 => X"02C0B02C0B02C0B02C0B02C4B12B312912831A27FCFE7FFB175B6FF800802594",
INIT_16 => X"2C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B",
INIT_17 => X"C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B0",
INIT_18 => X"EE7FFDF7FE783FFDFFEA0C00602FFFFFFFFFFFFFFFFFC0B02C0B02C0B02C0B02",
INIT_19 => X"BEFBEFBEFBEFBEFBEFBEFBEFBEEBAEBAEBAEBAEBBFFDF9FBEFFFFFFEBBCF9F96",
INIT_1A => X"FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFBEFBEFBEFBEF",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000FBFDFEFF7FBFDFEFF7FBFDFEFF7",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000",
INIT_22 => X"2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_26 => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFF",
INIT_2E => X"F5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA080402000000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"02000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_36 => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_37 => X"0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(29),        -- Port A data input
DOA(0)   => data_read_a_hi(29),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(29),        -- Port B data input
DOB(0)   => data_read_b_hi(29),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_30_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"FF9FE1F7FFBFFFFDFFD000000000000000000000000000000000000000000000",
INIT_19 => X"79E79E79E79E79E79E79E79E79E79E79E79E79E7AFBD75F5FDF7DF7FF7FFBFFE",
INIT_1A => X"3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE79E79E79E79E",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE000000000000000003F9FCFE7F3F9FCFE7F3F9FCFE7F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000",
INIT_22 => X"2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_26 => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFF",
INIT_2E => X"F5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA080402000000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"02000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_36 => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_37 => X"0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(30),        -- Port A data input
DOA(0)   => data_read_a_hi(30),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(30),        -- Port B data input
DOB(0)   => data_read_b_hi(30),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_31_7 : RAMB16_S1_S1
generic map (
INIT_00 => X"129000008004A00804A40000400800020000000C005FEA005800200400050100",
INIT_01 => X"A15FF18019700810180065FFFC0040801E80258CA2951C2200EC0906A0804140",
INIT_02 => X"146000808A0C060444692000402850040400408FF80000000010000000004000",
INIT_03 => X"000003F5D1202C70F654716A001A07F438184210960600000012108518004842",
INIT_04 => X"3E28FE3F6FE513703F70007472DA4128187B6DB530C1240A060C70580B439200",
INIT_05 => X"000F84040C088BE3E4AE40C1FD04CE38C0FC381FF8671FE01009048084C40010",
INIT_06 => X"0000000000000008000810200420620E00030BFE000181092CE7ED80DF800106",
INIT_07 => X"000000220FD1FF200040100540800000840200408002000C2244890200000200",
INIT_08 => X"0011F0780011E38004800E3CF3E0B1118C31747F000B33820209206FC9E80000",
INIT_09 => X"187FC301B124F2001600000000001A1F00110101092CE7ED81CF000401228800",
INIT_0A => X"0477330C4889CC012188310E08812982050800A91012494C31004124080886FE",
INIT_0B => X"9861D1403803800C1000C1000C1000C1000C1000C1000C1000C1800608006084",
INIT_0C => X"020400830602410901000D02D0002008012054040022102001017FE190022201",
INIT_0D => X"3A0000401E030B0C20C20188087FFA07FE203A80010002608030102008100408",
INIT_0E => X"3A000005E8010000004000F808000010100F02000008003A00000F0200000800",
INIT_0F => X"00000002006B80800000400003B80000000F02000008003A00000F0200000800",
INIT_10 => X"01E03200060000080405E8010000100000F600000081003740400000008000EE",
INIT_11 => X"201D0100000039000007404000000E1000001846282010A211AA000000000080",
INIT_12 => X"80000000E808000001C200003A0200000072000007E00080000007E0000000A0",
INIT_13 => X"0100000003E200000280800EE04000000000F8080000A02022AC04000000003D",
INIT_14 => X"9C06D082000A03200806A040019481D4000000000201E1A000040000A02022E8",
INIT_15 => X"0401004010040100401004010060C040040C200950402090128057C3FF800C60",
INIT_16 => X"4010040100401004010040100401004010040100401004010040100401004010",
INIT_17 => X"0100401004010040100401004010040100401004010040100401004010040100",
INIT_18 => X"000000000000000000001000802FFFFFFFFFFFFFFFFF81004010040100401004",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000",
INIT_22 => X"2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_26 => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFF",
INIT_2E => X"F5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA080402000000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"02000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_36 => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_37 => X"0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(31),        -- Port A data input
DOA(0)   => data_read_a_hi(31),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(31),        -- Port B data input
DOB(0)   => data_read_b_hi(31),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_0_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"ED39BA795990D275FB4A6E96ACC4731DEA4598B0AFB54867F6EE4618C3749803",
INIT_01 => X"58A0047C8607844847CA180001E4A2404042106208408208C2002069161734B3",
INIT_02 => X"8B1EC9562121F8051500147A0E5629A302CF28400615F5787B09FBF999BB1EFD",
INIT_03 => X"404EFC0A2AD6100F01A88E851CE47803C280110521898F6996088862C7B22221",
INIT_04 => X"C0D001C0100AEC83C008E7880D01A64661800002C21A52C590D2012194804844",
INIT_05 => X"650002C3F08754001B51981E007910070F01C1E003980015A204C22F32328BAF",
INIT_06 => X"BCDA4677CAEE7CF5BB870E1DDB9889C5FBFC440129A0604442180238203F70C1",
INIT_07 => X"7AAE0088B02000C2EC3A0E829836E0AF3325372E2AA8FDF3C18306758B24197A",
INIT_08 => X"D7E40002F7AE005FFB4730010411400A61080000F7F4C464B58294901606D5A5",
INIT_09 => X"C4801C40469B0CA9881A28C141118000C5A85A60444210123820B43B40804274",
INIT_0A => X"400800219010107ED453C041B13216656074EA560F0092A24856B05312226900",
INIT_0B => X"27122C3E04E03383E2781EA781E2781EA781E2781EA781E2781C33C0613C0E29",
INIT_0C => X"74EB1F50D0758A9650E520610A6A57A5529E2B439499CF96B086000000B09870",
INIT_0D => X"04F07E024108F4E28638EC57250004480155C1375A97A9121F8BA749D3A4E9D2",
INIT_0E => X"04F07E42177EFDF8570184071575970F8FC07D5BFF078004F07E007D5BFF0780",
INIT_0F => X"8F85ECB1FE047F5FB7B30E0700461E5AF8007D5BFF078004F07E007D5BFF0780",
INIT_10 => X"C0184D07C1DF15C7E3E2177EFDF8C3C03009C3CDD47C7F403FB3FDF89701C011",
INIT_11 => X"4F80FE659C6104C6D7103F9D1D064189B5924418D65FE45DEE55BBEDE34CF900",
INIT_12 => X"6395F64207F3A3A1483136B881FCCB38C2098DACA01FFF603F80001F80FDC81F",
INIT_13 => X"FED151E01015C3BB507D3F811FBEC32B81840714F8D91F4FC513F37C8AE07002",
INIT_14 => X"61692F293185D8D724E15D3FCC6B7C236FE0691A9500125C1F83F8CC1F4FC507",
INIT_15 => X"E93A4E93A4E93A4E93A4E93A4F942F90E9628540052090650525A0000066A00B",
INIT_16 => X"93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4",
INIT_17 => X"3A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E",
INIT_18 => X"09B56C74DAB15D1CF13501AA495000000000000000003A4E93A4E93A4E93A4E9",
INIT_19 => X"2082082082082082082082082082082082082082082084E41DC71C7155F3898E",
INIT_1A => X"3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F8208208208208",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE5294A5294A52800003E1F0F87C3E1F0F87C3E1F0F87C",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000030FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"A975EFFFAABDE00FFAEBDFFF5D2EAAAAAF7AEBDEBA0000000000000000000000",
INIT_22 => X"8000155087FC0155F7D168B55007BFDF45085168ABA002E82145085155545F7A",
INIT_23 => X"FFFD7545AA8028A00A2802AABAFF8028BEF5D7FFFE10005542145557FD5545FF",
INIT_24 => X"F7AEAAAAAA2FFFDF4500043FE105D2E954BAF7FFC0010080017555555568AAAF",
INIT_25 => X"A5D5168A00A2D142155005142010FFAE820AAFF842AABAA2AE95545FFD168ABA",
INIT_26 => X"FF5D2A821550000000BA007FD55FF5D7FC0145007FD7400550415410002E974B",
INIT_27 => X"F455D5142000082E82145FFD17DFEFFFD168BFFF780000BA007FE8AAAFF803FF",
INIT_28 => X"0000000000000000000000000000000000000000AAFBEAA00007BFDFFF082EBD",
INIT_29 => X"AABEA495FC716F002A975FFE3AA95E00EBAEBDFD75D2AA8A80EA8E2FE3F00000",
INIT_2A => X"56A16D557BC257D415E0216FA3F1E8FC0145B68B551475FAF6D1C556F0AA1C24",
INIT_2B => X"7FD24AFE3D02DAAAE12BD5545A2803AA0000542A0070071C50BAFEF1FAE0016D",
INIT_2C => X"A8B50F55A2F150005A3A438BD04AFAB8F550A8010E004924874825D7FEAA8548",
INIT_2D => X"A2A5504001C74BA42A1571E8028E3DB7816D0120155EA568E870BAEB8A05A2AE",
INIT_2E => X"2FFAFD2A82485FD2415A105C21451ED42A002545E055FFBE81D0BE8EA8A3AA05",
INIT_2F => X"100AA1D0F6F480B6A555A2A57A002A3D5FDB6A5C7E3DFFFE90B45B47ABA497A8",
INIT_30 => X"A0AFE80A8B0A000000000000000000000000000000000000000000000B55EAAA",
INIT_31 => X"ABEF5D557FEBA55022A3F70C6B405F4D2AE975EFAAAAB5E1AF3AABFF45592E88",
INIT_32 => X"411A8DED57CE1055555E5F58EFFC01FE2CACB65F520EBE9EF67D7BEA1FD5D556",
INIT_33 => X"A4AD0079C75D6070CC5CBB0280C029ABAA3EBC114728007521170821CE0FDE69",
INIT_34 => X"2A95E02A2AAB5EB0F280800EFAEE9F5D18F3142341D5DEEBEF55080034E0A592",
INIT_35 => X"B69C30E02116220415A9540AA854140A0A2047F353AAF6C77F7F20D968BF5781",
INIT_36 => X"ABEBE1B4D792A4AD1183454180DD3FDCAAAB7C91565455C141E41887D58AC448",
INIT_37 => X"F0000001FF01EABC4B8014174FF7DA80F52FEDE6BE93172D7D625B556EEAB157",
INIT_38 => X"FF0000001FF0000001FF0000001FF0000001FF0000001FF0000001FF0000001F",
INIT_39 => X"0000000000000000000000000001FF0000001FF0000001FF0000001FF0000001",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000100000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(0),        -- Port A data input
DOA(0)   => data_read_a_lo_256(0),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(0),        -- Port B data input
DOB(0)   => data_read_b_lo_256(0),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_1_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"212C001411984004084D000508C53810A03D1450E839B003342114428A000803",
INIT_01 => X"08000011400A100A81160000008C005400400002000000000000028001340000",
INIT_02 => X"C084484000002014400205851002007030450E0000A606C8C44CB4C6666C00E0",
INIT_03 => X"33DF380008164004000002000C80400002031943000101091608463061120118",
INIT_04 => X"4140008000000002000064000400004201000000000210458010070080100433",
INIT_05 => X"8500101040200000010009100000000508000100000000002010600100208D04",
INIT_06 => X"B5EDFDE24618AD433060C182BA860044204C000008A004100008000820280020",
INIT_07 => X"581E02100020000A81244890AA20263030517F122AA801F0983060AC564BF808",
INIT_08 => X"00820800C7A00045B103200000140A02234808000584000004808400020011A4",
INIT_09 => X"0000104000020082800808111008400000200204100000100820800144000414",
INIT_0A => X"12804062945211441E13C051156E800008402802060C94000040901102800000",
INIT_0B => X"24002006406401918C191AC191A4191A4191AC191AC191A4191A00C8560C8D29",
INIT_0C => X"0408010040050880383820080F105F05800302E0E08842422006000000041032",
INIT_0D => X"05000600000090C1841808172580000000008008020084082080204010200810",
INIT_0E => X"0500066210000178470184000000878402C000001E07800500062000001E0780",
INIT_0F => X"00003C404600000011A30E0700000009382000001E07800500062000001E0780",
INIT_10 => X"C0180000012010C20022100000F0C3C03000000055200340000000F88701C000",
INIT_11 => X"05800241186100004D100098190240001290002050068000001010486140F900",
INIT_12 => X"0000164A001303204800026880048230C2000094A0000F601F8000000001C908",
INIT_13 => X"12D051E01000000154200580003C030381840000004B08014401025480E07000",
INIT_14 => X"40082300218450C2800010094000482142E0601895001000000041C408014400",
INIT_15 => X"0802008020080200802008020080008208600500A82A15008000000000468000",
INIT_16 => X"8020080200802008020080200802008020080200802008020080200802008020",
INIT_17 => X"0200802008020080200802008020080200802008020080200802008020080200",
INIT_18 => X"BABEFC54A0810C7452B5420A1000000000000000000002008020080200802008",
INIT_19 => X"AAAAAAAAAAAAAAAAAAAAAAAAAAA28A28A28A28A2A8218D2C0C92492581328A46",
INIT_1A => X"2E974BA5D2E974BA5D2E974BA5D2E975BADD6EB75BADD6EB75BAAAAAAAAAAAAA",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFF6318C6318C63000002E974BA5D2E974BA5D2E974BA5D",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"00000000000000000000000C0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"002155557FFFFFF007FC21EFA2FFD74AAAAD5555550000000000000000000000",
INIT_22 => X"7FD75FFAAAA800AAF7AA974BAFFFBE8B45F7AEBDF455D2EAABEFF7FFE8BFF5D0",
INIT_23 => X"0557DF45AAD1400BAA2AE801550051555EFF7AA95400552AAAABAFFD1574105D",
INIT_24 => X"FFFBEAB55F780020AAAA80020AA082EAAB5500517DF555D2EAAA105500001550",
INIT_25 => X"AF7AE820AA0851574BAA2D1574AA5D7BFDEBAFFD540155557FD5400F78028BFF",
INIT_26 => X"FFFFD56AAAAFFFFD7555AAD168B45AAAEAAABAFF842ABEF5D517DF55552A974A",
INIT_27 => X"4BAF7AE80010082A97410557FEABFFAAFBE8BEFAAD1575EF557FFFE10557FFFF",
INIT_28 => X"00000000000000000000000000000000000000005D7FFDF4500043FE105D2E95",
INIT_29 => X"A8BC2EBDFEAF7F1F840017D4975D2FEF147FC51C7A2FBD5490BFD1C056A00000",
INIT_2A => X"AA8AAAE3D145410F7F1D55D71C002DABAEBAA974BAF7FFEFB45FFAABDF55492A",
INIT_2B => X"0E2AE85028B40155145F7AF6DBED5450AA1C2080BEF495FC71D54124924385FA",
INIT_2C => X"571D2E28E38E0216FA2D1E8E80140F45082B4002D082082AB8B6DBEDB7DF7F54",
INIT_2D => X"A97F7AF6D417E92482BF84020BA495557E3FF78E021FF1471FDEAAFFD56F16D5",
INIT_2E => X"7002FD74951D71EDFFABFD16FAAAE92BD5545A2DA3FB7DAAD4AAAAF487BC70BF",
INIT_2F => X"550A8010E00492487482FFFE82A85EBAE2FFC55554ADBD7A2FFC7BEFF6FFD7FC",
INIT_30 => X"400FBF9424F7000000000000000000000000000000000000000000000547AB8F",
INIT_31 => X"DF55F7AABFF55082CA8B4DF6C1E8F5E5400021EF005162BEF047FD5545AAFBF7",
INIT_32 => X"404547184164AA5D2EBEEB0A2D555410D3555714F8338AAAA1D0AE974AAF7FFF",
INIT_33 => X"AEABFFDF79DCBF755962010BDCBBC21455D7FEABEF75550ACBB7582225FF5843",
INIT_34 => X"D57D412F7D55F5E50C7F401BAAE8403CF5A3FFEAAEB083BC1000FF8409000512",
INIT_35 => X"2AA9FEAFDF7F431A9F7FFE81FF013A8001AFF801F8BA0C57740BDAA0688E5405",
INIT_36 => X"A2FBF7FED2C7F955445079E280A00C56145EF5D16BABAA3EBC3157ABD5FFE55F",
INIT_37 => X"0000000000596EBEF55080034E0A592A4AD00FB863550229BCABEB7DA403FFFD",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000100000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(1),        -- Port A data input
DOA(0)   => data_read_a_lo_256(1),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(1),        -- Port B data input
DOB(0)   => data_read_b_lo_256(1),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_2_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10E006600180111284380310006289800480032283E000A34301002001A0817",
INIT_01 => X"A14AC00A1079284D04A044A54E504368404000720885800802000006ECD10200",
INIT_02 => X"92250052A0348C310102048800A8507000040C8550200000480E0080001321E0",
INIT_03 => X"020204E4593C0824400C2220483042809292430400440180000890A4C9400242",
INIT_04 => X"486854B141002252142241502460480031B94420634850069A42241009610A04",
INIT_05 => X"800504244080892105AA6010A44882144840910A21220A8C820025E4A0000B00",
INIT_06 => X"A000442802280000340810209C444804206000AC800088096A0EA8C022208012",
INIT_07 => X"309820A848E0AA09826489A5CC49002001020112028201F8A20488260000108A",
INIT_08 => X"2400582881E0C1419D12041455509341A539C42A0D8208099002801700D10103",
INIT_09 => X"110D525861263100009200151409130A3C80C8C8096A06B8C12088400A9C2080",
INIT_0A => X"0451394CD0391A441583C04B580040089581001342801044877200D002A00DE0",
INIT_0B => X"144423040240450114901149013C9011C9013C9011C90134901144801A4808A5",
INIT_0C => X"D8A5345206D2C10082080A90C00000188150100C202A4640000E2B4081969420",
INIT_0D => X"050080400A0391A51240C480000AA902AA009028C83220008086952B4285A54A",
INIT_0E => X"05008021C00000000040000000020288000500000008000500802A0000000800",
INIT_0F => X"0002300000428000000040000000000D002A0000000800050080250000000800",
INIT_10 => X"0000000001204004000508000000100000000002054000130000000000800000",
INIT_11 => X"000C00000000000068144000000000001A000106200010021002000000000080",
INIT_12 => X"0002004A880000000000034098000000000000D024A000000000000001000900",
INIT_13 => X"00000000000000041400000A8000000000000000010A00000284000000000000",
INIT_14 => X"012100000002000280000000011080C000000000000000000000430000000260",
INIT_15 => X"A769DA769DA769DA368DA36CDA3A9A13A14801404134DA84A024024155000399",
INIT_16 => X"168DA769DA769DA769DA368DA368DA368DA769DA769DA769DA368DA368DA368D",
INIT_17 => X"68DA168DA169DA569DA569DA568DA168DA168DA169DA569DA569DA568DA168DA",
INIT_18 => X"138D70C030B51C50C7D000A2012F81F81F83F03F03F069DA569DA569DA568DA1",
INIT_19 => X"1041041041041041041041041041041041041041024860208165965975960040",
INIT_1A => X"25128944A25128944A25128944A25128944A25128944A2512894104104104104",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFF8421084210840703F25128944A25128944A25128944A",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"00000000000000000000000F0FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"415555087BFFF55A2AA800BAFFAE9540008002AA000000000000000000000000",
INIT_22 => X"7FE8B555551421455D0002145552EBFEBA007FC21EFA2FFD75EFAA8415410AA8",
INIT_23 => X"FFFE8B45552EBDF45FFAEAABFFF7FFE8B55F784155EFA2AEBDEAAA2FBEAABA5D",
INIT_24 => X"5D2AAAAAA5D2E820BAA2FBEAB5555557DF55A2AEBDF555D2E954BAA2AA974BAF",
INIT_25 => X"A5D04021EF557FC21FFAA8428BFFAAAA954AAAAAAAAAAAFFD1574105D7FFFF55",
INIT_26 => X"EFF7800215500557DF55AA80001FFAA80001550055575EFFF84021555D043DEA",
INIT_27 => X"B5500517DF555D042AA10A284154005D0015410085568A00FF80175FFA2D17DF",
INIT_28 => X"00000000000000000000000000000000000000005D00020AAAA80020AA082EAA",
INIT_29 => X"D55D2BE800042AFE8E1557D0075D2F45BEAA800AAFFAA9543A080038A2A00000",
INIT_2A => X"0BDEAAA2FBF8AAA557BE8B6D5D5FFABEF49040017D5D20B8EAA007FC51C7A2FB",
INIT_2B => X"0E174BFA02A974BAF7F5EFB455D2ABDF55492AA8BC7EBDFEAFEFFD00105FFBC2",
INIT_2C => X"3D155E105571D55D71C002DABA5524820BAB6FFEFB6D555578F7DB6A0BDF7D48",
INIT_2D => X"092A071555D5E3AE821D00001FF0871C016DBED1FDE90E3A497492B6AAADAAAE",
INIT_2E => X"0E3DA3DFD5E3DFFFBD5A38A021551C5F7AF6DBE8F401D7B6A0001470155C51D0",
INIT_2F => X"82B4002D082082AB8B6D1C5B7DF7FF78E075C5BE8555400550A38428007FED00",
INIT_30 => X"4AA00042AAA2000000000000000000000000000000000000000000000410F450",
INIT_31 => X"AAAA007FD5555AAFBD7545FBB8020A3F7AE975EF005560B55F7AA800AAF7AA95",
INIT_32 => X"E8F5EFF84165EFF7802BAB0A2FFEAABA557BEABEF057D68F5F5A00021EF55042",
INIT_33 => X"52ABFFFF841FFE75CA882108202E974AAF7D57DF55D7AABFF5428ACA8F45A6C1",
INIT_34 => X"84174A8FFAEBFEB0A2D55541051555694F002CA8AA80800020AAF7FBFFFEF045",
INIT_35 => X"7AAA155F595542455512A975455D3AA8A005500151FF0C57401E5F3D1E00A1A8",
INIT_36 => X"5D2A8A0B882FFFFE10AAAAAB755A66B6AF56A2AA801455D7FE8BFFF680800FFF",
INIT_37 => X"00000000000C3BC1000FF8409000512AEABFF5D79FCAF774AE005BE789555400",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000200000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(2),        -- Port A data input
DOA(0)   => data_read_a_lo_256(2),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(2),        -- Port B data input
DOB(0)   => data_read_b_lo_256(2),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_3_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"210C44A20020248B08431120001604B8156023104C4077133420400A02380202",
INIT_01 => X"015A2A424080216D3C2462C99E104B49404040028804A0080A000C16A0D90A0C",
INIT_02 => X"C0A4065000F0A95011000D1501005270B4045AB330860281CC08008222170060",
INIT_03 => X"AD22014098340394A4021320080841C40B411B4298042180002846B06900811A",
INIT_04 => X"244B32A86D20014A0D20403194904900071A24110F0BF400F85F92420E0C946E",
INIT_05 => X"80331030442898B4812840D0500008C528280B063006A64CA30004E5A4E40304",
INIT_06 => X"90016CA00E380042302040A0BC47160424428198C0038C89904E640023600816",
INIT_07 => X"1288020843A66620816049908AA0061011CA0142000009F0A810292E7402F088",
INIT_08 => X"20003C9984A0AC411102014D34EC2200214D5099048823019603A01A49410103",
INIT_09 => X"001CD74C4826220010A8891451284B661CA24A4C899046740121824004100080",
INIT_0A => X"44C9516DC0135C45159BE45F112B48804DC10203021290400772C0F402820D4C",
INIT_0B => X"B400624402404501A49018490184901A4901A4901849018C901A648056480C2D",
INIT_0C => X"D7A9B54000D7C10820680D08C420180381211081A022160000266723E1909021",
INIT_0D => X"400080200E199A4A2CA2994C0399981666409800CA52E4890806BD6B56BDAB52",
INIT_0E => X"40008008E00000000000000000024008000C8000000000400080028000000000",
INIT_0F => X"000A000000588000000000000000200400088000000000400080078000000000",
INIT_10 => X"0000001000004004000D800000000000000000022040000B4000000000000000",
INIT_11 => X"001A0000000000082006C000000000020804087220000122000A000000000000",
INIT_12 => X"00020800B8000000000041002E00000000001040466000000000000001020080",
INIT_13 => X"00000000000000048200004A600000000000000003008000320C000000000000",
INIT_14 => X"432900000222200871028000210400C4000000000000000000080200800030E0",
INIT_15 => X"AF6A5AF6A5AF6A5AF6A5AF6E5AFADA91AB68000101B4D20C08EC461733804A19",
INIT_16 => X"B6B5AF6A5AF6A5AF6A5AF6A5AF6A5AF6A5AB6B5AB6B5AB6B5AB6B5AB6B5AB6B5",
INIT_17 => X"6BDAB6B5A96ADAF6A5AD6ADAF6A5AD6ADAF6A5AD6BDAB6B5A96BDAB6B5A96BDA",
INIT_18 => X"C78C706428A14C586290008A044D54AAB556AA9556AAEBDAB6B5A96BDAB6B5A9",
INIT_19 => X"92492492492492492492492492410410410410412821600001249249015303C0",
INIT_1A => X"351A8D46A351A8D46A351A8D46A351A9D4EA753A9D4EA753A9D4924924924924",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000001543B351A8D46A351A8D46A351A8D46A",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"43DF55FFAA955EFA2D168B55557BEAA000055420000000000000000000000000",
INIT_22 => X"7BE8BFFA2D155410AA8415555087BFFF55A2AA800BAFFAE9554508002AA00AA8",
INIT_23 => X"52ABFEBA007FC21EF007FD75FFAA841541008002AB55AAAA955EF005568A0008",
INIT_24 => X"005168B455D042AB45F7FFD741000042AA10AAAABFF5508003FF555D00021455",
INIT_25 => X"0A2D1575FFF7AA975555D2E80145F78415545082EBDEAAA2FBEAABA5D7FC0155",
INIT_26 => X"55552A954BAFFFFE8B55552EBDE00F7AEAABFFF7FBEAB55F7AABDEBA5D7FC201",
INIT_27 => X"F55A2AEBDF555D2E954BA002EAAABA002A821EF5555554AA087BC01FFFFAAAAB",
INIT_28 => X"0000000000000000000000000000000000000000082E820BAA2FBEAB5555557D",
INIT_29 => X"95578080038A2AA28E3AF55E3A0BA5D7AADB6FB7D5D7FEAA3808554203A00000",
INIT_2A => X"0925D7085F6AA10087FEABD7AAD57AEBAB68E1557D1475FAF45BEAA800AAFFAA",
INIT_2B => X"04AAFFA41040017D5D20B8EAA007FC51C7A2FBD55D7BE80004AA1E8E2AB55B6A",
INIT_2C => X"2FBE80AA557BE8B6D5D5FFABEF49002FB55FFF5D0438140E2FA38B6AEBFF6D1D",
INIT_2D => X"AB8ABAE925D21C7010EADB525D7FFAE975C75D0A901FFFF801557D1C20B8EAAA",
INIT_2E => X"20875C21D5EB8AA8FFF012A954BAFFF5EFB455D20BDE00EBAAA8BC7EBDFEAFEF",
INIT_2F => X"BAB6FFEFB6D555578F7DB6A0BDF7DEB8E125FF002EADA921420871D74971D248",
INIT_30 => X"ABA0051400A20000000000000000000000000000000000000000000001C24820",
INIT_31 => X"8B55F7AA800BAF7AA955EF00042AAA2A2AEAAB55A28408145AAFFFFFFF5D7FEA",
INIT_32 => X"020A35D2ABEF55F7800015F087FEAA00007FEAB55FAD568AA2AFAE975EF55516",
INIT_33 => X"ABFEAAF7AE9DFF759A82AEF70800021EF55042AAAA007FD55558A7BD7145FBB8",
INIT_34 => X"84175EF55002AAB0A2FFEAABA557BEA3EF057968F575D003FF55F7D5420BA5D2",
INIT_35 => X"A8429F45A7D5EAF5FFBAEAAA10554155400AAFFD5145FBAC9755F05040255FFD",
INIT_36 => X"550415557085540000005156155FE90A8F5C082E974AAF7D57DF45552A3FF10A",
INIT_37 => X"00000000005500020AAF7FBFFFEF04552ABFFFF843FFE77C80825BC052ABFE10",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000100000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(3),        -- Port A data input
DOA(0)   => data_read_a_lo_256(3),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(3),        -- Port B data input
DOB(0)   => data_read_b_lo_256(3),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_4_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"A108400020612C80284210081034849800A000303100048B3432C82904204002",
INIT_01 => X"21066802000820491C00650E1E004360403008418984014902030906A8D10200",
INIT_02 => X"120404E00E4C0600000206100008402005040C00F104008040080080001310E0",
INIT_03 => X"DCA201514D1C0D706C5CF010083A0708BA0841945004010000080084C1000002",
INIT_04 => X"5C4CF21C48B133483C80417570D000083A62488074C1350EA60D785C0A6B0619",
INIT_05 => X"000F0400028083B381A60001E5546EB5C0E2B81E4166DE000139200004E50940",
INIT_06 => X"80004408020800023000102098000204A040038600018019004B800123208806",
INIT_07 => X"120C20204665E1008024188488800000001A01520000A1F08044892400001088",
INIT_08 => X"0801007AC0A1EB413102063CF3E0B3028D29F407059B0B000205A801C2200102",
INIT_09 => X"106052400922D00406BE1002C6150F41200280001900439001FD8A0004142000",
INIT_0A => X"047F2201D899BA503583504B58AB80804540001202805544314041B48A888EC5",
INIT_0B => X"1441E3443043410C5010C3010C1010C3010C1010C1010C3010C14086980861A5",
INIT_0C => X"020000A02600000805400502C0A0004A00625015000A12000026E1E180011220",
INIT_0D => X"400000000E43930C20C20188120782861E4004A800600401A030001008080400",
INIT_0E => X"40000021A8800000000000000000400800170024000000400000310024000000",
INIT_0F => X"0008000000AA80200800000000002000003400240000004000003B0024000000",
INIT_10 => X"00000010000000040004A080000000000000000020400006C008020000000000",
INIT_11 => X"002C008200000008001B4020200000020000090760000200110A040010000000",
INIT_12 => X"00000803E004040000004000E801040000001000086000000000000000020040",
INIT_13 => X"0000000000000000810000164001008000000000020040002240008020000000",
INIT_14 => X"04001040026026004000000002940040000410000000000000080000400000B8",
INIT_15 => X"040080201004008060000001806AC000004890015124D880100886D8F0014420",
INIT_16 => X"4010000180600000018020100400802010000080601000008020000401802000",
INIT_17 => X"0100000004008020180600000000000180600802010000000401802018020000",
INIT_18 => X"3807E05000140634504048820064B261934D964C326980004010000080600806",
INIT_19 => X"AAAAAAAAAAAAAAAAAAAAAAAAAAA28A28A28A28A2934C8D0CCD145144C0A28A06",
INIT_1A => X"068341A0D068341A0D068341A0D068351A8D46A351A8D46A351AAAAAAAAAAAAA",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000000173F068341A0D068341A0D068341A0D",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"57FE10FFFBEAA10007FD7410FFAA97555082A800AA0000000000000000000000",
INIT_22 => X"7FEAA00007BE8AAAAA843DF55FFAA955EFA2D168B55557BEAB45005542000005",
INIT_23 => X"87BFFF55A2AA800BAFFAE9555508002AA000055574105D2A800AA00043FEBA5D",
INIT_24 => X"A2D17DE1000517FE10AAAAA8AAA002E97545557BC00AAA2FFEAAAAAA84155550",
INIT_25 => X"0A2D157400AAAE974AAAAAA974BA08002AB55A2AA955EF005568A00087BE8BFF",
INIT_26 => X"BA080002145552ABFEAA007FC21EF007FD75FFAA8417410A2D140000F7FBC201",
INIT_27 => X"A10AAAABFF5508003FF55F7D568A00552EA8BEFA2AABDEAA087BEAAAAA2FBD54",
INIT_28 => X"000000000000000000000000000000000000000055042AB45F7FFD741000042A",
INIT_29 => X"EAB7808554203A145178E00FFFBE8A101475D5400F7A49057D0824850B800000",
INIT_2A => X"E8008200043FE925571EFA380871C7028A28E3AF55F7A0925D7AADB6FB7D5D7F",
INIT_2B => X"F5FDA38BE8E1557D1475FAF45BEAA800AAFFAA9557D080038AAA145157428492",
INIT_2C => X"85F6AA10087FEABD7AAD57AEBA08517DE00AAAEA8A9200249056D4175C5092AA",
INIT_2D => X"FEDB42028EBFBC2028BED152438AAA092492AAA4954281C0E2FB55B6A0925D70",
INIT_2E => X"A0875EDA80BEF1C743840040017D5520B8EAA007FC51C7007BD55D7BE80004AA",
INIT_2F => X"55FFF5D0438140E2FA38B6AEBFF6DBE84AAEBAF7DF6AA00412EAABFFAA803DEB",
INIT_30 => X"1EF0800154B200000000000000000000000000000000000000000000041002FB",
INIT_31 => X"0145AAFFFFFEF5D7FEABFF0051400A25D5568A00FFFFEAA105D5155410FF8402",
INIT_32 => X"2AAA25555410BA082E8201000043FE005D517DEBA0851574B2AAAEAAB55F7840",
INIT_33 => X"4001FF005575408AA557FEB2FFAE975EF555168B55F7AA800BAF7AA955EF0004",
INIT_34 => X"2ABFF55F7800015F087FEAA00007FEAB55FAD568AA200557DE00AAAAAAA00080",
INIT_35 => X"87BD6145FAAC000A2A6FBC00BAAAFBC00BAF7D1550AAAA8002010F2AC154B25F",
INIT_36 => X"082EA8BFFAA843FEBA08517DE00F3F9574B30800021EF55042AAAA007FD55550",
INIT_37 => X"000000000008003FF55F7D5420BA5D2ABFEAAF7AEBDFF779A82AA43F7FBE8A00",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000200000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(4),        -- Port A data input
DOA(0)   => data_read_a_lo_256(4),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(4),        -- Port B data input
DOB(0)   => data_read_b_lo_256(4),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_5_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50DF4A0791B3FCB694379283C81FD996A091832102004A337A20E07C0C1E006",
INIT_01 => X"294014468000A04D5C6A60000C34C24841280A00084000C8C212892EEAD53235",
INIT_02 => X"50AE41540CA1D9100002171C1F0A5171134E2A200D8633F8CD09DBFBBB970E7C",
INIT_03 => X"214E3C521D16021B64430CC51C45B8154689094241898749920842946B90010A",
INIT_04 => X"A2F20F7D7A314CB5C208E28A1BF0224A448920028A185340D0C20B2690000C22",
INIT_05 => X"7520B430B20B984809A8886E230C6106371146E1829941C58310402C600381CF",
INIT_06 => X"9CC96CD7C63A7495B9A356ACBC4601C57FD44F8549A46490261C4B39203F7080",
INIT_07 => X"12A88800B029E0C0A12C4B92AA36A2111167357C220095F3C8952A2E5D26F078",
INIT_08 => X"F3F00503B4AE105B534711820C0C0A1043080300F7E0E728B1829C2FEA0A95A1",
INIT_09 => X"C5184F084136848C9298A8560688F480C58858449026145B3830F40944906234",
INIT_0A => X"50EB4124D2B3902BF5C9700C1199DCA84DF46A974F92C7E28F1630D38088A438",
INIT_0B => X"B3144E5636E3178C86B8CC6B8CA6B8CE6B8C86B8CE6B8CA6B8CC15C6435C670C",
INIT_0C => X"79E51E70E070AA8132252008360A7E91504104C8948047D6B0AE1FE440B28A71",
INIT_0D => X"05F0FE40014090400400080329FF8089FF49611F589765923E139F09C78CE7C6",
INIT_0E => X"05F0FE64037FFD7857418407157797878F005F0DFF0F8005F0FE205F0DFF0F80",
INIT_0F => X"8F87FCB1F8053FDEB9B34E0700461E5FF8205F29FF0F8005F0FE205F29FF0F80",
INIT_10 => X"C0184D07C1FF55C3E3E0037FFCF8D3C03009C3CFD53C7E001FF2FAF89781C011",
INIT_11 => X"4E0CDF47186104C6FF177BD939024189BF900401165D645CEEF5BBCDF148F980",
INIT_12 => X"6397F64AEF7F2320483137F8A9BF8A30C2098DFCA06FFFE01F80001F81FDC94F",
INIT_13 => X"FFD051E01015C3BF553D3E0E5FFE838381840714F9DB4F4FA213F774A0E07002",
INIT_14 => X"8B652E2B3120C81284641D3E8DBF7D636FE070189500125C1F83FBCC4F4F80EF",
INIT_15 => X"E7394E339CE138CE5394E33D4E1E0E30E1208C251134921C12A44103F064014B",
INIT_16 => X"7384E3394E338CE538CE1394E3384E738CE139CE1394E7384E339CE139CE5384",
INIT_17 => X"38CE139CE1384E7384E7394E3384E738CE539CE139CE538CE5384E3394E7384E",
INIT_18 => X"7F7B9DB7FF3A1B6DB7ED438A9C3124B2DA6924965B4D384E7384E339CE138CE5",
INIT_19 => X"FBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEF9F7CFDFDDCF3CF3DF5E5BB4E",
INIT_1A => X"7BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEFBEFBEFBEFBE",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE000000000000118D27BBDDEEF77BBDDEEF77BBDDEEF7",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"E955450055421FFFFFBC0010AAD5574BA557FFDFFF0000000000000000000000",
INIT_22 => X"D5575EF55517FF5500557FE10FFFBEAA10007FD7410FFAA97410082A800AAAAA",
INIT_23 => X"FAA955EFA2D168B55557BEAB55005542000007FD74000055574BA5D7FD7555A2",
INIT_24 => X"007BC00AAAAAEBDF45A28428B45FFD168BFF00002AABA5D2ABFFFFAA843DF55F",
INIT_25 => X"AFF80174BAAAD1555EF5555555550055574105D2A800AA00043FEBA5D7FEAA00",
INIT_26 => X"FFAA8415555087BFFF55A2AA800BAFFAE95555080028A00A2FFFDE00F7D57FEB",
INIT_27 => X"545557BC00AAA2FFEAAAA082A97545F7D5420BA5D2E821FFA2D5554BA557BD75",
INIT_28 => X"000000000000000000000000000000000000000000517FE10AAAAA8AAA002E97",
INIT_29 => X"9043D0824850B8A2AE9756D145B401FFFFFFC7010BEDF524AA5571FDFEF00000",
INIT_2A => X"1524BA5571D757DB6D5525EF555178F6D145178E00EBFBE8A101475D5400F7A4",
INIT_2B => X"24BFFFFA28E3AF55F7A0925D7AADB6FB7D5D7FEAB7D0855420BA1471D7438085",
INIT_2C => X"0043FE925571EFA380871C7028B6AEBDF45B68A28B6DEBDF6DBEF1C0A28AAA55",
INIT_2D => X"A2FBF8E10EBD578EAAFF8415482BED1555EF55555057D145152428492E800820",
INIT_2E => X"FB6DF574A85575C55EFBE8E1557D1475FAF45BEAA800AAFFAA9557D080038AAA",
INIT_2F => X"00AAAEA8A9200249056D4175C50920875FDA381C209256DFFDF420BA552A821F",
INIT_30 => X"0BA55557DFF700000000000000000000000000000000000000000000008517DE",
INIT_31 => X"AA105D5155410FF84020AA0800154B2AAAA975FF5D7BC21EFF7FBD7400F7FBC0",
INIT_32 => X"400A25551554BA0051400BA5551575EFF7D1401FF5D5568BE7555568A00AAFFE",
INIT_33 => X"FFDFFF552EA8AAA55043DFF7AAAEAAB55F78400145AAFFFFFEF5D7FEABFF0051",
INIT_34 => X"55400BA082E8201000043FE005D517DEBA0851574B2FFAABFF45FFAAAABFFAAF",
INIT_35 => X"7AA955EF00002AAA2A2FBE8A00A2D16AAAAFF8002410FFD5575EF5555421E755",
INIT_36 => X"FFFFC00BA552A821EFFFFFD74BA5D51575F7FFAE975EF555168B55F7AA800BAF",
INIT_37 => X"000000000000557DE00AAAAAAA000804001FF0055554088A557FEB25D00021FF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000C00000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(5),        -- Port A data input
DOA(0)   => data_read_a_lo_256(5),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(5),        -- Port B data input
DOB(0)   => data_read_b_lo_256(5),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_6_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10800B0061A01002840002C03002818000402322520070B313301C4389B2082",
INIT_01 => X"274008482009404C18A160000C52424841000000090800090210000008510200",
INIT_02 => X"102430600C800110000006100009D070012408000000000648080000001210E0",
INIT_03 => X"000200501D1D02140C420200480140040608010040400104681A0084490C4802",
INIT_04 => X"404402820021000A00824002141000980500000808001114C000080624600600",
INIT_05 => X"120024204209981001A806500304610528000500000080000000300000012940",
INIT_06 => X"2000440832280002300010209C4400142061207A024008900008000220600220",
INIT_07 => X"130C8A220FF41F00902008808800182001020150000001F0800408264000100A",
INIT_08 => X"001BF002C4A01041B1120101000010128568837F04842B080020890008080342",
INIT_09 => X"011847140126805432A62A1596C8B5DF10000008900000100220C00084000008",
INIT_0A => X"44EB4104D09392053589F11C59898888454010830212C54081000410A0088C00",
INIT_0B => X"B0044245B25B456C0096C0096C4096C4096C2096C2096C6096C444B6004B600C",
INIT_0C => X"09040020280010000B3002820110101D0012402CC00802410C26800860070621",
INIT_0D => X"0500819D0000900208201040C4007920004884080000448C281018100C000200",
INIT_0E => X"05008182100000000000000000022AE800C00004000000050081A00004000000",
INIT_0F => X"0002330006000000080000000000000D07A00020000000050081A00020000000",
INIT_10 => X"0000000001204A340002100000000000000000020F4001400000020000000000",
INIT_11 => X"019300020000000068D08000200000001A692121000280000000000010000000",
INIT_12 => X"000201FA100400000000034696010000000000D3478000000000000001003F00",
INIT_13 => X"00000000000000043C0001C0A000008000000000012E000054AC000020000000",
INIT_14 => X"0200000040A410C2810800016000809400001000000000000000433300007600",
INIT_15 => X"060180400000008060180404002AC0200208940041309210B28048180F028000",
INIT_16 => X"2008000100601802000000100601800000000180600800000020180600000000",
INIT_17 => X"0180600000008040100200800000060100000802010040180200002018040100",
INIT_18 => X"7F8FF0F4FA955F7CF7F40A80907638C31C71C718638E00006018040080200004",
INIT_19 => X"38E38E38E38E38E38E38E38E38E38E38E38E38E39B6CEDECDDF7DF7DF5F78BCE",
INIT_1A => X"3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE38E38E38E38E",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFF000000000000196A03F9FCFE7F3F9FCFE7F3F9FCFE7F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"00000000000000000000000C0FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"BFDF45F7AA974AAAAAA97555F784174BAF7D5555FF0000000000000000000000",
INIT_22 => X"FBD7410AA8428AAAAAAE955450055421FFFFFBC0010AAD5574BA557FFDFFF087",
INIT_23 => X"FFBEAA10007FD7410FFAA97400082A800AA08515555508043FE00F7AA97555A2",
INIT_24 => X"55517FF55A2AA97400552AAAB45082E80155F7D1575EFFFAA9555500557FE10F",
INIT_25 => X"FF7AAA8A10082EAAB45A2FFC2000007FD74000055574BA5D7FD7555A2D5575EF",
INIT_26 => X"FFAA843DF55FFAA955EFA2D168B55557BEAB5500554200000003DE10FFD5401F",
INIT_27 => X"BFF00002AABA5D2ABFFFF087BD5545007BFDE10AA803FE105D516AABAFF843FF",
INIT_28 => X"0000000000000000000000000000000000000000AAAEBDF45A28428B45FFD168",
INIT_29 => X"524AA5571FDFEF1C7BFFF55FFA095482B6A49256DEB84104BAFFD1525FF00000",
INIT_2A => X"03DE28F7A49057DAAF5D2428A2842AAAAA2AE9756D145B401FFFFFFC7010BEDF",
INIT_2B => X"A49756D145178E00EBFBE8A101475D5400F7A4904380824850381C5B5057D1C0",
INIT_2C => X"571D757DB6D5525EF555178F6DAAA495428412AAFB451C2A8017DE3DF525FFFF",
INIT_2D => X"1C0E3FE00E3DB471EFE3AAAAA00082EA8B6DA2F1C50381471D74380851524BA5",
INIT_2E => X"049516AAB8FF8428FEFA28E3AF55F7A0925D7AADB6FB7D5D7FEAB7D0855420BA",
INIT_2F => X"45B68A28B6DEBDF6DBEF1C0A28AAA5524BFFFF1C7BD057D1C71FFE10A28038E1",
INIT_30 => X"0AAFFD1401E7000000000000000000000000000000000000000000000B6AEBDF",
INIT_31 => X"21EFF7FBD7400F7FBC00BA55557DFF7557BFDF55F78017400F780001FFAA8400",
INIT_32 => X"154B2557FC01EF55043FEAAFF80021EFA2D1420BAAA8428AA2AAAA975FF5D7BC",
INIT_33 => X"A821EFAAFBC01FFF780155F7555568A00AAFFEAA105D5155410FF84020AA0800",
INIT_34 => X"51554BA0051400BA5551575EFF7D1401FF5D5568BE7AA80174AA082ABDF555D2",
INIT_35 => X"D7FEABFF0051400A25D2EBFE10AAFFD55EFA2AEA8A10082EA8BEFAAD5554B255",
INIT_36 => X"55557DE00AA842AA0000516AABAFF8428BE7AAAEAAB55F78400145AAFFFFFEF5",
INIT_37 => X"0000000000FFAABFF45FFAAAABFFAAFFFDFFF552EA8AAA55043DFF7557BC01EF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000900000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(6),        -- Port A data input
DOA(0)   => data_read_a_lo_256(6),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(6),        -- Port B data input
DOB(0)   => data_read_b_lo_256(6),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_7_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10844B00482258A2842112C02450418800002300500030B313300C418992002",
INIT_01 => X"234008422008604D1C20E0000E11426840000000080000080200090000110204",
INIT_02 => X"1025207000B08910000206101188D03080144880010400044808000000122160",
INIT_03 => X"000200401914821004420000CA01000C0600010000605114291A008449484802",
INIT_04 => X"40440200002100080006500210101019040000000B085024D842080244000000",
INIT_05 => X"1A8024200009981001A8224001040104200204000000800CC2092CE4A0004900",
INIT_06 => X"A000440822280002340010209C040014A061200052500810000C490323208E28",
INIT_07 => X"128802020028000890240980A809102001020140000009F0800408264000100A",
INIT_08 => X"001A0602C4A01051B13281010408881203480200448423199046821008082351",
INIT_09 => X"336784144126811054809C1040140A001C8648481000045903318B80A400310A",
INIT_0A => X"000800009010100014114110312388984502148282A08415B032095048008100",
INIT_0B => X"20CDC1C483484D201192011920119201192051920519205192074C9018C90188",
INIT_0C => X"D8A5B44001D2C12901228F82F005310D293054048A2212004466000DA1908528",
INIT_0D => X"800F8108A0D09802082010408580008000000008C85264010816851B428DA146",
INIT_0E => X"800F81321000020000261900E28A204040E000A0000007800F814000A0000007",
INIT_0F => X"7072024807000020400000581C01C1A406400084000007800F81400084000007",
INIT_10 => X"060180E83800E820101210000200000CC3003C32080201C0000C000000160700",
INIT_11 => X"81DD00804086423120B74020023090644840A34000828800000004000420020B",
INIT_12 => X"1C6A0186E8000446120C8905BA0004810C84624237E00010001878007F0030C0",
INIT_13 => X"00080208E4083C44230201AEE0010040261900E30520C0806EAC0082000984C0",
INIT_14 => X"0121011088A600C032128201519480D40005802448160403E0700622C0806EE8",
INIT_15 => X"A1685A1685A168DA368DA36CDA30DA13A108810111349A943AA4401000928A19",
INIT_16 => X"368DA768DA1685A1685A5685A368DA368DA7685A1685A1685A768DA368DA368D",
INIT_17 => X"685A1685A169DA368DA1685A1695A368DA3685A1685A168DA368DA1685A1685A",
INIT_18 => X"00000000000000000000400A8448410400020820800069DA1685A168DA369DA3",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000003667B000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"0155EFAAAEA8ABAAAFBFDE0055556AA005D04155550000000000000000000000",
INIT_22 => X"556AA00FFAE95555087BFDF45F7AA974AAAAAA97555F784174BAF7D5555FFF78",
INIT_23 => X"055421FFFFFBC0010AAD5574BA557FFDFFF5555555EFAAFFFDFEFAAAAAAB455D",
INIT_24 => X"AA8428AAA557BFDFFF55003DFFFF7FBEAA00002EAAAAA082EA8A00AAAE955450",
INIT_25 => X"0552EBDE00007BEAAAAA2D14000008515555508043FE00F7AA97555A2FBD7410",
INIT_26 => X"FF00557FE10FFFBEAA10007FD7410FFAA97400082A800AAF7AE975FFA2800001",
INIT_27 => X"155F7D1575EFFFAA955555D51574AAAAFFD5545087FEAB455D516AB55557BD55",
INIT_28 => X"0000000000000000000000000000000000000000A2AA97400552AAAB45082E80",
INIT_29 => X"104BAFFD1525FFFF8E175C7A2AAAAA82A2F1FAE105D556AA10410E1755500000",
INIT_2A => X"1FFFD7AAAAAFB7D495F6AA10E3AE905551C7BFFF55FFA095482B6A49256DEB84",
INIT_2B => X"2EAAA00A2AE9756D145B401FFFFFFC7010BEDF524AA5571FDFEF415B575D7AAF",
INIT_2C => X"7A49057DAAF5D2428A2842AAAA497BFAFFF49003AFEFEBFBEAA001C2EA8A821C",
INIT_2D => X"F7A4905C7A28A070384120BDE100075EAA82BEDB470101C5B5057D1C003DE28F",
INIT_2E => X"D555F6AB57417BC05D7145178E00EBFBE8A101475D5400F7A490438082485038",
INIT_2F => X"28412AAFB451C2A8017DE3DF525FFFFA49756D495150492BEF1D2555087BE8B7",
INIT_30 => X"A10002E9754D000000000000000000000000000000000000000000000AAA4954",
INIT_31 => X"7400F780001FFAA84000AAFFD1401E7FFAA97555A2AEA8A10AAD568A00555168",
INIT_32 => X"7DFF7007BD5555AAD57DF55AAAEBDFEF007BE8A10AAAE8215D557BFDF55F7801",
INIT_33 => X"FEAA105D2EAAA005D2AAAA18AAAA975FF5D7BC21EFF7FBD7400F7FBC00BA5555",
INIT_34 => X"7FC01EF55043FEAAFF80021EFA2D1420BAAA8428AA2007FE8BFF080028BFFAAF",
INIT_35 => X"F84020AA0800154B2FF8402145A2AA954AA00043DE0000516AA10F7FBD740855",
INIT_36 => X"FFD140145007FE8BEF557BEAB55087FC215D555568A00AAFFEAA105D5155410F",
INIT_37 => X"0000000000AA80174AA082ABDF555D2A821EFAAFBC01FFF780155F7005140000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000000FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(7),        -- Port A data input
DOA(0)   => data_read_a_lo_256(7),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(7),        -- Port B data input
DOB(0)   => data_read_b_lo_256(7),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_8_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00000648E2840112C00000418000002700500030B3132000400812086",
INIT_01 => X"214009C21838284D042100000212026840000000180800080200080040510204",
INIT_02 => X"1021004000900110000006100088503000240800014400004808000000122160",
INIT_03 => X"0002004019110214044A82000121400C86000000000000860188008448400002",
INIT_04 => X"000402800031200A0000090214100889A5000000490090104800000224000400",
INIT_05 => X"10C025204289981000A820500344010428008500010080080909304040202004",
INIT_06 => X"8000440003280000340010208C04003420600000C6180810000C490703200010",
INIT_07 => X"130002000028000890240980A809012001020050000009F08004082640000082",
INIT_08 => X"20100402C4201041310041010008801201480200051023090024811008090A1A",
INIT_09 => X"0100001001248100308214528148A48008000008100004590711C04034000083",
INIT_0A => X"10804000801210140001C0103001088845010482004000008420041020008900",
INIT_0B => X"0004404002004400448000480004800048000480004800048000440022400200",
INIT_0C => X"880420000880204909004502D100A10C04205424010216010C26800805000004",
INIT_0D => X"8000801100509802082010400400018000488428800004082014000200010000",
INIT_0E => X"8000800A00000207A8BE7B00000200082040808000F07F80008000808000F07F",
INIT_0F => X"0002000402100000404CB1F8FC0000040000808000F07F80008000808000F07F",
INIT_10 => X"3E07800000004004080A000002072C3FCF0000020040804800040007687E3F00",
INIT_11 => X"10800018639EC00020100002C2F9B0000801016001008100000040120CB3067F",
INIT_12 => X"000200020000585EB6000100800030C73D8000402000001FC07FF80001000080",
INIT_13 => X"002EAE1FEC0000040200408000003C547E7B00000100801004000803551F8FC0",
INIT_14 => X"00000000440610C8000A808040000208901B86E568FE0C000000020080100400",
INIT_15 => X"0040100401004090240902449028D0230249850101349A98BAC0481000888810",
INIT_16 => X"0401004010040100401004010240902409024090240902409004010040100401",
INIT_17 => X"4010040100409024090240902409004010040100401004090240902409024090",
INIT_18 => X"543EBC57A10A1E75D6440A889050000000000000000040902409024010040100",
INIT_19 => X"79E79E79E79E79E79E79E79E79E79E79E79E79E7BF3CCD8DF5B2DB2CA4028A0A",
INIT_1A => X"4F87D3E1F4F87D3E1F4F87D3E1F4F87C3E1F0F87C3E1F0F87C3E79E79E79E79E",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000000D3E94F87D3E1F4F87D3E1F4F87D3E1F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"000000087BEAA10F7803DE00FFAEBFFFF0800155FF0000000000000000000000",
INIT_22 => X"7FC2145005155555F780155EFAAAEA8ABAAAFBFDE0055556AA005D0415555080",
INIT_23 => X"7AA974AAAAAA97555F784174BAF7D5555FF552AA8AAA557FC0010F780154105D",
INIT_24 => X"FFAE95555AAFFE8A00552EBFE00F7D17FF45F7FFFFF55AA80155FF087BFDF45F",
INIT_25 => X"5F7D140010552E821EFAAAABDF555555555EFAAFFFDFEFAAAAAAB455D556AA00",
INIT_26 => X"00AAAE955450055421FFFFFBC0010AAD5574BA557FFDFFF5504000AAAAAAA8B5",
INIT_27 => X"A00002EAAAAA082EA8A00002AA8A10F78402155AA8028A00A2D57FF45557BE8A",
INIT_28 => X"0000000000000000000000000000000000000000557BFDFFF55003DFFFF7FBEA",
INIT_29 => X"6AA10410E17555080E000280071E8A00EB8E3FE10F7AEBAFFF080A175D700000",
INIT_2A => X"1C2000FF8A17400557FC015514555757DFF8E175C7A2AAAAA82A2F1FAE105D55",
INIT_2B => X"8A105D71C7BFFF55FFA095482B6A49256DEB84104BAFFD1525FF492EA8AAA557",
INIT_2C => X"AAAAFB7D495F6AA10E3AE90555A2FBE8A38492ABDE10EBDF7AF6DE3FFF8F7DB6",
INIT_2D => X"550E00082B6A0AFB55F7D1420104124821D7AAA0BDF6D415B575D7AAF1FFFD7A",
INIT_2E => X"0B6D578F6D557FFDA00A2AE9756D145B401FFFFFFC7010BEDF524AA5571FDFEF",
INIT_2F => X"FF49003AFEFEBFBEAA001C2EA8A821C2EAAA001C2EA8A00F7800017DA2842FA0",
INIT_30 => X"BEF082E95545000000000000000000000000000000000000000000000497BFAF",
INIT_31 => X"8A10AAD568A00555168A10002E9754D082E820BA08556AA00AAAABFE00F7AEAA",
INIT_32 => X"401E7082EAAABA5D5140010F7AE974105D7BC21555D51575EFFFAA97555A2AEA",
INIT_33 => X"BEABFFAAFBEABFFF7AA80145557BFDF55F78017400F780001FFAA84000AAFFD1",
INIT_34 => X"7BD5555AAD57DF55AAAEBDFEF007BE8A10AAAE8215DA2FFE8ABA082ABFE00AAF",
INIT_35 => X"7FBC00BA55557DFF75D2E82010F7843DF45FFD540000000402145AA843FFFF00",
INIT_36 => X"F780021FFA2803DE10FFD16ABFF5D7BFDE10AAAA975FF5D7BC21EFF7FBD7400F",
INIT_37 => X"0000000000007FE8BFF080028BFFAAFFEAA105D2EAAA005D2AAAA185D2AAAA10",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000400000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(8),        -- Port A data input
DOA(0)   => data_read_a_lo_256(8),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(8),        -- Port B data input
DOB(0)   => data_read_b_lo_256(8),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_9_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000B0001800002840002C0000281800000030000000033022000000000002",
INIT_01 => X"8000098218302849180060000C004240413C0A61590001D90213C90008510200",
INIT_02 => X"000008700CB089100002061031200074810448800104008048080080001210E2",
INIT_03 => X"000200140C1822000A028010408100000628000140402080041A100040024840",
INIT_04 => X"41040000000400080002040200080800040000000B08D1055842080604600700",
INIT_05 => X"10002024000020102400010000026104200004000400800C8B0024E4E0010C40",
INIT_06 => X"8000440802280002700800008A840004A0610000C0000810000C590103600810",
INIT_07 => X"538600220028001890240980A80800200102025000000BF08200002440000883",
INIT_08 => X"00000402C220104131102101040810028528820005100003900E884000010007",
INIT_09 => X"00000005E000000600BCA284140200800C834948100004590111824404012080",
INIT_0A => X"04080000901012100A1141005922000245410002008880000032005080000800",
INIT_0B => X"2000020040044010440104401004010440100401044010040104400802008208",
INIT_0C => X"D1A1344420D2E100000808000000000481000000202002400006800825908402",
INIT_0D => X"0500000000109000000000000580008000080000C852240100068D0B4685A342",
INIT_0E => X"0500000A00000000000000000000028000408020000000050000208020000000",
INIT_0F => X"0000304002100020000000000000000900208004000000050000208004000000",
INIT_10 => X"0000000001200000000A00000000000000000000050000480008000000000000",
INIT_11 => X"009F0080000000004807C0200000000012000020000081000000040000000000",
INIT_12 => X"00000048F8000400000002403E0004000000009067E000000000000000000900",
INIT_13 => X"0000000000000000140000CEE001000000000000000A000036AC008000000000",
INIT_14 => X"03210000000400CA81000000619480D4000400000000000000004100000036E8",
INIT_15 => X"A368DA368DA3685A1685A1685A121A11A1419001512490040024001000008019",
INIT_16 => X"1685A1685A1685A1685A1685A368DA368DA368DA368DA368DA368DA368DA368D",
INIT_17 => X"685A1685A168DA368DA368DA368DA368DA368DA368DA3685A1685A1685A1685A",
INIT_18 => X"CCF48DE68A895C38E250080000000000000000000000685A1685A1685A1685A1",
INIT_19 => X"514514514514514514514514514D34D34D34D34D28E10040392482090157344C",
INIT_1A => X"4D268341A0D069349A0D069349A0D068341A0D068341A0D06834514514514514",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000001654D0D069349A0D068341A4D268341A",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"BE8B45002A974AAAA803DFFFAA843DF45FFFFEAABA0000000000000000000000",
INIT_22 => X"AEBDE00AAFBEAABA080000000087BEAA10F7803DE00FFAEBFFFF0800155FFAAF",
INIT_23 => X"AAEA8ABAAAFBFDE0055556AA005D0415555087BFDE00A2FBD7400F7FBFDFFFA2",
INIT_24 => X"005155555557BE8BEF007FFDEAAAAD1555EF0055401FFF7AEAAA10F780155EFA",
INIT_25 => X"0F7AA974AA082E80010A2AAAAA10552AA8AAA557FC0010F780154105D7FC2145",
INIT_26 => X"BA087BFDF45F7AA974AAAAAA97555F784174BAF7D5555FFF780154AA5D2AA8A1",
INIT_27 => X"F45F7FFFFF55AA80155FF080400145FFFBEAABAF7D17FEBAA2AEBDF45002EAAA",
INIT_28 => X"0000000000000000000000000000000000000000AAFFE8A00552EBFE00F7D17F",
INIT_29 => X"BAFFF080A175D7BEF1E8B6D002090482B68E38FC7BE8A3DF7DF7F5E8A9200000",
INIT_2A => X"BD0400FFF5FDFC7B6A0BDE38B6F5E8A92080E000280071E8A00EB8E3FE10F7AE",
INIT_2B => X"AAA8A38FF8E175C7A2AAAAA82A2F1FAE105D556AA10410E175550871FFE00A2F",
INIT_2C => X"F8A17400557FC015514555757D5D71E8BEF147BFAE82A2DB555C71C5B451D7FF",
INIT_2D => X"FF84174BA5D20AAA00E3AA904BA142A87010A2AEADA38492EA8AAA5571C2000F",
INIT_2E => X"AAAA0BFF7D0024ADA921C7BFFF55FFA095482B6A49256DEB84104BAFFD1525FF",
INIT_2F => X"38492ABDE10EBDF7AF6DE3FFF8F7DB68A105D7000400155FFFBEDA82FFD57DEB",
INIT_30 => X"FEFF7D16AA00000000000000000000000000000000000000000000000A2FBE8A",
INIT_31 => X"AA00AAAABFE00F7AEAABEF082E95545F7D568BEF080402000F7AAA8B55FFAABD",
INIT_32 => X"9754D00517DE00A2FFC2000F7D17FF55FF803FEAAFFD16AA00082E820BA08556",
INIT_33 => X"FD55555D7FD5555FFAAA8AAAFFAA97555A2AEA8A10AAD568A00555168A10002E",
INIT_34 => X"2EAAABA5D5140010F7AE974105D7BC21555D51575EF555568BEF5D7FE8A10AAF",
INIT_35 => X"A84000AAFFD1401E7FF80174AA5D0028A00AAAE800AA552A97400A2AEBDEAA08",
INIT_36 => X"F7FBFFE00FFD17FEAAA2803DFEF08043FE00557BFDF55F78017400F780001FFA",
INIT_37 => X"0000000000A2FFE8ABA082ABFE00AAFBEABFFAAFBEABFFF7AA80145080002145",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000800000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(9),        -- Port A data input
DOA(0)   => data_read_a_lo_256(9),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(9),        -- Port B data input
DOB(0)   => data_read_b_lo_256(9),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_10_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000B0001800002840002C0000281800020030000000033022000000180006",
INIT_01 => X"000008000000004C002000000010026840000000080000080200000000110200",
INIT_02 => X"0000004000800110000006100000003000040800010400004808000000120060",
INIT_03 => X"000200000810020000020000400100000600000000400000001A000040004800",
INIT_04 => X"0004000000000008000200020000000004000000080010004000000200000000",
INIT_05 => X"1000202000011010000000000000010520000400000080000000200000200004",
INIT_06 => X"80004408022800023000000088040004A061000040000810000C490103600000",
INIT_07 => X"120420020028000890240980A808002001020050000009F08000002440000082",
INIT_08 => X"00000402C0201051311001000000020201080200440400000000800000000000",
INIT_09 => X"0000105808000000000000000000008000008088100004590111800004000000",
INIT_0A => X"00804000801210440003C1411008800045000002000014000040009002800000",
INIT_0B => X"0400200000000000000004000040000000000000040000400000000000000221",
INIT_0C => X"0100802000000000000002802000000400100000000002000026000840011400",
INIT_0D => X"0500000000409002082010400400008000400008002044082000081004080204",
INIT_0E => X"0500000200000000000000000000028000400000000000050000200000000000",
INIT_0F => X"0000304002000000000000000000000900200000000000050000200000000000",
INIT_10 => X"0000000001200000000200000000000000000000050000400000000000000000",
INIT_11 => X"0082000000000000480080000000000012000101000080000000000000000000",
INIT_12 => X"0000004810000000000002400400000000000090400000000000000000000940",
INIT_13 => X"0000000000000000150000C00000000000000000000A40001400000000000000",
INIT_14 => X"02000000002400C2810000006000000000000000000000000000410040001400",
INIT_15 => X"020080200802008020080200800800220200840001309A08A848001000008000",
INIT_16 => X"0000000000000000000000000200802008020080200802008020080200802008",
INIT_17 => X"0080200802000000000000000000000000000000000000000000000000000000",
INIT_18 => X"940FE0D397124355520542821010000000000000000000802008020080200802",
INIT_19 => X"28A28A28A28A28A28A28A28A28A28A28A28A28A29554199854514514F546890A",
INIT_1A => X"32994CA6532995CAE572B94CA6532994CA6532994CA6532994CA28A28A28A28A",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000001867172B94CA6532994CA6572B95CAE5",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FC2155F7D155545AA80001EFAAFBEAB45557FFDE100000000000000000000000",
INIT_22 => X"FBE8BFFF78402155AAFBE8B45002A974AAAA803DFFFAA843DF45FFFFEAABA007",
INIT_23 => X"87BEAA10F7803DE00FFAEBFFFF0800155FF00042AB55FFD168B55AA8000010FF",
INIT_24 => X"AAFBEAABAA2FFD741055003DFEFF7AA801FFAAD16AABA002ABDE100800000000",
INIT_25 => X"FF7FBC0145F78028A00A2D142155087BFDE00A2FBD7400F7FBFDFFFA2AEBDE00",
INIT_26 => X"BAF780155EFAAAEA8ABAAAFBFDE0055556AA005D0415555007FD74105555555E",
INIT_27 => X"5EF0055401FFF7AEAAA105D042ABFF5D556AB55AAD168ABA002A975FFF7AEBDE",
INIT_28 => X"0000000000000000000000000000000000000000557BE8BEF007FFDEAAAAD155",
INIT_29 => X"3DF7DF7F5E8A92007BC217DEBDB55555AA8E071D7AAFBEFB455D71F8E0000000",
INIT_2A => X"B6DB55BE8E05000EBFFE8BC7E38E07145BEF1E8B6D002090482B68E38FC7BE8A",
INIT_2B => X"2EB8E00080E000280071E8A00EB8E3FE10F7AEBAFFF080A175D700042AB7DEBD",
INIT_2C => X"FF5FDFC7B6A0BDE38B6F5E8A92B6FBD5410490A3DFD7F7A4821D7A2D16FA8214",
INIT_2D => X"0071D54104951555D7EBF5C5155E3842AA00BED1421450871FFE00A2FBD0400F",
INIT_2E => X"20820955EFE3AEBDEAAFF8E175C7A2AAAAA82A2F1FAE105D556AA10410E17555",
INIT_2F => X"EF147BFAE82A2DB555C71C5B451D7FFAAA8A38410E2ABD749516FB55BED16FA8",
INIT_30 => X"F455D556AA000000000000000000000000000000000000000000000005D71E8B",
INIT_31 => X"2000F7AAA8B55FFAABDFEFF7D16AA00087FC01EFA2FFD7545AAAE97555A2FBFD",
INIT_32 => X"9554500042ABFFA2FFFFF45F7AE97400AAFFE8B45AAAA95545F7D568BEF08040",
INIT_33 => X"400155A2D57FE00552EA8A00082E820BA08556AA00AAAABFE00F7AEAABEF082E",
INIT_34 => X"517DE00A2FFC2000F7D17FF55FF803FEAAFFD16AA00FFFBD5400082EBFF45F78",
INIT_35 => X"55168A10002E9754D085155410085557555AAD557555A2802AA10FFD54214500",
INIT_36 => X"08557DF55F7D17FE000804155FFAAAABDEAAFFAA97555A2AEA8A10AAD568A005",
INIT_37 => X"0000000000555568BEF5D7FE8A10AAFFD55555D7FD5555FFAAA8AAA002AAAB45",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000008FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(10),        -- Port A data input
DOA(0)   => data_read_a_lo_256(10),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(10),        -- Port B data input
DOB(0)   => data_read_b_lo_256(10),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_11_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10180B05A0010402840602C2D001019000000300000000330A20080EC180002",
INIT_01 => X"AB400986B830284D1820E0000C3642484000000008000008820009080A512220",
INIT_02 => X"102A68440080011000000618062AD03502640800010410424908136019920868",
INIT_03 => X"004A0846191B22120642000442C110044600000101E9225CDC9A10844A9A4842",
INIT_04 => X"0094024000250808800216021138000B848000000800100040000102A0600200",
INIT_05 => X"7E4024242008A8102CA88A44010401042200444000888000000028000002A002",
INIT_06 => X"8088445712280000B18812288E0400253855200045C86810000C5B0503286A28",
INIT_07 => X"10008822A028004880200A80880208200122006C000015F0C20408264902C840",
INIT_08 => X"9390040280241041D1754100000018108728820024002B3A01A89540080824C8",
INIT_09 => X"A1001C41A1348498B080801010000080D00301081000045B0511D28D94012339",
INIT_0A => X"44080000901012428003414158230CBA4576708241C010908040341322008000",
INIT_0B => X"040464D280144050C72A0872A0C72A0872A0C72A0C72A0872A0C595043950421",
INIT_0C => X"0804001400000820110A42822204880CD81040442900021704E6000800001D54",
INIT_0D => X"80C62D0500409002082010404580018000404012004004192C10000000000000",
INIT_0E => X"80C62D5803161C526DB40506C120A806ABB0D808CC334A80A54B70D408CC32D2",
INIT_0F => X"2B5144D0DD903C54916D15458C0513005570D408CC334A80A54B70D808CC32D2",
INIT_10 => X"52148C4DB05621E363F813961C20EDA944016558C2347A080B10D8DD6422AA10",
INIT_11 => X"1880144D3345C65593800319C18BD1ECA1C9010112566F10AC4183C340DAE02D",
INIT_12 => X"5810503000633830DE3C2C9C00289A66AA8DE50E0800360614AC281430890600",
INIT_13 => X"0CD2A9CEA8199B6B082B55900314140365320485C4F00AD544407241C175C402",
INIT_14 => X"0000074044C4801832701A89D20A38093631425969020855A281844E00540404",
INIT_15 => X"0000000000000000000000000020C00200088101513492101280401000400200",
INIT_16 => X"2008020080200802008020080000000000000000000000000000000000000000",
INIT_17 => X"0080200802008020080200802008020080200802008020080200802008020080",
INIT_18 => X"804180C0B10A4210420140028400000000000000000000802008020080200802",
INIT_19 => X"000000000000000000000000000820820820820801C414947000000055062608",
INIT_1A => X"0000000004020000000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000001F87E000000000000010080000000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"ABDF5508557DF45002ABDFFFF7803DE10AA80000AA0000000000000000000000",
INIT_22 => X"FFE8A10A28000000007FC2155F7D155545AA80001EFAAFBEAB45557FFDE10082",
INIT_23 => X"02A974AAAA803DFFFAA843DF45FFFFEAABAA2AEBFF45FFAEBFEAA002A801FFF7",
INIT_24 => X"F78402155AAD155555A28428BFF002ABDE00A2AABFE10082ABFFEFAAFBE8B450",
INIT_25 => X"0002A80010A2842AAAA007BFFF4500042AB55FFD168B55AA8000010FFFBE8BFF",
INIT_26 => X"00080000000087BEAA10F7803DE00FFAEBFFFF0800155FF00557FF45557FC201",
INIT_27 => X"1FFAAD16AABA002ABDE10A2D168A10A284021FF5D00154BAF7FBE8BEFFFD5400",
INIT_28 => X"0000000000000000000000000000000000000000A2FFD741055003DFEFF7AA80",
INIT_29 => X"EFB455D71F8E00002EBDF6D005B78F7D142ABDFC7F78E3FE28B684070AA00000",
INIT_2A => X"0BDEAA1C2A801C7E3FFEFA10B68407038007BC217DEBDB55555AA8E071D7AAFB",
INIT_2B => X"20B8FEFBEF1E8B6D002090482B68E38FC7BE8A3DF7DF7F5E8A92BEAEBFF7DEBA",
INIT_2C => X"E8E05000EBFFE8BC7E38E07145B6D15756DA28A28BFF082ABAE10B6AAB8E2808",
INIT_2D => X"08517DF7D497BC5028142A87000A28A2AA92007FF8F7D00042AB7DEBDB6DB55B",
INIT_2E => X"2FFFFEFBC7E3DF42028080E000280071E8A00EB8E3FE10F7AEBAFFF080A175D7",
INIT_2F => X"10490A3DFD7F7A4821D7A2D16FA82142EB8E00B6DB6AA28A280001FF5D0A1048",
INIT_30 => X"EAAF784154BA000000000000000000000000000000000000000000000B6FBD54",
INIT_31 => X"7545AAAE97555A2FBFDF455D556AA00082EBFFEF007BE8BFF5D2ABDF55F7AABD",
INIT_32 => X"6AA00FFAEBFFEFAA803DEBA5D2E82155A2FBFDE00FF84154BA087FC01EFA2FFD",
INIT_33 => X"AAAA00FFAAA8AAA080028BFFF7D568BEF080402000F7AAA8B55FFAABDFEFF7D1",
INIT_34 => X"042ABFFA2FFFFF45F7AE97400AAFFE8B45AAAA95545F7D5555FFAAAAA8BFF002",
INIT_35 => X"7AEAABEF082E9554508557DFFF007BD54BA5D2E95400A2AEA8A00007FEABFF00",
INIT_36 => X"AA80001FF5D2E82000F7FFFFF45AAFFC20BA082E820BA08556AA00AAAABFE00F",
INIT_37 => X"0000000000FFFBD5400082EBFF45F78400155A2D57FE00552EA8A00FFFFE8AAA",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000800000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(11),        -- Port A data input
DOA(0)   => data_read_a_lo_256(11),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(11),        -- Port B data input
DOB(0)   => data_read_b_lo_256(11),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_12_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"A500C4B01BC0268A6940312C0DE045196A831A300500032B333287E4FC812006",
INIT_01 => X"AF400D869830E84D5823E0000C1742484000000008000008820009280A553235",
INIT_02 => X"502A7144008001100000171C022BD13412762A000586235ECC09C8423B960866",
INIT_03 => X"31863846191BA218064204000281200406A10843010022DEDF0852944A9C014A",
INIT_04 => X"0014030000250409000014821038080B840000400800102040000302F0600233",
INIT_05 => X"7FC034348008A8102CA88F48010601042400048000188000000938000002E088",
INIT_06 => X"9CC96CC6F63A5001F12B56A0AC8601F47AC06400D1F80C10020C493F03343A38",
INIT_07 => X"1020002030280098A12048908A16BA311177124C000003F08A94282E5C262861",
INIT_08 => X"827A0602902A10491165E10000049010C52882008600A73A01E8974008092CF8",
INIT_09 => X"47000001A1248008F000000000000080000F010C100204593F11A6CDF48023BF",
INIT_0A => X"040000208010120ACA01400058010CBA4D277C86CCE802B380003C1360008000",
INIT_0B => X"011C46D3C7BC1EF083AF0C3AF083AF083AF0C3AF083AF083AF0C1D7861D78400",
INIT_0C => X"08040014C9001AE91D17E50AD79FEFC87C2154745F82131FFCCE00080000095E",
INIT_0D => X"807BF7118180984004000803D40001880001001400C005031010000000000000",
INIT_0E => X"807BF76A109C944B5891BF06C5EEB14FCBF0D90076D61C807BF7D0D80876D49C",
INIT_0F => X"6DE38EB9FB10350C00A99F7CA80757365E50D80876D61C807BF7D0D90076D49C",
INIT_10 => X"841BCC69A0D8C6F7F0AA001C943A65756A0976EB5A7E7FC8951018186334F311",
INIT_11 => X"D5A014481991C6A737D80211912970CDCDD1864116D6C7080651CB4661F33615",
INIT_12 => X"349E929300423224AE19B9BEC0289033238D4E6EA805892946A9B011A7B152CF",
INIT_13 => X"6244CD7AC01CAAA56B3E6D9001068715D64006D2A961CF9B44512A2504532182",
INIT_14 => X"00000439FDC25C58067A9FAB46095A0B5289A0282D2E1444ACB12A17CF9B4414",
INIT_15 => X"0000000000000000000000040026C00000288401513492909280401000F70A00",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"088881360A95090CB05442029010000000000000000000000000000000000000",
INIT_19 => X"1041041041041041041041041049249249249249200100002D4514510051B946",
INIT_1A => X"592C964B2592C964B2592C964B2592C86432190C86432190C864104104104104",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000002007F592C964B2592C964B2592C964B2",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"43FE0008557DFFF0800020105D557FEAA00557DE100000000000000000000000",
INIT_22 => X"557DFFFF7AA80000082ABDF5508557DF45002ABDFFFF7803DE10AA80000AAAA8",
INIT_23 => X"7D155545AA80001EFAAFBEAB45557FFDE10AAD5420000051555FFA2AA8200000",
INIT_24 => X"A28000000A2D155410F7FFFFEBA08003FE00082AA8AAAAAFFC00BA007FC2155F",
INIT_25 => X"0A2AABFE1055516ABEF5D517DEAAA2AEBFF45FFAEBFEAA002A801FFF7FFE8A10",
INIT_26 => X"55AAFBE8B45002A974AAAA803DFFFAA843DF45FFFFEAABA000028A105D2ABFE1",
INIT_27 => X"E00A2AABFE10082ABFFEF085542000000417555002A820AA08557DFFFF7AA821",
INIT_28 => X"0000000000000000000000000000000000000000AAD155555A28428BFF002ABD",
INIT_29 => X"3FE28B684070AABE803AE38145B78FD7000005010495B7AE921C517DE1000000",
INIT_2A => X"B505FFB6A487000005F7AFD7F7A482038002EBDF6D005B78F7D142ABDFC7F78E",
INIT_2B => X"F5C2082007BC217DEBDB55555AA8E071D7AAFBEFB455D71F8E00BED547038145",
INIT_2C => X"C2A801C7E3FFEFA10B68407038B6D550428FFF1FDE821C003FE001C2EAAAAAB6",
INIT_2D => X"00002FA285D20BDE28A2A4B8E10555B68BEF5D517DEAABEAEBFF7DEBA0BDEAA1",
INIT_2E => X"2005F7DFD7F7A482155BEF1E8B6D002090482B68E38FC7BE8A3DF7DF7F5E8A92",
INIT_2F => X"6DA28A28BFF082ABAE10B6AAB8E280820B8FEF085F4703814001055514208208",
INIT_30 => X"A0055517DE00000000000000000000000000000000000000000000000B6D1575",
INIT_31 => X"8BFF5D2ABDF55F7AABDEAAF784154BAF7802AABA5D7FEAB45080015410007FEA",
INIT_32 => X"6AA00F7D1554BA5D7BC01FFFF8015410007FEAB45F780020BA082EBFFEF007BE",
INIT_33 => X"43FE10552EAAAAAFFD140000087FC01EFA2FFD7545AAAE97555A2FBFDF455D55",
INIT_34 => X"AEBFFEFAA803DEBA5D2E82155A2FBFDE00FF84154BAF7D1400BAFFD57FE005D0",
INIT_35 => X"FAABDFEFF7D16AA0008003FEBA55003DEBAA28428A105D7FEABEF55557DEBAFF",
INIT_36 => X"550402145550000010087FFFF45F78402145F7D568BEF080402000F7AAA8B55F",
INIT_37 => X"0000000000F7D5555FFAAAAA8BFF002AAAA00FFAAA8AAA080028BFF087BD54AA",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000000FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(12),        -- Port A data input
DOA(0)   => data_read_a_lo_256(12),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(12),        -- Port B data input
DOB(0)   => data_read_b_lo_256(12),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_13_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10110A0441812402840402822007818000E00700000000330A3000000008042",
INIT_01 => X"A1400984B830C848180260000C0042604001000008220008A200100802110200",
INIT_02 => X"10A00860009141100000C6180C285035000E0800010431004908135980120C60",
INIT_03 => X"004E20441910221B06420C85D5013804060000000040324C441A108468024842",
INIT_04 => X"0184034010250089C00EA8021938325B04800002091090014880080200000900",
INIT_05 => X"18002424B008881024A8004E01040104270004E0000080090500604840000481",
INIT_06 => X"80004414022A2490B00A142C8C840005794540015E006810001C4B01032C7E20",
INIT_07 => X"510200028028004880280A808816002101022468000011F082040A264006C000",
INIT_08 => X"D2B00402B220104B531001000008001041080200B660E30B200C8040080A9206",
INIT_09 => X"A1000809A93484D21000000000000080C90391881000145B0111A30404015000",
INIT_0A => X"000000008010102A82014100101118BA4510008241480290882400900000A000",
INIT_0B => X"0284484000000000400000000040000000000000040000000000000020000000",
INIT_0C => X"A944AA2000A02000212800020000000D80004084A0000390002E001843210400",
INIT_0D => X"859C1881A04090000000000021800180010341179065441356150A1285094284",
INIT_0E => X"859C188810C65A72A617520252781EA02520D589B9A260859C1840DD81B9A0E0",
INIT_0F => X"0E71F1052D942748C19484E39442D15961C0DD81B9A260859C1840D589B9A0E0",
INIT_10 => X"E60605C0C12CBD400B0810C65A61AA459D0047398500D5889D26907356533C00",
INIT_11 => X"8F60CA1562094650CA28398A42C051E0332181010109294C8E1160CB8C80A561",
INIT_12 => X"2645056D073148580A3C065141942AC4128CA199180C5232575138094450AD0A",
INIT_13 => X"84CA93A2FC008962142B17301A9A1A5196A80245208E0AC5C853C8028163B8C0",
INIT_14 => X"0240034000E4DC8A84000014982372011FC1E475F0F0084A3961F5A80AC5C816",
INIT_15 => X"4250942509425094250942509428D421420882020120981812C8403000088212",
INIT_16 => X"2509425094250942509425094250942509425094250942509425094250942509",
INIT_17 => X"5094250942509425094250942509425094250942509425094250942509425094",
INIT_18 => X"FF3F7DF7FF3E9F7DF7E24502A800000000000000000050942509425094250942",
INIT_19 => X"EBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBF7DFDFDDD555555F7EFBBEE",
INIT_1A => X"7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAEBAEBAEBAEBA",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000000007F7EBF5FAFD7EBF5FAFD7EBF5FAFD",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5554BA087FFFF55557BD54AAF7FBC01FFA2802ABEF0000000000000000000000",
INIT_22 => X"2E80155AA802AB45AA843FE0008557DFFF0800020105D557FEAA00557DE10AAD",
INIT_23 => X"8557DF45002ABDFFFF7803DE10AA80000AA087BD75EF087FFFFEF557BEAB4555",
INIT_24 => X"F7AA80000AAD1420AA087BD7555FFD168AAAFFAE820AA5D5557555082ABDF550",
INIT_25 => X"5FFD157555085140010F7AEAABFFAAD5420000051555FFA2AA8200000557DFFF",
INIT_26 => X"45007FC2155F7D155545AA80001EFAAFBEAB45557FFDE10AAAEA8BFFA2FBD754",
INIT_27 => X"E00082AA8AAAAAFFC00BA00002AAAAF7D5574BA557BE8A10A284154BAFFAAAAB",
INIT_28 => X"0000000000000000000000000000000000000000A2D155410F7FFFFEBA08003F",
INIT_29 => X"7AE921C517DE10A2DB50482147FFAF554971D0492E3F1C71C7BE8A2ABD700000",
INIT_2A => X"FFAFD7497BE8B5555208217DBE8A2AB45BE803AE38145B78FD7000005010495B",
INIT_2B => X"5F5056D002EBDF6D005B78F7D142ABDFC7F78E3FE28B684070AA1C71D25D7007",
INIT_2C => X"6A487000005F7AFD7F7A482038AADF47092147FD257DFFD568A82FFA4870BA55",
INIT_2D => X"A2A0ADBC7A2FFD257DE3DF52555085142000FFAAAFBFFBED547038145B505FFB",
INIT_2E => X"0B680124BAFFAAAFB45007BC217DEBDB55555AA8E071D7AAFBEFB455D71F8E00",
INIT_2F => X"28FFF1FDE821C003FE001C2EAAAAAB6F5C20821C002AA92FFDF574824171EAA1",
INIT_30 => X"545F7AEA8B55000000000000000000000000000000000000000000000B6D5504",
INIT_31 => X"AB45080015410007FEAA0055517DE00A2FFC00105D7BE8B55085142010AAD157",
INIT_32 => X"154BA5D5140145007BE8B55087BEAB555D04001EFF7AAA8B55F7802AABA5D7FE",
INIT_33 => X"16AA10FF80174AA557FC21EF082EBFFEF007BE8BFF5D2ABDF55F7AABDEAAF784",
INIT_34 => X"D1554BA5D7BC01FFFF8015410007FEAB45F780020BAA2FFD54105D7FC21EFFFD",
INIT_35 => X"2FBFDF455D556AA00A2803FF45AAFFC21EFAAFBC0155085540000FFAEBFFEFF7",
INIT_36 => X"F7FBD5410085568A10FF80020AAFFAABFF55087FC01EFA2FFD7545AAAE97555A",
INIT_37 => X"0000000000F7D1400BAFFD57FE005D043FE10552EAAAAAFFD1400005D042AA00",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000CFFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(13),        -- Port A data input
DOA(0)   => data_read_a_lo_256(13),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(13),        -- Port B data input
DOB(0)   => data_read_b_lo_256(13),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_14_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10020A000180000284008280000281800000030000000033022000000580002",
INIT_01 => X"A140098018300848184860000C20C24040000000084000084200000000110200",
INIT_02 => X"1020006000900110000006102028503400040800010400204908012018120E64",
INIT_03 => X"000200441910221006420000400100040600000000E9E401209A108448004842",
INIT_04 => X"0004020000250008000200021038000804000000090090004800080200000000",
INIT_05 => X"500024240008881024A800400104010420000400000080080100204040000000",
INIT_06 => X"8000440102282015B10A10288E0400042345400040006810000C5901033D7880",
INIT_07 => X"1100000200280048802008828812002001220064000005F1C2850A2649204070",
INIT_08 => X"00B00402802010411110010000080010010802000400230B000C804008080002",
INIT_09 => X"01000009A92480001000000000000080C8038188100004590111B68404010000",
INIT_0A => X"0000000080101000000141001001088A45000082400000008020009000008000",
INIT_0B => X"0004404000000000400004000000000000004000000000000004000000000000",
INIT_0C => X"8904A0200080200001080002000000088000400420000200002E000841010400",
INIT_0D => X"0500000C80409000000000000000018000000000806044010014081204090204",
INIT_0E => X"0500005813A0210D072E8D012001028402908004000587050000108004000707",
INIT_0F => X"9004300044900812386A280E5800088980108020000587050000108020000707",
INIT_10 => X"DE00482E19E30002007813A02096038AE200880405200308828062A68C0BC700",
INIT_11 => X"00000E5A08E6000048001292B83280001208A1011004011060049A1C59192055",
INIT_12 => X"492060480256530650000240001DB011CC00009000032C4C979E3806180C0900",
INIT_13 => X"5A3433EDE00154181400000007BCBD858F120120541A0000000033757465B2C0",
INIT_14 => X"02002C000024008A84001A0902000422E3E99681004802115652594000000001",
INIT_15 => X"0240902409024090240902409028D021020880000120901812C8401000000210",
INIT_16 => X"2409024090240902409024090240902409024090240902409024090240902409",
INIT_17 => X"4090240902409024090240902409024090240902409024090240902409024090",
INIT_18 => X"5C8FF0F7BE9D5F7DF65040028000000000000000000040902409024090240902",
INIT_19 => X"79E79E79E79E79E79E79E79E79E79E79E79E79E7BF7DDDDDFCF3CF3DF5579B4E",
INIT_1A => X"3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE79E79E79E79E",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000003FF803F9FCFE7F3F9FCFE7F3F9FCFE7F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"BE8B55A2AE80000F7D5555555D2AAAABAAAD1420BA0000000000000000000000",
INIT_22 => X"00155EF0804155EFAAD5554BA087FFFF55557BD54AAF7FBC01FFA2802ABEFA2F",
INIT_23 => X"8557DFFF0800020105D557FEAA00557DE10A2AA801FFA28402000AAAE9554555",
INIT_24 => X"AA802AB4500516AA00A2AE800BAFFFFC20BAF7AEA8B45080417400AA843FE000",
INIT_25 => X"0A2843FEBAFFFBD7410A2D168BFF087BD75EF087FFFFEF557BEAB45552E80155",
INIT_26 => X"AA082ABDF5508557DF45002ABDFFFF7803DE10AA80000AA005568ABAA2840201",
INIT_27 => X"AAAFFAE820AA5D5557555002E80155A280000005D7FFDF4555517DFEF00043FE",
INIT_28 => X"0000000000000000000000000000000000000000AAD1420AA087BD7555FFD168",
INIT_29 => X"C71C7BE8A2ABD7A2FFEDB55B6A080038E3DB50555412AA8ABAAADB4009200000",
INIT_2A => X"402038AAAA955554900105FF0800175D7A2DB50482147FFAF554971D0492E3F1",
INIT_2B => X"0A12410BE803AE38145B78FD7000005010495B7AE921C517DE10A2AE851FFB68",
INIT_2C => X"97BE8B5555208217DBE8A2AB451C556FA00A2A0800BAE3F1C0092EBAAADB6D08",
INIT_2D => X"00516DABAA28402038B6803DE82F7F5D5410A2D568BC71C71D25D7007FFAFD74",
INIT_2E => X"55D5F78FD7000E3FEAA002EBDF6D005B78F7D142ABDFC7F78E3FE28B684070AA",
INIT_2F => X"92147FD257DFFD568A82FFA4870BA555F5056D002A80155B680000105D7FF8F4",
INIT_30 => X"AAAAAFFC2000000000000000000000000000000000000000000000000AADF470",
INIT_31 => X"8B55085142010AAD157545F7AEA8B55A2FBFFF55FF84000AAAAFBC0145002AA8",
INIT_32 => X"7DE00A2AA955FFFF80020BAAAAA975450800001EF080417555A2FFC00105D7BE",
INIT_33 => X"140000A2AEBFFEF082A82010F7802AABA5D7FEAB45080015410007FEAA005551",
INIT_34 => X"5140145007BE8B55087BEAB555D04001EFF7AAA8B555D557FE00A280020BAAAD",
INIT_35 => X"7AABDEAAF784154BA08557FEAAA284000AAFF803DE00FFD557400AAD56AB455D",
INIT_36 => X"F780020105D7BEAB45557BE8B45082EBFEBA082EBFFEF007BE8BFF5D2ABDF55F",
INIT_37 => X"0000000000A2FFD54105D7FC21EFFFD16AA10FF80174AA557FC21EF082A80145",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000000FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(14),        -- Port A data input
DOA(0)   => data_read_a_lo_256(14),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(14),        -- Port B data input
DOB(0)   => data_read_b_lo_256(14),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_15_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000A000000000284000280000001800020030000000033022000000180002",
INIT_01 => X"A140098018300848180060000C00424040000000080000080200000000110200",
INIT_02 => X"102100400C8011100000061000A8503401044880010430004808000180122378",
INIT_03 => X"000200541D102210064200000045000546080000400020000008108448400042",
INIT_04 => X"8094020000254C880000028A1018000844000000880013504000002600000000",
INIT_05 => X"10002424000AA81024A82040010C61062001440002988000000024808001004B",
INIT_06 => X"80004400022A00003C8912248E0400042854400040006810000C4901032B1800",
INIT_07 => X"50200000B0280048A0280A828801002101020040000005F38204082640000000",
INIT_08 => X"01F00402802610411100110000000010010802000400230A0008884008080004",
INIT_09 => X"01000001A12481041000000000000080C0030108100004590111820404000000",
INIT_0A => X"0000000080101000004140001001088A45000082000000008000001080008000",
INIT_0B => X"0004404000000000400004000040000400000000000000000004000020000200",
INIT_0C => X"0804000020024100012808020000000981004004A0200310000C000800000000",
INIT_0D => X"0000001180009000000000002100018000000000004004010010000000000000",
INIT_0E => X"00000008000002000000000000000000000080A40000000000000080A4000000",
INIT_0F => X"00000000001000204800000000000000000080A40000000000000080A4000000",
INIT_10 => X"000000000000000000080000020000000000000000000008000C020000000000",
INIT_11 => X"000000824000000000000020220000000001800100020300000004003420480A",
INIT_12 => X"0000000000040440000000000001048000000000000000100800400000000000",
INIT_13 => X"000800000000000000000000000100C220050000000000000000008220884400",
INIT_14 => X"000000000000000830000000000000000016101C5C1400000000000000000000",
INIT_15 => X"0000000000000000000000000020C00000088000012090101280401000000200",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000040028000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"000010082A954BA00003DFEF085155400F78428BEF0000000000000000000000",
INIT_22 => X"8015400FF84001EFA2FBE8B55A2AE80000F7D5555555D2AAAABAAAD1420BAFF8",
INIT_23 => X"87FFFF55557BD54AAF7FBC01FFA2802ABEFF7AE95555A2FBE8BEFA2843DE00AA",
INIT_24 => X"0804155EFFFFBE8BFF0800174AA557BFDE10A2FBEAB45F7D56AABAAAD5554BA0",
INIT_25 => X"5FFD568BEF087FE8A1055003FE00A2AA801FFA28402000AAAE955455500155EF",
INIT_26 => X"45AA843FE0008557DFFF0800020105D557FEAA00557DE10F7D1574AAA2D16AB5",
INIT_27 => X"0BAF7AEA8B45080417400FFFFC2145080015400AA802AA00AAAE800BA5D00155",
INIT_28 => X"000000000000000000000000000000000000000000516AA00A2AE800BAFFFFC2",
INIT_29 => X"A8ABAAADB40092E38E070280024904AA1C0438FD7005150438F78A2DBFF00000",
INIT_2A => X"FE8BC7BE8E38E10A28017400E38A051FFA2FFEDB55B6A080038E3DB50555412A",
INIT_2B => X"D16AABAA2DB50482147FFAF554971D0492E3F1C71C7BE8A2ABD7E3AA9257DA2F",
INIT_2C => X"AAA955554900105FF0800175D7E3FFEFBD70000124AA557FFDE10A2FBEDB6DF7",
INIT_2D => X"FFDF50482A2DB6AB45FFD56DBD7087BEAA38410038E38A2AE851FFB68402038A",
INIT_2E => X"0AAA085082550A1057DBE803AE38145B78FD7000005010495B7AE921C517DE10",
INIT_2F => X"00A2A0800BAE3F1C0092EBAAADB6D080A12410FFF1C017D140410400BE8E28A1",
INIT_30 => X"0AAF7AEBDFEF0000000000000000000000000000000000000000000001C556FA",
INIT_31 => X"00AAAAFBC0145002AA8AAAAAFFC2000AAAA974AA0800020BA550028B55085540",
INIT_32 => X"A8B55AAAE821EFAAFBEAB55F7AAA8A00AA8417400AAAE975EFA2FBFFF55FF840",
INIT_33 => X"BFFE10A2FFFFFEFF7D568ABAA2FFC00105D7BE8B55085142010AAD157545F7AE",
INIT_34 => X"AA955FFFF80020BAAAAA975450800001EF080417555AAFFFDF450804020AA557",
INIT_35 => X"07FEAA0055517DE00FFFBC2000AAFBE8B55F7D17DF45007FE8AAA08002AAAAA2",
INIT_36 => X"5D0000010F7AAA8A10AA8017400552A801EFF7802AABA5D7FEAB450800154100",
INIT_37 => X"00000000005D557FE00A280020BAAAD140000A2AEBFFEF082A82010FFD5421EF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000C00000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(15),        -- Port A data input
DOA(0)   => data_read_a_lo_256(15),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(15),        -- Port B data input
DOB(0)   => data_read_b_lo_256(15),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_16_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"DA22C618B1000482B688B186588884862A400438255FC38381441205BA803003",
INIT_01 => X"264AC80028404C211203A952A90341080B173340412000E1005D628000820484",
INIT_02 => X"400034C206C405000001A48202084004003008255040826EE008B440200E2042",
INIT_03 => X"A459C1240181AB20AD27315B7F1983CA1C900040422A005762010010000C0400",
INIT_04 => X"296E542B6E3A825C15FB385321B4ADFE16AB45FD2C400002E205231201290A28",
INIT_05 => X"B9E5815006028179808C00A0D2152B90707A1E0BD423CAC0000D610000000710",
INIT_06 => X"81F104A1415C292164280081C6AB88742086ACACDE240000A80090CE82A803B9",
INIT_07 => X"400800000ACCAA280940580400A37B8896CA4D000A80C1102A00001C14028009",
INIT_08 => X"0015452880C8D90409A02D965965200100104F2B00822512000000231520A024",
INIT_09 => X"A5AA80018120E00066000000000012C9000A0000D0A80000BF8028E87C1B9927",
INIT_0A => X"00520228080108039501200848002912300208092B940192D1000000000000A8",
INIT_0B => X"03561180063DB4F6110001100011000110001100011000110001080008800080",
INIT_0C => X"080200854409418B02ED0000502A02972000040BB401100010012B4C90000100",
INIT_0D => X"6D061A1F8D60D80820500101244AA8A2AA242E80000009200120000000000000",
INIT_0E => X"6D066210E5001DB4A5B400C7D553847165A99000C6564CDD051DC99000C65555",
INIT_0F => X"21D0C48F254946148107354292673D1F72C99000C6564CDD0565C99000C65555",
INIT_10 => X"952D2058F33225787810F5001D6121A9559224D1FF97D0272F04D89441A56D8A",
INIT_11 => X"6C1C74485B81E31306C71D1093AB8A64811BADC00992180D58033B1172F2A025",
INIT_12 => X"7B86DED8E3A212748F0E0CA638E890B7A8546120C0AFF5B548AC431FB1C7DB07",
INIT_13 => X"EFCE9B26DECA1AD36A2E4F40DF6AAAF260AF88899E8B8B93D12A877178DD0032",
INIT_14 => X"A8009F8B108C80A1021B9A8BB8056662CA1951596800FC01A38D4D4B072B922F",
INIT_15 => X"00000000000000000000000000044000102A0001148442A1108103595580A840",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"4C690DA64C1C4F68A36040000000000000000000000000000000000000000000",
INIT_19 => X"D14D14D14D14D14D14D14D14D14514514514514529E5F87869E79E78558D1154",
INIT_1A => X"3D1E8F47A7D3E9F4FA7D3E9F4FA7D3E9F47A7D1E9F47A7D1E9F4D14D14D14D14",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE000000000000000007D3E9F4FA7D3E8F47A3D1E8F47A",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFEFF7D168B55AAD17FFFF552EBFE00007FC00AA0000000000000000000000",
INIT_22 => X"04000BA552A821FFFF8000010082A954BA00003DFEF085155400F78428BEF087",
INIT_23 => X"2AE80000F7D5555555D2AAAABAAAD1420BA5D2E975EFF7D568BFFFF80175EF00",
INIT_24 => X"FF84001EF0000020AA5D00154005D043FF45555540000082EAABFFA2FBE8B55A",
INIT_25 => X"0087FD74BAAAAEBFFEF557FC00AAF7AE95555A2FBE8BEFA2843DE00AA8015400",
INIT_26 => X"FFAAD5554BA087FFFF55557BD54AAF7FBC01FFA2802ABEF557BEABEF5D041541",
INIT_27 => X"E10A2FBEAB45F7D56AABA082A97545F7D16ABFFFFAABFEAAFF84001FF002A821",
INIT_28 => X"0000000000000000000000000000000000000000FFFBE8BFF0800174AA557BFD",
INIT_29 => X"50438F78A2DBFF0871F8FC7E3D56AB6DBEDB7FFEF552AB8E38087FC209200000",
INIT_2A => X"16ABFFE38E175EF1400000BA412E871FFE38E070280024904AA1C0438FD70051",
INIT_2B => X"2EAFBD7A2FFEDB55B6A080038E3DB50555412AA8ABAAADB400924920925EFF7D",
INIT_2C => X"E8E38E10A28017400E38A051FF0804050BA410A1240055003FF6D5551420101C",
INIT_2D => X"4975EDBC7550E12410087FD74AAB6AABFFC7557FC00BAE3AA9257DA2FFE8BC7B",
INIT_2E => X"AF780051C70824851D7A2DB50482147FFAF554971D0492E3F1C71C7BE8A2ABD7",
INIT_2F => X"D70000124AA557FFDE10A2FBEDB6DF7D16AABA08249756DF7D168BC7F7AABAEA",
INIT_30 => X"AAA007BC0000000000000000000000000000000000000000000000000E3FFEFB",
INIT_31 => X"20BA550028B550855400AAF7AEBDFEF08516AB55A2D16ABEFFFFBFDFFF552AAA",
INIT_32 => X"C20000000021EFF7D568BFFA2AA955FF5D04020AA002A955EFAAAA974AA08000",
INIT_33 => X"03DFEF5D51420005D2ABFF45A2FBFFF55FF84000AAAAFBC0145002AA8AAAAAFF",
INIT_34 => X"AE821EFAAFBEAB55F7AAA8A00AA8417400AAAE975EF0800174BA002E820105D0",
INIT_35 => X"AD157545F7AEA8B5500557DF45552A82000007BD74AAF7AEBDF455D7BC20BAAA",
INIT_36 => X"F7D568B55FFAAAAABAFF8415545000015555A2FFC00105D7BE8B55085142010A",
INIT_37 => X"0000000000AAFFFDF450804020AA557BFFE10A2FFFFFEFF7D568ABA0804155FF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000400000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(16),        -- Port A data input
DOA(0)   => data_read_a_lo_256(16),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(16),        -- Port B data input
DOB(0)   => data_read_b_lo_256(16),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_17_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"5284CE4FB7BD2C8994A13392DBD02E14006B82AC7E800D44D3DD2FD5F9B961C0",
INIT_01 => X"F9BA301F7E03FC6793F2199B39FC233C11D93AE6F3BB92B32091DBC339B24542",
INIT_02 => X"1D5FC0C08F040404446965C0607FB8A217C400C33A908078551BD04222186338",
INIT_03 => X"8504930A37F65820CB24111B7F08014A0AB84A52B6D2AFF97C1B5AC757F06D6B",
INIT_04 => X"250834336D1E81500FDB38302292ADFE103B6DBD204037F202042075E2B1D00A",
INIT_05 => X"8F039786062C6CE092F5FE005236781C402A0807B4070670083DC68206D7E6D0",
INIT_06 => X"0CD26803C3582408962C58B183F8AEF42045919B30E085DD2ED57D4EED08CA6A",
INIT_07 => X"700000B30380670B8142500448E3E01E94EF1340A28AC1AC8156044D1400AA00",
INIT_08 => X"009F3A1B0120A1C51DFFC40C30E5F0182D0950190C0810BE00E9A76E4C6FFBE4",
INIT_09 => X"8FCCC200A59BDD2FFE3F3EC7C7DEF207000F00059D2ED56D7EED2ED3C9A867DC",
INIT_0A => X"0617112E46F05D02DD814102F800633F1D0A7CC9AE7A08BFF0001D35682AC0CE",
INIT_0B => X"8A3F06ABD73DBCF4FBCF4FBCF4FBCF4FBCF4FBCF4FBCF4FBCF4FBE7A7DE7A780",
INIT_0C => X"001000974F08518F5AFFC94B533FADA7FDE97D6BFF329E1B50FF99F086000D9E",
INIT_0D => X"F50B018F95EA3DED1652EC0B27E67F419E2E1E8000C0036340B8000000000000",
INIT_0E => X"F50B01C8DF7F96197DB4AFC8C8886AF672A1537F759299F50B03C1537F759199",
INIT_0F => X"6068331C5103E7EF0FBEED6BB6A9412007C1537F759299F50B03C1537F759199",
INIT_10 => X"21F2CD7F252CDABB3CE8CF7F963AB9FD6AD434201AA68B837FFD1F7B7125B68C",
INIT_11 => X"BD055EB6D555CB2949C15BA7270FF256526BBFD55BBE71D79F73C7AC6DB9BF37",
INIT_12 => X"94080BF82B74E4E1FE4ACA4E0ABD6DAAAB965293036FF6B652A99A6026027FBE",
INIT_13 => X"EF5CBA7A43482800FEFAFD06B8CFCCAB7550D0C2022EAEBD438697AD2EBA9168",
INIT_14 => X"AC00A8BBFC8B501CF7A0FED9A548FA19752C4A4EADAE42FCBC38C3B7BEBF42CF",
INIT_15 => X"0000000000000000000000000026E100002F382DBD9ECFE117805F20CFDAAB00",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"09EDCC4052E917114F981800C000000000000000000000000000000000000000",
INIT_19 => X"EBA69AEBA69A69AEBA69AEBA69A69A69A69A69A68698686981D75D7443720030",
INIT_1A => X"46A351A8D068341A0D068341A0D068341A0D46A341A0D46A341A69AEBA69A69A",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000000000046A351A8D46A351A8D46A351A8D",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFEFF7FBEAB450804001EFAAD57FEAA0000000000000000000000",
INIT_22 => X"51401EF087FD74AA087FFFFEFF7D168B55AAD17FFFF552EBFE00007FC00AA087",
INIT_23 => X"82A954BA00003DFEF085155400F78428BEFAAD168A000004020AA5D7BE8B4500",
INIT_24 => X"552A821FF5D00020BA552A82000552A821555D7FEAB55FF80175EFFF80000100",
INIT_25 => X"FAAFBC01EF5D0015555557BFDEBA5D2E975EFF7D568BFFFF80175EF0004000BA",
INIT_26 => X"BAA2FBE8B55A2AE80000F7D5555555D2AAAABAAAD1420BAFFFFFDF45AAD17FFF",
INIT_27 => X"F45555540000082EAABFF00516AA10552E820BA007FEABEF005555555A2D1554",
INIT_28 => X"00000000000000000000000000000000000000000000020AA5D00154005D043F",
INIT_29 => X"B8E38087FC2092147FFFFFFFFFBFDFC7EBF5E8B550000071EFB6DF7AE9200000",
INIT_2A => X"A07082497FEFB6D1451471EF007BD04920871F8FC7E3D56AB6DBEDB7FFEF552A",
INIT_2B => X"8E175FFE38E070280024904AA1C0438FD7005150438F78A2DBFFBED16AA381C0",
INIT_2C => X"38E175EF1400000BA412E871FF550A00092492A850105D2A80155417BEFB6DEB",
INIT_2D => X"FFF5FFF6DAADF7FFD7B6F1C71EF55001756D5D7BFAEBA4920925EFF7D16ABFFE",
INIT_2E => X"700515556DA2DF50492A2FFEDB55B6A080038E3DB50555412AA8ABAAADB40092",
INIT_2F => X"BA410A1240055003FF6D5551420101C2EAFBD7145B6AA28492487082007FEDBD",
INIT_30 => X"5EFFFFBEAA000000000000000000000000000000000000000000000000804050",
INIT_31 => X"ABEFFFFBFDFFF552AAAAAA007BC0000557FFDFEFF7FBFFF55A2D16AB55000017",
INIT_32 => X"BDFEFF7D568AAA5D2A97410007BFFFFF5551555EF087FC200008516AB55A2D16",
INIT_33 => X"A82155087FFFFEFAAAA975EFAAAA974AA0800020BA550028B550855400AAF7AE",
INIT_34 => X"00021EFF7D568BFFA2AA955FF5D04020AA002A955EF5D2E80010002A954005D2",
INIT_35 => X"02AA8AAAAAFFC2000FFD57DFFFAAFFFDF55FFD1575FF5504175EF5D7FEAAAA00",
INIT_36 => X"000415410007BFFF450051555EFA2FBC0000A2FBFFF55FF84000AAAAFBC01450",
INIT_37 => X"00000000000800174BA002E820105D003DFEF5D51420005D2ABFF45557FE8AAA",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000CFFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(17),        -- Port A data input
DOA(0)   => data_read_a_lo_256(17),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(17),        -- Port B data input
DOB(0)   => data_read_b_lo_256(17),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_18_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"69844019080000A21A611406840014122A641074155FC28A2024001001801003",
INIT_01 => X"01067920034004180005E9E3C90360C0041C0181002001602025800008440084",
INIT_02 => X"40AC3CAA22D605200000856E2481902400344A20F802C22054001000021E2379",
INIT_03 => X"A54C23B34C81EB2076471000800981140C010101750D1007E58040102B0E0100",
INIT_04 => X"22660C1C0065003C04040013236E105016A028402D618803EB092B9201490B2A",
INIT_05 => X"B8E080000000005889AC41E04508A99070200E010001C1CA11803850C8000100",
INIT_06 => X"800A4CE301545001F40050216C09950004C2047BCF1C8090C02800C0120886B3",
INIT_07 => X"814A0080064C1F300020080182001A9E02C03400082002700000217294007101",
INIT_08 => X"000117088080990419002D86184A01018030430700802541420440022030041A",
INIT_09 => X"7030C30B885200D274004008080003C32A10A19090C02010E102294406168800",
INIT_0A => X"00602A01880980037109700C04C44C92A88DCC2211E44174112840880000060D",
INIT_0B => X"11C0D95C20C2030A003080030800308003080030800308003080018400184004",
INIT_0C => X"8304E02809832E6021002020404042000F00008400811824AD4007ECD9436261",
INIT_0D => X"0AFCE5D22A82B20000520100C801F8A07E103000A1285C84000418360C1B060D",
INIT_0E => X"0AFCFD8CB17E5B4F045557575E6EFBE3942C1040A41D660AFCE1CC1040A41E66",
INIT_0F => X"8E7FFBB385661C08D1455ABA91E6FF5FDFCC1040A41D660AFCF9CC1040A41E66",
INIT_10 => X"015F82C006C3AF31E64CB17E5A9655017F1FC73FAF1D61B1040294C58AD1FF5F",
INIT_11 => X"B95454005BAA36DCF8E519001BF80DEB3EE2020EA678189C6EC32881F7F75648",
INIT_12 => X"67D7EDFCA320037E81BD77D728A800B7546DBDFF12904747A351145FC53ABF8D",
INIT_13 => X"92B764225C57C97EBE76E1254F0C0D4514A84F5573FE9DBA4A38E247C522CC0E",
INIT_14 => X"BE84370001B6922070440556B15F7FABBC40151D7C747D8220673C3B9DB84B20",
INIT_15 => X"06C1B06C1B06C1B06C1B06C1B0491069068000004060300A005A01183F240014",
INIT_16 => X"6C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B",
INIT_17 => X"C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B0",
INIT_18 => X"B80EE173C2300F7DF16000000000000000000000000041B06C1B06C1B06C1B06",
INIT_19 => X"AAAAAA28A28A28AAAAAAA28A28A28A28A28A28A2910591505C104104B28BBECE",
INIT_1A => X"128944A25128944A25128944A25128944A2552A954AA5128944AAAA28A28A28A",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000128944A25128944A25128944A25",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFDFEF5D2A974BA082E954000000000000000000000000",
INIT_22 => X"0028B55002E82000087FFFFFFFFFFFFFEFF7FBEAB450804001EFAAD57FEAA087",
INIT_23 => X"7D168B55AAD17FFFF552EBFE00007FC00AA087FFFFFFFFFBFDF45AAD568B5508",
INIT_24 => X"087FD74AAAAFFFDF45A2D16AB55F7FFFFFFF00043DE10AA843DE00087FFFFEFF",
INIT_25 => X"A55042ABEF5D7FD75FFAAD540145AAD168A000004020AA5D7BE8B450051401EF",
INIT_26 => X"45FF8000010082A954BA00003DFEF085155400F78428BEFAA80000000804154B",
INIT_27 => X"1555D7FEAB55FF80175EF5D00020105D2A97400082E95555085168A10557FD75",
INIT_28 => X"00000000000000000000000000000000000000005D00020BA552A82000552A82",
INIT_29 => X"071EFB6DF7AE921C7FFFFFFFFFFFFFFFF7FBFDFFF5D2A954AA082A9242800000",
INIT_2A => X"1FAF55A2DF6DB7D1C002AB7D002A82028147FFFFFFFFFBFDFC7EBF5E8B550000",
INIT_2B => X"8E38E280871F8FC7E3D56AB6DBEDB7FFEF552AB8E38087FC2092087FFDFC7E3F",
INIT_2C => X"97FEFB6D1451471EF007BD0492B6F1F8F55AADF6DB7DE3F5FAFC708003DE28B6",
INIT_2D => X"A28407038140410492550A2ABC7497BD25FFAADF4516DBED16AA381C0A070824",
INIT_2E => X"D1C516FA28417BD5545E38E070280024904AA1C0438FD7005150438F78A2DBFF",
INIT_2F => X"92492A850105D2A80155417BEFB6DEB8E175FF5D0E05000492097428002E9557",
INIT_30 => X"4AA082A820AA000000000000000000000000000000000000000000000550A000",
INIT_31 => X"FF55A2D16AB550000175EFFFFBEAA00557FFFFFFFFFFFDFEFF7FBFFFEF552E97",
INIT_32 => X"C0000087BFDF45AAD568B55AAFBFDFEF55042ABEF002A800AA557FFDFEFF7FBF",
INIT_33 => X"16AB4500043DEAAFFAEAAAAA08516AB55A2D16ABEFFFFBFDFFF552AAAAAA007B",
INIT_34 => X"D568AAA5D2A97410007BFFFFF5551555EF087FC2000FFD56AB45A2FFFDFFFAAD",
INIT_35 => X"855400AAF7AEBDFEFA280154BA550400000552AA8B45087FC01EFA2FFD55EFF7",
INIT_36 => X"0804154BA082A975EF5D517DEAA007BD5545AAAA974AA0800020BA550028B550",
INIT_37 => X"00000000005D2E80010002A954005D2A82155087FFFFEFAAAA975EF5D2E97400",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000400000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(18),        -- Port A data input
DOA(0)   => data_read_a_lo_256(18),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(18),        -- Port B data input
DOB(0)   => data_read_b_lo_256(18),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_19_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"042200000000000041088001001AA00000000000000000000000500802000003",
INIT_01 => X"074018000024000000000404000000000A22000800000800004A200000000001",
INIT_02 => X"0000048002C405000000000006A84000000000200893C246A20000000020031A",
INIT_03 => X"082A58E411004B2000071000000981000C000000002045000200000000000000",
INIT_04 => X"200604000000001C0400001320000000162000002C4000026201201200090800",
INIT_05 => X"1020800000000058840200204000099070200E010001C0400000000000000000",
INIT_06 => X"0012048037805421402850001402498820022802400480405008901100A00102",
INIT_07 => X"00000000020C0130481204919200010C82000000000006002A548902A0020109",
INIT_08 => X"0001150800009900000005861840000000004301000B000000000001C1C00000",
INIT_09 => X"001F00002024B20002000000000002C300000000405000103010204000000000",
INIT_0A => X"00000000000000000000000000000040002000044000000000000000000002F0",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000420003B00000000000000000040012C80000000",
INIT_0D => X"45001A03C0825A0D20800000000018A006001000000000000000000000000000",
INIT_0E => X"450002131E01A1F6EA0A0020211146E069C2ACC01AE80045001D82ACC01AE800",
INIT_0F => X"1188340C3E1CFAD27CC2E004481020892282ACC01AE80045000582ACC01AE800",
INIT_10 => X"DEA03228D810007019931E01A1E5BA02802008C06F029D4C7B76639CEC0A0020",
INIT_11 => X"428AA3592000000206C2A4DAC00000008113C246A181C03FE4662A84575768DF",
INIT_12 => X"08201090549B5800000000261546B24000000000C53807E7CC06618018C51210",
INIT_13 => X"13F6A185A0A0168128411ACB800C0E108A0720288C011046B5986247C5452291",
INIT_14 => X"0000C220010808C10D9A92A74CD7CF4A080031B1515B212143D841431046B58A",
INIT_15 => X"00000000000000000000000000000000000000000000000000000118030004E0",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"3F0C7010C660C744192000000000000000000000000000000000000000000000",
INIT_19 => X"1861861861869A61861861861861861861861861A8208C4C1534D34C07208BBA",
INIT_1A => X"0984C26130984C26130984C26130984D26930984C26130984C261861861869A6",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE000000000000000000984C26130984C26130984C2613",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF552A974AA0004174BA0000000000000000000000",
INIT_22 => X"2E974BAA2FFFFE10087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974BA082E95400F7F",
INIT_23 => X"FFFFFFEFF7FBEAB450804001EFAAD57FEAAF7FFFFFFFFFFFFFFFFF7FBFDFFF55",
INIT_24 => X"002E82000F7FFFFFFFFFFFFDFEFA2D568B550004001EFAAAEA8ABA087FFFFFFF",
INIT_25 => X"5AAD16ABEF5D2ABFF55080402010087FFFFFFFFFBFDF45AAD568B55080028B55",
INIT_26 => X"BA087FFFFEFF7D168B55AAD17FFFF552EBFE00007FC00AAF7FFFFFFFF7FBE8B5",
INIT_27 => X"FFF00043DE10AA843DE00557FFDFEFA2D16AB55A2FFFDFEF5D2EBFE00AAFFFFE",
INIT_28 => X"0000000000000000000000000000000000000000AAFFFDF45A2D16AB55F7FFFF",
INIT_29 => X"954AA082A92428E3FFFFFFFFFFFFFFFFFFFFFFFEF552A974AA0000104AA00000",
INIT_2A => X"FFDFEFF7F5FAFC7492A974AAB6F5F8E101C7FFFFFFFFFFFFFFFF7FBFDFFF5D2A",
INIT_2B => X"A4A8AAA147FFFFFFFFFBFDFC7EBF5E8B550000071EFB6DF7AE92EBFFFFFFFFFF",
INIT_2C => X"2DF6DB7D1C002AB7D002A82028FFFFFFFEFF7F1F8FD7AAD16AB450000001FFBE",
INIT_2D => X"F7FBF8FC7E3F5EAB45B6DF6FBEF5D2AB8F7D000000010087FFDFC7E3F1FAF55A",
INIT_2E => X"7412ABFE28B6F5F8E820871F8FC7E3D56AB6DBEDB7FFEF552AB8E38087FC2092",
INIT_2F => X"55AADF6DB7DE3F5FAFC708003DE28B68E38E284971F8FC7AAD56DB6DBEF5F8FD",
INIT_30 => X"4AA0004000AA000000000000000000000000000000000000000000000B6F1F8F",
INIT_31 => X"DFEFF7FBFFFEF552E974AA082A820AAA2FFFFFFFFFFFFFFFFFFFFFDFEF552E95",
INIT_32 => X"EAA00A2FFFFFFFF7FBFDFFFFFD568B55002A954AAF7D568A00557FFFFFFFFFFF",
INIT_33 => X"56AB450004001EFFF842AAAA557FFDFEFF7FBFFF55A2D16AB550000175EFFFFB",
INIT_34 => X"7BFDF45AAD568B55AAFBFDFEF55042ABEF002A800AAF7FBFDFEFF7D56AB45AAD",
INIT_35 => X"52AAAAAA007BC0000FFFBE8B55AAD168B55F7FFFFFFF552AA8BEF08040200008",
INIT_36 => X"A2D57FFFFF7D568B45002ABDEAAFFD16AA0008516AB55A2D16ABEFFFFBFDFFF5",
INIT_37 => X"0000000000FFD56AB45A2FFFDFFFAAD16AB4500043DEAAFFAEAAAAA08556AB55",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000800000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(19),        -- Port A data input
DOA(0)   => data_read_a_lo_256(19),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(19),        -- Port B data input
DOB(0)   => data_read_b_lo_256(19),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_20_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000003",
INIT_01 => X"A65FF80000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000048002CC070000000000000000000000002FF86100200000000220002362",
INIT_03 => X"0000000000080F6000977060009B87A03C000000000000000000000000000000",
INIT_04 => X"3F2EFC040388137C3E20C477600142019E6000003CC0000A6601601A000B0000",
INIT_05 => X"102F91D10802ABFB80000021C8010FB0F0F43E1FE867DFC04400390210000220",
INIT_06 => X"90492261000080003400000010008000004203FE400580000000803000200006",
INIT_07 => X"401000004FFDFF28C4300C0010200100004000002AA001F00000000014000000",
INIT_08 => X"0801F5780259FB00000007BEFBC010002008FF7F00000000010018A81000041C",
INIT_09 => X"00000000020000000000000000000ADF00000020000000800000802830011023",
INIT_0A => X"0000000000000200020000000000000000000000000000000200200290000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"08120000B9090A700000200000004000000400000080002000407FED80000000",
INIT_0D => X"000079804000F00000000000C01FF8A7FE003000000004008100000000000000",
INIT_0E => X"0000798201000000100000000135386000401000010000000079801000010000",
INIT_0F => X"0185C300020004000010000000000252C7801000010000000079801000010000",
INIT_10 => X"00000010C1F30F300002010000080000000000CD8A0000400400000010000000",
INIT_11 => X"008040000000000292C0080000000000A5604000000284000818505200080000",
INIT_12 => X"0015E1B00100000000001496008000000000052B000048080000000000FC3600",
INIT_13 => X"80000000000002BA280000800830300000000000B8B400000401881010000000",
INIT_14 => X"00000000020020020001000040283024E6FB8604020080000383383B00000400",
INIT_15 => X"000000000000000000000004010201001003020200000000000127DBFF004000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"038200010089120104D204002000000000000000000000000000000000000000",
INIT_19 => X"B2CB2CB2CB2CB2CB2CB2CB2CB2C30C30C30C30C306982121A1E79E79A0700030",
INIT_1A => X"432190C86432190C86432190C86432190C86432190C86432190CB2CB2CB2CB2C",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000432190C86432190C86432190C86",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA0804020100000000000000000000000",
INIT_22 => X"2E954AA000400000F7FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0004174BAFFF",
INIT_23 => X"FFFFFFFFFFFFFDFEF5D2A974BA082E95400007FFFFFFFFFFFFFFFFFFFFFFEF55",
INIT_24 => X"A2FFFFE10FFFFFFFFFFFFFFFFFFFFFBFDFFF5D2E954BA007FC00BA087FFFFFFF",
INIT_25 => X"FF7FBFFF550800020BAAAD56AAAAF7FFFFFFFFFFFFFFFFF7FBFDFFF552E974BA",
INIT_26 => X"10087FFFFFFFFFFFFFEFF7FBEAB450804001EFAAD57FEAA007FFFFFFFFFFFFFE",
INIT_27 => X"B550004001EFAAAEA8ABA5D7FFFFFFFFFFFDFEFF7D56AB450000021EFA2D57DE",
INIT_28 => X"0000000000000000000000000000000000000000F7FFFFFFFFFFFFDFEFA2D568",
INIT_29 => X"974AA0000104AAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA08000500000000",
INIT_2A => X"FFFFFFFFFBFDFEF5D2E974AA000A07000E3FFFFFFFFFFFFFFFFFFFFFFFEF552A",
INIT_2B => X"71C50BA1C7FFFFFFFFFFFFFFFF7FBFDFFF5D2A954AA082A92428087FFFFFFFFF",
INIT_2C => X"7F5FAFC7492A974AAB6F5F8E10E3FFFFFFFFFFFFFFEFF7FBFFFFF552E974AA00",
INIT_2D => X"1C7FFFFFFFFFBFDFEFE3F5F8F450004050AABEDF6FABAEBFFFFFFFFFFFFDFEFF",
INIT_2E => X"50804021FFB6D57DE28147FFFFFFFFFBFDFC7EBF5E8B550000071EFB6DF7AE92",
INIT_2F => X"EFF7F1F8FD7AAD16AB450000001FFBEA4A8AAA497FFFFFFF7FBF8FC7EBD168B4",
INIT_30 => X"4AA080017410000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFDFEF552E954AA0004000AAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A95",
INIT_32 => X"820AA087FFFFFFFFFFFFFEFF7FBFDFFF5D2A974AA002E95410A2FFFFFFFFFFFF",
INIT_33 => X"FFDFEF5D2E954AA0051554BA557FFFFFFFFFFFDFEFF7FBFFFEF552E974AA082A",
INIT_34 => X"FFFFFFFF7FBFDFFFFFD568B55002A954AAF7D568A00AAFFFFFFFFFFBFDFEFFFF",
INIT_35 => X"000175EFFFFBEAA005D7FFFFEFF7FBFDFFFAAD16AB450804174AAFFFFFFEBAA2",
INIT_36 => X"F7FFEAB45A2D568B550804001EFF7D57DEBA557FFDFEFF7FBFFF55A2D16AB550",
INIT_37 => X"0000000000F7FBFDFEFF7D56AB45AAD56AB450004001EFFF842AAAA087BFDFEF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000000FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(20),        -- Port A data input
DOA(0)   => data_read_a_lo_256(20),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(20),        -- Port B data input
DOB(0)   => data_read_b_lo_256(20),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_21_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"4A302428B824900A128C090A5C1800261500213C005FE812D10420054085A202",
INIT_01 => X"081FFE3440B609703B0427F801A40B8115BC4F655300340288A40D30040E4DD8",
INIT_02 => X"04CA478082CC1740002019824E0203100640303FF8C0B31061096E21A1840814",
INIT_03 => X"8C329E9204020FE002577800405B87047D5042129D8D0248903200013290C800",
INIT_04 => X"3E7FFE02482553FC3C020277E128080A1E6000003CC0000A6601E03A8B0F0008",
INIT_05 => X"F43F8140000203FFC806C8A1C1048FF0F0E07E1F00F7FFC00024010000468310",
INIT_06 => X"08710C10015E083D01A24404786BE0014114C3FE4187A009A663A680100B3096",
INIT_07 => X"200800008FDFFF00290000100211019812E210488228000000900260026C6058",
INIT_08 => X"0EF1F5FA0041FF080AC707FEFBC110008420F7FF388B70A20389346FE8000580",
INIT_09 => X"917FC30010107688862A28C54518DBFF00020004C0A6044901112A0908AA0A30",
INIT_0A => X"006309044081A001B188300E20806520398C6021569249C4B3007127080806FF",
INIT_0B => X"904595123203040D9228D9228D9228D9228D9228D9228D9228D99146C9146C84",
INIT_0C => X"88042090068008003120000806001402504110C48002403601887FEF80022A51",
INIT_0D => X"26C0AC404E43032CA0C205880A7FFAB7FE01409400400C0594A4002200110008",
INIT_0E => X"26C0AC086A170250454004C6012280129B034A080C0B0016A0D20346080C0A80",
INIT_0F => X"0B064092D85938C0112144050224120C500346080C0B0016A0D2034A080C0A80",
INIT_10 => X"40702E058355458967E86A170220D1800093414B0414782E4B5000D81480809A",
INIT_11 => X"081B1545104135443306C35901024F88A88049062A747512B76783C5D040E080",
INIT_12 => X"40160040D86B202049B22198362A8A208279854400A036801480031401900800",
INIT_13 => X"0DD001C002D38334000914028354008301008C0CF1480245108C7640A0604032",
INIT_14 => X"AC0496022300233104662848808E191526205018030060540284FA0C0044022C",
INIT_15 => X"004010040100401004010040102090010008000001C0E010020007DFFFC06E60",
INIT_16 => X"0401004010040100401004010040100401004010040100401004010040100401",
INIT_17 => X"4010040100401004010040100401004010040100401004010040100401004010",
INIT_18 => X"FF7FFDF7FF3E3DFDF7E000000000000000000000000040100401004010040100",
INIT_19 => X"FBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBFFDFDFFFCF3CF3FFFEF9FEE",
INIT_1A => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFEFF7FBFDFEFF7FBFDFEFBEFBEFBEFBE",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0004000100000000000000000000000",
INIT_22 => X"2A954BA0004154BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080402010FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF552A974AA0004174BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"000400000007FFFFFFFFFFFFFFFFFFFFFFEF552E974BA0804000AAF7FFFFFFFF",
INIT_25 => X"FFFFFFDFEF5D2E974BA002E97400007FFFFFFFFFFFFFFFFFFFFFFEF552E954AA",
INIT_26 => X"BA087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974BA082E95400007FFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2E954BA007FC00BA5D7FFFFFFFFFFFFFFFFFFBFDFEF5D2A954AA002E974",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFBFD",
INIT_29 => X"954AA080005000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA00000200000000",
INIT_2A => X"FFFFFFFFFFFFFFF552A974BA0000174AAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0A000AAE3FFFFFFFFFFFFFFFFFFFFFFFEF552A974AA0000104AAF7FFFFFFFFFF",
INIT_2C => X"FFBFDFEF5D2E974AA000A07000007FFFFFFFFFFFFFFFFFFFFDFEF552E954BA08",
INIT_2D => X"1C7FFFFFFFFFFFFFFFFFFBFDFEF5D2A974BA002A95400087FFFFFFFFFFFFFFFF",
INIT_2E => X"F552E974BA0020924BA1C7FFFFFFFFFFFFFFFF7FBFDFFF5D2A954AA082A92428",
INIT_2F => X"FFFFFFFFFEFF7FBFFFFF552E974AA0071C50BA557FFFFFFFFFFFFFFFF7FBFDFF",
INIT_30 => X"4BA000002000000000000000000000000000000000000000000000000E3FFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2A954AA080017410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"000AAF7FFFFFFFFFFFFFFFFFFFFFFFEF552A974BA0000174BAFFFFFFFFFFFFFF",
INIT_33 => X"BFDFEF5D2A954BA082E800AAA2FFFFFFFFFFFFFFFFFFFFFDFEF552E954AA0004",
INIT_34 => X"7FFFFFFFFFFFFFEFF7FBFDFFF5D2A974AA002E95410087FFFFFFFFFFFFFFFF7F",
INIT_35 => X"52E974AA082A820AA557FFFFFFFFFFFFFEFF7FBFFFFF552E954BA002E9741008",
INIT_36 => X"FFFBFDFEFF7FFFFFEF5D2A974BA0000020AA557FFFFFFFFFFFDFEFF7FBFFFEF5",
INIT_37 => X"0000000000AAFFFFFFFFFFBFDFEFFFFFFDFEF5D2E954AA0051554BA5D7FFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(21),        -- Port A data input
DOA(0)   => data_read_a_lo_256(21),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(21),        -- Port B data input
DOB(0)   => data_read_b_lo_256(21),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_22_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"5290F4CDE914905A14A43D33F488243E17122300F55FEB189B343A1140548380",
INIT_01 => X"A94007B259F6A975386262000C344BA9573C6FF57B18A5FB0ABFCD3C2C5F4F0C",
INIT_02 => X"D56B4302AC01005111011BD506AA5205274056900596A539584E2E6DFE4B2418",
INIT_03 => X"6B03F2F6151A2081F24001E8400008F401CB10C6594423C8923AD6B55AD0EB5A",
INIT_04 => X"8001023D37E50880436200808BC8492A0089249600101100008087248B64426E",
INIT_05 => X"A51035B41C0A88046CAEE8C23C08E040011C0020F8882001102D620A06D68301",
INIT_06 => X"B93FF975CF7889D085E997A2144E8FC2060B880081A26DCD4047EFF9EF018980",
INIT_07 => X"283800AA500200E8024AD03546A3262FB5AA5542A882040C7A64CBD64065F028",
INIT_08 => X"141008801018040E48D500400015805060040080A2A0F4A82381B4000A0905A0",
INIT_09 => X"4D0000002126F30C902A29C54539C020E11810098D4067EFF9FF284D483E2AB4",
INIT_0A => X"1400006100003202D040050220103D2A512C6A8C4F0008AA800470370000A000",
INIT_0B => X"013456520CA09281C2A81C2A81C2A81C2A81C2A81C2A81C2A81C9540E1540E00",
INIT_0C => X"A1402A13C0A10A893165281A1C2A7283516344C594A85536B1AD800214202C50",
INIT_0D => X"3C70FC20515808A0100820112300011000287B071105034406950A0285014280",
INIT_0E => X"3C70FC48E11CFC48400184CE0D6783139B0959A41606003C70FA0958AC160480",
INIT_0F => X"0D87E8B3B811B52048B10E0402AE1606D80958AC1606003C70FA0959A4160480",
INIT_10 => X"80F84E0185594581E088E11CFC38414020DD42CF909D7E0A551C02180300C0DD",
INIT_11 => X"441154C258012D86F3044A3133004A99BD8455300654458A1D588C4061403000",
INIT_12 => X"A096A240894626600953379822A984B0025B0DEC0345C9200680027181B44887",
INIT_13 => X"E2404160035482BE521C2C04A90783C18000D610B9D8070B12B1A2A62040202A",
INIT_14 => X"304244A91102C93A2D608D2A258DF8034284200C050070E40C80620C870B02C4",
INIT_15 => X"4411044110441104411044110466C440446CA06951D4EA801000980400646002",
INIT_16 => X"0100441104411044110441104411044110441104411044110441104411044110",
INIT_17 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_18 => X"FE8FF1F7DEBDDF7DF7D05122890000000003FFFFFFFF90040100401004010040",
INIT_19 => X"79E79E79E79E79E79E79E79E79E79E79E79E79E7BFFDFD7DDDF7DF7DF7DFBFDE",
INIT_1A => X"3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE79E79E79E79E",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE000000000000000003F9FCFE7F3F9FCFE7F3F9FCFE7F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0800000000000000000000000000000",
INIT_22 => X"2E974AA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000400010FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E954AA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"0004154BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA000015400FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF552A974AA0800154AAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA",
INIT_26 => X"BAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0004174BAFFFFFFFFFFFFFFFFF",
INIT_27 => X"FEF552E974BA0804000AAA2FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0000174",
INIT_28 => X"0000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040001000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E954AA000402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0417410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080005000FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF552A974BA0000174AAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA00",
INIT_2D => X"E3FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0804154BAF7FFFFFFFFFFFFFFFFF",
INIT_2E => X"F552E954BA000E124BAE3FFFFFFFFFFFFFFFFFFFFFFFEF552A974AA0000104AA",
INIT_2F => X"FFFFFFFFFFFFFFFFDFEF552E954BA080A000AAA2FFFFFFFFFFFFFFFFFFFFFFFE",
INIT_30 => X"4BA080400010000000000000000000000000000000000000000000000007FFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"17410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000400010FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF552A954BA000415400FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954AA0800",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFEF552A974BA0000174BAF7FFFFFFFFFFFFFFFFFFF",
INIT_35 => X"52E954AA0004000AAA2FFFFFFFFFFFFFFFFFFFFFDFEF552E974AA0804174AAF7",
INIT_36 => X"FFFFFFFFFFFFBFDFEF5D2E954BA002A820BAA2FFFFFFFFFFFFFFFFFFFFFDFEF5",
INIT_37 => X"0000000000087FFFFFFFFFFFFFFFF7FBFDFEF5D2A954BA082E800AAAAFFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000000FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(22),        -- Port A data input
DOA(0)   => data_read_a_lo_256(22),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(22),        -- Port B data input
DOB(0)   => data_read_b_lo_256(22),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_23_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"EF20906D902424807BC8241BC81801B97D38AD3C0800103362A6741C80A12A02",
INIT_01 => X"001FFF8409F089003B4422000D80C80106804A7951C5B9D1C828043EA28838F9",
INIT_02 => X"028406A002DC176444683862400003111001303FFC00F240D50146013B300500",
INIT_03 => X"001B243004080FE000177003145F87017D584B10D804034800200200A1008008",
INIT_04 => X"BEFFFC0248005FFC3C18A2FFE12222425E600000BDC0800AEE01E81A100F0A00",
INIT_05 => X"D03F8000000003FF810640A1C0008FF2F0E17E1F02FFFFC80100004044800080",
INIT_06 => X"800264B4854650040123428C204BF40F439647FF4807E189A477EF81DF0AF116",
INIT_07 => X"01000000FFDFFFE800401005C0A0008F86C60840AAAA100C68D1810C9F4A0020",
INIT_08 => X"1BE1F5F80003FF0002021FFEFBC80000000077FF184B03010004002FE1F29002",
INIT_09 => X"907FC308181204800600000000001BFFA800808189A657EF81DD0C00079CC800",
INIT_0A => X"0063090442A18001B188300C48907120AC810033149249C433200180082A06FF",
INIT_0B => X"9A41C1443243050C1010C1010C1010C1010C1010C1010C1010C1008608086084",
INIT_0C => X"000082A00600200080000500C000400800601200000254A000007FEFC1030221",
INIT_0D => X"0A9080400E0BF30C20CA858E087FFABFFE01409780214EE49620001000080004",
INIT_0E => X"0A908044294700701641005218521210150E5789F90A000A90800E5F81F90880",
INIT_0F => X"0E0220036864A7DCA190440301E2105C000E5F81F90A000A90800E5789F90880",
INIT_10 => X"C1400500C6CE5400032429470068924010164302048156305D66F8701681000E",
INIT_11 => X"2E0CCB0500013440600339C800004D8018000857A82920CE8CB220C81400A180",
INIT_12 => X"220344406739000009B0030019960A00026880C0422C52B01700044901488822",
INIT_13 => X"85C811A010428104128996465ADA020180804A040108A2658217C4008060300C",
INIT_14 => X"BE0692020328CA0028042054A92771C50FC070109000C1C819078280A265920E",
INIT_15 => X"020080200802008020080200800800200200000000000008004807DFFF000470",
INIT_16 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_17 => X"0080200802008020080200802008020080200802008020080200802008020080",
INIT_18 => X"0000000000000000000000000000000000000000000000802008020080200802",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000",
INIT_22 => X"2E974BA080002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E974BA000400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000400000FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF5D2E954AA080000010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA",
INIT_26 => X"10FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080402010FFFFFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2A954BA000015400FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA0804000",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E974BA080002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF5D2E954AA000402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA00",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080002010FFFFFFFFFFFFFFFFFFF",
INIT_2E => X"F5D2A954BA080407000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080005000",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF5D2A954BA000417410FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA080402000000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"02000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000010FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF5D2E974AA000402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0000",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000400010FFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"D2A954AA080017410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954AA080002000FF",
INIT_36 => X"FFFFFFFFFFFFFFFFFF552A954BA080015410FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_37 => X"0000000000F7FFFFFFFFFFFFFFFFFFFFFFFFF552A954BA000415400F7FFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000000FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(23),        -- Port A data input
DOA(0)   => data_read_a_lo_256(23),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(23),        -- Port B data input
DOB(0)   => data_read_b_lo_256(23),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_24_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100600007FFF000080108004000800020000840041000080808",
INIT_02 => X"0000068002CC07400000090C080002000000103FF811F150231000520ABE4404",
INIT_03 => X"8428180000080FE000177000001B87003D4000000E8B84010020000000008000",
INIT_04 => X"3E2FFC024800137C3C000077E00000001E6000003CC0000A6601E01A000F0200",
INIT_05 => X"103F8000000003FF80000021C0000FF0F0E03E1F0067FFC00000000000000000",
INIT_06 => X"00132412079001AD00810005E8000001401643FE4007E5501AA00000DC8C3006",
INIT_07 => X"000000000FDFFF62695A5685C094831D966000008002100C2040A178B600C240",
INIT_08 => X"08E1F5F80001FF00000007FEFBC00000000077FF000B00000000002FE0000000",
INIT_09 => X"107FC300000000000600000000001BFFA0000005501AA00000CE200000940000",
INIT_0A => X"00630104408180012188300C00814080008000010012414433000100080806FD",
INIT_0B => X"904181003003000C1000C1000C1000C1000C1000C1000C1000C1000608006084",
INIT_0C => X"00000080060000000000000012002C00000000000000000000007FEF80020201",
INIT_0D => X"440082404E0B332CA2C20188087FFAB7FE000082000000008220000000000000",
INIT_0E => X"4400824903210308074084210002460402009280010D80440084009280010F00",
INIT_0F => X"800A2400401A0C82183248060010280C20009280010D80440084009280010F00",
INIT_10 => X"C0A078160000404A0469032102981380202080026420020D06C002A08481C020",
INIT_11 => X"00164F400860000824059AD01802000208104817B00011306B2D9B0DD5082080",
INIT_12 => X"41021800B35A0300400041202C9E8010C0001040C5836CC01780018601030088",
INIT_13 => X"DB1011E000A140058220004AEFFC8101810021084301880030A8B77400603011",
INIT_14 => X"8C063C0220002201490418082010A57263E010000201033016085A40880030A1",
INIT_15 => X"000000000000000000000000000000000000000000000000000007DFFF0006E0",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"F6E7CC1132CDB444199000000000000000000000000000000000000000000000",
INIT_19 => X"79E79E79E79EFBEFBEFBEFBEFBEF9EF9EF9EF9EFA69861219575D75FF2D0AEEA",
INIT_1A => X"0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1EFBEFBEFBE79E",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE000000000000000000783C1E0F0783C1E0F0783C1E0F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020100000000000000000000000",
INIT_22 => X"2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"080002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_26 => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000400010FFFFFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2E974AA000400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0004000",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040201000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF5D2E974BA080002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFF",
INIT_2E => X"F5D2E974AA000400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF5D2E974AA000400000FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA080402010000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"00010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000010FFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002010FF",
INIT_36 => X"FFFFFFFFFFFFFFFFFF5D2E974AA000002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_37 => X"0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000402010FFFFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(24),        -- Port A data input
DOA(0)   => data_read_a_lo_256(24),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(24),        -- Port B data input
DOB(0)   => data_read_b_lo_256(24),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_25_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100200002000000080100004000000020000800041000080808",
INIT_02 => X"0000068002CC474000000800000002000000103FFCE302008000000880844A04",
INIT_03 => X"00000101C0200FF004177800081B87003D400000080000000020000000008000",
INIT_04 => X"3E2FFE024820137C3C004077F01000001E7249213CC1264A660DF05A000F9000",
INIT_05 => X"103F81C1002203FF80000021C1140FF8F0E03E1F0067FFE04800258280010052",
INIT_06 => X"80480AE20000000100000001C8608001401643FE4007C00000000000CC083006",
INIT_07 => X"280800000FDFFFEA4050140540B00100840000080002A00C2040810000000010",
INIT_08 => X"C8E1F5FA21C9FF80040007FEFBE031018C31F7FFBAEBC0020008086FE0000100",
INIT_09 => X"107FC301800000000600000000001BFFE00301000000000000CC020000140000",
INIT_0A => X"0077330C4889CC292588300C0080400000800001001243443B000100880806FD",
INIT_0B => X"904189003003000C1000C1000C1000C1000C1000C1000C1000C1000608006084",
INIT_0C => X"8B04228026824100000000000000000000000000000004A000007FEF80020201",
INIT_0D => X"400000400E03C30C20C2818C087FFAB7FE01409700C10007962418220C110608",
INIT_0E => X"4000000001010000004000000000400400001200000800400000001200000800",
INIT_0F => X"0008000000000480000040000000200000001200000800400000001200000800",
INIT_10 => X"0000001001000002000001010000100000000000202000000440000000800000",
INIT_11 => X"0000410000000008000008400000000200000806300400000820000020004880",
INIT_12 => X"0000080001080000000040000082000000001000000040800800000000020008",
INIT_13 => X"8100000000000000802000000840000200040000020008000000840000804000",
INIT_14 => X"8C04100200000200000610000000210000000018140000000008000008000000",
INIT_15 => X"04411044110441104411044510629041040D180400000010028047DFFF800C60",
INIT_16 => X"4411044110441104411044110441104411044110441104411044110441104411",
INIT_17 => X"4110441104411044110441104411044110441104411044110441104411044110",
INIT_18 => X"196A8C5A2932EC15DA080800002FFFFFFFFFFFFFFFFFC1104411044110441104",
INIT_19 => X"92492492492410410410410410410492410492412000531215A69A6BFBA2894A",
INIT_1A => X"B158AC562B158AC562B158AC562B1588C46231188C46231188C4924924924924",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000B158AC562B158AC562B158AC562",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000",
INIT_22 => X"2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF5D2E974BA080400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_26 => X"10FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0800000",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400000FFFFFFFFFFFFFFFFFFF",
INIT_2E => X"F5D2E974BA080000010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA080402000000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"02000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400000FF",
INIT_36 => X"FFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_37 => X"0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000000FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(25),        -- Port A data input
DOA(0)   => data_read_a_lo_256(25),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(25),        -- Port B data input
DOB(0)   => data_read_b_lo_256(25),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_26_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"E9264EAB20190CA3BA4997AA9002AE9C001006B0778015CFA17E0811039879C7",
INIT_01 => X"F1FFF9BB1F773C7F9BB07DFFFDD863FC5FFF3FEFFBBF9FFB22FFFBC7B9F30686",
INIT_02 => X"9B3184F8AFDEAF300029E4E300FC78A6258548EFFA71C00172082400003A2161",
INIT_03 => X"0213C3FDFFFC7F74FFBF737A603B87FEBE1A5294F65628A0001B9CE6CC606E73",
INIT_04 => X"7E2EFEBF6FFEB37C3FF3017776FFCDA43E7B6DFD7DEBFD8E6F5F78DF0BFBD644",
INIT_05 => X"902F87C74E8CCFFBB6FF70E1FE61FFBDF0FEBE1FFD67DFFEFFBDA7F7FED50870",
INIT_06 => X"213246200BCC8920360C1831CD7DF60A244B9BFEE00589DDBCEFEDC1DFA08957",
INIT_07 => X"B1D4223B4FFDFF21CC721C85DCE1458E8782484020A2C1FCA3468D77E0000300",
INIT_08 => X"2C05FD7BC471FBD13D980FBEFBEBF30B8D79FF7F451F33CFD60FE8FFFDF54003",
INIT_09 => X"19FFC71FEFED7B251E35768E8ED6BFDF3EB3EBF9DDBCE7FDC1DF8A760F3EACC0",
INIT_0A => X"56F7730ECCDBDF152199F51EDDCDEBCFF589807B7096CD4CF73AC1FC98884FFF",
INIT_0B => X"B867D3683A03A40F78C0D78C0D78C0D78C0D78C0D78C0D78C0D7A606BC606B8C",
INIT_0C => X"DFBFF5EB36DFE51FC3A80D73D840303983EE7F0EA03BDA680137FFFDFFD7E681",
INIT_0D => X"3F0080425E6BFF8DB0DAE19C09FFFFE7FE3EBEA8EB7AFEE5C9AEBD7F5EBFAF5F",
INIT_0E => X"3F00800DEC010280004000F808020290100FA2F60008003F00800FA2F6000800",
INIT_0F => X"00023002007BC0A14E00400003B8000D000FA2F60008003F00800FA2F6000800",
INIT_10 => X"01E0320007204008040DEC010300100000F600020581003F604D0700008000EE",
INIT_11 => X"201F21A2C40039006807C46426040E101A0259DFE82011A311AA042016040080",
INIT_12 => X"80020048F88C84C101C203403E434588007200D047F00090200007E0010009B0",
INIT_13 => X"0109000003E2000416C0804FE04140E80000F808010AB02033AC048A2A00003D",
INIT_14 => X"FFAFD082003B032FB987E04021D481D4000419060201E1A000044300B02033E8",
INIT_15 => X"AFEBFAFEBFAFEBFAFEBFAFEFFBFBFBFBBFCFBB0FFDFEFFEF2DFFFFFBFF802FFD",
INIT_16 => X"FEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBF",
INIT_17 => X"EBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFA",
INIT_18 => X"F491E166CC8553F86EDB5C88646FFFFFFFFFFFFFFFFFEBFAFEBFAFEBFAFEBFAF",
INIT_19 => X"1861861861861861861861861861869A69A61861AFBD54D5F871C71D475B15BC",
INIT_1A => X"0984C26130984C26130984C26130984C26130984C26130984C26186186186186",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE000000000000000000984C26130984C26130984C2613",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000",
INIT_22 => X"2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_26 => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFF",
INIT_2E => X"F5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA080402000000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"02010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_36 => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_37 => X"0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(26),        -- Port A data input
DOA(0)   => data_read_a_lo_256(26),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(26),        -- Port B data input
DOB(0)   => data_read_b_lo_256(26),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_27_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"00080A40000A41248002029000050A088000008242A0004404480002000A1155",
INIT_01 => X"F1FFF1C11F781C129C107DFFFE0860941E81258CA2B71C2220EC1B86E1A00002",
INIT_02 => X"183080988B2EAE00002BE001117C78C6848140CFFA0000800042008000011081",
INIT_03 => X"000003FDF3E47C74F7BCF36A203A47F6B8184210B6160820001318C60C204C63",
INIT_04 => X"7E28FEBF6FEEB3723F71017476DFC524397B6DF572EB6C8E175E70D90F539600",
INIT_05 => X"000F86064C8DDFE3B6FF50D1FC61DE39C8FCB91FF9671FE6B68984B5BCE40834",
INIT_06 => X"0000000800000042020C18300520620A80231BFE200181092CE7ED80DFC00147",
INIT_07 => X"8AC4AA3B0FD1FF201044110560884000840200520002080C23468D0300000282",
INIT_08 => X"2005F0784411E390A4880E3DF7E2FB0B8E717C7F411F3BC6D60B60FFDDE44001",
INIT_09 => X"18FFD757E7ED7A211E81C09818109E1F16B16B71092CE7ED81CF403601228C40",
INIT_0A => X"46FF730E5CCBCD55219AB55F0DEFABC7054880693016DD4C755AC16C1A884FFE",
INIT_0B => X"BC63F1683803C00E3440C3440C3440C3440C3440C3440C3440C3C2061A2061AD",
INIT_0C => X"56BF55CB165EC51D41880FA3F040202883B475062033186801137FF1BAD6F281",
INIT_0D => X"3B0000421E2B0F2E2AE215C808FFFA47FE62BAA86B1AB268E92AB56D5AB6AD5B",
INIT_0E => X"3B000025EC010080004000F808000098100F22520008003B00002F2252000800",
INIT_0F => X"00001042006BC0810600400003B80001002F22520008003B00002F2252000800",
INIT_10 => X"01E032000620000C0405EC010100100000F6000001C1003760410500008000EE",
INIT_11 => X"201D2120840039000817444404040E10020218DE282010A311AA002002040080",
INIT_12 => X"8000000AE888808101C20040BA4241080072001027F00080200007E0000001F0",
INIT_13 => X"0101000003E2000007C0800FE04040280000F8080002F02023AC04080A00003D",
INIT_14 => X"DDAFD082001B03249887E04001D481D4000009020201E1A000040100F02023E8",
INIT_15 => X"ADAB6ADAB6ADAB6ADAB6ADAB6BF1EBDABD8E270BF84A25C6ACB777E3FF800C6D",
INIT_16 => X"DAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6",
INIT_17 => X"AB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6A",
INIT_18 => X"100481CA860402104A471688747FFFFFFFFFFFFFFFFFAB6ADAB6ADAB6ADAB6AD",
INIT_19 => X"0000000000000000000000000008200000000000200072F210000001490E2168",
INIT_1A => X"A05028140A05028140A05028140A050080402010080402010080000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000A05028140A05028140A05028140",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000",
INIT_22 => X"2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_26 => X"10FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFF",
INIT_2E => X"F5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA080402000000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"02000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FF",
INIT_36 => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_37 => X"0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000000FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(27),        -- Port A data input
DOA(0)   => data_read_a_lo_256(27),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(27),        -- Port B data input
DOB(0)   => data_read_b_lo_256(27),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_28_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"02200AA400180030808802A900002A08001280A08A801044104A1000001818C3",
INIT_01 => X"50A00011460214428114180000882214413D0A71592A01D92213D28005210202",
INIT_02 => X"8A54800A210200111100C2110054289220810440030404010844000444410001",
INIT_03 => X"4200040822D4500001E0000028000002000211842010092000018C6295200631",
INIT_04 => X"00400000000B8000000140000005840C00000040002008808100048100100044",
INIT_05 => X"0000222200244400135110000135100000000000000000024CA0A01018000320",
INIT_06 => X"A004912008208040024489121144080400081000200008104000000020000041",
INIT_07 => X"A85800994000000A0200802004204420210001022AA8A0001122448142491008",
INIT_08 => X"0414000201800004080A000000124058200408000880004440004080160C4100",
INIT_09 => X"0080000206CB0821082B694D4D29400002002038104000000020003204000440",
INIT_0A => X"12000843066021001400040024440245400082D022040000400800081022C000",
INIT_0B => X"0002002C004001036050160501605016050160501605016050160280B0280B00",
INIT_0C => X"0012400810080414C0A800310840102182C62302A0194C08001680100E4040A0",
INIT_0D => X"05000002003004208208841401800040000A0000200814004198000400020001",
INIT_0E => X"0500000004000080000000000000028000002052000000050000002052000000",
INIT_0F => X"0000300000004001060000000000000900002052000000050000002052000000",
INIT_10 => X"0000000001200000000004000100000000000000050000002001050000000000",
INIT_11 => X"00002020840000004800040404040000120200A9000000010000002002040000",
INIT_12 => X"0000004800808081000002400040410800000090001000002000000000000910",
INIT_13 => X"0001000000000000144000010000402800000000000A1000010000080A000000",
INIT_14 => X"0080000000110006B08140000040000000000902000000000000410010000100",
INIT_15 => X"0080200802008020080200802101210810C39A66A90A85420413A82000000204",
INIT_16 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_17 => X"8020080200802008020080200802008020080200802008020080200802008020",
INIT_18 => X"110A00246972BD89A40A0C22E100000000000000000000200802008020080200",
INIT_19 => X"82082082082082082082082082082082082082080D35050758C30C31DE21102C",
INIT_1A => X"B0582C160B0582C160B0582C160B0580C06030180C06030180C0820820820820",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000B0582C160B0582C160B0582C160",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000",
INIT_22 => X"2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_26 => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFF",
INIT_2E => X"F5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA080402000000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"02000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_36 => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_37 => X"0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000000FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(28),        -- Port A data input
DOA(0)   => data_read_a_lo_256(28),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(28),        -- Port B data input
DOB(0)   => data_read_b_lo_256(28),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_29_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"79964E4BA01DACAB9E659792D00AAE160002829C7FDFEFCEE97C2815039D70C3",
INIT_01 => X"50BFF9AB0775343F9AB01DF80D5821FC0FFF3FEFD1AF9FF1207FFBC7B9720586",
INIT_02 => X"0D15846807D207200021C4E200D428A2018408600271C000720A0000003A2161",
INIT_03 => X"0002C009EEFC5F10F9B70178681B80FA3E000100765029A00019084345606421",
INIT_04 => X"3E6E023D27DA937C03E3407712E5CDA41E0924DC3D20B98AE905189F0BF8C000",
INIT_05 => X"902003C30E0447F877F930203E213F8CF01E3E00FC67C03A4D9C87525E510160",
INIT_06 => X"0012460003CC002036040811D919F402244293FEE00400CCB46BA4C164A08857",
INIT_07 => X"914800110FFC0001CC320C81D841418E82800100000041FCA1428575A0001108",
INIT_08 => X"0805FD0180E1F8C1111A0782082B50080508FF00048B124D4005C8AFF4154102",
INIT_09 => X"0180000ABFEF89250815568A8AD6ABC02A02A0B0CCB463B4C0748A720B1EA4C0",
INIT_0A => X"021410028450530014014002D445624DB481806A62840800C22800B8900042FF",
INIT_0B => X"0806522C0A40A50268D0068D0068D0068D0068D0068D0068D006A68034680300",
INIT_0C => X"8912E0A83289641F42A80561D040203182AC3D0AA0118A080036FFFC4F4164A0",
INIT_0D => X"050080424069F5A51250648801BFFFE0003E3E00A0685A85410C0816040B0205",
INIT_0E => X"050080080400028000000000000202900000A0F600000005008000A0F6000000",
INIT_0F => X"00023000001040214E0000000000000D0000A0F600000005008000A0F6000000",
INIT_10 => X"000000000120400800080400030000000000000205800008200D070000000000",
INIT_11 => X"000220A2C400000068008424260400001A0241DAC80001010000042016040000",
INIT_12 => X"00020048108484C10000034004414588000000D04010001020000000010009B0",
INIT_13 => X"000900000000000416C00041000140E800000000010AB0001100008A2A000000",
INIT_14 => X"A282C0000033010FB181E00020400000000419060000000000004300B0001100",
INIT_15 => X"02C0B02C0B02C0B02C0B02C4B12B312912831A27FCFE7FFB175B6FF800802594",
INIT_16 => X"2C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B",
INIT_17 => X"C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B0",
INIT_18 => X"EE7FFDF7FE783FFDFFEA0C00602FFFFFFFFFFFFFFFFFC0B02C0B02C0B02C0B02",
INIT_19 => X"BEFBEFBEFBEFBEFBEFBEFBEFBEEBAEBAEBAEBAEBBFFDF9FBEFFFFFFEBBCF9F96",
INIT_1A => X"FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFBEFBEFBEFBEF",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000FBFDFEFF7FBFDFEFF7FBFDFEFF7",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000",
INIT_22 => X"2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_26 => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFF",
INIT_2E => X"F5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA080402000000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"02000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_36 => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_37 => X"0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(29),        -- Port A data input
DOA(0)   => data_read_a_lo_256(29),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(29),        -- Port B data input
DOB(0)   => data_read_b_lo_256(29),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_30_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"FF9FE1F7FFBFFFFDFFD000000000000000000000000000000000000000000000",
INIT_19 => X"79E79E79E79E79E79E79E79E79E79E79E79E79E7AFBD75F5FDF7DF7FF7FFBFFE",
INIT_1A => X"3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE79E79E79E79E",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE000000000000000003F9FCFE7F3F9FCFE7F3F9FCFE7F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000",
INIT_22 => X"2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_26 => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFF",
INIT_2E => X"F5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA080402000000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"02000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_36 => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_37 => X"0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(30),        -- Port A data input
DOA(0)   => data_read_a_lo_256(30),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(30),        -- Port B data input
DOB(0)   => data_read_b_lo_256(30),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_31_6 : RAMB16_S1_S1
generic map (
INIT_00 => X"129000008004A00804A40000400800020000000C005FEA005800200400050100",
INIT_01 => X"A15FF18019700810180065FFFC0040801E80258CA2951C2200EC0906A0804140",
INIT_02 => X"146000808A0C060444692000402850040400408FF80000000010000000004000",
INIT_03 => X"000003F5D1202C70F654716A001A07F438184210960600000012108518004842",
INIT_04 => X"3E28FE3F6FE513703F70007472DA4128187B6DB530C1240A060C70580B439200",
INIT_05 => X"000F84040C088BE3E4AE40C1FD04CE38C0FC381FF8671FE01009048084C40010",
INIT_06 => X"0000000000000008000810200420620E00030BFE000181092CE7ED80DF800106",
INIT_07 => X"000000220FD1FF200040100540800000840200408002000C2244890200000200",
INIT_08 => X"0011F0780011E38004800E3CF3E0B1118C31747F000B33820209206FC9E80000",
INIT_09 => X"187FC301B124F2001600000000001A1F00110101092CE7ED81CF000401228800",
INIT_0A => X"0477330C4889CC012188310E08812982050800A91012494C31004124080886FE",
INIT_0B => X"9861D1403803800C1000C1000C1000C1000C1000C1000C1000C1800608006084",
INIT_0C => X"020400830602410901000D02D0002008012054040022102001017FE190022201",
INIT_0D => X"3A0000401E030B0C20C20188087FFA07FE203A80010002608030102008100408",
INIT_0E => X"3A000005E8010000004000F808000010100F02000008003A00000F0200000800",
INIT_0F => X"00000002006B80800000400003B80000000F02000008003A00000F0200000800",
INIT_10 => X"01E03200060000080405E8010000100000F600000081003740400000008000EE",
INIT_11 => X"201D0100000039000007404000000E1000001846282010A211AA000000000080",
INIT_12 => X"80000000E808000001C200003A0200000072000007E00080000007E0000000A0",
INIT_13 => X"0100000003E200000280800EE04000000000F8080000A02022AC04000000003D",
INIT_14 => X"9C06D082000A03200806A040019481D4000000000201E1A000040000A02022E8",
INIT_15 => X"0401004010040100401004010060C040040C200950402090128057C3FF800C60",
INIT_16 => X"4010040100401004010040100401004010040100401004010040100401004010",
INIT_17 => X"0100401004010040100401004010040100401004010040100401004010040100",
INIT_18 => X"000000000000000000001000802FFFFFFFFFFFFFFFFF81004010040100401004",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000",
INIT_22 => X"2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_26 => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFF",
INIT_2E => X"F5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA080402000000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"02000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_36 => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_37 => X"0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(31),        -- Port A data input
DOA(0)   => data_read_a_lo_256(31),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(31),        -- Port B data input
DOB(0)   => data_read_b_lo_256(31),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_0_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"ED39BA795990D275FB4A6E96ACC4731DEA4598B0AFB54867F6EE4618C3749803",
INIT_01 => X"58A0047C8607844847CA180001E4A2404042106208408208C2002069161734B3",
INIT_02 => X"8B1EC9562121F8051500147A0E5629A302CF28400615F5787B09FBF999BB1EFD",
INIT_03 => X"404EFC0A2AD6100F01A88E851CE47803C280110521898F6996088862C7B22221",
INIT_04 => X"C0D001C0100AEC83C008E7880D01A64661800002C21A52C590D2012194804844",
INIT_05 => X"650002C3F08754001B51981E007910070F01C1E003980015A204C22F32328BAF",
INIT_06 => X"BCDA4677CAEE7CF5BB870E1DDB9889C5FBFC440129A0604442180238203F70C1",
INIT_07 => X"7AAE0088B02000C2EC3A0E829836E0AF3325372E2AA8FDF3C18306758B24197A",
INIT_08 => X"D7E40002F7AE005FFB4730010411400A61080000F7F4C464B58294901606D5A5",
INIT_09 => X"C4801C40469B0CA9881A28C141118000C5A85A60444210123820B43B40804274",
INIT_0A => X"400800219010107ED453C041B13216656074EA560F0092A24856B05312226900",
INIT_0B => X"27122C3E04E03383E2781EA781E2781EA781E2781EA781E2781C33C0613C0E29",
INIT_0C => X"74EB1F50D0758A9650E520610A6A57A5529E2B439499CF96B086000000B09870",
INIT_0D => X"04F07E024108F4E28638EC57250004480155C1375A97A9121F8BA749D3A4E9D2",
INIT_0E => X"04F07E42177EFDF8570184071575970F8FC07D5BFF078004F07E007D5BFF0780",
INIT_0F => X"8F85ECB1FE047F5FB7B30E0700461E5AF8007D5BFF078004F07E007D5BFF0780",
INIT_10 => X"C0184D07C1DF15C7E3E2177EFDF8C3C03009C3CDD47C7F403FB3FDF89701C011",
INIT_11 => X"4F80FE659C6104C6D7103F9D1D064189B5924418D65FE45DEE55BBEDE34CF900",
INIT_12 => X"6395F64207F3A3A1483136B881FCCB38C2098DACA01FFF603F80001F80FDC81F",
INIT_13 => X"FED151E01015C3BB507D3F811FBEC32B81840714F8D91F4FC513F37C8AE07002",
INIT_14 => X"61692F293185D8D724E15D3FCC6B7C236FE0691A9500125C1F83F8CC1F4FC507",
INIT_15 => X"E93A4E93A4E93A4E93A4E93A4F942F90E9628540052090650525A0000066A00B",
INIT_16 => X"93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4",
INIT_17 => X"3A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E",
INIT_18 => X"09B56C74DAB15D1CF13501AA495000000000000000003A4E93A4E93A4E93A4E9",
INIT_19 => X"2082082082082082082082082082082082082082082084E41DC71C7155F3898E",
INIT_1A => X"3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F8208208208208",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE5294A5294A52800003E1F0F87C3E1F0F87C3E1F0F87C",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000030FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"A975EFFFAABDE00FFAEBDFFF5D2EAAAAAF7AEBDEBA0000000000000000000000",
INIT_22 => X"8000155087FC0155F7D168B55007BFDF45085168ABA002E82145085155545F7A",
INIT_23 => X"FFFD7545AA8028A00A2802AABAFF8028BEF5D7FFFE10005542145557FD5545FF",
INIT_24 => X"F7AEAAAAAA2FFFDF4500043FE105D2E954BAF7FFC0010080017555555568AAAF",
INIT_25 => X"A5D5168A00A2D142155005142010FFAE820AAFF842AABAA2AE95545FFD168ABA",
INIT_26 => X"FF5D2A821550000000BA007FD55FF5D7FC0145007FD7400550415410002E974B",
INIT_27 => X"F455D5142000082E82145FFD17DFEFFFD168BFFF780000BA007FE8AAAFF803FF",
INIT_28 => X"0000000000000000000000000000000000000000AAFBEAA00007BFDFFF082EBD",
INIT_29 => X"AABEA495FC716F002A975FFE3AA95E00EBAEBDFD75D2AA8A80EA8E2FE3F00000",
INIT_2A => X"56A16D557BC257D415E0216FA3F1E8FC0145B68B551475FAF6D1C556F0AA1C24",
INIT_2B => X"7FD24AFE3D02DAAAE12BD5545A2803AA0000542A0070071C50BAFEF1FAE0016D",
INIT_2C => X"A8B50F55A2F150005A3A438BD04AFAB8F550A8010E004924874825D7FEAA8548",
INIT_2D => X"A2A5504001C74BA42A1571E8028E3DB7816D0120155EA568E870BAEB8A05A2AE",
INIT_2E => X"2FFAFD2A82485FD2415A105C21451ED42A002545E055FFBE81D0BE8EA8A3AA05",
INIT_2F => X"100AA1D0F6F480B6A555A2A57A002A3D5FDB6A5C7E3DFFFE90B45B47ABA497A8",
INIT_30 => X"A0AFE80A8B0A000000000000000000000000000000000000000000000B55EAAA",
INIT_31 => X"ABEF5D557FEBA55022A3F70C6B405F4D2AE975EFAAAAB5E1AF3AABFF45592E88",
INIT_32 => X"411A8DED57CE1055555E5F58EFFC01FE2CACB65F520EBE9EF67D7BEA1FD5D556",
INIT_33 => X"A4AD0079C75D6070CC5CBB0280C029ABAA3EBC114728007521170821CE0FDE69",
INIT_34 => X"2A95E02A2AAB5EB0F280800EFAEE9F5D18F3142341D5DEEBEF55080034E0A592",
INIT_35 => X"B69C30E02116220415A9540AA854140A0A2047F353AAF6C77F7F20D968BF5781",
INIT_36 => X"ABEBE1B4D792A4AD1183454180DD3FDCAAAB7C91565455C141E41887D58AC448",
INIT_37 => X"F0000001FF01EABC4B8014174FF7DA80F52FEDE6BE93172D7D625B556EEAB157",
INIT_38 => X"FF0000001FF0000001FF0000001FF0000001FF0000001FF0000001FF0000001F",
INIT_39 => X"0000000000000000000000000001FF0000001FF0000001FF0000001FF0000001",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000100000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(0),        -- Port A data input
DOA(0)   => data_read_a_hi_256(0),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(0),        -- Port B data input
DOB(0)   => data_read_b_hi_256(0),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_1_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"212C001411984004084D000508C53810A03D1450E839B003342114428A000803",
INIT_01 => X"08000011400A100A81160000008C005400400002000000000000028001340000",
INIT_02 => X"C084484000002014400205851002007030450E0000A606C8C44CB4C6666C00E0",
INIT_03 => X"33DF380008164004000002000C80400002031943000101091608463061120118",
INIT_04 => X"4140008000000002000064000400004201000000000210458010070080100433",
INIT_05 => X"8500101040200000010009100000000508000100000000002010600100208D04",
INIT_06 => X"B5EDFDE24618AD433060C182BA860044204C000008A004100008000820280020",
INIT_07 => X"581E02100020000A81244890AA20263030517F122AA801F0983060AC564BF808",
INIT_08 => X"00820800C7A00045B103200000140A02234808000584000004808400020011A4",
INIT_09 => X"0000104000020082800808111008400000200204100000100820800144000414",
INIT_0A => X"12804062945211441E13C051156E800008402802060C94000040901102800000",
INIT_0B => X"24002006406401918C191AC191A4191A4191AC191AC191A4191A00C8560C8D29",
INIT_0C => X"0408010040050880383820080F105F05800302E0E08842422006000000041032",
INIT_0D => X"05000600000090C1841808172580000000008008020084082080204010200810",
INIT_0E => X"0500066210000178470184000000878402C000001E07800500062000001E0780",
INIT_0F => X"00003C404600000011A30E0700000009382000001E07800500062000001E0780",
INIT_10 => X"C0180000012010C20022100000F0C3C03000000055200340000000F88701C000",
INIT_11 => X"05800241186100004D100098190240001290002050068000001010486140F900",
INIT_12 => X"0000164A001303204800026880048230C2000094A0000F601F8000000001C908",
INIT_13 => X"12D051E01000000154200580003C030381840000004B08014401025480E07000",
INIT_14 => X"40082300218450C2800010094000482142E0601895001000000041C408014400",
INIT_15 => X"0802008020080200802008020080008208600500A82A15008000000000468000",
INIT_16 => X"8020080200802008020080200802008020080200802008020080200802008020",
INIT_17 => X"0200802008020080200802008020080200802008020080200802008020080200",
INIT_18 => X"BABEFC54A0810C7452B5420A1000000000000000000002008020080200802008",
INIT_19 => X"AAAAAAAAAAAAAAAAAAAAAAAAAAA28A28A28A28A2A8218D2C0C92492581328A46",
INIT_1A => X"2E974BA5D2E974BA5D2E974BA5D2E975BADD6EB75BADD6EB75BAAAAAAAAAAAAA",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFF6318C6318C63000002E974BA5D2E974BA5D2E974BA5D",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"00000000000000000000000C0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"002155557FFFFFF007FC21EFA2FFD74AAAAD5555550000000000000000000000",
INIT_22 => X"7FD75FFAAAA800AAF7AA974BAFFFBE8B45F7AEBDF455D2EAABEFF7FFE8BFF5D0",
INIT_23 => X"0557DF45AAD1400BAA2AE801550051555EFF7AA95400552AAAABAFFD1574105D",
INIT_24 => X"FFFBEAB55F780020AAAA80020AA082EAAB5500517DF555D2EAAA105500001550",
INIT_25 => X"AF7AE820AA0851574BAA2D1574AA5D7BFDEBAFFD540155557FD5400F78028BFF",
INIT_26 => X"FFFFD56AAAAFFFFD7555AAD168B45AAAEAAABAFF842ABEF5D517DF55552A974A",
INIT_27 => X"4BAF7AE80010082A97410557FEABFFAAFBE8BEFAAD1575EF557FFFE10557FFFF",
INIT_28 => X"00000000000000000000000000000000000000005D7FFDF4500043FE105D2E95",
INIT_29 => X"A8BC2EBDFEAF7F1F840017D4975D2FEF147FC51C7A2FBD5490BFD1C056A00000",
INIT_2A => X"AA8AAAE3D145410F7F1D55D71C002DABAEBAA974BAF7FFEFB45FFAABDF55492A",
INIT_2B => X"0E2AE85028B40155145F7AF6DBED5450AA1C2080BEF495FC71D54124924385FA",
INIT_2C => X"571D2E28E38E0216FA2D1E8E80140F45082B4002D082082AB8B6DBEDB7DF7F54",
INIT_2D => X"A97F7AF6D417E92482BF84020BA495557E3FF78E021FF1471FDEAAFFD56F16D5",
INIT_2E => X"7002FD74951D71EDFFABFD16FAAAE92BD5545A2DA3FB7DAAD4AAAAF487BC70BF",
INIT_2F => X"550A8010E00492487482FFFE82A85EBAE2FFC55554ADBD7A2FFC7BEFF6FFD7FC",
INIT_30 => X"400FBF9424F7000000000000000000000000000000000000000000000547AB8F",
INIT_31 => X"DF55F7AABFF55082CA8B4DF6C1E8F5E5400021EF005162BEF047FD5545AAFBF7",
INIT_32 => X"404547184164AA5D2EBEEB0A2D555410D3555714F8338AAAA1D0AE974AAF7FFF",
INIT_33 => X"AEABFFDF79DCBF755962010BDCBBC21455D7FEABEF75550ACBB7582225FF5843",
INIT_34 => X"D57D412F7D55F5E50C7F401BAAE8403CF5A3FFEAAEB083BC1000FF8409000512",
INIT_35 => X"2AA9FEAFDF7F431A9F7FFE81FF013A8001AFF801F8BA0C57740BDAA0688E5405",
INIT_36 => X"A2FBF7FED2C7F955445079E280A00C56145EF5D16BABAA3EBC3157ABD5FFE55F",
INIT_37 => X"0000000000596EBEF55080034E0A592A4AD00FB863550229BCABEB7DA403FFFD",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000100000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(1),        -- Port A data input
DOA(0)   => data_read_a_hi_256(1),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(1),        -- Port B data input
DOB(0)   => data_read_b_hi_256(1),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_2_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10E006600180111284380310006289800480032283E000A34301002001A0817",
INIT_01 => X"A14AC00A1079284D04A044A54E504368404000720885800802000006ECD10200",
INIT_02 => X"92250052A0348C310102048800A8507000040C8550200000480E0080001321E0",
INIT_03 => X"020204E4593C0824400C2220483042809292430400440180000890A4C9400242",
INIT_04 => X"486854B141002252142241502460480031B94420634850069A42241009610A04",
INIT_05 => X"800504244080892105AA6010A44882144840910A21220A8C820025E4A0000B00",
INIT_06 => X"A000442802280000340810209C444804206000AC800088096A0EA8C022208012",
INIT_07 => X"309820A848E0AA09826489A5CC49002001020112028201F8A20488260000108A",
INIT_08 => X"2400582881E0C1419D12041455509341A539C42A0D8208099002801700D10103",
INIT_09 => X"110D525861263100009200151409130A3C80C8C8096A06B8C12088400A9C2080",
INIT_0A => X"0451394CD0391A441583C04B580040089581001342801044877200D002A00DE0",
INIT_0B => X"144423040240450114901149013C9011C9013C9011C90134901144801A4808A5",
INIT_0C => X"D8A5345206D2C10082080A90C00000188150100C202A4640000E2B4081969420",
INIT_0D => X"050080400A0391A51240C480000AA902AA009028C83220008086952B4285A54A",
INIT_0E => X"05008021C00000000040000000020288000500000008000500802A0000000800",
INIT_0F => X"0002300000428000000040000000000D002A0000000800050080250000000800",
INIT_10 => X"0000000001204004000508000000100000000002054000130000000000800000",
INIT_11 => X"000C00000000000068144000000000001A000106200010021002000000000080",
INIT_12 => X"0002004A880000000000034098000000000000D024A000000000000001000900",
INIT_13 => X"00000000000000041400000A8000000000000000010A00000284000000000000",
INIT_14 => X"012100000002000280000000011080C000000000000000000000430000000260",
INIT_15 => X"A769DA769DA769DA368DA36CDA3A9A13A14801404134DA84A024024155000399",
INIT_16 => X"168DA769DA769DA769DA368DA368DA368DA769DA769DA769DA368DA368DA368D",
INIT_17 => X"68DA168DA169DA569DA569DA568DA168DA168DA169DA569DA569DA568DA168DA",
INIT_18 => X"138D70C030B51C50C7D000A2012F81F81F83F03F03F069DA569DA569DA568DA1",
INIT_19 => X"1041041041041041041041041041041041041041024860208165965975960040",
INIT_1A => X"25128944A25128944A25128944A25128944A25128944A2512894104104104104",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFF8421084210840703F25128944A25128944A25128944A",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"00000000000000000000000F0FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"415555087BFFF55A2AA800BAFFAE9540008002AA000000000000000000000000",
INIT_22 => X"7FE8B555551421455D0002145552EBFEBA007FC21EFA2FFD75EFAA8415410AA8",
INIT_23 => X"FFFE8B45552EBDF45FFAEAABFFF7FFE8B55F784155EFA2AEBDEAAA2FBEAABA5D",
INIT_24 => X"5D2AAAAAA5D2E820BAA2FBEAB5555557DF55A2AEBDF555D2E954BAA2AA974BAF",
INIT_25 => X"A5D04021EF557FC21FFAA8428BFFAAAA954AAAAAAAAAAAFFD1574105D7FFFF55",
INIT_26 => X"EFF7800215500557DF55AA80001FFAA80001550055575EFFF84021555D043DEA",
INIT_27 => X"B5500517DF555D042AA10A284154005D0015410085568A00FF80175FFA2D17DF",
INIT_28 => X"00000000000000000000000000000000000000005D00020AAAA80020AA082EAA",
INIT_29 => X"D55D2BE800042AFE8E1557D0075D2F45BEAA800AAFFAA9543A080038A2A00000",
INIT_2A => X"0BDEAAA2FBF8AAA557BE8B6D5D5FFABEF49040017D5D20B8EAA007FC51C7A2FB",
INIT_2B => X"0E174BFA02A974BAF7F5EFB455D2ABDF55492AA8BC7EBDFEAFEFFD00105FFBC2",
INIT_2C => X"3D155E105571D55D71C002DABA5524820BAB6FFEFB6D555578F7DB6A0BDF7D48",
INIT_2D => X"092A071555D5E3AE821D00001FF0871C016DBED1FDE90E3A497492B6AAADAAAE",
INIT_2E => X"0E3DA3DFD5E3DFFFBD5A38A021551C5F7AF6DBE8F401D7B6A0001470155C51D0",
INIT_2F => X"82B4002D082082AB8B6D1C5B7DF7FF78E075C5BE8555400550A38428007FED00",
INIT_30 => X"4AA00042AAA2000000000000000000000000000000000000000000000410F450",
INIT_31 => X"AAAA007FD5555AAFBD7545FBB8020A3F7AE975EF005560B55F7AA800AAF7AA95",
INIT_32 => X"E8F5EFF84165EFF7802BAB0A2FFEAABA557BEABEF057D68F5F5A00021EF55042",
INIT_33 => X"52ABFFFF841FFE75CA882108202E974AAF7D57DF55D7AABFF5428ACA8F45A6C1",
INIT_34 => X"84174A8FFAEBFEB0A2D55541051555694F002CA8AA80800020AAF7FBFFFEF045",
INIT_35 => X"7AAA155F595542455512A975455D3AA8A005500151FF0C57401E5F3D1E00A1A8",
INIT_36 => X"5D2A8A0B882FFFFE10AAAAAB755A66B6AF56A2AA801455D7FE8BFFF680800FFF",
INIT_37 => X"00000000000C3BC1000FF8409000512AEABFF5D79FCAF774AE005BE789555400",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000200000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(2),        -- Port A data input
DOA(0)   => data_read_a_hi_256(2),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(2),        -- Port B data input
DOB(0)   => data_read_b_hi_256(2),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_3_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"210C44A20020248B08431120001604B8156023104C4077133420400A02380202",
INIT_01 => X"015A2A424080216D3C2462C99E104B49404040028804A0080A000C16A0D90A0C",
INIT_02 => X"C0A4065000F0A95011000D1501005270B4045AB330860281CC08008222170060",
INIT_03 => X"AD22014098340394A4021320080841C40B411B4298042180002846B06900811A",
INIT_04 => X"244B32A86D20014A0D20403194904900071A24110F0BF400F85F92420E0C946E",
INIT_05 => X"80331030442898B4812840D0500008C528280B063006A64CA30004E5A4E40304",
INIT_06 => X"90016CA00E380042302040A0BC47160424428198C0038C89904E640023600816",
INIT_07 => X"1288020843A66620816049908AA0061011CA0142000009F0A810292E7402F088",
INIT_08 => X"20003C9984A0AC411102014D34EC2200214D5099048823019603A01A49410103",
INIT_09 => X"001CD74C4826220010A8891451284B661CA24A4C899046740121824004100080",
INIT_0A => X"44C9516DC0135C45159BE45F112B48804DC10203021290400772C0F402820D4C",
INIT_0B => X"B400624402404501A49018490184901A4901A4901849018C901A648056480C2D",
INIT_0C => X"D7A9B54000D7C10820680D08C420180381211081A022160000266723E1909021",
INIT_0D => X"400080200E199A4A2CA2994C0399981666409800CA52E4890806BD6B56BDAB52",
INIT_0E => X"40008008E00000000000000000024008000C8000000000400080028000000000",
INIT_0F => X"000A000000588000000000000000200400088000000000400080078000000000",
INIT_10 => X"0000001000004004000D800000000000000000022040000B4000000000000000",
INIT_11 => X"001A0000000000082006C000000000020804087220000122000A000000000000",
INIT_12 => X"00020800B8000000000041002E00000000001040466000000000000001020080",
INIT_13 => X"00000000000000048200004A600000000000000003008000320C000000000000",
INIT_14 => X"432900000222200871028000210400C4000000000000000000080200800030E0",
INIT_15 => X"AF6A5AF6A5AF6A5AF6A5AF6E5AFADA91AB68000101B4D20C08EC461733804A19",
INIT_16 => X"B6B5AF6A5AF6A5AF6A5AF6A5AF6A5AF6A5AB6B5AB6B5AB6B5AB6B5AB6B5AB6B5",
INIT_17 => X"6BDAB6B5A96ADAF6A5AD6ADAF6A5AD6ADAF6A5AD6BDAB6B5A96BDAB6B5A96BDA",
INIT_18 => X"C78C706428A14C586290008A044D54AAB556AA9556AAEBDAB6B5A96BDAB6B5A9",
INIT_19 => X"92492492492492492492492492410410410410412821600001249249015303C0",
INIT_1A => X"351A8D46A351A8D46A351A8D46A351A9D4EA753A9D4EA753A9D4924924924924",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000001543B351A8D46A351A8D46A351A8D46A",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"43DF55FFAA955EFA2D168B55557BEAA000055420000000000000000000000000",
INIT_22 => X"7BE8BFFA2D155410AA8415555087BFFF55A2AA800BAFFAE9554508002AA00AA8",
INIT_23 => X"52ABFEBA007FC21EF007FD75FFAA841541008002AB55AAAA955EF005568A0008",
INIT_24 => X"005168B455D042AB45F7FFD741000042AA10AAAABFF5508003FF555D00021455",
INIT_25 => X"0A2D1575FFF7AA975555D2E80145F78415545082EBDEAAA2FBEAABA5D7FC0155",
INIT_26 => X"55552A954BAFFFFE8B55552EBDE00F7AEAABFFF7FBEAB55F7AABDEBA5D7FC201",
INIT_27 => X"F55A2AEBDF555D2E954BA002EAAABA002A821EF5555554AA087BC01FFFFAAAAB",
INIT_28 => X"0000000000000000000000000000000000000000082E820BAA2FBEAB5555557D",
INIT_29 => X"95578080038A2AA28E3AF55E3A0BA5D7AADB6FB7D5D7FEAA3808554203A00000",
INIT_2A => X"0925D7085F6AA10087FEABD7AAD57AEBAB68E1557D1475FAF45BEAA800AAFFAA",
INIT_2B => X"04AAFFA41040017D5D20B8EAA007FC51C7A2FBD55D7BE80004AA1E8E2AB55B6A",
INIT_2C => X"2FBE80AA557BE8B6D5D5FFABEF49002FB55FFF5D0438140E2FA38B6AEBFF6D1D",
INIT_2D => X"AB8ABAE925D21C7010EADB525D7FFAE975C75D0A901FFFF801557D1C20B8EAAA",
INIT_2E => X"20875C21D5EB8AA8FFF012A954BAFFF5EFB455D20BDE00EBAAA8BC7EBDFEAFEF",
INIT_2F => X"BAB6FFEFB6D555578F7DB6A0BDF7DEB8E125FF002EADA921420871D74971D248",
INIT_30 => X"ABA0051400A20000000000000000000000000000000000000000000001C24820",
INIT_31 => X"8B55F7AA800BAF7AA955EF00042AAA2A2AEAAB55A28408145AAFFFFFFF5D7FEA",
INIT_32 => X"020A35D2ABEF55F7800015F087FEAA00007FEAB55FAD568AA2AFAE975EF55516",
INIT_33 => X"ABFEAAF7AE9DFF759A82AEF70800021EF55042AAAA007FD55558A7BD7145FBB8",
INIT_34 => X"84175EF55002AAB0A2FFEAABA557BEA3EF057968F575D003FF55F7D5420BA5D2",
INIT_35 => X"A8429F45A7D5EAF5FFBAEAAA10554155400AAFFD5145FBAC9755F05040255FFD",
INIT_36 => X"550415557085540000005156155FE90A8F5C082E974AAF7D57DF45552A3FF10A",
INIT_37 => X"00000000005500020AAF7FBFFFEF04552ABFFFF843FFE77C80825BC052ABFE10",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000100000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(3),        -- Port A data input
DOA(0)   => data_read_a_hi_256(3),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(3),        -- Port B data input
DOB(0)   => data_read_b_hi_256(3),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_4_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"A108400020612C80284210081034849800A000303100048B3432C82904204002",
INIT_01 => X"21066802000820491C00650E1E004360403008418984014902030906A8D10200",
INIT_02 => X"120404E00E4C0600000206100008402005040C00F104008040080080001310E0",
INIT_03 => X"DCA201514D1C0D706C5CF010083A0708BA0841945004010000080084C1000002",
INIT_04 => X"5C4CF21C48B133483C80417570D000083A62488074C1350EA60D785C0A6B0619",
INIT_05 => X"000F0400028083B381A60001E5546EB5C0E2B81E4166DE000139200004E50940",
INIT_06 => X"80004408020800023000102098000204A040038600018019004B800123208806",
INIT_07 => X"120C20204665E1008024188488800000001A01520000A1F08044892400001088",
INIT_08 => X"0801007AC0A1EB413102063CF3E0B3028D29F407059B0B000205A801C2200102",
INIT_09 => X"106052400922D00406BE1002C6150F41200280001900439001FD8A0004142000",
INIT_0A => X"047F2201D899BA503583504B58AB80804540001202805544314041B48A888EC5",
INIT_0B => X"1441E3443043410C5010C3010C1010C3010C1010C1010C3010C14086980861A5",
INIT_0C => X"020000A02600000805400502C0A0004A00625015000A12000026E1E180011220",
INIT_0D => X"400000000E43930C20C20188120782861E4004A800600401A030001008080400",
INIT_0E => X"40000021A8800000000000000000400800170024000000400000310024000000",
INIT_0F => X"0008000000AA80200800000000002000003400240000004000003B0024000000",
INIT_10 => X"00000010000000040004A080000000000000000020400006C008020000000000",
INIT_11 => X"002C008200000008001B4020200000020000090760000200110A040010000000",
INIT_12 => X"00000803E004040000004000E801040000001000086000000000000000020040",
INIT_13 => X"0000000000000000810000164001008000000000020040002240008020000000",
INIT_14 => X"04001040026026004000000002940040000410000000000000080000400000B8",
INIT_15 => X"040080201004008060000001806AC000004890015124D880100886D8F0014420",
INIT_16 => X"4010000180600000018020100400802010000080601000008020000401802000",
INIT_17 => X"0100000004008020180600000000000180600802010000000401802018020000",
INIT_18 => X"3807E05000140634504048820064B261934D964C326980004010000080600806",
INIT_19 => X"AAAAAAAAAAAAAAAAAAAAAAAAAAA28A28A28A28A2934C8D0CCD145144C0A28A06",
INIT_1A => X"068341A0D068341A0D068341A0D068351A8D46A351A8D46A351AAAAAAAAAAAAA",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000000173F068341A0D068341A0D068341A0D",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"57FE10FFFBEAA10007FD7410FFAA97555082A800AA0000000000000000000000",
INIT_22 => X"7FEAA00007BE8AAAAA843DF55FFAA955EFA2D168B55557BEAB45005542000005",
INIT_23 => X"87BFFF55A2AA800BAFFAE9555508002AA000055574105D2A800AA00043FEBA5D",
INIT_24 => X"A2D17DE1000517FE10AAAAA8AAA002E97545557BC00AAA2FFEAAAAAA84155550",
INIT_25 => X"0A2D157400AAAE974AAAAAA974BA08002AB55A2AA955EF005568A00087BE8BFF",
INIT_26 => X"BA080002145552ABFEAA007FC21EF007FD75FFAA8417410A2D140000F7FBC201",
INIT_27 => X"A10AAAABFF5508003FF55F7D568A00552EA8BEFA2AABDEAA087BEAAAAA2FBD54",
INIT_28 => X"000000000000000000000000000000000000000055042AB45F7FFD741000042A",
INIT_29 => X"EAB7808554203A145178E00FFFBE8A101475D5400F7A49057D0824850B800000",
INIT_2A => X"E8008200043FE925571EFA380871C7028A28E3AF55F7A0925D7AADB6FB7D5D7F",
INIT_2B => X"F5FDA38BE8E1557D1475FAF45BEAA800AAFFAA9557D080038AAA145157428492",
INIT_2C => X"85F6AA10087FEABD7AAD57AEBA08517DE00AAAEA8A9200249056D4175C5092AA",
INIT_2D => X"FEDB42028EBFBC2028BED152438AAA092492AAA4954281C0E2FB55B6A0925D70",
INIT_2E => X"A0875EDA80BEF1C743840040017D5520B8EAA007FC51C7007BD55D7BE80004AA",
INIT_2F => X"55FFF5D0438140E2FA38B6AEBFF6DBE84AAEBAF7DF6AA00412EAABFFAA803DEB",
INIT_30 => X"1EF0800154B200000000000000000000000000000000000000000000041002FB",
INIT_31 => X"0145AAFFFFFEF5D7FEABFF0051400A25D5568A00FFFFEAA105D5155410FF8402",
INIT_32 => X"2AAA25555410BA082E8201000043FE005D517DEBA0851574B2AAAEAAB55F7840",
INIT_33 => X"4001FF005575408AA557FEB2FFAE975EF555168B55F7AA800BAF7AA955EF0004",
INIT_34 => X"2ABFF55F7800015F087FEAA00007FEAB55FAD568AA200557DE00AAAAAAA00080",
INIT_35 => X"87BD6145FAAC000A2A6FBC00BAAAFBC00BAF7D1550AAAA8002010F2AC154B25F",
INIT_36 => X"082EA8BFFAA843FEBA08517DE00F3F9574B30800021EF55042AAAA007FD55550",
INIT_37 => X"000000000008003FF55F7D5420BA5D2ABFEAAF7AEBDFF779A82AA43F7FBE8A00",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000200000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(4),        -- Port A data input
DOA(0)   => data_read_a_hi_256(4),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(4),        -- Port B data input
DOB(0)   => data_read_b_hi_256(4),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_5_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50DF4A0791B3FCB694379283C81FD996A091832102004A337A20E07C0C1E006",
INIT_01 => X"294014468000A04D5C6A60000C34C24841280A00084000C8C212892EEAD53235",
INIT_02 => X"50AE41540CA1D9100002171C1F0A5171134E2A200D8633F8CD09DBFBBB970E7C",
INIT_03 => X"214E3C521D16021B64430CC51C45B8154689094241898749920842946B90010A",
INIT_04 => X"A2F20F7D7A314CB5C208E28A1BF0224A448920028A185340D0C20B2690000C22",
INIT_05 => X"7520B430B20B984809A8886E230C6106371146E1829941C58310402C600381CF",
INIT_06 => X"9CC96CD7C63A7495B9A356ACBC4601C57FD44F8549A46490261C4B39203F7080",
INIT_07 => X"12A88800B029E0C0A12C4B92AA36A2111167357C220095F3C8952A2E5D26F078",
INIT_08 => X"F3F00503B4AE105B534711820C0C0A1043080300F7E0E728B1829C2FEA0A95A1",
INIT_09 => X"C5184F084136848C9298A8560688F480C58858449026145B3830F40944906234",
INIT_0A => X"50EB4124D2B3902BF5C9700C1199DCA84DF46A974F92C7E28F1630D38088A438",
INIT_0B => X"B3144E5636E3178C86B8CC6B8CA6B8CE6B8C86B8CE6B8CA6B8CC15C6435C670C",
INIT_0C => X"79E51E70E070AA8132252008360A7E91504104C8948047D6B0AE1FE440B28A71",
INIT_0D => X"05F0FE40014090400400080329FF8089FF49611F589765923E139F09C78CE7C6",
INIT_0E => X"05F0FE64037FFD7857418407157797878F005F0DFF0F8005F0FE205F0DFF0F80",
INIT_0F => X"8F87FCB1F8053FDEB9B34E0700461E5FF8205F29FF0F8005F0FE205F29FF0F80",
INIT_10 => X"C0184D07C1FF55C3E3E0037FFCF8D3C03009C3CFD53C7E001FF2FAF89781C011",
INIT_11 => X"4E0CDF47186104C6FF177BD939024189BF900401165D645CEEF5BBCDF148F980",
INIT_12 => X"6397F64AEF7F2320483137F8A9BF8A30C2098DFCA06FFFE01F80001F81FDC94F",
INIT_13 => X"FFD051E01015C3BF553D3E0E5FFE838381840714F9DB4F4FA213F774A0E07002",
INIT_14 => X"8B652E2B3120C81284641D3E8DBF7D636FE070189500125C1F83FBCC4F4F80EF",
INIT_15 => X"E7394E339CE138CE5394E33D4E1E0E30E1208C251134921C12A44103F064014B",
INIT_16 => X"7384E3394E338CE538CE1394E3384E738CE139CE1394E7384E339CE139CE5384",
INIT_17 => X"38CE139CE1384E7384E7394E3384E738CE539CE139CE538CE5384E3394E7384E",
INIT_18 => X"7F7B9DB7FF3A1B6DB7ED438A9C3124B2DA6924965B4D384E7384E339CE138CE5",
INIT_19 => X"FBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEF9F7CFDFDDCF3CF3DF5E5BB4E",
INIT_1A => X"7BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEFBEFBEFBEFBE",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE000000000000118D27BBDDEEF77BBDDEEF77BBDDEEF7",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"E955450055421FFFFFBC0010AAD5574BA557FFDFFF0000000000000000000000",
INIT_22 => X"D5575EF55517FF5500557FE10FFFBEAA10007FD7410FFAA97410082A800AAAAA",
INIT_23 => X"FAA955EFA2D168B55557BEAB55005542000007FD74000055574BA5D7FD7555A2",
INIT_24 => X"007BC00AAAAAEBDF45A28428B45FFD168BFF00002AABA5D2ABFFFFAA843DF55F",
INIT_25 => X"AFF80174BAAAD1555EF5555555550055574105D2A800AA00043FEBA5D7FEAA00",
INIT_26 => X"FFAA8415555087BFFF55A2AA800BAFFAE95555080028A00A2FFFDE00F7D57FEB",
INIT_27 => X"545557BC00AAA2FFEAAAA082A97545F7D5420BA5D2E821FFA2D5554BA557BD75",
INIT_28 => X"000000000000000000000000000000000000000000517FE10AAAAA8AAA002E97",
INIT_29 => X"9043D0824850B8A2AE9756D145B401FFFFFFC7010BEDF524AA5571FDFEF00000",
INIT_2A => X"1524BA5571D757DB6D5525EF555178F6D145178E00EBFBE8A101475D5400F7A4",
INIT_2B => X"24BFFFFA28E3AF55F7A0925D7AADB6FB7D5D7FEAB7D0855420BA1471D7438085",
INIT_2C => X"0043FE925571EFA380871C7028B6AEBDF45B68A28B6DEBDF6DBEF1C0A28AAA55",
INIT_2D => X"A2FBF8E10EBD578EAAFF8415482BED1555EF55555057D145152428492E800820",
INIT_2E => X"FB6DF574A85575C55EFBE8E1557D1475FAF45BEAA800AAFFAA9557D080038AAA",
INIT_2F => X"00AAAEA8A9200249056D4175C50920875FDA381C209256DFFDF420BA552A821F",
INIT_30 => X"0BA55557DFF700000000000000000000000000000000000000000000008517DE",
INIT_31 => X"AA105D5155410FF84020AA0800154B2AAAA975FF5D7BC21EFF7FBD7400F7FBC0",
INIT_32 => X"400A25551554BA0051400BA5551575EFF7D1401FF5D5568BE7555568A00AAFFE",
INIT_33 => X"FFDFFF552EA8AAA55043DFF7AAAEAAB55F78400145AAFFFFFEF5D7FEABFF0051",
INIT_34 => X"55400BA082E8201000043FE005D517DEBA0851574B2FFAABFF45FFAAAABFFAAF",
INIT_35 => X"7AA955EF00002AAA2A2FBE8A00A2D16AAAAFF8002410FFD5575EF5555421E755",
INIT_36 => X"FFFFC00BA552A821EFFFFFD74BA5D51575F7FFAE975EF555168B55F7AA800BAF",
INIT_37 => X"000000000000557DE00AAAAAAA000804001FF0055554088A557FEB25D00021FF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000C00000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(5),        -- Port A data input
DOA(0)   => data_read_a_hi_256(5),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(5),        -- Port B data input
DOB(0)   => data_read_b_hi_256(5),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_6_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10800B0061A01002840002C03002818000402322520070B313301C4389B2082",
INIT_01 => X"274008482009404C18A160000C52424841000000090800090210000008510200",
INIT_02 => X"102430600C800110000006100009D070012408000000000648080000001210E0",
INIT_03 => X"000200501D1D02140C420200480140040608010040400104681A0084490C4802",
INIT_04 => X"404402820021000A00824002141000980500000808001114C000080624600600",
INIT_05 => X"120024204209981001A806500304610528000500000080000000300000012940",
INIT_06 => X"2000440832280002300010209C4400142061207A024008900008000220600220",
INIT_07 => X"130C8A220FF41F00902008808800182001020150000001F0800408264000100A",
INIT_08 => X"001BF002C4A01041B1120101000010128568837F04842B080020890008080342",
INIT_09 => X"011847140126805432A62A1596C8B5DF10000008900000100220C00084000008",
INIT_0A => X"44EB4104D09392053589F11C59898888454010830212C54081000410A0088C00",
INIT_0B => X"B0044245B25B456C0096C0096C4096C4096C2096C2096C6096C444B6004B600C",
INIT_0C => X"09040020280010000B3002820110101D0012402CC00802410C26800860070621",
INIT_0D => X"0500819D0000900208201040C4007920004884080000448C281018100C000200",
INIT_0E => X"05008182100000000000000000022AE800C00004000000050081A00004000000",
INIT_0F => X"0002330006000000080000000000000D07A00020000000050081A00020000000",
INIT_10 => X"0000000001204A340002100000000000000000020F4001400000020000000000",
INIT_11 => X"019300020000000068D08000200000001A692121000280000000000010000000",
INIT_12 => X"000201FA100400000000034696010000000000D3478000000000000001003F00",
INIT_13 => X"00000000000000043C0001C0A000008000000000012E000054AC000020000000",
INIT_14 => X"0200000040A410C2810800016000809400001000000000000000433300007600",
INIT_15 => X"060180400000008060180404002AC0200208940041309210B28048180F028000",
INIT_16 => X"2008000100601802000000100601800000000180600800000020180600000000",
INIT_17 => X"0180600000008040100200800000060100000802010040180200002018040100",
INIT_18 => X"7F8FF0F4FA955F7CF7F40A80907638C31C71C718638E00006018040080200004",
INIT_19 => X"38E38E38E38E38E38E38E38E38E38E38E38E38E39B6CEDECDDF7DF7DF5F78BCE",
INIT_1A => X"3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE38E38E38E38E",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFF000000000000196A03F9FCFE7F3F9FCFE7F3F9FCFE7F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"00000000000000000000000C0FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"BFDF45F7AA974AAAAAA97555F784174BAF7D5555FF0000000000000000000000",
INIT_22 => X"FBD7410AA8428AAAAAAE955450055421FFFFFBC0010AAD5574BA557FFDFFF087",
INIT_23 => X"FFBEAA10007FD7410FFAA97400082A800AA08515555508043FE00F7AA97555A2",
INIT_24 => X"55517FF55A2AA97400552AAAB45082E80155F7D1575EFFFAA9555500557FE10F",
INIT_25 => X"FF7AAA8A10082EAAB45A2FFC2000007FD74000055574BA5D7FD7555A2D5575EF",
INIT_26 => X"FFAA843DF55FFAA955EFA2D168B55557BEAB5500554200000003DE10FFD5401F",
INIT_27 => X"BFF00002AABA5D2ABFFFF087BD5545007BFDE10AA803FE105D516AABAFF843FF",
INIT_28 => X"0000000000000000000000000000000000000000AAAEBDF45A28428B45FFD168",
INIT_29 => X"524AA5571FDFEF1C7BFFF55FFA095482B6A49256DEB84104BAFFD1525FF00000",
INIT_2A => X"03DE28F7A49057DAAF5D2428A2842AAAAA2AE9756D145B401FFFFFFC7010BEDF",
INIT_2B => X"A49756D145178E00EBFBE8A101475D5400F7A4904380824850381C5B5057D1C0",
INIT_2C => X"571D757DB6D5525EF555178F6DAAA495428412AAFB451C2A8017DE3DF525FFFF",
INIT_2D => X"1C0E3FE00E3DB471EFE3AAAAA00082EA8B6DA2F1C50381471D74380851524BA5",
INIT_2E => X"049516AAB8FF8428FEFA28E3AF55F7A0925D7AADB6FB7D5D7FEAB7D0855420BA",
INIT_2F => X"45B68A28B6DEBDF6DBEF1C0A28AAA5524BFFFF1C7BD057D1C71FFE10A28038E1",
INIT_30 => X"0AAFFD1401E7000000000000000000000000000000000000000000000B6AEBDF",
INIT_31 => X"21EFF7FBD7400F7FBC00BA55557DFF7557BFDF55F78017400F780001FFAA8400",
INIT_32 => X"154B2557FC01EF55043FEAAFF80021EFA2D1420BAAA8428AA2AAAA975FF5D7BC",
INIT_33 => X"A821EFAAFBC01FFF780155F7555568A00AAFFEAA105D5155410FF84020AA0800",
INIT_34 => X"51554BA0051400BA5551575EFF7D1401FF5D5568BE7AA80174AA082ABDF555D2",
INIT_35 => X"D7FEABFF0051400A25D2EBFE10AAFFD55EFA2AEA8A10082EA8BEFAAD5554B255",
INIT_36 => X"55557DE00AA842AA0000516AABAFF8428BE7AAAEAAB55F78400145AAFFFFFEF5",
INIT_37 => X"0000000000FFAABFF45FFAAAABFFAAFFFDFFF552EA8AAA55043DFF7557BC01EF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000900000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(6),        -- Port A data input
DOA(0)   => data_read_a_hi_256(6),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(6),        -- Port B data input
DOB(0)   => data_read_b_hi_256(6),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_7_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10844B00482258A2842112C02450418800002300500030B313300C418992002",
INIT_01 => X"234008422008604D1C20E0000E11426840000000080000080200090000110204",
INIT_02 => X"1025207000B08910000206101188D03080144880010400044808000000122160",
INIT_03 => X"000200401914821004420000CA01000C0600010000605114291A008449484802",
INIT_04 => X"40440200002100080006500210101019040000000B085024D842080244000000",
INIT_05 => X"1A8024200009981001A8224001040104200204000000800CC2092CE4A0004900",
INIT_06 => X"A000440822280002340010209C040014A061200052500810000C490323208E28",
INIT_07 => X"128802020028000890240980A809102001020140000009F0800408264000100A",
INIT_08 => X"001A0602C4A01051B13281010408881203480200448423199046821008082351",
INIT_09 => X"336784144126811054809C1040140A001C8648481000045903318B80A400310A",
INIT_0A => X"000800009010100014114110312388984502148282A08415B032095048008100",
INIT_0B => X"20CDC1C483484D201192011920119201192051920519205192074C9018C90188",
INIT_0C => X"D8A5B44001D2C12901228F82F005310D293054048A2212004466000DA1908528",
INIT_0D => X"800F8108A0D09802082010408580008000000008C85264010816851B428DA146",
INIT_0E => X"800F81321000020000261900E28A204040E000A0000007800F814000A0000007",
INIT_0F => X"7072024807000020400000581C01C1A406400084000007800F81400084000007",
INIT_10 => X"060180E83800E820101210000200000CC3003C32080201C0000C000000160700",
INIT_11 => X"81DD00804086423120B74020023090644840A34000828800000004000420020B",
INIT_12 => X"1C6A0186E8000446120C8905BA0004810C84624237E00010001878007F0030C0",
INIT_13 => X"00080208E4083C44230201AEE0010040261900E30520C0806EAC0082000984C0",
INIT_14 => X"0121011088A600C032128201519480D40005802448160403E0700622C0806EE8",
INIT_15 => X"A1685A1685A168DA368DA36CDA30DA13A108810111349A943AA4401000928A19",
INIT_16 => X"368DA768DA1685A1685A5685A368DA368DA7685A1685A1685A768DA368DA368D",
INIT_17 => X"685A1685A169DA368DA1685A1695A368DA3685A1685A168DA368DA1685A1685A",
INIT_18 => X"00000000000000000000400A8448410400020820800069DA1685A168DA369DA3",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000003667B000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"0155EFAAAEA8ABAAAFBFDE0055556AA005D04155550000000000000000000000",
INIT_22 => X"556AA00FFAE95555087BFDF45F7AA974AAAAAA97555F784174BAF7D5555FFF78",
INIT_23 => X"055421FFFFFBC0010AAD5574BA557FFDFFF5555555EFAAFFFDFEFAAAAAAB455D",
INIT_24 => X"AA8428AAA557BFDFFF55003DFFFF7FBEAA00002EAAAAA082EA8A00AAAE955450",
INIT_25 => X"0552EBDE00007BEAAAAA2D14000008515555508043FE00F7AA97555A2FBD7410",
INIT_26 => X"FF00557FE10FFFBEAA10007FD7410FFAA97400082A800AAF7AE975FFA2800001",
INIT_27 => X"155F7D1575EFFFAA955555D51574AAAAFFD5545087FEAB455D516AB55557BD55",
INIT_28 => X"0000000000000000000000000000000000000000A2AA97400552AAAB45082E80",
INIT_29 => X"104BAFFD1525FFFF8E175C7A2AAAAA82A2F1FAE105D556AA10410E1755500000",
INIT_2A => X"1FFFD7AAAAAFB7D495F6AA10E3AE905551C7BFFF55FFA095482B6A49256DEB84",
INIT_2B => X"2EAAA00A2AE9756D145B401FFFFFFC7010BEDF524AA5571FDFEF415B575D7AAF",
INIT_2C => X"7A49057DAAF5D2428A2842AAAA497BFAFFF49003AFEFEBFBEAA001C2EA8A821C",
INIT_2D => X"F7A4905C7A28A070384120BDE100075EAA82BEDB470101C5B5057D1C003DE28F",
INIT_2E => X"D555F6AB57417BC05D7145178E00EBFBE8A101475D5400F7A490438082485038",
INIT_2F => X"28412AAFB451C2A8017DE3DF525FFFFA49756D495150492BEF1D2555087BE8B7",
INIT_30 => X"A10002E9754D000000000000000000000000000000000000000000000AAA4954",
INIT_31 => X"7400F780001FFAA84000AAFFD1401E7FFAA97555A2AEA8A10AAD568A00555168",
INIT_32 => X"7DFF7007BD5555AAD57DF55AAAEBDFEF007BE8A10AAAE8215D557BFDF55F7801",
INIT_33 => X"FEAA105D2EAAA005D2AAAA18AAAA975FF5D7BC21EFF7FBD7400F7FBC00BA5555",
INIT_34 => X"7FC01EF55043FEAAFF80021EFA2D1420BAAA8428AA2007FE8BFF080028BFFAAF",
INIT_35 => X"F84020AA0800154B2FF8402145A2AA954AA00043DE0000516AA10F7FBD740855",
INIT_36 => X"FFD140145007FE8BEF557BEAB55087FC215D555568A00AAFFEAA105D5155410F",
INIT_37 => X"0000000000AA80174AA082ABDF555D2A821EFAAFBC01FFF780155F7005140000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000000FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(7),        -- Port A data input
DOA(0)   => data_read_a_hi_256(7),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(7),        -- Port B data input
DOB(0)   => data_read_b_hi_256(7),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_8_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00000648E2840112C00000418000002700500030B3132000400812086",
INIT_01 => X"214009C21838284D042100000212026840000000180800080200080040510204",
INIT_02 => X"1021004000900110000006100088503000240800014400004808000000122160",
INIT_03 => X"0002004019110214044A82000121400C86000000000000860188008448400002",
INIT_04 => X"000402800031200A0000090214100889A5000000490090104800000224000400",
INIT_05 => X"10C025204289981000A820500344010428008500010080080909304040202004",
INIT_06 => X"8000440003280000340010208C04003420600000C6180810000C490703200010",
INIT_07 => X"130002000028000890240980A809012001020050000009F08004082640000082",
INIT_08 => X"20100402C4201041310041010008801201480200051023090024811008090A1A",
INIT_09 => X"0100001001248100308214528148A48008000008100004590711C04034000083",
INIT_0A => X"10804000801210140001C0103001088845010482004000008420041020008900",
INIT_0B => X"0004404002004400448000480004800048000480004800048000440022400200",
INIT_0C => X"880420000880204909004502D100A10C04205424010216010C26800805000004",
INIT_0D => X"8000801100509802082010400400018000488428800004082014000200010000",
INIT_0E => X"8000800A00000207A8BE7B00000200082040808000F07F80008000808000F07F",
INIT_0F => X"0002000402100000404CB1F8FC0000040000808000F07F80008000808000F07F",
INIT_10 => X"3E07800000004004080A000002072C3FCF0000020040804800040007687E3F00",
INIT_11 => X"10800018639EC00020100002C2F9B0000801016001008100000040120CB3067F",
INIT_12 => X"000200020000585EB6000100800030C73D8000402000001FC07FF80001000080",
INIT_13 => X"002EAE1FEC0000040200408000003C547E7B00000100801004000803551F8FC0",
INIT_14 => X"00000000440610C8000A808040000208901B86E568FE0C000000020080100400",
INIT_15 => X"0040100401004090240902449028D0230249850101349A98BAC0481000888810",
INIT_16 => X"0401004010040100401004010240902409024090240902409004010040100401",
INIT_17 => X"4010040100409024090240902409004010040100401004090240902409024090",
INIT_18 => X"543EBC57A10A1E75D6440A889050000000000000000040902409024010040100",
INIT_19 => X"79E79E79E79E79E79E79E79E79E79E79E79E79E7BF3CCD8DF5B2DB2CA4028A0A",
INIT_1A => X"4F87D3E1F4F87D3E1F4F87D3E1F4F87C3E1F0F87C3E1F0F87C3E79E79E79E79E",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000000D3E94F87D3E1F4F87D3E1F4F87D3E1F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"000000087BEAA10F7803DE00FFAEBFFFF0800155FF0000000000000000000000",
INIT_22 => X"7FC2145005155555F780155EFAAAEA8ABAAAFBFDE0055556AA005D0415555080",
INIT_23 => X"7AA974AAAAAA97555F784174BAF7D5555FF552AA8AAA557FC0010F780154105D",
INIT_24 => X"FFAE95555AAFFE8A00552EBFE00F7D17FF45F7FFFFF55AA80155FF087BFDF45F",
INIT_25 => X"5F7D140010552E821EFAAAABDF555555555EFAAFFFDFEFAAAAAAB455D556AA00",
INIT_26 => X"00AAAE955450055421FFFFFBC0010AAD5574BA557FFDFFF5504000AAAAAAA8B5",
INIT_27 => X"A00002EAAAAA082EA8A00002AA8A10F78402155AA8028A00A2D57FF45557BE8A",
INIT_28 => X"0000000000000000000000000000000000000000557BFDFFF55003DFFFF7FBEA",
INIT_29 => X"6AA10410E17555080E000280071E8A00EB8E3FE10F7AEBAFFF080A175D700000",
INIT_2A => X"1C2000FF8A17400557FC015514555757DFF8E175C7A2AAAAA82A2F1FAE105D55",
INIT_2B => X"8A105D71C7BFFF55FFA095482B6A49256DEB84104BAFFD1525FF492EA8AAA557",
INIT_2C => X"AAAAFB7D495F6AA10E3AE90555A2FBE8A38492ABDE10EBDF7AF6DE3FFF8F7DB6",
INIT_2D => X"550E00082B6A0AFB55F7D1420104124821D7AAA0BDF6D415B575D7AAF1FFFD7A",
INIT_2E => X"0B6D578F6D557FFDA00A2AE9756D145B401FFFFFFC7010BEDF524AA5571FDFEF",
INIT_2F => X"FF49003AFEFEBFBEAA001C2EA8A821C2EAAA001C2EA8A00F7800017DA2842FA0",
INIT_30 => X"BEF082E95545000000000000000000000000000000000000000000000497BFAF",
INIT_31 => X"8A10AAD568A00555168A10002E9754D082E820BA08556AA00AAAABFE00F7AEAA",
INIT_32 => X"401E7082EAAABA5D5140010F7AE974105D7BC21555D51575EFFFAA97555A2AEA",
INIT_33 => X"BEABFFAAFBEABFFF7AA80145557BFDF55F78017400F780001FFAA84000AAFFD1",
INIT_34 => X"7BD5555AAD57DF55AAAEBDFEF007BE8A10AAAE8215DA2FFE8ABA082ABFE00AAF",
INIT_35 => X"7FBC00BA55557DFF75D2E82010F7843DF45FFD540000000402145AA843FFFF00",
INIT_36 => X"F780021FFA2803DE10FFD16ABFF5D7BFDE10AAAA975FF5D7BC21EFF7FBD7400F",
INIT_37 => X"0000000000007FE8BFF080028BFFAAFFEAA105D2EAAA005D2AAAA185D2AAAA10",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000400000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(8),        -- Port A data input
DOA(0)   => data_read_a_hi_256(8),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(8),        -- Port B data input
DOB(0)   => data_read_b_hi_256(8),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_9_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000B0001800002840002C0000281800000030000000033022000000000002",
INIT_01 => X"8000098218302849180060000C004240413C0A61590001D90213C90008510200",
INIT_02 => X"000008700CB089100002061031200074810448800104008048080080001210E2",
INIT_03 => X"000200140C1822000A028010408100000628000140402080041A100040024840",
INIT_04 => X"41040000000400080002040200080800040000000B08D1055842080604600700",
INIT_05 => X"10002024000020102400010000026104200004000400800C8B0024E4E0010C40",
INIT_06 => X"8000440802280002700800008A840004A0610000C0000810000C590103600810",
INIT_07 => X"538600220028001890240980A80800200102025000000BF08200002440000883",
INIT_08 => X"00000402C220104131102101040810028528820005100003900E884000010007",
INIT_09 => X"00000005E000000600BCA284140200800C834948100004590111824404012080",
INIT_0A => X"04080000901012100A1141005922000245410002008880000032005080000800",
INIT_0B => X"2000020040044010440104401004010440100401044010040104400802008208",
INIT_0C => X"D1A1344420D2E100000808000000000481000000202002400006800825908402",
INIT_0D => X"0500000000109000000000000580008000080000C852240100068D0B4685A342",
INIT_0E => X"0500000A00000000000000000000028000408020000000050000208020000000",
INIT_0F => X"0000304002100020000000000000000900208004000000050000208004000000",
INIT_10 => X"0000000001200000000A00000000000000000000050000480008000000000000",
INIT_11 => X"009F0080000000004807C0200000000012000020000081000000040000000000",
INIT_12 => X"00000048F8000400000002403E0004000000009067E000000000000000000900",
INIT_13 => X"0000000000000000140000CEE001000000000000000A000036AC008000000000",
INIT_14 => X"03210000000400CA81000000619480D4000400000000000000004100000036E8",
INIT_15 => X"A368DA368DA3685A1685A1685A121A11A1419001512490040024001000008019",
INIT_16 => X"1685A1685A1685A1685A1685A368DA368DA368DA368DA368DA368DA368DA368D",
INIT_17 => X"685A1685A168DA368DA368DA368DA368DA368DA368DA3685A1685A1685A1685A",
INIT_18 => X"CCF48DE68A895C38E250080000000000000000000000685A1685A1685A1685A1",
INIT_19 => X"514514514514514514514514514D34D34D34D34D28E10040392482090157344C",
INIT_1A => X"4D268341A0D069349A0D069349A0D068341A0D068341A0D06834514514514514",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000001654D0D069349A0D068341A4D268341A",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"BE8B45002A974AAAA803DFFFAA843DF45FFFFEAABA0000000000000000000000",
INIT_22 => X"AEBDE00AAFBEAABA080000000087BEAA10F7803DE00FFAEBFFFF0800155FFAAF",
INIT_23 => X"AAEA8ABAAAFBFDE0055556AA005D0415555087BFDE00A2FBD7400F7FBFDFFFA2",
INIT_24 => X"005155555557BE8BEF007FFDEAAAAD1555EF0055401FFF7AEAAA10F780155EFA",
INIT_25 => X"0F7AA974AA082E80010A2AAAAA10552AA8AAA557FC0010F780154105D7FC2145",
INIT_26 => X"BA087BFDF45F7AA974AAAAAA97555F784174BAF7D5555FFF780154AA5D2AA8A1",
INIT_27 => X"F45F7FFFFF55AA80155FF080400145FFFBEAABAF7D17FEBAA2AEBDF45002EAAA",
INIT_28 => X"0000000000000000000000000000000000000000AAFFE8A00552EBFE00F7D17F",
INIT_29 => X"BAFFF080A175D7BEF1E8B6D002090482B68E38FC7BE8A3DF7DF7F5E8A9200000",
INIT_2A => X"BD0400FFF5FDFC7B6A0BDE38B6F5E8A92080E000280071E8A00EB8E3FE10F7AE",
INIT_2B => X"AAA8A38FF8E175C7A2AAAAA82A2F1FAE105D556AA10410E175550871FFE00A2F",
INIT_2C => X"F8A17400557FC015514555757D5D71E8BEF147BFAE82A2DB555C71C5B451D7FF",
INIT_2D => X"FF84174BA5D20AAA00E3AA904BA142A87010A2AEADA38492EA8AAA5571C2000F",
INIT_2E => X"AAAA0BFF7D0024ADA921C7BFFF55FFA095482B6A49256DEB84104BAFFD1525FF",
INIT_2F => X"38492ABDE10EBDF7AF6DE3FFF8F7DB68A105D7000400155FFFBEDA82FFD57DEB",
INIT_30 => X"FEFF7D16AA00000000000000000000000000000000000000000000000A2FBE8A",
INIT_31 => X"AA00AAAABFE00F7AEAABEF082E95545F7D568BEF080402000F7AAA8B55FFAABD",
INIT_32 => X"9754D00517DE00A2FFC2000F7D17FF55FF803FEAAFFD16AA00082E820BA08556",
INIT_33 => X"FD55555D7FD5555FFAAA8AAAFFAA97555A2AEA8A10AAD568A00555168A10002E",
INIT_34 => X"2EAAABA5D5140010F7AE974105D7BC21555D51575EF555568BEF5D7FE8A10AAF",
INIT_35 => X"A84000AAFFD1401E7FF80174AA5D0028A00AAAE800AA552A97400A2AEBDEAA08",
INIT_36 => X"F7FBFFE00FFD17FEAAA2803DFEF08043FE00557BFDF55F78017400F780001FFA",
INIT_37 => X"0000000000A2FFE8ABA082ABFE00AAFBEABFFAAFBEABFFF7AA80145080002145",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000800000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(9),        -- Port A data input
DOA(0)   => data_read_a_hi_256(9),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(9),        -- Port B data input
DOB(0)   => data_read_b_hi_256(9),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_10_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000B0001800002840002C0000281800020030000000033022000000180006",
INIT_01 => X"000008000000004C002000000010026840000000080000080200000000110200",
INIT_02 => X"0000004000800110000006100000003000040800010400004808000000120060",
INIT_03 => X"000200000810020000020000400100000600000000400000001A000040004800",
INIT_04 => X"0004000000000008000200020000000004000000080010004000000200000000",
INIT_05 => X"1000202000011010000000000000010520000400000080000000200000200004",
INIT_06 => X"80004408022800023000000088040004A061000040000810000C490103600000",
INIT_07 => X"120420020028000890240980A808002001020050000009F08000002440000082",
INIT_08 => X"00000402C0201051311001000000020201080200440400000000800000000000",
INIT_09 => X"0000105808000000000000000000008000008088100004590111800004000000",
INIT_0A => X"00804000801210440003C1411008800045000002000014000040009002800000",
INIT_0B => X"0400200000000000000004000040000000000000040000400000000000000221",
INIT_0C => X"0100802000000000000002802000000400100000000002000026000840011400",
INIT_0D => X"0500000000409002082010400400008000400008002044082000081004080204",
INIT_0E => X"0500000200000000000000000000028000400000000000050000200000000000",
INIT_0F => X"0000304002000000000000000000000900200000000000050000200000000000",
INIT_10 => X"0000000001200000000200000000000000000000050000400000000000000000",
INIT_11 => X"0082000000000000480080000000000012000101000080000000000000000000",
INIT_12 => X"0000004810000000000002400400000000000090400000000000000000000940",
INIT_13 => X"0000000000000000150000C00000000000000000000A40001400000000000000",
INIT_14 => X"02000000002400C2810000006000000000000000000000000000410040001400",
INIT_15 => X"020080200802008020080200800800220200840001309A08A848001000008000",
INIT_16 => X"0000000000000000000000000200802008020080200802008020080200802008",
INIT_17 => X"0080200802000000000000000000000000000000000000000000000000000000",
INIT_18 => X"940FE0D397124355520542821010000000000000000000802008020080200802",
INIT_19 => X"28A28A28A28A28A28A28A28A28A28A28A28A28A29554199854514514F546890A",
INIT_1A => X"32994CA6532995CAE572B94CA6532994CA6532994CA6532994CA28A28A28A28A",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000001867172B94CA6532994CA6572B95CAE5",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FC2155F7D155545AA80001EFAAFBEAB45557FFDE100000000000000000000000",
INIT_22 => X"FBE8BFFF78402155AAFBE8B45002A974AAAA803DFFFAA843DF45FFFFEAABA007",
INIT_23 => X"87BEAA10F7803DE00FFAEBFFFF0800155FF00042AB55FFD168B55AA8000010FF",
INIT_24 => X"AAFBEAABAA2FFD741055003DFEFF7AA801FFAAD16AABA002ABDE100800000000",
INIT_25 => X"FF7FBC0145F78028A00A2D142155087BFDE00A2FBD7400F7FBFDFFFA2AEBDE00",
INIT_26 => X"BAF780155EFAAAEA8ABAAAFBFDE0055556AA005D0415555007FD74105555555E",
INIT_27 => X"5EF0055401FFF7AEAAA105D042ABFF5D556AB55AAD168ABA002A975FFF7AEBDE",
INIT_28 => X"0000000000000000000000000000000000000000557BE8BEF007FFDEAAAAD155",
INIT_29 => X"3DF7DF7F5E8A92007BC217DEBDB55555AA8E071D7AAFBEFB455D71F8E0000000",
INIT_2A => X"B6DB55BE8E05000EBFFE8BC7E38E07145BEF1E8B6D002090482B68E38FC7BE8A",
INIT_2B => X"2EB8E00080E000280071E8A00EB8E3FE10F7AEBAFFF080A175D700042AB7DEBD",
INIT_2C => X"FF5FDFC7B6A0BDE38B6F5E8A92B6FBD5410490A3DFD7F7A4821D7A2D16FA8214",
INIT_2D => X"0071D54104951555D7EBF5C5155E3842AA00BED1421450871FFE00A2FBD0400F",
INIT_2E => X"20820955EFE3AEBDEAAFF8E175C7A2AAAAA82A2F1FAE105D556AA10410E17555",
INIT_2F => X"EF147BFAE82A2DB555C71C5B451D7FFAAA8A38410E2ABD749516FB55BED16FA8",
INIT_30 => X"F455D556AA000000000000000000000000000000000000000000000005D71E8B",
INIT_31 => X"2000F7AAA8B55FFAABDFEFF7D16AA00087FC01EFA2FFD7545AAAE97555A2FBFD",
INIT_32 => X"9554500042ABFFA2FFFFF45F7AE97400AAFFE8B45AAAA95545F7D568BEF08040",
INIT_33 => X"400155A2D57FE00552EA8A00082E820BA08556AA00AAAABFE00F7AEAABEF082E",
INIT_34 => X"517DE00A2FFC2000F7D17FF55FF803FEAAFFD16AA00FFFBD5400082EBFF45F78",
INIT_35 => X"55168A10002E9754D085155410085557555AAD557555A2802AA10FFD54214500",
INIT_36 => X"08557DF55F7D17FE000804155FFAAAABDEAAFFAA97555A2AEA8A10AAD568A005",
INIT_37 => X"0000000000555568BEF5D7FE8A10AAFFD55555D7FD5555FFAAA8AAA002AAAB45",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000008FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(10),        -- Port A data input
DOA(0)   => data_read_a_hi_256(10),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(10),        -- Port B data input
DOB(0)   => data_read_b_hi_256(10),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_11_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10180B05A0010402840602C2D001019000000300000000330A20080EC180002",
INIT_01 => X"AB400986B830284D1820E0000C3642484000000008000008820009080A512220",
INIT_02 => X"102A68440080011000000618062AD03502640800010410424908136019920868",
INIT_03 => X"004A0846191B22120642000442C110044600000101E9225CDC9A10844A9A4842",
INIT_04 => X"0094024000250808800216021138000B848000000800100040000102A0600200",
INIT_05 => X"7E4024242008A8102CA88A44010401042200444000888000000028000002A002",
INIT_06 => X"8088445712280000B18812288E0400253855200045C86810000C5B0503286A28",
INIT_07 => X"10008822A028004880200A80880208200122006C000015F0C20408264902C840",
INIT_08 => X"9390040280241041D1754100000018108728820024002B3A01A89540080824C8",
INIT_09 => X"A1001C41A1348498B080801010000080D00301081000045B0511D28D94012339",
INIT_0A => X"44080000901012428003414158230CBA4576708241C010908040341322008000",
INIT_0B => X"040464D280144050C72A0872A0C72A0872A0C72A0C72A0872A0C595043950421",
INIT_0C => X"0804001400000820110A42822204880CD81040442900021704E6000800001D54",
INIT_0D => X"80C62D0500409002082010404580018000404012004004192C10000000000000",
INIT_0E => X"80C62D5803161C526DB40506C120A806ABB0D808CC334A80A54B70D408CC32D2",
INIT_0F => X"2B5144D0DD903C54916D15458C0513005570D408CC334A80A54B70D808CC32D2",
INIT_10 => X"52148C4DB05621E363F813961C20EDA944016558C2347A080B10D8DD6422AA10",
INIT_11 => X"1880144D3345C65593800319C18BD1ECA1C9010112566F10AC4183C340DAE02D",
INIT_12 => X"5810503000633830DE3C2C9C00289A66AA8DE50E0800360614AC281430890600",
INIT_13 => X"0CD2A9CEA8199B6B082B55900314140365320485C4F00AD544407241C175C402",
INIT_14 => X"0000074044C4801832701A89D20A38093631425969020855A281844E00540404",
INIT_15 => X"0000000000000000000000000020C00200088101513492101280401000400200",
INIT_16 => X"2008020080200802008020080000000000000000000000000000000000000000",
INIT_17 => X"0080200802008020080200802008020080200802008020080200802008020080",
INIT_18 => X"804180C0B10A4210420140028400000000000000000000802008020080200802",
INIT_19 => X"000000000000000000000000000820820820820801C414947000000055062608",
INIT_1A => X"0000000004020000000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000001F87E000000000000010080000000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"ABDF5508557DF45002ABDFFFF7803DE10AA80000AA0000000000000000000000",
INIT_22 => X"FFE8A10A28000000007FC2155F7D155545AA80001EFAAFBEAB45557FFDE10082",
INIT_23 => X"02A974AAAA803DFFFAA843DF45FFFFEAABAA2AEBFF45FFAEBFEAA002A801FFF7",
INIT_24 => X"F78402155AAD155555A28428BFF002ABDE00A2AABFE10082ABFFEFAAFBE8B450",
INIT_25 => X"0002A80010A2842AAAA007BFFF4500042AB55FFD168B55AA8000010FFFBE8BFF",
INIT_26 => X"00080000000087BEAA10F7803DE00FFAEBFFFF0800155FF00557FF45557FC201",
INIT_27 => X"1FFAAD16AABA002ABDE10A2D168A10A284021FF5D00154BAF7FBE8BEFFFD5400",
INIT_28 => X"0000000000000000000000000000000000000000A2FFD741055003DFEFF7AA80",
INIT_29 => X"EFB455D71F8E00002EBDF6D005B78F7D142ABDFC7F78E3FE28B684070AA00000",
INIT_2A => X"0BDEAA1C2A801C7E3FFEFA10B68407038007BC217DEBDB55555AA8E071D7AAFB",
INIT_2B => X"20B8FEFBEF1E8B6D002090482B68E38FC7BE8A3DF7DF7F5E8A92BEAEBFF7DEBA",
INIT_2C => X"E8E05000EBFFE8BC7E38E07145B6D15756DA28A28BFF082ABAE10B6AAB8E2808",
INIT_2D => X"08517DF7D497BC5028142A87000A28A2AA92007FF8F7D00042AB7DEBDB6DB55B",
INIT_2E => X"2FFFFEFBC7E3DF42028080E000280071E8A00EB8E3FE10F7AEBAFFF080A175D7",
INIT_2F => X"10490A3DFD7F7A4821D7A2D16FA82142EB8E00B6DB6AA28A280001FF5D0A1048",
INIT_30 => X"EAAF784154BA000000000000000000000000000000000000000000000B6FBD54",
INIT_31 => X"7545AAAE97555A2FBFDF455D556AA00082EBFFEF007BE8BFF5D2ABDF55F7AABD",
INIT_32 => X"6AA00FFAEBFFEFAA803DEBA5D2E82155A2FBFDE00FF84154BA087FC01EFA2FFD",
INIT_33 => X"AAAA00FFAAA8AAA080028BFFF7D568BEF080402000F7AAA8B55FFAABDFEFF7D1",
INIT_34 => X"042ABFFA2FFFFF45F7AE97400AAFFE8B45AAAA95545F7D5555FFAAAAA8BFF002",
INIT_35 => X"7AEAABEF082E9554508557DFFF007BD54BA5D2E95400A2AEA8A00007FEABFF00",
INIT_36 => X"AA80001FF5D2E82000F7FFFFF45AAFFC20BA082E820BA08556AA00AAAABFE00F",
INIT_37 => X"0000000000FFFBD5400082EBFF45F78400155A2D57FE00552EA8A00FFFFE8AAA",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000800000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(11),        -- Port A data input
DOA(0)   => data_read_a_hi_256(11),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(11),        -- Port B data input
DOB(0)   => data_read_b_hi_256(11),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_12_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"A500C4B01BC0268A6940312C0DE045196A831A300500032B333287E4FC812006",
INIT_01 => X"AF400D869830E84D5823E0000C1742484000000008000008820009280A553235",
INIT_02 => X"502A7144008001100000171C022BD13412762A000586235ECC09C8423B960866",
INIT_03 => X"31863846191BA218064204000281200406A10843010022DEDF0852944A9C014A",
INIT_04 => X"0014030000250409000014821038080B840000400800102040000302F0600233",
INIT_05 => X"7FC034348008A8102CA88F48010601042400048000188000000938000002E088",
INIT_06 => X"9CC96CC6F63A5001F12B56A0AC8601F47AC06400D1F80C10020C493F03343A38",
INIT_07 => X"1020002030280098A12048908A16BA311177124C000003F08A94282E5C262861",
INIT_08 => X"827A0602902A10491165E10000049010C52882008600A73A01E8974008092CF8",
INIT_09 => X"47000001A1248008F000000000000080000F010C100204593F11A6CDF48023BF",
INIT_0A => X"040000208010120ACA01400058010CBA4D277C86CCE802B380003C1360008000",
INIT_0B => X"011C46D3C7BC1EF083AF0C3AF083AF083AF0C3AF083AF083AF0C1D7861D78400",
INIT_0C => X"08040014C9001AE91D17E50AD79FEFC87C2154745F82131FFCCE00080000095E",
INIT_0D => X"807BF7118180984004000803D40001880001001400C005031010000000000000",
INIT_0E => X"807BF76A109C944B5891BF06C5EEB14FCBF0D90076D61C807BF7D0D80876D49C",
INIT_0F => X"6DE38EB9FB10350C00A99F7CA80757365E50D80876D61C807BF7D0D90076D49C",
INIT_10 => X"841BCC69A0D8C6F7F0AA001C943A65756A0976EB5A7E7FC8951018186334F311",
INIT_11 => X"D5A014481991C6A737D80211912970CDCDD1864116D6C7080651CB4661F33615",
INIT_12 => X"349E929300423224AE19B9BEC0289033238D4E6EA805892946A9B011A7B152CF",
INIT_13 => X"6244CD7AC01CAAA56B3E6D9001068715D64006D2A961CF9B44512A2504532182",
INIT_14 => X"00000439FDC25C58067A9FAB46095A0B5289A0282D2E1444ACB12A17CF9B4414",
INIT_15 => X"0000000000000000000000040026C00000288401513492909280401000F70A00",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"088881360A95090CB05442029010000000000000000000000000000000000000",
INIT_19 => X"1041041041041041041041041049249249249249200100002D4514510051B946",
INIT_1A => X"592C964B2592C964B2592C964B2592C86432190C86432190C864104104104104",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000002007F592C964B2592C964B2592C964B2",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"43FE0008557DFFF0800020105D557FEAA00557DE100000000000000000000000",
INIT_22 => X"557DFFFF7AA80000082ABDF5508557DF45002ABDFFFF7803DE10AA80000AAAA8",
INIT_23 => X"7D155545AA80001EFAAFBEAB45557FFDE10AAD5420000051555FFA2AA8200000",
INIT_24 => X"A28000000A2D155410F7FFFFEBA08003FE00082AA8AAAAAFFC00BA007FC2155F",
INIT_25 => X"0A2AABFE1055516ABEF5D517DEAAA2AEBFF45FFAEBFEAA002A801FFF7FFE8A10",
INIT_26 => X"55AAFBE8B45002A974AAAA803DFFFAA843DF45FFFFEAABA000028A105D2ABFE1",
INIT_27 => X"E00A2AABFE10082ABFFEF085542000000417555002A820AA08557DFFFF7AA821",
INIT_28 => X"0000000000000000000000000000000000000000AAD155555A28428BFF002ABD",
INIT_29 => X"3FE28B684070AABE803AE38145B78FD7000005010495B7AE921C517DE1000000",
INIT_2A => X"B505FFB6A487000005F7AFD7F7A482038002EBDF6D005B78F7D142ABDFC7F78E",
INIT_2B => X"F5C2082007BC217DEBDB55555AA8E071D7AAFBEFB455D71F8E00BED547038145",
INIT_2C => X"C2A801C7E3FFEFA10B68407038B6D550428FFF1FDE821C003FE001C2EAAAAAB6",
INIT_2D => X"00002FA285D20BDE28A2A4B8E10555B68BEF5D517DEAABEAEBFF7DEBA0BDEAA1",
INIT_2E => X"2005F7DFD7F7A482155BEF1E8B6D002090482B68E38FC7BE8A3DF7DF7F5E8A92",
INIT_2F => X"6DA28A28BFF082ABAE10B6AAB8E280820B8FEF085F4703814001055514208208",
INIT_30 => X"A0055517DE00000000000000000000000000000000000000000000000B6D1575",
INIT_31 => X"8BFF5D2ABDF55F7AABDEAAF784154BAF7802AABA5D7FEAB45080015410007FEA",
INIT_32 => X"6AA00F7D1554BA5D7BC01FFFF8015410007FEAB45F780020BA082EBFFEF007BE",
INIT_33 => X"43FE10552EAAAAAFFD140000087FC01EFA2FFD7545AAAE97555A2FBFDF455D55",
INIT_34 => X"AEBFFEFAA803DEBA5D2E82155A2FBFDE00FF84154BAF7D1400BAFFD57FE005D0",
INIT_35 => X"FAABDFEFF7D16AA0008003FEBA55003DEBAA28428A105D7FEABEF55557DEBAFF",
INIT_36 => X"550402145550000010087FFFF45F78402145F7D568BEF080402000F7AAA8B55F",
INIT_37 => X"0000000000F7D5555FFAAAAA8BFF002AAAA00FFAAA8AAA080028BFF087BD54AA",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000000FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(12),        -- Port A data input
DOA(0)   => data_read_a_hi_256(12),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(12),        -- Port B data input
DOB(0)   => data_read_b_hi_256(12),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_13_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10110A0441812402840402822007818000E00700000000330A3000000008042",
INIT_01 => X"A1400984B830C848180260000C0042604001000008220008A200100802110200",
INIT_02 => X"10A00860009141100000C6180C285035000E0800010431004908135980120C60",
INIT_03 => X"004E20441910221B06420C85D5013804060000000040324C441A108468024842",
INIT_04 => X"0184034010250089C00EA8021938325B04800002091090014880080200000900",
INIT_05 => X"18002424B008881024A8004E01040104270004E0000080090500604840000481",
INIT_06 => X"80004414022A2490B00A142C8C840005794540015E006810001C4B01032C7E20",
INIT_07 => X"510200028028004880280A808816002101022468000011F082040A264006C000",
INIT_08 => X"D2B00402B220104B531001000008001041080200B660E30B200C8040080A9206",
INIT_09 => X"A1000809A93484D21000000000000080C90391881000145B0111A30404015000",
INIT_0A => X"000000008010102A82014100101118BA4510008241480290882400900000A000",
INIT_0B => X"0284484000000000400000000040000000000000040000000000000020000000",
INIT_0C => X"A944AA2000A02000212800020000000D80004084A0000390002E001843210400",
INIT_0D => X"859C1881A04090000000000021800180010341179065441356150A1285094284",
INIT_0E => X"859C188810C65A72A617520252781EA02520D589B9A260859C1840DD81B9A0E0",
INIT_0F => X"0E71F1052D942748C19484E39442D15961C0DD81B9A260859C1840D589B9A0E0",
INIT_10 => X"E60605C0C12CBD400B0810C65A61AA459D0047398500D5889D26907356533C00",
INIT_11 => X"8F60CA1562094650CA28398A42C051E0332181010109294C8E1160CB8C80A561",
INIT_12 => X"2645056D073148580A3C065141942AC4128CA199180C5232575138094450AD0A",
INIT_13 => X"84CA93A2FC008962142B17301A9A1A5196A80245208E0AC5C853C8028163B8C0",
INIT_14 => X"0240034000E4DC8A84000014982372011FC1E475F0F0084A3961F5A80AC5C816",
INIT_15 => X"4250942509425094250942509428D421420882020120981812C8403000088212",
INIT_16 => X"2509425094250942509425094250942509425094250942509425094250942509",
INIT_17 => X"5094250942509425094250942509425094250942509425094250942509425094",
INIT_18 => X"FF3F7DF7FF3E9F7DF7E24502A800000000000000000050942509425094250942",
INIT_19 => X"EBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBF7DFDFDDD555555F7EFBBEE",
INIT_1A => X"7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAEBAEBAEBAEBA",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000000007F7EBF5FAFD7EBF5FAFD7EBF5FAFD",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5554BA087FFFF55557BD54AAF7FBC01FFA2802ABEF0000000000000000000000",
INIT_22 => X"2E80155AA802AB45AA843FE0008557DFFF0800020105D557FEAA00557DE10AAD",
INIT_23 => X"8557DF45002ABDFFFF7803DE10AA80000AA087BD75EF087FFFFEF557BEAB4555",
INIT_24 => X"F7AA80000AAD1420AA087BD7555FFD168AAAFFAE820AA5D5557555082ABDF550",
INIT_25 => X"5FFD157555085140010F7AEAABFFAAD5420000051555FFA2AA8200000557DFFF",
INIT_26 => X"45007FC2155F7D155545AA80001EFAAFBEAB45557FFDE10AAAEA8BFFA2FBD754",
INIT_27 => X"E00082AA8AAAAAFFC00BA00002AAAAF7D5574BA557BE8A10A284154BAFFAAAAB",
INIT_28 => X"0000000000000000000000000000000000000000A2D155410F7FFFFEBA08003F",
INIT_29 => X"7AE921C517DE10A2DB50482147FFAF554971D0492E3F1C71C7BE8A2ABD700000",
INIT_2A => X"FFAFD7497BE8B5555208217DBE8A2AB45BE803AE38145B78FD7000005010495B",
INIT_2B => X"5F5056D002EBDF6D005B78F7D142ABDFC7F78E3FE28B684070AA1C71D25D7007",
INIT_2C => X"6A487000005F7AFD7F7A482038AADF47092147FD257DFFD568A82FFA4870BA55",
INIT_2D => X"A2A0ADBC7A2FFD257DE3DF52555085142000FFAAAFBFFBED547038145B505FFB",
INIT_2E => X"0B680124BAFFAAAFB45007BC217DEBDB55555AA8E071D7AAFBEFB455D71F8E00",
INIT_2F => X"28FFF1FDE821C003FE001C2EAAAAAB6F5C20821C002AA92FFDF574824171EAA1",
INIT_30 => X"545F7AEA8B55000000000000000000000000000000000000000000000B6D5504",
INIT_31 => X"AB45080015410007FEAA0055517DE00A2FFC00105D7BE8B55085142010AAD157",
INIT_32 => X"154BA5D5140145007BE8B55087BEAB555D04001EFF7AAA8B55F7802AABA5D7FE",
INIT_33 => X"16AA10FF80174AA557FC21EF082EBFFEF007BE8BFF5D2ABDF55F7AABDEAAF784",
INIT_34 => X"D1554BA5D7BC01FFFF8015410007FEAB45F780020BAA2FFD54105D7FC21EFFFD",
INIT_35 => X"2FBFDF455D556AA00A2803FF45AAFFC21EFAAFBC0155085540000FFAEBFFEFF7",
INIT_36 => X"F7FBD5410085568A10FF80020AAFFAABFF55087FC01EFA2FFD7545AAAE97555A",
INIT_37 => X"0000000000F7D1400BAFFD57FE005D043FE10552EAAAAAFFD1400005D042AA00",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000CFFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(13),        -- Port A data input
DOA(0)   => data_read_a_hi_256(13),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(13),        -- Port B data input
DOB(0)   => data_read_b_hi_256(13),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_14_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10020A000180000284008280000281800000030000000033022000000580002",
INIT_01 => X"A140098018300848184860000C20C24040000000084000084200000000110200",
INIT_02 => X"1020006000900110000006102028503400040800010400204908012018120E64",
INIT_03 => X"000200441910221006420000400100040600000000E9E401209A108448004842",
INIT_04 => X"0004020000250008000200021038000804000000090090004800080200000000",
INIT_05 => X"500024240008881024A800400104010420000400000080080100204040000000",
INIT_06 => X"8000440102282015B10A10288E0400042345400040006810000C5901033D7880",
INIT_07 => X"1100000200280048802008828812002001220064000005F1C2850A2649204070",
INIT_08 => X"00B00402802010411110010000080010010802000400230B000C804008080002",
INIT_09 => X"01000009A92480001000000000000080C8038188100004590111B68404010000",
INIT_0A => X"0000000080101000000141001001088A45000082400000008020009000008000",
INIT_0B => X"0004404000000000400004000000000000004000000000000004000000000000",
INIT_0C => X"8904A0200080200001080002000000088000400420000200002E000841010400",
INIT_0D => X"0500000C80409000000000000000018000000000806044010014081204090204",
INIT_0E => X"0500005813A0210D072E8D012001028402908004000587050000108004000707",
INIT_0F => X"9004300044900812386A280E5800088980108020000587050000108020000707",
INIT_10 => X"DE00482E19E30002007813A02096038AE200880405200308828062A68C0BC700",
INIT_11 => X"00000E5A08E6000048001292B83280001208A1011004011060049A1C59192055",
INIT_12 => X"492060480256530650000240001DB011CC00009000032C4C979E3806180C0900",
INIT_13 => X"5A3433EDE00154181400000007BCBD858F120120541A0000000033757465B2C0",
INIT_14 => X"02002C000024008A84001A0902000422E3E99681004802115652594000000001",
INIT_15 => X"0240902409024090240902409028D021020880000120901812C8401000000210",
INIT_16 => X"2409024090240902409024090240902409024090240902409024090240902409",
INIT_17 => X"4090240902409024090240902409024090240902409024090240902409024090",
INIT_18 => X"5C8FF0F7BE9D5F7DF65040028000000000000000000040902409024090240902",
INIT_19 => X"79E79E79E79E79E79E79E79E79E79E79E79E79E7BF7DDDDDFCF3CF3DF5579B4E",
INIT_1A => X"3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE79E79E79E79E",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000003FF803F9FCFE7F3F9FCFE7F3F9FCFE7F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"BE8B55A2AE80000F7D5555555D2AAAABAAAD1420BA0000000000000000000000",
INIT_22 => X"00155EF0804155EFAAD5554BA087FFFF55557BD54AAF7FBC01FFA2802ABEFA2F",
INIT_23 => X"8557DFFF0800020105D557FEAA00557DE10A2AA801FFA28402000AAAE9554555",
INIT_24 => X"AA802AB4500516AA00A2AE800BAFFFFC20BAF7AEA8B45080417400AA843FE000",
INIT_25 => X"0A2843FEBAFFFBD7410A2D168BFF087BD75EF087FFFFEF557BEAB45552E80155",
INIT_26 => X"AA082ABDF5508557DF45002ABDFFFF7803DE10AA80000AA005568ABAA2840201",
INIT_27 => X"AAAFFAE820AA5D5557555002E80155A280000005D7FFDF4555517DFEF00043FE",
INIT_28 => X"0000000000000000000000000000000000000000AAD1420AA087BD7555FFD168",
INIT_29 => X"C71C7BE8A2ABD7A2FFEDB55B6A080038E3DB50555412AA8ABAAADB4009200000",
INIT_2A => X"402038AAAA955554900105FF0800175D7A2DB50482147FFAF554971D0492E3F1",
INIT_2B => X"0A12410BE803AE38145B78FD7000005010495B7AE921C517DE10A2AE851FFB68",
INIT_2C => X"97BE8B5555208217DBE8A2AB451C556FA00A2A0800BAE3F1C0092EBAAADB6D08",
INIT_2D => X"00516DABAA28402038B6803DE82F7F5D5410A2D568BC71C71D25D7007FFAFD74",
INIT_2E => X"55D5F78FD7000E3FEAA002EBDF6D005B78F7D142ABDFC7F78E3FE28B684070AA",
INIT_2F => X"92147FD257DFFD568A82FFA4870BA555F5056D002A80155B680000105D7FF8F4",
INIT_30 => X"AAAAAFFC2000000000000000000000000000000000000000000000000AADF470",
INIT_31 => X"8B55085142010AAD157545F7AEA8B55A2FBFFF55FF84000AAAAFBC0145002AA8",
INIT_32 => X"7DE00A2AA955FFFF80020BAAAAA975450800001EF080417555A2FFC00105D7BE",
INIT_33 => X"140000A2AEBFFEF082A82010F7802AABA5D7FEAB45080015410007FEAA005551",
INIT_34 => X"5140145007BE8B55087BEAB555D04001EFF7AAA8B555D557FE00A280020BAAAD",
INIT_35 => X"7AABDEAAF784154BA08557FEAAA284000AAFF803DE00FFD557400AAD56AB455D",
INIT_36 => X"F780020105D7BEAB45557BE8B45082EBFEBA082EBFFEF007BE8BFF5D2ABDF55F",
INIT_37 => X"0000000000A2FFD54105D7FC21EFFFD16AA10FF80174AA557FC21EF082A80145",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000000FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(14),        -- Port A data input
DOA(0)   => data_read_a_hi_256(14),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(14),        -- Port B data input
DOB(0)   => data_read_b_hi_256(14),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_15_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000A000000000284000280000001800020030000000033022000000180002",
INIT_01 => X"A140098018300848180060000C00424040000000080000080200000000110200",
INIT_02 => X"102100400C8011100000061000A8503401044880010430004808000180122378",
INIT_03 => X"000200541D102210064200000045000546080000400020000008108448400042",
INIT_04 => X"8094020000254C880000028A1018000844000000880013504000002600000000",
INIT_05 => X"10002424000AA81024A82040010C61062001440002988000000024808001004B",
INIT_06 => X"80004400022A00003C8912248E0400042854400040006810000C4901032B1800",
INIT_07 => X"50200000B0280048A0280A828801002101020040000005F38204082640000000",
INIT_08 => X"01F00402802610411100110000000010010802000400230A0008884008080004",
INIT_09 => X"01000001A12481041000000000000080C0030108100004590111820404000000",
INIT_0A => X"0000000080101000004140001001088A45000082000000008000001080008000",
INIT_0B => X"0004404000000000400004000040000400000000000000000004000020000200",
INIT_0C => X"0804000020024100012808020000000981004004A0200310000C000800000000",
INIT_0D => X"0000001180009000000000002100018000000000004004010010000000000000",
INIT_0E => X"00000008000002000000000000000000000080A40000000000000080A4000000",
INIT_0F => X"00000000001000204800000000000000000080A40000000000000080A4000000",
INIT_10 => X"000000000000000000080000020000000000000000000008000C020000000000",
INIT_11 => X"000000824000000000000020220000000001800100020300000004003420480A",
INIT_12 => X"0000000000040440000000000001048000000000000000100800400000000000",
INIT_13 => X"000800000000000000000000000100C220050000000000000000008220884400",
INIT_14 => X"000000000000000830000000000000000016101C5C1400000000000000000000",
INIT_15 => X"0000000000000000000000000020C00000088000012090101280401000000200",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000040028000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"000010082A954BA00003DFEF085155400F78428BEF0000000000000000000000",
INIT_22 => X"8015400FF84001EFA2FBE8B55A2AE80000F7D5555555D2AAAABAAAD1420BAFF8",
INIT_23 => X"87FFFF55557BD54AAF7FBC01FFA2802ABEFF7AE95555A2FBE8BEFA2843DE00AA",
INIT_24 => X"0804155EFFFFBE8BFF0800174AA557BFDE10A2FBEAB45F7D56AABAAAD5554BA0",
INIT_25 => X"5FFD568BEF087FE8A1055003FE00A2AA801FFA28402000AAAE955455500155EF",
INIT_26 => X"45AA843FE0008557DFFF0800020105D557FEAA00557DE10F7D1574AAA2D16AB5",
INIT_27 => X"0BAF7AEA8B45080417400FFFFC2145080015400AA802AA00AAAE800BA5D00155",
INIT_28 => X"000000000000000000000000000000000000000000516AA00A2AE800BAFFFFC2",
INIT_29 => X"A8ABAAADB40092E38E070280024904AA1C0438FD7005150438F78A2DBFF00000",
INIT_2A => X"FE8BC7BE8E38E10A28017400E38A051FFA2FFEDB55B6A080038E3DB50555412A",
INIT_2B => X"D16AABAA2DB50482147FFAF554971D0492E3F1C71C7BE8A2ABD7E3AA9257DA2F",
INIT_2C => X"AAA955554900105FF0800175D7E3FFEFBD70000124AA557FFDE10A2FBEDB6DF7",
INIT_2D => X"FFDF50482A2DB6AB45FFD56DBD7087BEAA38410038E38A2AE851FFB68402038A",
INIT_2E => X"0AAA085082550A1057DBE803AE38145B78FD7000005010495B7AE921C517DE10",
INIT_2F => X"00A2A0800BAE3F1C0092EBAAADB6D080A12410FFF1C017D140410400BE8E28A1",
INIT_30 => X"0AAF7AEBDFEF0000000000000000000000000000000000000000000001C556FA",
INIT_31 => X"00AAAAFBC0145002AA8AAAAAFFC2000AAAA974AA0800020BA550028B55085540",
INIT_32 => X"A8B55AAAE821EFAAFBEAB55F7AAA8A00AA8417400AAAE975EFA2FBFFF55FF840",
INIT_33 => X"BFFE10A2FFFFFEFF7D568ABAA2FFC00105D7BE8B55085142010AAD157545F7AE",
INIT_34 => X"AA955FFFF80020BAAAAA975450800001EF080417555AAFFFDF450804020AA557",
INIT_35 => X"07FEAA0055517DE00FFFBC2000AAFBE8B55F7D17DF45007FE8AAA08002AAAAA2",
INIT_36 => X"5D0000010F7AAA8A10AA8017400552A801EFF7802AABA5D7FEAB450800154100",
INIT_37 => X"00000000005D557FE00A280020BAAAD140000A2AEBFFEF082A82010FFD5421EF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000C00000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(15),        -- Port A data input
DOA(0)   => data_read_a_hi_256(15),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(15),        -- Port B data input
DOB(0)   => data_read_b_hi_256(15),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_16_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"DA22C618B1000482B688B186588884862A400438255FC38381441205BA803003",
INIT_01 => X"264AC80028404C211203A952A90341080B173340412000E1005D628000820484",
INIT_02 => X"400034C206C405000001A48202084004003008255040826EE008B440200E2042",
INIT_03 => X"A459C1240181AB20AD27315B7F1983CA1C900040422A005762010010000C0400",
INIT_04 => X"296E542B6E3A825C15FB385321B4ADFE16AB45FD2C400002E205231201290A28",
INIT_05 => X"B9E5815006028179808C00A0D2152B90707A1E0BD423CAC0000D610000000710",
INIT_06 => X"81F104A1415C292164280081C6AB88742086ACACDE240000A80090CE82A803B9",
INIT_07 => X"400800000ACCAA280940580400A37B8896CA4D000A80C1102A00001C14028009",
INIT_08 => X"0015452880C8D90409A02D965965200100104F2B00822512000000231520A024",
INIT_09 => X"A5AA80018120E00066000000000012C9000A0000D0A80000BF8028E87C1B9927",
INIT_0A => X"00520228080108039501200848002912300208092B940192D1000000000000A8",
INIT_0B => X"03561180063DB4F6110001100011000110001100011000110001080008800080",
INIT_0C => X"080200854409418B02ED0000502A02972000040BB401100010012B4C90000100",
INIT_0D => X"6D061A1F8D60D80820500101244AA8A2AA242E80000009200120000000000000",
INIT_0E => X"6D066210E5001DB4A5B400C7D553847165A99000C6564CDD051DC99000C65555",
INIT_0F => X"21D0C48F254946148107354292673D1F72C99000C6564CDD0565C99000C65555",
INIT_10 => X"952D2058F33225787810F5001D6121A9559224D1FF97D0272F04D89441A56D8A",
INIT_11 => X"6C1C74485B81E31306C71D1093AB8A64811BADC00992180D58033B1172F2A025",
INIT_12 => X"7B86DED8E3A212748F0E0CA638E890B7A8546120C0AFF5B548AC431FB1C7DB07",
INIT_13 => X"EFCE9B26DECA1AD36A2E4F40DF6AAAF260AF88899E8B8B93D12A877178DD0032",
INIT_14 => X"A8009F8B108C80A1021B9A8BB8056662CA1951596800FC01A38D4D4B072B922F",
INIT_15 => X"00000000000000000000000000044000102A0001148442A1108103595580A840",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"4C690DA64C1C4F68A36040000000000000000000000000000000000000000000",
INIT_19 => X"D14D14D14D14D14D14D14D14D14514514514514529E5F87869E79E78558D1154",
INIT_1A => X"3D1E8F47A7D3E9F4FA7D3E9F4FA7D3E9F47A7D1E9F47A7D1E9F4D14D14D14D14",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE000000000000000007D3E9F4FA7D3E8F47A3D1E8F47A",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFEFF7D168B55AAD17FFFF552EBFE00007FC00AA0000000000000000000000",
INIT_22 => X"04000BA552A821FFFF8000010082A954BA00003DFEF085155400F78428BEF087",
INIT_23 => X"2AE80000F7D5555555D2AAAABAAAD1420BA5D2E975EFF7D568BFFFF80175EF00",
INIT_24 => X"FF84001EF0000020AA5D00154005D043FF45555540000082EAABFFA2FBE8B55A",
INIT_25 => X"0087FD74BAAAAEBFFEF557FC00AAF7AE95555A2FBE8BEFA2843DE00AA8015400",
INIT_26 => X"FFAAD5554BA087FFFF55557BD54AAF7FBC01FFA2802ABEF557BEABEF5D041541",
INIT_27 => X"E10A2FBEAB45F7D56AABA082A97545F7D16ABFFFFAABFEAAFF84001FF002A821",
INIT_28 => X"0000000000000000000000000000000000000000FFFBE8BFF0800174AA557BFD",
INIT_29 => X"50438F78A2DBFF0871F8FC7E3D56AB6DBEDB7FFEF552AB8E38087FC209200000",
INIT_2A => X"16ABFFE38E175EF1400000BA412E871FFE38E070280024904AA1C0438FD70051",
INIT_2B => X"2EAFBD7A2FFEDB55B6A080038E3DB50555412AA8ABAAADB400924920925EFF7D",
INIT_2C => X"E8E38E10A28017400E38A051FF0804050BA410A1240055003FF6D5551420101C",
INIT_2D => X"4975EDBC7550E12410087FD74AAB6AABFFC7557FC00BAE3AA9257DA2FFE8BC7B",
INIT_2E => X"AF780051C70824851D7A2DB50482147FFAF554971D0492E3F1C71C7BE8A2ABD7",
INIT_2F => X"D70000124AA557FFDE10A2FBEDB6DF7D16AABA08249756DF7D168BC7F7AABAEA",
INIT_30 => X"AAA007BC0000000000000000000000000000000000000000000000000E3FFEFB",
INIT_31 => X"20BA550028B550855400AAF7AEBDFEF08516AB55A2D16ABEFFFFBFDFFF552AAA",
INIT_32 => X"C20000000021EFF7D568BFFA2AA955FF5D04020AA002A955EFAAAA974AA08000",
INIT_33 => X"03DFEF5D51420005D2ABFF45A2FBFFF55FF84000AAAAFBC0145002AA8AAAAAFF",
INIT_34 => X"AE821EFAAFBEAB55F7AAA8A00AA8417400AAAE975EF0800174BA002E820105D0",
INIT_35 => X"AD157545F7AEA8B5500557DF45552A82000007BD74AAF7AEBDF455D7BC20BAAA",
INIT_36 => X"F7D568B55FFAAAAABAFF8415545000015555A2FFC00105D7BE8B55085142010A",
INIT_37 => X"0000000000AAFFFDF450804020AA557BFFE10A2FFFFFEFF7D568ABA0804155FF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000400000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(16),        -- Port A data input
DOA(0)   => data_read_a_hi_256(16),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(16),        -- Port B data input
DOB(0)   => data_read_b_hi_256(16),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_17_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"5284CE4FB7BD2C8994A13392DBD02E14006B82AC7E800D44D3DD2FD5F9B961C0",
INIT_01 => X"F9BA301F7E03FC6793F2199B39FC233C11D93AE6F3BB92B32091DBC339B24542",
INIT_02 => X"1D5FC0C08F040404446965C0607FB8A217C400C33A908078551BD04222186338",
INIT_03 => X"8504930A37F65820CB24111B7F08014A0AB84A52B6D2AFF97C1B5AC757F06D6B",
INIT_04 => X"250834336D1E81500FDB38302292ADFE103B6DBD204037F202042075E2B1D00A",
INIT_05 => X"8F039786062C6CE092F5FE005236781C402A0807B4070670083DC68206D7E6D0",
INIT_06 => X"0CD26803C3582408962C58B183F8AEF42045919B30E085DD2ED57D4EED08CA6A",
INIT_07 => X"700000B30380670B8142500448E3E01E94EF1340A28AC1AC8156044D1400AA00",
INIT_08 => X"009F3A1B0120A1C51DFFC40C30E5F0182D0950190C0810BE00E9A76E4C6FFBE4",
INIT_09 => X"8FCCC200A59BDD2FFE3F3EC7C7DEF207000F00059D2ED56D7EED2ED3C9A867DC",
INIT_0A => X"0617112E46F05D02DD814102F800633F1D0A7CC9AE7A08BFF0001D35682AC0CE",
INIT_0B => X"8A3F06ABD73DBCF4FBCF4FBCF4FBCF4FBCF4FBCF4FBCF4FBCF4FBE7A7DE7A780",
INIT_0C => X"001000974F08518F5AFFC94B533FADA7FDE97D6BFF329E1B50FF99F086000D9E",
INIT_0D => X"F50B018F95EA3DED1652EC0B27E67F419E2E1E8000C0036340B8000000000000",
INIT_0E => X"F50B01C8DF7F96197DB4AFC8C8886AF672A1537F759299F50B03C1537F759199",
INIT_0F => X"6068331C5103E7EF0FBEED6BB6A9412007C1537F759299F50B03C1537F759199",
INIT_10 => X"21F2CD7F252CDABB3CE8CF7F963AB9FD6AD434201AA68B837FFD1F7B7125B68C",
INIT_11 => X"BD055EB6D555CB2949C15BA7270FF256526BBFD55BBE71D79F73C7AC6DB9BF37",
INIT_12 => X"94080BF82B74E4E1FE4ACA4E0ABD6DAAAB965293036FF6B652A99A6026027FBE",
INIT_13 => X"EF5CBA7A43482800FEFAFD06B8CFCCAB7550D0C2022EAEBD438697AD2EBA9168",
INIT_14 => X"AC00A8BBFC8B501CF7A0FED9A548FA19752C4A4EADAE42FCBC38C3B7BEBF42CF",
INIT_15 => X"0000000000000000000000000026E100002F382DBD9ECFE117805F20CFDAAB00",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"09EDCC4052E917114F981800C000000000000000000000000000000000000000",
INIT_19 => X"EBA69AEBA69A69AEBA69AEBA69A69A69A69A69A68698686981D75D7443720030",
INIT_1A => X"46A351A8D068341A0D068341A0D068341A0D46A341A0D46A341A69AEBA69A69A",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000000000046A351A8D46A351A8D46A351A8D",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFEFF7FBEAB450804001EFAAD57FEAA0000000000000000000000",
INIT_22 => X"51401EF087FD74AA087FFFFEFF7D168B55AAD17FFFF552EBFE00007FC00AA087",
INIT_23 => X"82A954BA00003DFEF085155400F78428BEFAAD168A000004020AA5D7BE8B4500",
INIT_24 => X"552A821FF5D00020BA552A82000552A821555D7FEAB55FF80175EFFF80000100",
INIT_25 => X"FAAFBC01EF5D0015555557BFDEBA5D2E975EFF7D568BFFFF80175EF0004000BA",
INIT_26 => X"BAA2FBE8B55A2AE80000F7D5555555D2AAAABAAAD1420BAFFFFFDF45AAD17FFF",
INIT_27 => X"F45555540000082EAABFF00516AA10552E820BA007FEABEF005555555A2D1554",
INIT_28 => X"00000000000000000000000000000000000000000000020AA5D00154005D043F",
INIT_29 => X"B8E38087FC2092147FFFFFFFFFBFDFC7EBF5E8B550000071EFB6DF7AE9200000",
INIT_2A => X"A07082497FEFB6D1451471EF007BD04920871F8FC7E3D56AB6DBEDB7FFEF552A",
INIT_2B => X"8E175FFE38E070280024904AA1C0438FD7005150438F78A2DBFFBED16AA381C0",
INIT_2C => X"38E175EF1400000BA412E871FF550A00092492A850105D2A80155417BEFB6DEB",
INIT_2D => X"FFF5FFF6DAADF7FFD7B6F1C71EF55001756D5D7BFAEBA4920925EFF7D16ABFFE",
INIT_2E => X"700515556DA2DF50492A2FFEDB55B6A080038E3DB50555412AA8ABAAADB40092",
INIT_2F => X"BA410A1240055003FF6D5551420101C2EAFBD7145B6AA28492487082007FEDBD",
INIT_30 => X"5EFFFFBEAA000000000000000000000000000000000000000000000000804050",
INIT_31 => X"ABEFFFFBFDFFF552AAAAAA007BC0000557FFDFEFF7FBFFF55A2D16AB55000017",
INIT_32 => X"BDFEFF7D568AAA5D2A97410007BFFFFF5551555EF087FC200008516AB55A2D16",
INIT_33 => X"A82155087FFFFEFAAAA975EFAAAA974AA0800020BA550028B550855400AAF7AE",
INIT_34 => X"00021EFF7D568BFFA2AA955FF5D04020AA002A955EF5D2E80010002A954005D2",
INIT_35 => X"02AA8AAAAAFFC2000FFD57DFFFAAFFFDF55FFD1575FF5504175EF5D7FEAAAA00",
INIT_36 => X"000415410007BFFF450051555EFA2FBC0000A2FBFFF55FF84000AAAAFBC01450",
INIT_37 => X"00000000000800174BA002E820105D003DFEF5D51420005D2ABFF45557FE8AAA",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000CFFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(17),        -- Port A data input
DOA(0)   => data_read_a_hi_256(17),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(17),        -- Port B data input
DOB(0)   => data_read_b_hi_256(17),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_18_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"69844019080000A21A611406840014122A641074155FC28A2024001001801003",
INIT_01 => X"01067920034004180005E9E3C90360C0041C0181002001602025800008440084",
INIT_02 => X"40AC3CAA22D605200000856E2481902400344A20F802C22054001000021E2379",
INIT_03 => X"A54C23B34C81EB2076471000800981140C010101750D1007E58040102B0E0100",
INIT_04 => X"22660C1C0065003C04040013236E105016A028402D618803EB092B9201490B2A",
INIT_05 => X"B8E080000000005889AC41E04508A99070200E010001C1CA11803850C8000100",
INIT_06 => X"800A4CE301545001F40050216C09950004C2047BCF1C8090C02800C0120886B3",
INIT_07 => X"814A0080064C1F300020080182001A9E02C03400082002700000217294007101",
INIT_08 => X"000117088080990419002D86184A01018030430700802541420440022030041A",
INIT_09 => X"7030C30B885200D274004008080003C32A10A19090C02010E102294406168800",
INIT_0A => X"00602A01880980037109700C04C44C92A88DCC2211E44174112840880000060D",
INIT_0B => X"11C0D95C20C2030A003080030800308003080030800308003080018400184004",
INIT_0C => X"8304E02809832E6021002020404042000F00008400811824AD4007ECD9436261",
INIT_0D => X"0AFCE5D22A82B20000520100C801F8A07E103000A1285C84000418360C1B060D",
INIT_0E => X"0AFCFD8CB17E5B4F045557575E6EFBE3942C1040A41D660AFCE1CC1040A41E66",
INIT_0F => X"8E7FFBB385661C08D1455ABA91E6FF5FDFCC1040A41D660AFCF9CC1040A41E66",
INIT_10 => X"015F82C006C3AF31E64CB17E5A9655017F1FC73FAF1D61B1040294C58AD1FF5F",
INIT_11 => X"B95454005BAA36DCF8E519001BF80DEB3EE2020EA678189C6EC32881F7F75648",
INIT_12 => X"67D7EDFCA320037E81BD77D728A800B7546DBDFF12904747A351145FC53ABF8D",
INIT_13 => X"92B764225C57C97EBE76E1254F0C0D4514A84F5573FE9DBA4A38E247C522CC0E",
INIT_14 => X"BE84370001B6922070440556B15F7FABBC40151D7C747D8220673C3B9DB84B20",
INIT_15 => X"06C1B06C1B06C1B06C1B06C1B0491069068000004060300A005A01183F240014",
INIT_16 => X"6C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B",
INIT_17 => X"C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B0",
INIT_18 => X"B80EE173C2300F7DF16000000000000000000000000041B06C1B06C1B06C1B06",
INIT_19 => X"AAAAAA28A28A28AAAAAAA28A28A28A28A28A28A2910591505C104104B28BBECE",
INIT_1A => X"128944A25128944A25128944A25128944A2552A954AA5128944AAAA28A28A28A",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000128944A25128944A25128944A25",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFDFEF5D2A974BA082E954000000000000000000000000",
INIT_22 => X"0028B55002E82000087FFFFFFFFFFFFFEFF7FBEAB450804001EFAAD57FEAA087",
INIT_23 => X"7D168B55AAD17FFFF552EBFE00007FC00AA087FFFFFFFFFBFDF45AAD568B5508",
INIT_24 => X"087FD74AAAAFFFDF45A2D16AB55F7FFFFFFF00043DE10AA843DE00087FFFFEFF",
INIT_25 => X"A55042ABEF5D7FD75FFAAD540145AAD168A000004020AA5D7BE8B450051401EF",
INIT_26 => X"45FF8000010082A954BA00003DFEF085155400F78428BEFAA80000000804154B",
INIT_27 => X"1555D7FEAB55FF80175EF5D00020105D2A97400082E95555085168A10557FD75",
INIT_28 => X"00000000000000000000000000000000000000005D00020BA552A82000552A82",
INIT_29 => X"071EFB6DF7AE921C7FFFFFFFFFFFFFFFF7FBFDFFF5D2A954AA082A9242800000",
INIT_2A => X"1FAF55A2DF6DB7D1C002AB7D002A82028147FFFFFFFFFBFDFC7EBF5E8B550000",
INIT_2B => X"8E38E280871F8FC7E3D56AB6DBEDB7FFEF552AB8E38087FC2092087FFDFC7E3F",
INIT_2C => X"97FEFB6D1451471EF007BD0492B6F1F8F55AADF6DB7DE3F5FAFC708003DE28B6",
INIT_2D => X"A28407038140410492550A2ABC7497BD25FFAADF4516DBED16AA381C0A070824",
INIT_2E => X"D1C516FA28417BD5545E38E070280024904AA1C0438FD7005150438F78A2DBFF",
INIT_2F => X"92492A850105D2A80155417BEFB6DEB8E175FF5D0E05000492097428002E9557",
INIT_30 => X"4AA082A820AA000000000000000000000000000000000000000000000550A000",
INIT_31 => X"FF55A2D16AB550000175EFFFFBEAA00557FFFFFFFFFFFDFEFF7FBFFFEF552E97",
INIT_32 => X"C0000087BFDF45AAD568B55AAFBFDFEF55042ABEF002A800AA557FFDFEFF7FBF",
INIT_33 => X"16AB4500043DEAAFFAEAAAAA08516AB55A2D16ABEFFFFBFDFFF552AAAAAA007B",
INIT_34 => X"D568AAA5D2A97410007BFFFFF5551555EF087FC2000FFD56AB45A2FFFDFFFAAD",
INIT_35 => X"855400AAF7AEBDFEFA280154BA550400000552AA8B45087FC01EFA2FFD55EFF7",
INIT_36 => X"0804154BA082A975EF5D517DEAA007BD5545AAAA974AA0800020BA550028B550",
INIT_37 => X"00000000005D2E80010002A954005D2A82155087FFFFEFAAAA975EF5D2E97400",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000400000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(18),        -- Port A data input
DOA(0)   => data_read_a_hi_256(18),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(18),        -- Port B data input
DOB(0)   => data_read_b_hi_256(18),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_19_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"042200000000000041088001001AA00000000000000000000000500802000003",
INIT_01 => X"074018000024000000000404000000000A22000800000800004A200000000001",
INIT_02 => X"0000048002C405000000000006A84000000000200893C246A20000000020031A",
INIT_03 => X"082A58E411004B2000071000000981000C000000002045000200000000000000",
INIT_04 => X"200604000000001C0400001320000000162000002C4000026201201200090800",
INIT_05 => X"1020800000000058840200204000099070200E010001C0400000000000000000",
INIT_06 => X"0012048037805421402850001402498820022802400480405008901100A00102",
INIT_07 => X"00000000020C0130481204919200010C82000000000006002A548902A0020109",
INIT_08 => X"0001150800009900000005861840000000004301000B000000000001C1C00000",
INIT_09 => X"001F00002024B20002000000000002C300000000405000103010204000000000",
INIT_0A => X"00000000000000000000000000000040002000044000000000000000000002F0",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000420003B00000000000000000040012C80000000",
INIT_0D => X"45001A03C0825A0D20800000000018A006001000000000000000000000000000",
INIT_0E => X"450002131E01A1F6EA0A0020211146E069C2ACC01AE80045001D82ACC01AE800",
INIT_0F => X"1188340C3E1CFAD27CC2E004481020892282ACC01AE80045000582ACC01AE800",
INIT_10 => X"DEA03228D810007019931E01A1E5BA02802008C06F029D4C7B76639CEC0A0020",
INIT_11 => X"428AA3592000000206C2A4DAC00000008113C246A181C03FE4662A84575768DF",
INIT_12 => X"08201090549B5800000000261546B24000000000C53807E7CC06618018C51210",
INIT_13 => X"13F6A185A0A0168128411ACB800C0E108A0720288C011046B5986247C5452291",
INIT_14 => X"0000C220010808C10D9A92A74CD7CF4A080031B1515B212143D841431046B58A",
INIT_15 => X"00000000000000000000000000000000000000000000000000000118030004E0",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"3F0C7010C660C744192000000000000000000000000000000000000000000000",
INIT_19 => X"1861861861869A61861861861861861861861861A8208C4C1534D34C07208BBA",
INIT_1A => X"0984C26130984C26130984C26130984D26930984C26130984C261861861869A6",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE000000000000000000984C26130984C26130984C2613",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF552A974AA0004174BA0000000000000000000000",
INIT_22 => X"2E974BAA2FFFFE10087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974BA082E95400F7F",
INIT_23 => X"FFFFFFEFF7FBEAB450804001EFAAD57FEAAF7FFFFFFFFFFFFFFFFF7FBFDFFF55",
INIT_24 => X"002E82000F7FFFFFFFFFFFFDFEFA2D568B550004001EFAAAEA8ABA087FFFFFFF",
INIT_25 => X"5AAD16ABEF5D2ABFF55080402010087FFFFFFFFFBFDF45AAD568B55080028B55",
INIT_26 => X"BA087FFFFEFF7D168B55AAD17FFFF552EBFE00007FC00AAF7FFFFFFFF7FBE8B5",
INIT_27 => X"FFF00043DE10AA843DE00557FFDFEFA2D16AB55A2FFFDFEF5D2EBFE00AAFFFFE",
INIT_28 => X"0000000000000000000000000000000000000000AAFFFDF45A2D16AB55F7FFFF",
INIT_29 => X"954AA082A92428E3FFFFFFFFFFFFFFFFFFFFFFFEF552A974AA0000104AA00000",
INIT_2A => X"FFDFEFF7F5FAFC7492A974AAB6F5F8E101C7FFFFFFFFFFFFFFFF7FBFDFFF5D2A",
INIT_2B => X"A4A8AAA147FFFFFFFFFBFDFC7EBF5E8B550000071EFB6DF7AE92EBFFFFFFFFFF",
INIT_2C => X"2DF6DB7D1C002AB7D002A82028FFFFFFFEFF7F1F8FD7AAD16AB450000001FFBE",
INIT_2D => X"F7FBF8FC7E3F5EAB45B6DF6FBEF5D2AB8F7D000000010087FFDFC7E3F1FAF55A",
INIT_2E => X"7412ABFE28B6F5F8E820871F8FC7E3D56AB6DBEDB7FFEF552AB8E38087FC2092",
INIT_2F => X"55AADF6DB7DE3F5FAFC708003DE28B68E38E284971F8FC7AAD56DB6DBEF5F8FD",
INIT_30 => X"4AA0004000AA000000000000000000000000000000000000000000000B6F1F8F",
INIT_31 => X"DFEFF7FBFFFEF552E974AA082A820AAA2FFFFFFFFFFFFFFFFFFFFFDFEF552E95",
INIT_32 => X"EAA00A2FFFFFFFF7FBFDFFFFFD568B55002A954AAF7D568A00557FFFFFFFFFFF",
INIT_33 => X"56AB450004001EFFF842AAAA557FFDFEFF7FBFFF55A2D16AB550000175EFFFFB",
INIT_34 => X"7BFDF45AAD568B55AAFBFDFEF55042ABEF002A800AAF7FBFDFEFF7D56AB45AAD",
INIT_35 => X"52AAAAAA007BC0000FFFBE8B55AAD168B55F7FFFFFFF552AA8BEF08040200008",
INIT_36 => X"A2D57FFFFF7D568B45002ABDEAAFFD16AA0008516AB55A2D16ABEFFFFBFDFFF5",
INIT_37 => X"0000000000FFD56AB45A2FFFDFFFAAD16AB4500043DEAAFFAEAAAAA08556AB55",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000800000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(19),        -- Port A data input
DOA(0)   => data_read_a_hi_256(19),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(19),        -- Port B data input
DOB(0)   => data_read_b_hi_256(19),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_20_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000003",
INIT_01 => X"A65FF80000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000048002CC070000000000000000000000002FF86100200000000220002362",
INIT_03 => X"0000000000080F6000977060009B87A03C000000000000000000000000000000",
INIT_04 => X"3F2EFC040388137C3E20C477600142019E6000003CC0000A6601601A000B0000",
INIT_05 => X"102F91D10802ABFB80000021C8010FB0F0F43E1FE867DFC04400390210000220",
INIT_06 => X"90492261000080003400000010008000004203FE400580000000803000200006",
INIT_07 => X"401000004FFDFF28C4300C0010200100004000002AA001F00000000014000000",
INIT_08 => X"0801F5780259FB00000007BEFBC010002008FF7F00000000010018A81000041C",
INIT_09 => X"00000000020000000000000000000ADF00000020000000800000802830011023",
INIT_0A => X"0000000000000200020000000000000000000000000000000200200290000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"08120000B9090A700000200000004000000400000080002000407FED80000000",
INIT_0D => X"000079804000F00000000000C01FF8A7FE003000000004008100000000000000",
INIT_0E => X"0000798201000000100000000135386000401000010000000079801000010000",
INIT_0F => X"0185C300020004000010000000000252C7801000010000000079801000010000",
INIT_10 => X"00000010C1F30F300002010000080000000000CD8A0000400400000010000000",
INIT_11 => X"008040000000000292C0080000000000A5604000000284000818505200080000",
INIT_12 => X"0015E1B00100000000001496008000000000052B000048080000000000FC3600",
INIT_13 => X"80000000000002BA280000800830300000000000B8B400000401881010000000",
INIT_14 => X"00000000020020020001000040283024E6FB8604020080000383383B00000400",
INIT_15 => X"000000000000000000000004010201001003020200000000000127DBFF004000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"038200010089120104D204002000000000000000000000000000000000000000",
INIT_19 => X"B2CB2CB2CB2CB2CB2CB2CB2CB2C30C30C30C30C306982121A1E79E79A0700030",
INIT_1A => X"432190C86432190C86432190C86432190C86432190C86432190CB2CB2CB2CB2C",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000432190C86432190C86432190C86",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA0804020100000000000000000000000",
INIT_22 => X"2E954AA000400000F7FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0004174BAFFF",
INIT_23 => X"FFFFFFFFFFFFFDFEF5D2A974BA082E95400007FFFFFFFFFFFFFFFFFFFFFFEF55",
INIT_24 => X"A2FFFFE10FFFFFFFFFFFFFFFFFFFFFBFDFFF5D2E954BA007FC00BA087FFFFFFF",
INIT_25 => X"FF7FBFFF550800020BAAAD56AAAAF7FFFFFFFFFFFFFFFFF7FBFDFFF552E974BA",
INIT_26 => X"10087FFFFFFFFFFFFFEFF7FBEAB450804001EFAAD57FEAA007FFFFFFFFFFFFFE",
INIT_27 => X"B550004001EFAAAEA8ABA5D7FFFFFFFFFFFDFEFF7D56AB450000021EFA2D57DE",
INIT_28 => X"0000000000000000000000000000000000000000F7FFFFFFFFFFFFDFEFA2D568",
INIT_29 => X"974AA0000104AAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA08000500000000",
INIT_2A => X"FFFFFFFFFBFDFEF5D2E974AA000A07000E3FFFFFFFFFFFFFFFFFFFFFFFEF552A",
INIT_2B => X"71C50BA1C7FFFFFFFFFFFFFFFF7FBFDFFF5D2A954AA082A92428087FFFFFFFFF",
INIT_2C => X"7F5FAFC7492A974AAB6F5F8E10E3FFFFFFFFFFFFFFEFF7FBFFFFF552E974AA00",
INIT_2D => X"1C7FFFFFFFFFBFDFEFE3F5F8F450004050AABEDF6FABAEBFFFFFFFFFFFFDFEFF",
INIT_2E => X"50804021FFB6D57DE28147FFFFFFFFFBFDFC7EBF5E8B550000071EFB6DF7AE92",
INIT_2F => X"EFF7F1F8FD7AAD16AB450000001FFBEA4A8AAA497FFFFFFF7FBF8FC7EBD168B4",
INIT_30 => X"4AA080017410000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFDFEF552E954AA0004000AAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A95",
INIT_32 => X"820AA087FFFFFFFFFFFFFEFF7FBFDFFF5D2A974AA002E95410A2FFFFFFFFFFFF",
INIT_33 => X"FFDFEF5D2E954AA0051554BA557FFFFFFFFFFFDFEFF7FBFFFEF552E974AA082A",
INIT_34 => X"FFFFFFFF7FBFDFFFFFD568B55002A954AAF7D568A00AAFFFFFFFFFFBFDFEFFFF",
INIT_35 => X"000175EFFFFBEAA005D7FFFFEFF7FBFDFFFAAD16AB450804174AAFFFFFFEBAA2",
INIT_36 => X"F7FFEAB45A2D568B550804001EFF7D57DEBA557FFDFEFF7FBFFF55A2D16AB550",
INIT_37 => X"0000000000F7FBFDFEFF7D56AB45AAD56AB450004001EFFF842AAAA087BFDFEF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000000FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(20),        -- Port A data input
DOA(0)   => data_read_a_hi_256(20),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(20),        -- Port B data input
DOB(0)   => data_read_b_hi_256(20),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_21_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"4A302428B824900A128C090A5C1800261500213C005FE812D10420054085A202",
INIT_01 => X"081FFE3440B609703B0427F801A40B8115BC4F655300340288A40D30040E4DD8",
INIT_02 => X"04CA478082CC1740002019824E0203100640303FF8C0B31061096E21A1840814",
INIT_03 => X"8C329E9204020FE002577800405B87047D5042129D8D0248903200013290C800",
INIT_04 => X"3E7FFE02482553FC3C020277E128080A1E6000003CC0000A6601E03A8B0F0008",
INIT_05 => X"F43F8140000203FFC806C8A1C1048FF0F0E07E1F00F7FFC00024010000468310",
INIT_06 => X"08710C10015E083D01A24404786BE0014114C3FE4187A009A663A680100B3096",
INIT_07 => X"200800008FDFFF00290000100211019812E210488228000000900260026C6058",
INIT_08 => X"0EF1F5FA0041FF080AC707FEFBC110008420F7FF388B70A20389346FE8000580",
INIT_09 => X"917FC30010107688862A28C54518DBFF00020004C0A6044901112A0908AA0A30",
INIT_0A => X"006309044081A001B188300E20806520398C6021569249C4B3007127080806FF",
INIT_0B => X"904595123203040D9228D9228D9228D9228D9228D9228D9228D99146C9146C84",
INIT_0C => X"88042090068008003120000806001402504110C48002403601887FEF80022A51",
INIT_0D => X"26C0AC404E43032CA0C205880A7FFAB7FE01409400400C0594A4002200110008",
INIT_0E => X"26C0AC086A170250454004C6012280129B034A080C0B0016A0D20346080C0A80",
INIT_0F => X"0B064092D85938C0112144050224120C500346080C0B0016A0D2034A080C0A80",
INIT_10 => X"40702E058355458967E86A170220D1800093414B0414782E4B5000D81480809A",
INIT_11 => X"081B1545104135443306C35901024F88A88049062A747512B76783C5D040E080",
INIT_12 => X"40160040D86B202049B22198362A8A208279854400A036801480031401900800",
INIT_13 => X"0DD001C002D38334000914028354008301008C0CF1480245108C7640A0604032",
INIT_14 => X"AC0496022300233104662848808E191526205018030060540284FA0C0044022C",
INIT_15 => X"004010040100401004010040102090010008000001C0E010020007DFFFC06E60",
INIT_16 => X"0401004010040100401004010040100401004010040100401004010040100401",
INIT_17 => X"4010040100401004010040100401004010040100401004010040100401004010",
INIT_18 => X"FF7FFDF7FF3E3DFDF7E000000000000000000000000040100401004010040100",
INIT_19 => X"FBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBFFDFDFFFCF3CF3FFFEF9FEE",
INIT_1A => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFEFF7FBFDFEFF7FBFDFEFBEFBEFBEFBE",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0004000100000000000000000000000",
INIT_22 => X"2A954BA0004154BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080402010FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF552A974AA0004174BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"000400000007FFFFFFFFFFFFFFFFFFFFFFEF552E974BA0804000AAF7FFFFFFFF",
INIT_25 => X"FFFFFFDFEF5D2E974BA002E97400007FFFFFFFFFFFFFFFFFFFFFFEF552E954AA",
INIT_26 => X"BA087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974BA082E95400007FFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2E954BA007FC00BA5D7FFFFFFFFFFFFFFFFFFBFDFEF5D2A954AA002E974",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFBFD",
INIT_29 => X"954AA080005000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA00000200000000",
INIT_2A => X"FFFFFFFFFFFFFFF552A974BA0000174AAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0A000AAE3FFFFFFFFFFFFFFFFFFFFFFFEF552A974AA0000104AAF7FFFFFFFFFF",
INIT_2C => X"FFBFDFEF5D2E974AA000A07000007FFFFFFFFFFFFFFFFFFFFDFEF552E954BA08",
INIT_2D => X"1C7FFFFFFFFFFFFFFFFFFBFDFEF5D2A974BA002A95400087FFFFFFFFFFFFFFFF",
INIT_2E => X"F552E974BA0020924BA1C7FFFFFFFFFFFFFFFF7FBFDFFF5D2A954AA082A92428",
INIT_2F => X"FFFFFFFFFEFF7FBFFFFF552E974AA0071C50BA557FFFFFFFFFFFFFFFF7FBFDFF",
INIT_30 => X"4BA000002000000000000000000000000000000000000000000000000E3FFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2A954AA080017410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"000AAF7FFFFFFFFFFFFFFFFFFFFFFFEF552A974BA0000174BAFFFFFFFFFFFFFF",
INIT_33 => X"BFDFEF5D2A954BA082E800AAA2FFFFFFFFFFFFFFFFFFFFFDFEF552E954AA0004",
INIT_34 => X"7FFFFFFFFFFFFFEFF7FBFDFFF5D2A974AA002E95410087FFFFFFFFFFFFFFFF7F",
INIT_35 => X"52E974AA082A820AA557FFFFFFFFFFFFFEFF7FBFFFFF552E954BA002E9741008",
INIT_36 => X"FFFBFDFEFF7FFFFFEF5D2A974BA0000020AA557FFFFFFFFFFFDFEFF7FBFFFEF5",
INIT_37 => X"0000000000AAFFFFFFFFFFBFDFEFFFFFFDFEF5D2E954AA0051554BA5D7FFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(21),        -- Port A data input
DOA(0)   => data_read_a_hi_256(21),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(21),        -- Port B data input
DOB(0)   => data_read_b_hi_256(21),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_22_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"5290F4CDE914905A14A43D33F488243E17122300F55FEB189B343A1140548380",
INIT_01 => X"A94007B259F6A975386262000C344BA9573C6FF57B18A5FB0ABFCD3C2C5F4F0C",
INIT_02 => X"D56B4302AC01005111011BD506AA5205274056900596A539584E2E6DFE4B2418",
INIT_03 => X"6B03F2F6151A2081F24001E8400008F401CB10C6594423C8923AD6B55AD0EB5A",
INIT_04 => X"8001023D37E50880436200808BC8492A0089249600101100008087248B64426E",
INIT_05 => X"A51035B41C0A88046CAEE8C23C08E040011C0020F8882001102D620A06D68301",
INIT_06 => X"B93FF975CF7889D085E997A2144E8FC2060B880081A26DCD4047EFF9EF018980",
INIT_07 => X"283800AA500200E8024AD03546A3262FB5AA5542A882040C7A64CBD64065F028",
INIT_08 => X"141008801018040E48D500400015805060040080A2A0F4A82381B4000A0905A0",
INIT_09 => X"4D0000002126F30C902A29C54539C020E11810098D4067EFF9FF284D483E2AB4",
INIT_0A => X"1400006100003202D040050220103D2A512C6A8C4F0008AA800470370000A000",
INIT_0B => X"013456520CA09281C2A81C2A81C2A81C2A81C2A81C2A81C2A81C9540E1540E00",
INIT_0C => X"A1402A13C0A10A893165281A1C2A7283516344C594A85536B1AD800214202C50",
INIT_0D => X"3C70FC20515808A0100820112300011000287B071105034406950A0285014280",
INIT_0E => X"3C70FC48E11CFC48400184CE0D6783139B0959A41606003C70FA0958AC160480",
INIT_0F => X"0D87E8B3B811B52048B10E0402AE1606D80958AC1606003C70FA0959A4160480",
INIT_10 => X"80F84E0185594581E088E11CFC38414020DD42CF909D7E0A551C02180300C0DD",
INIT_11 => X"441154C258012D86F3044A3133004A99BD8455300654458A1D588C4061403000",
INIT_12 => X"A096A240894626600953379822A984B0025B0DEC0345C9200680027181B44887",
INIT_13 => X"E2404160035482BE521C2C04A90783C18000D610B9D8070B12B1A2A62040202A",
INIT_14 => X"304244A91102C93A2D608D2A258DF8034284200C050070E40C80620C870B02C4",
INIT_15 => X"4411044110441104411044110466C440446CA06951D4EA801000980400646002",
INIT_16 => X"0100441104411044110441104411044110441104411044110441104411044110",
INIT_17 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_18 => X"FE8FF1F7DEBDDF7DF7D05122890000000003FFFFFFFF90040100401004010040",
INIT_19 => X"79E79E79E79E79E79E79E79E79E79E79E79E79E7BFFDFD7DDDF7DF7DF7DFBFDE",
INIT_1A => X"3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE79E79E79E79E",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE000000000000000003F9FCFE7F3F9FCFE7F3F9FCFE7F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0800000000000000000000000000000",
INIT_22 => X"2E974AA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000400010FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E954AA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"0004154BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA000015400FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF552A974AA0800154AAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA",
INIT_26 => X"BAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0004174BAFFFFFFFFFFFFFFFFF",
INIT_27 => X"FEF552E974BA0804000AAA2FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0000174",
INIT_28 => X"0000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040001000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E954AA000402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0417410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080005000FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF552A974BA0000174AAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA00",
INIT_2D => X"E3FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0804154BAF7FFFFFFFFFFFFFFFFF",
INIT_2E => X"F552E954BA000E124BAE3FFFFFFFFFFFFFFFFFFFFFFFEF552A974AA0000104AA",
INIT_2F => X"FFFFFFFFFFFFFFFFDFEF552E954BA080A000AAA2FFFFFFFFFFFFFFFFFFFFFFFE",
INIT_30 => X"4BA080400010000000000000000000000000000000000000000000000007FFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"17410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000400010FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF552A954BA000415400FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954AA0800",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFEF552A974BA0000174BAF7FFFFFFFFFFFFFFFFFFF",
INIT_35 => X"52E954AA0004000AAA2FFFFFFFFFFFFFFFFFFFFFDFEF552E974AA0804174AAF7",
INIT_36 => X"FFFFFFFFFFFFBFDFEF5D2E954BA002A820BAA2FFFFFFFFFFFFFFFFFFFFFDFEF5",
INIT_37 => X"0000000000087FFFFFFFFFFFFFFFF7FBFDFEF5D2A954BA082E800AAAAFFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000000FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(22),        -- Port A data input
DOA(0)   => data_read_a_hi_256(22),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(22),        -- Port B data input
DOB(0)   => data_read_b_hi_256(22),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_23_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"EF20906D902424807BC8241BC81801B97D38AD3C0800103362A6741C80A12A02",
INIT_01 => X"001FFF8409F089003B4422000D80C80106804A7951C5B9D1C828043EA28838F9",
INIT_02 => X"028406A002DC176444683862400003111001303FFC00F240D50146013B300500",
INIT_03 => X"001B243004080FE000177003145F87017D584B10D804034800200200A1008008",
INIT_04 => X"BEFFFC0248005FFC3C18A2FFE12222425E600000BDC0800AEE01E81A100F0A00",
INIT_05 => X"D03F8000000003FF810640A1C0008FF2F0E17E1F02FFFFC80100004044800080",
INIT_06 => X"800264B4854650040123428C204BF40F439647FF4807E189A477EF81DF0AF116",
INIT_07 => X"01000000FFDFFFE800401005C0A0008F86C60840AAAA100C68D1810C9F4A0020",
INIT_08 => X"1BE1F5F80003FF0002021FFEFBC80000000077FF184B03010004002FE1F29002",
INIT_09 => X"907FC308181204800600000000001BFFA800808189A657EF81DD0C00079CC800",
INIT_0A => X"0063090442A18001B188300C48907120AC810033149249C433200180082A06FF",
INIT_0B => X"9A41C1443243050C1010C1010C1010C1010C1010C1010C1010C1008608086084",
INIT_0C => X"000082A00600200080000500C000400800601200000254A000007FEFC1030221",
INIT_0D => X"0A9080400E0BF30C20CA858E087FFABFFE01409780214EE49620001000080004",
INIT_0E => X"0A908044294700701641005218521210150E5789F90A000A90800E5F81F90880",
INIT_0F => X"0E0220036864A7DCA190440301E2105C000E5F81F90A000A90800E5789F90880",
INIT_10 => X"C1400500C6CE5400032429470068924010164302048156305D66F8701681000E",
INIT_11 => X"2E0CCB0500013440600339C800004D8018000857A82920CE8CB220C81400A180",
INIT_12 => X"220344406739000009B0030019960A00026880C0422C52B01700044901488822",
INIT_13 => X"85C811A010428104128996465ADA020180804A040108A2658217C4008060300C",
INIT_14 => X"BE0692020328CA0028042054A92771C50FC070109000C1C819078280A265920E",
INIT_15 => X"020080200802008020080200800800200200000000000008004807DFFF000470",
INIT_16 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_17 => X"0080200802008020080200802008020080200802008020080200802008020080",
INIT_18 => X"0000000000000000000000000000000000000000000000802008020080200802",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000",
INIT_22 => X"2E974BA080002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E974BA000400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000400000FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF5D2E954AA080000010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA",
INIT_26 => X"10FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080402010FFFFFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2A954BA000015400FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA0804000",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E974BA080002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF5D2E954AA000402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA00",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080002010FFFFFFFFFFFFFFFFFFF",
INIT_2E => X"F5D2A954BA080407000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080005000",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF5D2A954BA000417410FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA080402000000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"02000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000010FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF5D2E974AA000402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0000",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000400010FFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"D2A954AA080017410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954AA080002000FF",
INIT_36 => X"FFFFFFFFFFFFFFFFFF552A954BA080015410FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_37 => X"0000000000F7FFFFFFFFFFFFFFFFFFFFFFFFF552A954BA000415400F7FFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000000FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(23),        -- Port A data input
DOA(0)   => data_read_a_hi_256(23),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(23),        -- Port B data input
DOB(0)   => data_read_b_hi_256(23),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_24_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100600007FFF000080108004000800020000840041000080808",
INIT_02 => X"0000068002CC07400000090C080002000000103FF811F150231000520ABE4404",
INIT_03 => X"8428180000080FE000177000001B87003D4000000E8B84010020000000008000",
INIT_04 => X"3E2FFC024800137C3C000077E00000001E6000003CC0000A6601E01A000F0200",
INIT_05 => X"103F8000000003FF80000021C0000FF0F0E03E1F0067FFC00000000000000000",
INIT_06 => X"00132412079001AD00810005E8000001401643FE4007E5501AA00000DC8C3006",
INIT_07 => X"000000000FDFFF62695A5685C094831D966000008002100C2040A178B600C240",
INIT_08 => X"08E1F5F80001FF00000007FEFBC00000000077FF000B00000000002FE0000000",
INIT_09 => X"107FC300000000000600000000001BFFA0000005501AA00000CE200000940000",
INIT_0A => X"00630104408180012188300C00814080008000010012414433000100080806FD",
INIT_0B => X"904181003003000C1000C1000C1000C1000C1000C1000C1000C1000608006084",
INIT_0C => X"00000080060000000000000012002C00000000000000000000007FEF80020201",
INIT_0D => X"440082404E0B332CA2C20188087FFAB7FE000082000000008220000000000000",
INIT_0E => X"4400824903210308074084210002460402009280010D80440084009280010F00",
INIT_0F => X"800A2400401A0C82183248060010280C20009280010D80440084009280010F00",
INIT_10 => X"C0A078160000404A0469032102981380202080026420020D06C002A08481C020",
INIT_11 => X"00164F400860000824059AD01802000208104817B00011306B2D9B0DD5082080",
INIT_12 => X"41021800B35A0300400041202C9E8010C0001040C5836CC01780018601030088",
INIT_13 => X"DB1011E000A140058220004AEFFC8101810021084301880030A8B77400603011",
INIT_14 => X"8C063C0220002201490418082010A57263E010000201033016085A40880030A1",
INIT_15 => X"000000000000000000000000000000000000000000000000000007DFFF0006E0",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"F6E7CC1132CDB444199000000000000000000000000000000000000000000000",
INIT_19 => X"79E79E79E79EFBEFBEFBEFBEFBEF9EF9EF9EF9EFA69861219575D75FF2D0AEEA",
INIT_1A => X"0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1EFBEFBEFBE79E",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE000000000000000000783C1E0F0783C1E0F0783C1E0F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020100000000000000000000000",
INIT_22 => X"2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"080002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_26 => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000400010FFFFFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2E974AA000400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0004000",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040201000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF5D2E974BA080002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFF",
INIT_2E => X"F5D2E974AA000400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF5D2E974AA000400000FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA080402010000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"00010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000010FFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002010FF",
INIT_36 => X"FFFFFFFFFFFFFFFFFF5D2E974AA000002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_37 => X"0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000402010FFFFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(24),        -- Port A data input
DOA(0)   => data_read_a_hi_256(24),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(24),        -- Port B data input
DOB(0)   => data_read_b_hi_256(24),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_25_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100200002000000080100004000000020000800041000080808",
INIT_02 => X"0000068002CC474000000800000002000000103FFCE302008000000880844A04",
INIT_03 => X"00000101C0200FF004177800081B87003D400000080000000020000000008000",
INIT_04 => X"3E2FFE024820137C3C004077F01000001E7249213CC1264A660DF05A000F9000",
INIT_05 => X"103F81C1002203FF80000021C1140FF8F0E03E1F0067FFE04800258280010052",
INIT_06 => X"80480AE20000000100000001C8608001401643FE4007C00000000000CC083006",
INIT_07 => X"280800000FDFFFEA4050140540B00100840000080002A00C2040810000000010",
INIT_08 => X"C8E1F5FA21C9FF80040007FEFBE031018C31F7FFBAEBC0020008086FE0000100",
INIT_09 => X"107FC301800000000600000000001BFFE00301000000000000CC020000140000",
INIT_0A => X"0077330C4889CC292588300C0080400000800001001243443B000100880806FD",
INIT_0B => X"904189003003000C1000C1000C1000C1000C1000C1000C1000C1000608006084",
INIT_0C => X"8B04228026824100000000000000000000000000000004A000007FEF80020201",
INIT_0D => X"400000400E03C30C20C2818C087FFAB7FE01409700C10007962418220C110608",
INIT_0E => X"4000000001010000004000000000400400001200000800400000001200000800",
INIT_0F => X"0008000000000480000040000000200000001200000800400000001200000800",
INIT_10 => X"0000001001000002000001010000100000000000202000000440000000800000",
INIT_11 => X"0000410000000008000008400000000200000806300400000820000020004880",
INIT_12 => X"0000080001080000000040000082000000001000000040800800000000020008",
INIT_13 => X"8100000000000000802000000840000200040000020008000000840000804000",
INIT_14 => X"8C04100200000200000610000000210000000018140000000008000008000000",
INIT_15 => X"04411044110441104411044510629041040D180400000010028047DFFF800C60",
INIT_16 => X"4411044110441104411044110441104411044110441104411044110441104411",
INIT_17 => X"4110441104411044110441104411044110441104411044110441104411044110",
INIT_18 => X"196A8C5A2932EC15DA080800002FFFFFFFFFFFFFFFFFC1104411044110441104",
INIT_19 => X"92492492492410410410410410410492410492412000531215A69A6BFBA2894A",
INIT_1A => X"B158AC562B158AC562B158AC562B1588C46231188C46231188C4924924924924",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000B158AC562B158AC562B158AC562",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000",
INIT_22 => X"2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF5D2E974BA080400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_26 => X"10FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0800000",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400000FFFFFFFFFFFFFFFFFFF",
INIT_2E => X"F5D2E974BA080000010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA080402000000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"02000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400000FF",
INIT_36 => X"FFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_37 => X"0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000000FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(25),        -- Port A data input
DOA(0)   => data_read_a_hi_256(25),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(25),        -- Port B data input
DOB(0)   => data_read_b_hi_256(25),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_26_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"E9264EAB20190CA3BA4997AA9002AE9C001006B0778015CFA17E0811039879C7",
INIT_01 => X"F1FFF9BB1F773C7F9BB07DFFFDD863FC5FFF3FEFFBBF9FFB22FFFBC7B9F30686",
INIT_02 => X"9B3184F8AFDEAF300029E4E300FC78A6258548EFFA71C00172082400003A2161",
INIT_03 => X"0213C3FDFFFC7F74FFBF737A603B87FEBE1A5294F65628A0001B9CE6CC606E73",
INIT_04 => X"7E2EFEBF6FFEB37C3FF3017776FFCDA43E7B6DFD7DEBFD8E6F5F78DF0BFBD644",
INIT_05 => X"902F87C74E8CCFFBB6FF70E1FE61FFBDF0FEBE1FFD67DFFEFFBDA7F7FED50870",
INIT_06 => X"213246200BCC8920360C1831CD7DF60A244B9BFEE00589DDBCEFEDC1DFA08957",
INIT_07 => X"B1D4223B4FFDFF21CC721C85DCE1458E8782484020A2C1FCA3468D77E0000300",
INIT_08 => X"2C05FD7BC471FBD13D980FBEFBEBF30B8D79FF7F451F33CFD60FE8FFFDF54003",
INIT_09 => X"19FFC71FEFED7B251E35768E8ED6BFDF3EB3EBF9DDBCE7FDC1DF8A760F3EACC0",
INIT_0A => X"56F7730ECCDBDF152199F51EDDCDEBCFF589807B7096CD4CF73AC1FC98884FFF",
INIT_0B => X"B867D3683A03A40F78C0D78C0D78C0D78C0D78C0D78C0D78C0D7A606BC606B8C",
INIT_0C => X"DFBFF5EB36DFE51FC3A80D73D840303983EE7F0EA03BDA680137FFFDFFD7E681",
INIT_0D => X"3F0080425E6BFF8DB0DAE19C09FFFFE7FE3EBEA8EB7AFEE5C9AEBD7F5EBFAF5F",
INIT_0E => X"3F00800DEC010280004000F808020290100FA2F60008003F00800FA2F6000800",
INIT_0F => X"00023002007BC0A14E00400003B8000D000FA2F60008003F00800FA2F6000800",
INIT_10 => X"01E0320007204008040DEC010300100000F600020581003F604D0700008000EE",
INIT_11 => X"201F21A2C40039006807C46426040E101A0259DFE82011A311AA042016040080",
INIT_12 => X"80020048F88C84C101C203403E434588007200D047F00090200007E0010009B0",
INIT_13 => X"0109000003E2000416C0804FE04140E80000F808010AB02033AC048A2A00003D",
INIT_14 => X"FFAFD082003B032FB987E04021D481D4000419060201E1A000044300B02033E8",
INIT_15 => X"AFEBFAFEBFAFEBFAFEBFAFEFFBFBFBFBBFCFBB0FFDFEFFEF2DFFFFFBFF802FFD",
INIT_16 => X"FEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBF",
INIT_17 => X"EBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFA",
INIT_18 => X"F491E166CC8553F86EDB5C88646FFFFFFFFFFFFFFFFFEBFAFEBFAFEBFAFEBFAF",
INIT_19 => X"1861861861861861861861861861869A69A61861AFBD54D5F871C71D475B15BC",
INIT_1A => X"0984C26130984C26130984C26130984C26130984C26130984C26186186186186",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE000000000000000000984C26130984C26130984C2613",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000",
INIT_22 => X"2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_26 => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFF",
INIT_2E => X"F5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA080402000000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"02010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_36 => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_37 => X"0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(26),        -- Port A data input
DOA(0)   => data_read_a_hi_256(26),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(26),        -- Port B data input
DOB(0)   => data_read_b_hi_256(26),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_27_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"00080A40000A41248002029000050A088000008242A0004404480002000A1155",
INIT_01 => X"F1FFF1C11F781C129C107DFFFE0860941E81258CA2B71C2220EC1B86E1A00002",
INIT_02 => X"183080988B2EAE00002BE001117C78C6848140CFFA0000800042008000011081",
INIT_03 => X"000003FDF3E47C74F7BCF36A203A47F6B8184210B6160820001318C60C204C63",
INIT_04 => X"7E28FEBF6FEEB3723F71017476DFC524397B6DF572EB6C8E175E70D90F539600",
INIT_05 => X"000F86064C8DDFE3B6FF50D1FC61DE39C8FCB91FF9671FE6B68984B5BCE40834",
INIT_06 => X"0000000800000042020C18300520620A80231BFE200181092CE7ED80DFC00147",
INIT_07 => X"8AC4AA3B0FD1FF201044110560884000840200520002080C23468D0300000282",
INIT_08 => X"2005F0784411E390A4880E3DF7E2FB0B8E717C7F411F3BC6D60B60FFDDE44001",
INIT_09 => X"18FFD757E7ED7A211E81C09818109E1F16B16B71092CE7ED81CF403601228C40",
INIT_0A => X"46FF730E5CCBCD55219AB55F0DEFABC7054880693016DD4C755AC16C1A884FFE",
INIT_0B => X"BC63F1683803C00E3440C3440C3440C3440C3440C3440C3440C3C2061A2061AD",
INIT_0C => X"56BF55CB165EC51D41880FA3F040202883B475062033186801137FF1BAD6F281",
INIT_0D => X"3B0000421E2B0F2E2AE215C808FFFA47FE62BAA86B1AB268E92AB56D5AB6AD5B",
INIT_0E => X"3B000025EC010080004000F808000098100F22520008003B00002F2252000800",
INIT_0F => X"00001042006BC0810600400003B80001002F22520008003B00002F2252000800",
INIT_10 => X"01E032000620000C0405EC010100100000F6000001C1003760410500008000EE",
INIT_11 => X"201D2120840039000817444404040E10020218DE282010A311AA002002040080",
INIT_12 => X"8000000AE888808101C20040BA4241080072001027F00080200007E0000001F0",
INIT_13 => X"0101000003E2000007C0800FE04040280000F8080002F02023AC04080A00003D",
INIT_14 => X"DDAFD082001B03249887E04001D481D4000009020201E1A000040100F02023E8",
INIT_15 => X"ADAB6ADAB6ADAB6ADAB6ADAB6BF1EBDABD8E270BF84A25C6ACB777E3FF800C6D",
INIT_16 => X"DAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6",
INIT_17 => X"AB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6A",
INIT_18 => X"100481CA860402104A471688747FFFFFFFFFFFFFFFFFAB6ADAB6ADAB6ADAB6AD",
INIT_19 => X"0000000000000000000000000008200000000000200072F210000001490E2168",
INIT_1A => X"A05028140A05028140A05028140A050080402010080402010080000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000A05028140A05028140A05028140",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000",
INIT_22 => X"2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_26 => X"10FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFF",
INIT_2E => X"F5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA080402000000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"02000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FF",
INIT_36 => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_37 => X"0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000000FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(27),        -- Port A data input
DOA(0)   => data_read_a_hi_256(27),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(27),        -- Port B data input
DOB(0)   => data_read_b_hi_256(27),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_28_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"02200AA400180030808802A900002A08001280A08A801044104A1000001818C3",
INIT_01 => X"50A00011460214428114180000882214413D0A71592A01D92213D28005210202",
INIT_02 => X"8A54800A210200111100C2110054289220810440030404010844000444410001",
INIT_03 => X"4200040822D4500001E0000028000002000211842010092000018C6295200631",
INIT_04 => X"00400000000B8000000140000005840C00000040002008808100048100100044",
INIT_05 => X"0000222200244400135110000135100000000000000000024CA0A01018000320",
INIT_06 => X"A004912008208040024489121144080400081000200008104000000020000041",
INIT_07 => X"A85800994000000A0200802004204420210001022AA8A0001122448142491008",
INIT_08 => X"0414000201800004080A000000124058200408000880004440004080160C4100",
INIT_09 => X"0080000206CB0821082B694D4D29400002002038104000000020003204000440",
INIT_0A => X"12000843066021001400040024440245400082D022040000400800081022C000",
INIT_0B => X"0002002C004001036050160501605016050160501605016050160280B0280B00",
INIT_0C => X"0012400810080414C0A800310840102182C62302A0194C08001680100E4040A0",
INIT_0D => X"05000002003004208208841401800040000A0000200814004198000400020001",
INIT_0E => X"0500000004000080000000000000028000002052000000050000002052000000",
INIT_0F => X"0000300000004001060000000000000900002052000000050000002052000000",
INIT_10 => X"0000000001200000000004000100000000000000050000002001050000000000",
INIT_11 => X"00002020840000004800040404040000120200A9000000010000002002040000",
INIT_12 => X"0000004800808081000002400040410800000090001000002000000000000910",
INIT_13 => X"0001000000000000144000010000402800000000000A1000010000080A000000",
INIT_14 => X"0080000000110006B08140000040000000000902000000000000410010000100",
INIT_15 => X"0080200802008020080200802101210810C39A66A90A85420413A82000000204",
INIT_16 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_17 => X"8020080200802008020080200802008020080200802008020080200802008020",
INIT_18 => X"110A00246972BD89A40A0C22E100000000000000000000200802008020080200",
INIT_19 => X"82082082082082082082082082082082082082080D35050758C30C31DE21102C",
INIT_1A => X"B0582C160B0582C160B0582C160B0580C06030180C06030180C0820820820820",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000B0582C160B0582C160B0582C160",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000",
INIT_22 => X"2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_26 => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFF",
INIT_2E => X"F5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA080402000000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"02000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_36 => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_37 => X"0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000000FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(28),        -- Port A data input
DOA(0)   => data_read_a_hi_256(28),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(28),        -- Port B data input
DOB(0)   => data_read_b_hi_256(28),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_29_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"79964E4BA01DACAB9E659792D00AAE160002829C7FDFEFCEE97C2815039D70C3",
INIT_01 => X"50BFF9AB0775343F9AB01DF80D5821FC0FFF3FEFD1AF9FF1207FFBC7B9720586",
INIT_02 => X"0D15846807D207200021C4E200D428A2018408600271C000720A0000003A2161",
INIT_03 => X"0002C009EEFC5F10F9B70178681B80FA3E000100765029A00019084345606421",
INIT_04 => X"3E6E023D27DA937C03E3407712E5CDA41E0924DC3D20B98AE905189F0BF8C000",
INIT_05 => X"902003C30E0447F877F930203E213F8CF01E3E00FC67C03A4D9C87525E510160",
INIT_06 => X"0012460003CC002036040811D919F402244293FEE00400CCB46BA4C164A08857",
INIT_07 => X"914800110FFC0001CC320C81D841418E82800100000041FCA1428575A0001108",
INIT_08 => X"0805FD0180E1F8C1111A0782082B50080508FF00048B124D4005C8AFF4154102",
INIT_09 => X"0180000ABFEF89250815568A8AD6ABC02A02A0B0CCB463B4C0748A720B1EA4C0",
INIT_0A => X"021410028450530014014002D445624DB481806A62840800C22800B8900042FF",
INIT_0B => X"0806522C0A40A50268D0068D0068D0068D0068D0068D0068D006A68034680300",
INIT_0C => X"8912E0A83289641F42A80561D040203182AC3D0AA0118A080036FFFC4F4164A0",
INIT_0D => X"050080424069F5A51250648801BFFFE0003E3E00A0685A85410C0816040B0205",
INIT_0E => X"050080080400028000000000000202900000A0F600000005008000A0F6000000",
INIT_0F => X"00023000001040214E0000000000000D0000A0F600000005008000A0F6000000",
INIT_10 => X"000000000120400800080400030000000000000205800008200D070000000000",
INIT_11 => X"000220A2C400000068008424260400001A0241DAC80001010000042016040000",
INIT_12 => X"00020048108484C10000034004414588000000D04010001020000000010009B0",
INIT_13 => X"000900000000000416C00041000140E800000000010AB0001100008A2A000000",
INIT_14 => X"A282C0000033010FB181E00020400000000419060000000000004300B0001100",
INIT_15 => X"02C0B02C0B02C0B02C0B02C4B12B312912831A27FCFE7FFB175B6FF800802594",
INIT_16 => X"2C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B",
INIT_17 => X"C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B0",
INIT_18 => X"EE7FFDF7FE783FFDFFEA0C00602FFFFFFFFFFFFFFFFFC0B02C0B02C0B02C0B02",
INIT_19 => X"BEFBEFBEFBEFBEFBEFBEFBEFBEEBAEBAEBAEBAEBBFFDF9FBEFFFFFFEBBCF9F96",
INIT_1A => X"FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFBEFBEFBEFBEF",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000FBFDFEFF7FBFDFEFF7FBFDFEFF7",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000",
INIT_22 => X"2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_26 => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFF",
INIT_2E => X"F5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA080402000000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"02000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_36 => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_37 => X"0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(29),        -- Port A data input
DOA(0)   => data_read_a_hi_256(29),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(29),        -- Port B data input
DOB(0)   => data_read_b_hi_256(29),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_30_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"FF9FE1F7FFBFFFFDFFD000000000000000000000000000000000000000000000",
INIT_19 => X"79E79E79E79E79E79E79E79E79E79E79E79E79E7AFBD75F5FDF7DF7FF7FFBFFE",
INIT_1A => X"3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE79E79E79E79E",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE000000000000000003F9FCFE7F3F9FCFE7F3F9FCFE7F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000",
INIT_22 => X"2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_26 => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFF",
INIT_2E => X"F5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA080402000000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"02000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_36 => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_37 => X"0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(30),        -- Port A data input
DOA(0)   => data_read_a_hi_256(30),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(30),        -- Port B data input
DOB(0)   => data_read_b_hi_256(30),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_31_5 : RAMB16_S1_S1
generic map (
INIT_00 => X"129000008004A00804A40000400800020000000C005FEA005800200400050100",
INIT_01 => X"A15FF18019700810180065FFFC0040801E80258CA2951C2200EC0906A0804140",
INIT_02 => X"146000808A0C060444692000402850040400408FF80000000010000000004000",
INIT_03 => X"000003F5D1202C70F654716A001A07F438184210960600000012108518004842",
INIT_04 => X"3E28FE3F6FE513703F70007472DA4128187B6DB530C1240A060C70580B439200",
INIT_05 => X"000F84040C088BE3E4AE40C1FD04CE38C0FC381FF8671FE01009048084C40010",
INIT_06 => X"0000000000000008000810200420620E00030BFE000181092CE7ED80DF800106",
INIT_07 => X"000000220FD1FF200040100540800000840200408002000C2244890200000200",
INIT_08 => X"0011F0780011E38004800E3CF3E0B1118C31747F000B33820209206FC9E80000",
INIT_09 => X"187FC301B124F2001600000000001A1F00110101092CE7ED81CF000401228800",
INIT_0A => X"0477330C4889CC012188310E08812982050800A91012494C31004124080886FE",
INIT_0B => X"9861D1403803800C1000C1000C1000C1000C1000C1000C1000C1800608006084",
INIT_0C => X"020400830602410901000D02D0002008012054040022102001017FE190022201",
INIT_0D => X"3A0000401E030B0C20C20188087FFA07FE203A80010002608030102008100408",
INIT_0E => X"3A000005E8010000004000F808000010100F02000008003A00000F0200000800",
INIT_0F => X"00000002006B80800000400003B80000000F02000008003A00000F0200000800",
INIT_10 => X"01E03200060000080405E8010000100000F600000081003740400000008000EE",
INIT_11 => X"201D0100000039000007404000000E1000001846282010A211AA000000000080",
INIT_12 => X"80000000E808000001C200003A0200000072000007E00080000007E0000000A0",
INIT_13 => X"0100000003E200000280800EE04000000000F8080000A02022AC04000000003D",
INIT_14 => X"9C06D082000A03200806A040019481D4000000000201E1A000040000A02022E8",
INIT_15 => X"0401004010040100401004010060C040040C200950402090128057C3FF800C60",
INIT_16 => X"4010040100401004010040100401004010040100401004010040100401004010",
INIT_17 => X"0100401004010040100401004010040100401004010040100401004010040100",
INIT_18 => X"000000000000000000001000802FFFFFFFFFFFFFFFFF81004010040100401004",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000",
INIT_22 => X"2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_26 => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFF",
INIT_2E => X"F5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA080402000000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"02000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_36 => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_37 => X"0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(31),        -- Port A data input
DOA(0)   => data_read_a_hi_256(31),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(31),        -- Port B data input
DOB(0)   => data_read_b_hi_256(31),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_0_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"ED39BA795990D275FB4A6E96ACC4731DEA4598B0AFB54867F6EE4618C3749803",
INIT_01 => X"58A0047C8607844847CA180001E4A2404042106208408208C2002069161734B3",
INIT_02 => X"8B1EC9562121F8051500147A0E5629A302CF28400615F5787B09FBF999BB1EFD",
INIT_03 => X"404EFC0A2AD6100F01A88E851CE47803C280110521898F6996088862C7B22221",
INIT_04 => X"C0D001C0100AEC83C008E7880D01A64661800002C21A52C590D2012194804844",
INIT_05 => X"650002C3F08754001B51981E007910070F01C1E003980015A204C22F32328BAF",
INIT_06 => X"BCDA4677CAEE7CF5BB870E1DDB9889C5FBFC440129A0604442180238203F70C1",
INIT_07 => X"7AAE0088B02000C2EC3A0E829836E0AF3325372E2AA8FDF3C18306758B24197A",
INIT_08 => X"D7E40002F7AE005FFB4730010411400A61080000F7F4C464B58294901606D5A5",
INIT_09 => X"C4801C40469B0CA9881A28C141118000C5A85A60444210123820B43B40804274",
INIT_0A => X"400800219010107ED453C041B13216656074EA560F0092A24856B05312226900",
INIT_0B => X"27122C3E04E03383E2781EA781E2781EA781E2781EA781E2781C33C0613C0E29",
INIT_0C => X"74EB1F50D0758A9650E520610A6A57A5529E2B439499CF96B086000000B09870",
INIT_0D => X"04F07E024108F4E28638EC57250004480155C1375A97A9121F8BA749D3A4E9D2",
INIT_0E => X"04F07E42177EFDF8570184071575970F8FC07D5BFF078004F07E007D5BFF0780",
INIT_0F => X"8F85ECB1FE047F5FB7B30E0700461E5AF8007D5BFF078004F07E007D5BFF0780",
INIT_10 => X"C0184D07C1DF15C7E3E2177EFDF8C3C03009C3CDD47C7F403FB3FDF89701C011",
INIT_11 => X"4F80FE659C6104C6D7103F9D1D064189B5924418D65FE45DEE55BBEDE34CF900",
INIT_12 => X"6395F64207F3A3A1483136B881FCCB38C2098DACA01FFF603F80001F80FDC81F",
INIT_13 => X"FED151E01015C3BB507D3F811FBEC32B81840714F8D91F4FC513F37C8AE07002",
INIT_14 => X"61692F293185D8D724E15D3FCC6B7C236FE0691A9500125C1F83F8CC1F4FC507",
INIT_15 => X"E93A4E93A4E93A4E93A4E93A4F942F90E9628540052090650525A0000066A00B",
INIT_16 => X"93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4",
INIT_17 => X"3A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E",
INIT_18 => X"09B56C74DAB15D1CF13501AA495000000000000000003A4E93A4E93A4E93A4E9",
INIT_19 => X"2082082082082082082082082082082082082082082084E41DC71C7155F3898E",
INIT_1A => X"3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F8208208208208",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE5294A5294A52800003E1F0F87C3E1F0F87C3E1F0F87C",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000030FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"A975EFFFAABDE00FFAEBDFFF5D2EAAAAAF7AEBDEBA0000000000000000000000",
INIT_22 => X"8000155087FC0155F7D168B55007BFDF45085168ABA002E82145085155545F7A",
INIT_23 => X"FFFD7545AA8028A00A2802AABAFF8028BEF5D7FFFE10005542145557FD5545FF",
INIT_24 => X"F7AEAAAAAA2FFFDF4500043FE105D2E954BAF7FFC0010080017555555568AAAF",
INIT_25 => X"A5D5168A00A2D142155005142010FFAE820AAFF842AABAA2AE95545FFD168ABA",
INIT_26 => X"FF5D2A821550000000BA007FD55FF5D7FC0145007FD7400550415410002E974B",
INIT_27 => X"F455D5142000082E82145FFD17DFEFFFD168BFFF780000BA007FE8AAAFF803FF",
INIT_28 => X"0000000000000000000000000000000000000000AAFBEAA00007BFDFFF082EBD",
INIT_29 => X"AABEA495FC716F002A975FFE3AA95E00EBAEBDFD75D2AA8A80EA8E2FE3F00000",
INIT_2A => X"56A16D557BC257D415E0216FA3F1E8FC0145B68B551475FAF6D1C556F0AA1C24",
INIT_2B => X"7FD24AFE3D02DAAAE12BD5545A2803AA0000542A0070071C50BAFEF1FAE0016D",
INIT_2C => X"A8B50F55A2F150005A3A438BD04AFAB8F550A8010E004924874825D7FEAA8548",
INIT_2D => X"A2A5504001C74BA42A1571E8028E3DB7816D0120155EA568E870BAEB8A05A2AE",
INIT_2E => X"2FFAFD2A82485FD2415A105C21451ED42A002545E055FFBE81D0BE8EA8A3AA05",
INIT_2F => X"100AA1D0F6F480B6A555A2A57A002A3D5FDB6A5C7E3DFFFE90B45B47ABA497A8",
INIT_30 => X"A0AFE80A8B0A000000000000000000000000000000000000000000000B55EAAA",
INIT_31 => X"ABEF5D557FEBA55022A3F70C6B405F4D2AE975EFAAAAB5E1AF3AABFF45592E88",
INIT_32 => X"411A8DED57CE1055555E5F58EFFC01FE2CACB65F520EBE9EF67D7BEA1FD5D556",
INIT_33 => X"A4AD0079C75D6070CC5CBB0280C029ABAA3EBC114728007521170821CE0FDE69",
INIT_34 => X"2A95E02A2AAB5EB0F280800EFAEE9F5D18F3142341D5DEEBEF55080034E0A592",
INIT_35 => X"B69C30E02116220415A9540AA854140A0A2047F353AAF6C77F7F20D968BF5781",
INIT_36 => X"ABEBE1B4D792A4AD1183454180DD3FDCAAAB7C91565455C141E41887D58AC448",
INIT_37 => X"F0000001FF01EABC4B8014174FF7DA80F52FEDE6BE93172D7D625B556EEAB157",
INIT_38 => X"FF0000001FF0000001FF0000001FF0000001FF0000001FF0000001FF0000001F",
INIT_39 => X"0000000000000000000000000001FF0000001FF0000001FF0000001FF0000001",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000100000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(0),               -- Port A write enable input
DIA(0)   => data_write_a(0),        -- Port A data input
DOA(0)   => data_read_a_lo_512(0),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(0),               -- Port B write enable input
DIB(0)   => data_write_b(0),        -- Port B data input
DOB(0)   => data_read_b_lo_512(0),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_1_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"212C001411984004084D000508C53810A03D1450E839B003342114428A000803",
INIT_01 => X"08000011400A100A81160000008C005400400002000000000000028001340000",
INIT_02 => X"C084484000002014400205851002007030450E0000A606C8C44CB4C6666C00E0",
INIT_03 => X"33DF380008164004000002000C80400002031943000101091608463061120118",
INIT_04 => X"4140008000000002000064000400004201000000000210458010070080100433",
INIT_05 => X"8500101040200000010009100000000508000100000000002010600100208D04",
INIT_06 => X"B5EDFDE24618AD433060C182BA860044204C000008A004100008000820280020",
INIT_07 => X"581E02100020000A81244890AA20263030517F122AA801F0983060AC564BF808",
INIT_08 => X"00820800C7A00045B103200000140A02234808000584000004808400020011A4",
INIT_09 => X"0000104000020082800808111008400000200204100000100820800144000414",
INIT_0A => X"12804062945211441E13C051156E800008402802060C94000040901102800000",
INIT_0B => X"24002006406401918C191AC191A4191A4191AC191AC191A4191A00C8560C8D29",
INIT_0C => X"0408010040050880383820080F105F05800302E0E08842422006000000041032",
INIT_0D => X"05000600000090C1841808172580000000008008020084082080204010200810",
INIT_0E => X"0500066210000178470184000000878402C000001E07800500062000001E0780",
INIT_0F => X"00003C404600000011A30E0700000009382000001E07800500062000001E0780",
INIT_10 => X"C0180000012010C20022100000F0C3C03000000055200340000000F88701C000",
INIT_11 => X"05800241186100004D100098190240001290002050068000001010486140F900",
INIT_12 => X"0000164A001303204800026880048230C2000094A0000F601F8000000001C908",
INIT_13 => X"12D051E01000000154200580003C030381840000004B08014401025480E07000",
INIT_14 => X"40082300218450C2800010094000482142E0601895001000000041C408014400",
INIT_15 => X"0802008020080200802008020080008208600500A82A15008000000000468000",
INIT_16 => X"8020080200802008020080200802008020080200802008020080200802008020",
INIT_17 => X"0200802008020080200802008020080200802008020080200802008020080200",
INIT_18 => X"BABEFC54A0810C7452B5420A1000000000000000000002008020080200802008",
INIT_19 => X"AAAAAAAAAAAAAAAAAAAAAAAAAAA28A28A28A28A2A8218D2C0C92492581328A46",
INIT_1A => X"2E974BA5D2E974BA5D2E974BA5D2E975BADD6EB75BADD6EB75BAAAAAAAAAAAAA",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFF6318C6318C63000002E974BA5D2E974BA5D2E974BA5D",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"00000000000000000000000C0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"002155557FFFFFF007FC21EFA2FFD74AAAAD5555550000000000000000000000",
INIT_22 => X"7FD75FFAAAA800AAF7AA974BAFFFBE8B45F7AEBDF455D2EAABEFF7FFE8BFF5D0",
INIT_23 => X"0557DF45AAD1400BAA2AE801550051555EFF7AA95400552AAAABAFFD1574105D",
INIT_24 => X"FFFBEAB55F780020AAAA80020AA082EAAB5500517DF555D2EAAA105500001550",
INIT_25 => X"AF7AE820AA0851574BAA2D1574AA5D7BFDEBAFFD540155557FD5400F78028BFF",
INIT_26 => X"FFFFD56AAAAFFFFD7555AAD168B45AAAEAAABAFF842ABEF5D517DF55552A974A",
INIT_27 => X"4BAF7AE80010082A97410557FEABFFAAFBE8BEFAAD1575EF557FFFE10557FFFF",
INIT_28 => X"00000000000000000000000000000000000000005D7FFDF4500043FE105D2E95",
INIT_29 => X"A8BC2EBDFEAF7F1F840017D4975D2FEF147FC51C7A2FBD5490BFD1C056A00000",
INIT_2A => X"AA8AAAE3D145410F7F1D55D71C002DABAEBAA974BAF7FFEFB45FFAABDF55492A",
INIT_2B => X"0E2AE85028B40155145F7AF6DBED5450AA1C2080BEF495FC71D54124924385FA",
INIT_2C => X"571D2E28E38E0216FA2D1E8E80140F45082B4002D082082AB8B6DBEDB7DF7F54",
INIT_2D => X"A97F7AF6D417E92482BF84020BA495557E3FF78E021FF1471FDEAAFFD56F16D5",
INIT_2E => X"7002FD74951D71EDFFABFD16FAAAE92BD5545A2DA3FB7DAAD4AAAAF487BC70BF",
INIT_2F => X"550A8010E00492487482FFFE82A85EBAE2FFC55554ADBD7A2FFC7BEFF6FFD7FC",
INIT_30 => X"400FBF9424F7000000000000000000000000000000000000000000000547AB8F",
INIT_31 => X"DF55F7AABFF55082CA8B4DF6C1E8F5E5400021EF005162BEF047FD5545AAFBF7",
INIT_32 => X"404547184164AA5D2EBEEB0A2D555410D3555714F8338AAAA1D0AE974AAF7FFF",
INIT_33 => X"AEABFFDF79DCBF755962010BDCBBC21455D7FEABEF75550ACBB7582225FF5843",
INIT_34 => X"D57D412F7D55F5E50C7F401BAAE8403CF5A3FFEAAEB083BC1000FF8409000512",
INIT_35 => X"2AA9FEAFDF7F431A9F7FFE81FF013A8001AFF801F8BA0C57740BDAA0688E5405",
INIT_36 => X"A2FBF7FED2C7F955445079E280A00C56145EF5D16BABAA3EBC3157ABD5FFE55F",
INIT_37 => X"0000000000596EBEF55080034E0A592A4AD00FB863550229BCABEB7DA403FFFD",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000100000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(0),               -- Port A write enable input
DIA(0)   => data_write_a(1),        -- Port A data input
DOA(0)   => data_read_a_lo_512(1),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(0),               -- Port B write enable input
DIB(0)   => data_write_b(1),        -- Port B data input
DOB(0)   => data_read_b_lo_512(1),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_2_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10E006600180111284380310006289800480032283E000A34301002001A0817",
INIT_01 => X"A14AC00A1079284D04A044A54E504368404000720885800802000006ECD10200",
INIT_02 => X"92250052A0348C310102048800A8507000040C8550200000480E0080001321E0",
INIT_03 => X"020204E4593C0824400C2220483042809292430400440180000890A4C9400242",
INIT_04 => X"486854B141002252142241502460480031B94420634850069A42241009610A04",
INIT_05 => X"800504244080892105AA6010A44882144840910A21220A8C820025E4A0000B00",
INIT_06 => X"A000442802280000340810209C444804206000AC800088096A0EA8C022208012",
INIT_07 => X"309820A848E0AA09826489A5CC49002001020112028201F8A20488260000108A",
INIT_08 => X"2400582881E0C1419D12041455509341A539C42A0D8208099002801700D10103",
INIT_09 => X"110D525861263100009200151409130A3C80C8C8096A06B8C12088400A9C2080",
INIT_0A => X"0451394CD0391A441583C04B580040089581001342801044877200D002A00DE0",
INIT_0B => X"144423040240450114901149013C9011C9013C9011C90134901144801A4808A5",
INIT_0C => X"D8A5345206D2C10082080A90C00000188150100C202A4640000E2B4081969420",
INIT_0D => X"050080400A0391A51240C480000AA902AA009028C83220008086952B4285A54A",
INIT_0E => X"05008021C00000000040000000020288000500000008000500802A0000000800",
INIT_0F => X"0002300000428000000040000000000D002A0000000800050080250000000800",
INIT_10 => X"0000000001204004000508000000100000000002054000130000000000800000",
INIT_11 => X"000C00000000000068144000000000001A000106200010021002000000000080",
INIT_12 => X"0002004A880000000000034098000000000000D024A000000000000001000900",
INIT_13 => X"00000000000000041400000A8000000000000000010A00000284000000000000",
INIT_14 => X"012100000002000280000000011080C000000000000000000000430000000260",
INIT_15 => X"A769DA769DA769DA368DA36CDA3A9A13A14801404134DA84A024024155000399",
INIT_16 => X"168DA769DA769DA769DA368DA368DA368DA769DA769DA769DA368DA368DA368D",
INIT_17 => X"68DA168DA169DA569DA569DA568DA168DA168DA169DA569DA569DA568DA168DA",
INIT_18 => X"138D70C030B51C50C7D000A2012F81F81F83F03F03F069DA569DA569DA568DA1",
INIT_19 => X"1041041041041041041041041041041041041041024860208165965975960040",
INIT_1A => X"25128944A25128944A25128944A25128944A25128944A2512894104104104104",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFF8421084210840703F25128944A25128944A25128944A",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"00000000000000000000000F0FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"415555087BFFF55A2AA800BAFFAE9540008002AA000000000000000000000000",
INIT_22 => X"7FE8B555551421455D0002145552EBFEBA007FC21EFA2FFD75EFAA8415410AA8",
INIT_23 => X"FFFE8B45552EBDF45FFAEAABFFF7FFE8B55F784155EFA2AEBDEAAA2FBEAABA5D",
INIT_24 => X"5D2AAAAAA5D2E820BAA2FBEAB5555557DF55A2AEBDF555D2E954BAA2AA974BAF",
INIT_25 => X"A5D04021EF557FC21FFAA8428BFFAAAA954AAAAAAAAAAAFFD1574105D7FFFF55",
INIT_26 => X"EFF7800215500557DF55AA80001FFAA80001550055575EFFF84021555D043DEA",
INIT_27 => X"B5500517DF555D042AA10A284154005D0015410085568A00FF80175FFA2D17DF",
INIT_28 => X"00000000000000000000000000000000000000005D00020AAAA80020AA082EAA",
INIT_29 => X"D55D2BE800042AFE8E1557D0075D2F45BEAA800AAFFAA9543A080038A2A00000",
INIT_2A => X"0BDEAAA2FBF8AAA557BE8B6D5D5FFABEF49040017D5D20B8EAA007FC51C7A2FB",
INIT_2B => X"0E174BFA02A974BAF7F5EFB455D2ABDF55492AA8BC7EBDFEAFEFFD00105FFBC2",
INIT_2C => X"3D155E105571D55D71C002DABA5524820BAB6FFEFB6D555578F7DB6A0BDF7D48",
INIT_2D => X"092A071555D5E3AE821D00001FF0871C016DBED1FDE90E3A497492B6AAADAAAE",
INIT_2E => X"0E3DA3DFD5E3DFFFBD5A38A021551C5F7AF6DBE8F401D7B6A0001470155C51D0",
INIT_2F => X"82B4002D082082AB8B6D1C5B7DF7FF78E075C5BE8555400550A38428007FED00",
INIT_30 => X"4AA00042AAA2000000000000000000000000000000000000000000000410F450",
INIT_31 => X"AAAA007FD5555AAFBD7545FBB8020A3F7AE975EF005560B55F7AA800AAF7AA95",
INIT_32 => X"E8F5EFF84165EFF7802BAB0A2FFEAABA557BEABEF057D68F5F5A00021EF55042",
INIT_33 => X"52ABFFFF841FFE75CA882108202E974AAF7D57DF55D7AABFF5428ACA8F45A6C1",
INIT_34 => X"84174A8FFAEBFEB0A2D55541051555694F002CA8AA80800020AAF7FBFFFEF045",
INIT_35 => X"7AAA155F595542455512A975455D3AA8A005500151FF0C57401E5F3D1E00A1A8",
INIT_36 => X"5D2A8A0B882FFFFE10AAAAAB755A66B6AF56A2AA801455D7FE8BFFF680800FFF",
INIT_37 => X"00000000000C3BC1000FF8409000512AEABFF5D79FCAF774AE005BE789555400",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000200000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(0),               -- Port A write enable input
DIA(0)   => data_write_a(2),        -- Port A data input
DOA(0)   => data_read_a_lo_512(2),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(0),               -- Port B write enable input
DIB(0)   => data_write_b(2),        -- Port B data input
DOB(0)   => data_read_b_lo_512(2),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_3_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"210C44A20020248B08431120001604B8156023104C4077133420400A02380202",
INIT_01 => X"015A2A424080216D3C2462C99E104B49404040028804A0080A000C16A0D90A0C",
INIT_02 => X"C0A4065000F0A95011000D1501005270B4045AB330860281CC08008222170060",
INIT_03 => X"AD22014098340394A4021320080841C40B411B4298042180002846B06900811A",
INIT_04 => X"244B32A86D20014A0D20403194904900071A24110F0BF400F85F92420E0C946E",
INIT_05 => X"80331030442898B4812840D0500008C528280B063006A64CA30004E5A4E40304",
INIT_06 => X"90016CA00E380042302040A0BC47160424428198C0038C89904E640023600816",
INIT_07 => X"1288020843A66620816049908AA0061011CA0142000009F0A810292E7402F088",
INIT_08 => X"20003C9984A0AC411102014D34EC2200214D5099048823019603A01A49410103",
INIT_09 => X"001CD74C4826220010A8891451284B661CA24A4C899046740121824004100080",
INIT_0A => X"44C9516DC0135C45159BE45F112B48804DC10203021290400772C0F402820D4C",
INIT_0B => X"B400624402404501A49018490184901A4901A4901849018C901A648056480C2D",
INIT_0C => X"D7A9B54000D7C10820680D08C420180381211081A022160000266723E1909021",
INIT_0D => X"400080200E199A4A2CA2994C0399981666409800CA52E4890806BD6B56BDAB52",
INIT_0E => X"40008008E00000000000000000024008000C8000000000400080028000000000",
INIT_0F => X"000A000000588000000000000000200400088000000000400080078000000000",
INIT_10 => X"0000001000004004000D800000000000000000022040000B4000000000000000",
INIT_11 => X"001A0000000000082006C000000000020804087220000122000A000000000000",
INIT_12 => X"00020800B8000000000041002E00000000001040466000000000000001020080",
INIT_13 => X"00000000000000048200004A600000000000000003008000320C000000000000",
INIT_14 => X"432900000222200871028000210400C4000000000000000000080200800030E0",
INIT_15 => X"AF6A5AF6A5AF6A5AF6A5AF6E5AFADA91AB68000101B4D20C08EC461733804A19",
INIT_16 => X"B6B5AF6A5AF6A5AF6A5AF6A5AF6A5AF6A5AB6B5AB6B5AB6B5AB6B5AB6B5AB6B5",
INIT_17 => X"6BDAB6B5A96ADAF6A5AD6ADAF6A5AD6ADAF6A5AD6BDAB6B5A96BDAB6B5A96BDA",
INIT_18 => X"C78C706428A14C586290008A044D54AAB556AA9556AAEBDAB6B5A96BDAB6B5A9",
INIT_19 => X"92492492492492492492492492410410410410412821600001249249015303C0",
INIT_1A => X"351A8D46A351A8D46A351A8D46A351A9D4EA753A9D4EA753A9D4924924924924",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000001543B351A8D46A351A8D46A351A8D46A",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"43DF55FFAA955EFA2D168B55557BEAA000055420000000000000000000000000",
INIT_22 => X"7BE8BFFA2D155410AA8415555087BFFF55A2AA800BAFFAE9554508002AA00AA8",
INIT_23 => X"52ABFEBA007FC21EF007FD75FFAA841541008002AB55AAAA955EF005568A0008",
INIT_24 => X"005168B455D042AB45F7FFD741000042AA10AAAABFF5508003FF555D00021455",
INIT_25 => X"0A2D1575FFF7AA975555D2E80145F78415545082EBDEAAA2FBEAABA5D7FC0155",
INIT_26 => X"55552A954BAFFFFE8B55552EBDE00F7AEAABFFF7FBEAB55F7AABDEBA5D7FC201",
INIT_27 => X"F55A2AEBDF555D2E954BA002EAAABA002A821EF5555554AA087BC01FFFFAAAAB",
INIT_28 => X"0000000000000000000000000000000000000000082E820BAA2FBEAB5555557D",
INIT_29 => X"95578080038A2AA28E3AF55E3A0BA5D7AADB6FB7D5D7FEAA3808554203A00000",
INIT_2A => X"0925D7085F6AA10087FEABD7AAD57AEBAB68E1557D1475FAF45BEAA800AAFFAA",
INIT_2B => X"04AAFFA41040017D5D20B8EAA007FC51C7A2FBD55D7BE80004AA1E8E2AB55B6A",
INIT_2C => X"2FBE80AA557BE8B6D5D5FFABEF49002FB55FFF5D0438140E2FA38B6AEBFF6D1D",
INIT_2D => X"AB8ABAE925D21C7010EADB525D7FFAE975C75D0A901FFFF801557D1C20B8EAAA",
INIT_2E => X"20875C21D5EB8AA8FFF012A954BAFFF5EFB455D20BDE00EBAAA8BC7EBDFEAFEF",
INIT_2F => X"BAB6FFEFB6D555578F7DB6A0BDF7DEB8E125FF002EADA921420871D74971D248",
INIT_30 => X"ABA0051400A20000000000000000000000000000000000000000000001C24820",
INIT_31 => X"8B55F7AA800BAF7AA955EF00042AAA2A2AEAAB55A28408145AAFFFFFFF5D7FEA",
INIT_32 => X"020A35D2ABEF55F7800015F087FEAA00007FEAB55FAD568AA2AFAE975EF55516",
INIT_33 => X"ABFEAAF7AE9DFF759A82AEF70800021EF55042AAAA007FD55558A7BD7145FBB8",
INIT_34 => X"84175EF55002AAB0A2FFEAABA557BEA3EF057968F575D003FF55F7D5420BA5D2",
INIT_35 => X"A8429F45A7D5EAF5FFBAEAAA10554155400AAFFD5145FBAC9755F05040255FFD",
INIT_36 => X"550415557085540000005156155FE90A8F5C082E974AAF7D57DF45552A3FF10A",
INIT_37 => X"00000000005500020AAF7FBFFFEF04552ABFFFF843FFE77C80825BC052ABFE10",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000100000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(0),               -- Port A write enable input
DIA(0)   => data_write_a(3),        -- Port A data input
DOA(0)   => data_read_a_lo_512(3),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(0),               -- Port B write enable input
DIB(0)   => data_write_b(3),        -- Port B data input
DOB(0)   => data_read_b_lo_512(3),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_4_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A108400020612C80284210081034849800A000303100048B3432C82904204002",
INIT_01 => X"21066802000820491C00650E1E004360403008418984014902030906A8D10200",
INIT_02 => X"120404E00E4C0600000206100008402005040C00F104008040080080001310E0",
INIT_03 => X"DCA201514D1C0D706C5CF010083A0708BA0841945004010000080084C1000002",
INIT_04 => X"5C4CF21C48B133483C80417570D000083A62488074C1350EA60D785C0A6B0619",
INIT_05 => X"000F0400028083B381A60001E5546EB5C0E2B81E4166DE000139200004E50940",
INIT_06 => X"80004408020800023000102098000204A040038600018019004B800123208806",
INIT_07 => X"120C20204665E1008024188488800000001A01520000A1F08044892400001088",
INIT_08 => X"0801007AC0A1EB413102063CF3E0B3028D29F407059B0B000205A801C2200102",
INIT_09 => X"106052400922D00406BE1002C6150F41200280001900439001FD8A0004142000",
INIT_0A => X"047F2201D899BA503583504B58AB80804540001202805544314041B48A888EC5",
INIT_0B => X"1441E3443043410C5010C3010C1010C3010C1010C1010C3010C14086980861A5",
INIT_0C => X"020000A02600000805400502C0A0004A00625015000A12000026E1E180011220",
INIT_0D => X"400000000E43930C20C20188120782861E4004A800600401A030001008080400",
INIT_0E => X"40000021A8800000000000000000400800170024000000400000310024000000",
INIT_0F => X"0008000000AA80200800000000002000003400240000004000003B0024000000",
INIT_10 => X"00000010000000040004A080000000000000000020400006C008020000000000",
INIT_11 => X"002C008200000008001B4020200000020000090760000200110A040010000000",
INIT_12 => X"00000803E004040000004000E801040000001000086000000000000000020040",
INIT_13 => X"0000000000000000810000164001008000000000020040002240008020000000",
INIT_14 => X"04001040026026004000000002940040000410000000000000080000400000B8",
INIT_15 => X"040080201004008060000001806AC000004890015124D880100886D8F0014420",
INIT_16 => X"4010000180600000018020100400802010000080601000008020000401802000",
INIT_17 => X"0100000004008020180600000000000180600802010000000401802018020000",
INIT_18 => X"3807E05000140634504048820064B261934D964C326980004010000080600806",
INIT_19 => X"AAAAAAAAAAAAAAAAAAAAAAAAAAA28A28A28A28A2934C8D0CCD145144C0A28A06",
INIT_1A => X"068341A0D068341A0D068341A0D068351A8D46A351A8D46A351AAAAAAAAAAAAA",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000000173F068341A0D068341A0D068341A0D",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"57FE10FFFBEAA10007FD7410FFAA97555082A800AA0000000000000000000000",
INIT_22 => X"7FEAA00007BE8AAAAA843DF55FFAA955EFA2D168B55557BEAB45005542000005",
INIT_23 => X"87BFFF55A2AA800BAFFAE9555508002AA000055574105D2A800AA00043FEBA5D",
INIT_24 => X"A2D17DE1000517FE10AAAAA8AAA002E97545557BC00AAA2FFEAAAAAA84155550",
INIT_25 => X"0A2D157400AAAE974AAAAAA974BA08002AB55A2AA955EF005568A00087BE8BFF",
INIT_26 => X"BA080002145552ABFEAA007FC21EF007FD75FFAA8417410A2D140000F7FBC201",
INIT_27 => X"A10AAAABFF5508003FF55F7D568A00552EA8BEFA2AABDEAA087BEAAAAA2FBD54",
INIT_28 => X"000000000000000000000000000000000000000055042AB45F7FFD741000042A",
INIT_29 => X"EAB7808554203A145178E00FFFBE8A101475D5400F7A49057D0824850B800000",
INIT_2A => X"E8008200043FE925571EFA380871C7028A28E3AF55F7A0925D7AADB6FB7D5D7F",
INIT_2B => X"F5FDA38BE8E1557D1475FAF45BEAA800AAFFAA9557D080038AAA145157428492",
INIT_2C => X"85F6AA10087FEABD7AAD57AEBA08517DE00AAAEA8A9200249056D4175C5092AA",
INIT_2D => X"FEDB42028EBFBC2028BED152438AAA092492AAA4954281C0E2FB55B6A0925D70",
INIT_2E => X"A0875EDA80BEF1C743840040017D5520B8EAA007FC51C7007BD55D7BE80004AA",
INIT_2F => X"55FFF5D0438140E2FA38B6AEBFF6DBE84AAEBAF7DF6AA00412EAABFFAA803DEB",
INIT_30 => X"1EF0800154B200000000000000000000000000000000000000000000041002FB",
INIT_31 => X"0145AAFFFFFEF5D7FEABFF0051400A25D5568A00FFFFEAA105D5155410FF8402",
INIT_32 => X"2AAA25555410BA082E8201000043FE005D517DEBA0851574B2AAAEAAB55F7840",
INIT_33 => X"4001FF005575408AA557FEB2FFAE975EF555168B55F7AA800BAF7AA955EF0004",
INIT_34 => X"2ABFF55F7800015F087FEAA00007FEAB55FAD568AA200557DE00AAAAAAA00080",
INIT_35 => X"87BD6145FAAC000A2A6FBC00BAAAFBC00BAF7D1550AAAA8002010F2AC154B25F",
INIT_36 => X"082EA8BFFAA843FEBA08517DE00F3F9574B30800021EF55042AAAA007FD55550",
INIT_37 => X"000000000008003FF55F7D5420BA5D2ABFEAAF7AEBDFF779A82AA43F7FBE8A00",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000200000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(0),               -- Port A write enable input
DIA(0)   => data_write_a(4),        -- Port A data input
DOA(0)   => data_read_a_lo_512(4),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(0),               -- Port B write enable input
DIB(0)   => data_write_b(4),        -- Port B data input
DOB(0)   => data_read_b_lo_512(4),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_5_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50DF4A0791B3FCB694379283C81FD996A091832102004A337A20E07C0C1E006",
INIT_01 => X"294014468000A04D5C6A60000C34C24841280A00084000C8C212892EEAD53235",
INIT_02 => X"50AE41540CA1D9100002171C1F0A5171134E2A200D8633F8CD09DBFBBB970E7C",
INIT_03 => X"214E3C521D16021B64430CC51C45B8154689094241898749920842946B90010A",
INIT_04 => X"A2F20F7D7A314CB5C208E28A1BF0224A448920028A185340D0C20B2690000C22",
INIT_05 => X"7520B430B20B984809A8886E230C6106371146E1829941C58310402C600381CF",
INIT_06 => X"9CC96CD7C63A7495B9A356ACBC4601C57FD44F8549A46490261C4B39203F7080",
INIT_07 => X"12A88800B029E0C0A12C4B92AA36A2111167357C220095F3C8952A2E5D26F078",
INIT_08 => X"F3F00503B4AE105B534711820C0C0A1043080300F7E0E728B1829C2FEA0A95A1",
INIT_09 => X"C5184F084136848C9298A8560688F480C58858449026145B3830F40944906234",
INIT_0A => X"50EB4124D2B3902BF5C9700C1199DCA84DF46A974F92C7E28F1630D38088A438",
INIT_0B => X"B3144E5636E3178C86B8CC6B8CA6B8CE6B8C86B8CE6B8CA6B8CC15C6435C670C",
INIT_0C => X"79E51E70E070AA8132252008360A7E91504104C8948047D6B0AE1FE440B28A71",
INIT_0D => X"05F0FE40014090400400080329FF8089FF49611F589765923E139F09C78CE7C6",
INIT_0E => X"05F0FE64037FFD7857418407157797878F005F0DFF0F8005F0FE205F0DFF0F80",
INIT_0F => X"8F87FCB1F8053FDEB9B34E0700461E5FF8205F29FF0F8005F0FE205F29FF0F80",
INIT_10 => X"C0184D07C1FF55C3E3E0037FFCF8D3C03009C3CFD53C7E001FF2FAF89781C011",
INIT_11 => X"4E0CDF47186104C6FF177BD939024189BF900401165D645CEEF5BBCDF148F980",
INIT_12 => X"6397F64AEF7F2320483137F8A9BF8A30C2098DFCA06FFFE01F80001F81FDC94F",
INIT_13 => X"FFD051E01015C3BF553D3E0E5FFE838381840714F9DB4F4FA213F774A0E07002",
INIT_14 => X"8B652E2B3120C81284641D3E8DBF7D636FE070189500125C1F83FBCC4F4F80EF",
INIT_15 => X"E7394E339CE138CE5394E33D4E1E0E30E1208C251134921C12A44103F064014B",
INIT_16 => X"7384E3394E338CE538CE1394E3384E738CE139CE1394E7384E339CE139CE5384",
INIT_17 => X"38CE139CE1384E7384E7394E3384E738CE539CE139CE538CE5384E3394E7384E",
INIT_18 => X"7F7B9DB7FF3A1B6DB7ED438A9C3124B2DA6924965B4D384E7384E339CE138CE5",
INIT_19 => X"FBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEF9F7CFDFDDCF3CF3DF5E5BB4E",
INIT_1A => X"7BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEFBEFBEFBEFBE",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE000000000000118D27BBDDEEF77BBDDEEF77BBDDEEF7",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"E955450055421FFFFFBC0010AAD5574BA557FFDFFF0000000000000000000000",
INIT_22 => X"D5575EF55517FF5500557FE10FFFBEAA10007FD7410FFAA97410082A800AAAAA",
INIT_23 => X"FAA955EFA2D168B55557BEAB55005542000007FD74000055574BA5D7FD7555A2",
INIT_24 => X"007BC00AAAAAEBDF45A28428B45FFD168BFF00002AABA5D2ABFFFFAA843DF55F",
INIT_25 => X"AFF80174BAAAD1555EF5555555550055574105D2A800AA00043FEBA5D7FEAA00",
INIT_26 => X"FFAA8415555087BFFF55A2AA800BAFFAE95555080028A00A2FFFDE00F7D57FEB",
INIT_27 => X"545557BC00AAA2FFEAAAA082A97545F7D5420BA5D2E821FFA2D5554BA557BD75",
INIT_28 => X"000000000000000000000000000000000000000000517FE10AAAAA8AAA002E97",
INIT_29 => X"9043D0824850B8A2AE9756D145B401FFFFFFC7010BEDF524AA5571FDFEF00000",
INIT_2A => X"1524BA5571D757DB6D5525EF555178F6D145178E00EBFBE8A101475D5400F7A4",
INIT_2B => X"24BFFFFA28E3AF55F7A0925D7AADB6FB7D5D7FEAB7D0855420BA1471D7438085",
INIT_2C => X"0043FE925571EFA380871C7028B6AEBDF45B68A28B6DEBDF6DBEF1C0A28AAA55",
INIT_2D => X"A2FBF8E10EBD578EAAFF8415482BED1555EF55555057D145152428492E800820",
INIT_2E => X"FB6DF574A85575C55EFBE8E1557D1475FAF45BEAA800AAFFAA9557D080038AAA",
INIT_2F => X"00AAAEA8A9200249056D4175C50920875FDA381C209256DFFDF420BA552A821F",
INIT_30 => X"0BA55557DFF700000000000000000000000000000000000000000000008517DE",
INIT_31 => X"AA105D5155410FF84020AA0800154B2AAAA975FF5D7BC21EFF7FBD7400F7FBC0",
INIT_32 => X"400A25551554BA0051400BA5551575EFF7D1401FF5D5568BE7555568A00AAFFE",
INIT_33 => X"FFDFFF552EA8AAA55043DFF7AAAEAAB55F78400145AAFFFFFEF5D7FEABFF0051",
INIT_34 => X"55400BA082E8201000043FE005D517DEBA0851574B2FFAABFF45FFAAAABFFAAF",
INIT_35 => X"7AA955EF00002AAA2A2FBE8A00A2D16AAAAFF8002410FFD5575EF5555421E755",
INIT_36 => X"FFFFC00BA552A821EFFFFFD74BA5D51575F7FFAE975EF555168B55F7AA800BAF",
INIT_37 => X"000000000000557DE00AAAAAAA000804001FF0055554088A557FEB25D00021FF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000C00000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(0),               -- Port A write enable input
DIA(0)   => data_write_a(5),        -- Port A data input
DOA(0)   => data_read_a_lo_512(5),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(0),               -- Port B write enable input
DIB(0)   => data_write_b(5),        -- Port B data input
DOB(0)   => data_read_b_lo_512(5),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_6_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10800B0061A01002840002C03002818000402322520070B313301C4389B2082",
INIT_01 => X"274008482009404C18A160000C52424841000000090800090210000008510200",
INIT_02 => X"102430600C800110000006100009D070012408000000000648080000001210E0",
INIT_03 => X"000200501D1D02140C420200480140040608010040400104681A0084490C4802",
INIT_04 => X"404402820021000A00824002141000980500000808001114C000080624600600",
INIT_05 => X"120024204209981001A806500304610528000500000080000000300000012940",
INIT_06 => X"2000440832280002300010209C4400142061207A024008900008000220600220",
INIT_07 => X"130C8A220FF41F00902008808800182001020150000001F0800408264000100A",
INIT_08 => X"001BF002C4A01041B1120101000010128568837F04842B080020890008080342",
INIT_09 => X"011847140126805432A62A1596C8B5DF10000008900000100220C00084000008",
INIT_0A => X"44EB4104D09392053589F11C59898888454010830212C54081000410A0088C00",
INIT_0B => X"B0044245B25B456C0096C0096C4096C4096C2096C2096C6096C444B6004B600C",
INIT_0C => X"09040020280010000B3002820110101D0012402CC00802410C26800860070621",
INIT_0D => X"0500819D0000900208201040C4007920004884080000448C281018100C000200",
INIT_0E => X"05008182100000000000000000022AE800C00004000000050081A00004000000",
INIT_0F => X"0002330006000000080000000000000D07A00020000000050081A00020000000",
INIT_10 => X"0000000001204A340002100000000000000000020F4001400000020000000000",
INIT_11 => X"019300020000000068D08000200000001A692121000280000000000010000000",
INIT_12 => X"000201FA100400000000034696010000000000D3478000000000000001003F00",
INIT_13 => X"00000000000000043C0001C0A000008000000000012E000054AC000020000000",
INIT_14 => X"0200000040A410C2810800016000809400001000000000000000433300007600",
INIT_15 => X"060180400000008060180404002AC0200208940041309210B28048180F028000",
INIT_16 => X"2008000100601802000000100601800000000180600800000020180600000000",
INIT_17 => X"0180600000008040100200800000060100000802010040180200002018040100",
INIT_18 => X"7F8FF0F4FA955F7CF7F40A80907638C31C71C718638E00006018040080200004",
INIT_19 => X"38E38E38E38E38E38E38E38E38E38E38E38E38E39B6CEDECDDF7DF7DF5F78BCE",
INIT_1A => X"3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE38E38E38E38E",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFF000000000000196A03F9FCFE7F3F9FCFE7F3F9FCFE7F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"00000000000000000000000C0FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"BFDF45F7AA974AAAAAA97555F784174BAF7D5555FF0000000000000000000000",
INIT_22 => X"FBD7410AA8428AAAAAAE955450055421FFFFFBC0010AAD5574BA557FFDFFF087",
INIT_23 => X"FFBEAA10007FD7410FFAA97400082A800AA08515555508043FE00F7AA97555A2",
INIT_24 => X"55517FF55A2AA97400552AAAB45082E80155F7D1575EFFFAA9555500557FE10F",
INIT_25 => X"FF7AAA8A10082EAAB45A2FFC2000007FD74000055574BA5D7FD7555A2D5575EF",
INIT_26 => X"FFAA843DF55FFAA955EFA2D168B55557BEAB5500554200000003DE10FFD5401F",
INIT_27 => X"BFF00002AABA5D2ABFFFF087BD5545007BFDE10AA803FE105D516AABAFF843FF",
INIT_28 => X"0000000000000000000000000000000000000000AAAEBDF45A28428B45FFD168",
INIT_29 => X"524AA5571FDFEF1C7BFFF55FFA095482B6A49256DEB84104BAFFD1525FF00000",
INIT_2A => X"03DE28F7A49057DAAF5D2428A2842AAAAA2AE9756D145B401FFFFFFC7010BEDF",
INIT_2B => X"A49756D145178E00EBFBE8A101475D5400F7A4904380824850381C5B5057D1C0",
INIT_2C => X"571D757DB6D5525EF555178F6DAAA495428412AAFB451C2A8017DE3DF525FFFF",
INIT_2D => X"1C0E3FE00E3DB471EFE3AAAAA00082EA8B6DA2F1C50381471D74380851524BA5",
INIT_2E => X"049516AAB8FF8428FEFA28E3AF55F7A0925D7AADB6FB7D5D7FEAB7D0855420BA",
INIT_2F => X"45B68A28B6DEBDF6DBEF1C0A28AAA5524BFFFF1C7BD057D1C71FFE10A28038E1",
INIT_30 => X"0AAFFD1401E7000000000000000000000000000000000000000000000B6AEBDF",
INIT_31 => X"21EFF7FBD7400F7FBC00BA55557DFF7557BFDF55F78017400F780001FFAA8400",
INIT_32 => X"154B2557FC01EF55043FEAAFF80021EFA2D1420BAAA8428AA2AAAA975FF5D7BC",
INIT_33 => X"A821EFAAFBC01FFF780155F7555568A00AAFFEAA105D5155410FF84020AA0800",
INIT_34 => X"51554BA0051400BA5551575EFF7D1401FF5D5568BE7AA80174AA082ABDF555D2",
INIT_35 => X"D7FEABFF0051400A25D2EBFE10AAFFD55EFA2AEA8A10082EA8BEFAAD5554B255",
INIT_36 => X"55557DE00AA842AA0000516AABAFF8428BE7AAAEAAB55F78400145AAFFFFFEF5",
INIT_37 => X"0000000000FFAABFF45FFAAAABFFAAFFFDFFF552EA8AAA55043DFF7557BC01EF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000900000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(0),               -- Port A write enable input
DIA(0)   => data_write_a(6),        -- Port A data input
DOA(0)   => data_read_a_lo_512(6),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(0),               -- Port B write enable input
DIB(0)   => data_write_b(6),        -- Port B data input
DOB(0)   => data_read_b_lo_512(6),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_7_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10844B00482258A2842112C02450418800002300500030B313300C418992002",
INIT_01 => X"234008422008604D1C20E0000E11426840000000080000080200090000110204",
INIT_02 => X"1025207000B08910000206101188D03080144880010400044808000000122160",
INIT_03 => X"000200401914821004420000CA01000C0600010000605114291A008449484802",
INIT_04 => X"40440200002100080006500210101019040000000B085024D842080244000000",
INIT_05 => X"1A8024200009981001A8224001040104200204000000800CC2092CE4A0004900",
INIT_06 => X"A000440822280002340010209C040014A061200052500810000C490323208E28",
INIT_07 => X"128802020028000890240980A809102001020140000009F0800408264000100A",
INIT_08 => X"001A0602C4A01051B13281010408881203480200448423199046821008082351",
INIT_09 => X"336784144126811054809C1040140A001C8648481000045903318B80A400310A",
INIT_0A => X"000800009010100014114110312388984502148282A08415B032095048008100",
INIT_0B => X"20CDC1C483484D201192011920119201192051920519205192074C9018C90188",
INIT_0C => X"D8A5B44001D2C12901228F82F005310D293054048A2212004466000DA1908528",
INIT_0D => X"800F8108A0D09802082010408580008000000008C85264010816851B428DA146",
INIT_0E => X"800F81321000020000261900E28A204040E000A0000007800F814000A0000007",
INIT_0F => X"7072024807000020400000581C01C1A406400084000007800F81400084000007",
INIT_10 => X"060180E83800E820101210000200000CC3003C32080201C0000C000000160700",
INIT_11 => X"81DD00804086423120B74020023090644840A34000828800000004000420020B",
INIT_12 => X"1C6A0186E8000446120C8905BA0004810C84624237E00010001878007F0030C0",
INIT_13 => X"00080208E4083C44230201AEE0010040261900E30520C0806EAC0082000984C0",
INIT_14 => X"0121011088A600C032128201519480D40005802448160403E0700622C0806EE8",
INIT_15 => X"A1685A1685A168DA368DA36CDA30DA13A108810111349A943AA4401000928A19",
INIT_16 => X"368DA768DA1685A1685A5685A368DA368DA7685A1685A1685A768DA368DA368D",
INIT_17 => X"685A1685A169DA368DA1685A1695A368DA3685A1685A168DA368DA1685A1685A",
INIT_18 => X"00000000000000000000400A8448410400020820800069DA1685A168DA369DA3",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000003667B000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"0155EFAAAEA8ABAAAFBFDE0055556AA005D04155550000000000000000000000",
INIT_22 => X"556AA00FFAE95555087BFDF45F7AA974AAAAAA97555F784174BAF7D5555FFF78",
INIT_23 => X"055421FFFFFBC0010AAD5574BA557FFDFFF5555555EFAAFFFDFEFAAAAAAB455D",
INIT_24 => X"AA8428AAA557BFDFFF55003DFFFF7FBEAA00002EAAAAA082EA8A00AAAE955450",
INIT_25 => X"0552EBDE00007BEAAAAA2D14000008515555508043FE00F7AA97555A2FBD7410",
INIT_26 => X"FF00557FE10FFFBEAA10007FD7410FFAA97400082A800AAF7AE975FFA2800001",
INIT_27 => X"155F7D1575EFFFAA955555D51574AAAAFFD5545087FEAB455D516AB55557BD55",
INIT_28 => X"0000000000000000000000000000000000000000A2AA97400552AAAB45082E80",
INIT_29 => X"104BAFFD1525FFFF8E175C7A2AAAAA82A2F1FAE105D556AA10410E1755500000",
INIT_2A => X"1FFFD7AAAAAFB7D495F6AA10E3AE905551C7BFFF55FFA095482B6A49256DEB84",
INIT_2B => X"2EAAA00A2AE9756D145B401FFFFFFC7010BEDF524AA5571FDFEF415B575D7AAF",
INIT_2C => X"7A49057DAAF5D2428A2842AAAA497BFAFFF49003AFEFEBFBEAA001C2EA8A821C",
INIT_2D => X"F7A4905C7A28A070384120BDE100075EAA82BEDB470101C5B5057D1C003DE28F",
INIT_2E => X"D555F6AB57417BC05D7145178E00EBFBE8A101475D5400F7A490438082485038",
INIT_2F => X"28412AAFB451C2A8017DE3DF525FFFFA49756D495150492BEF1D2555087BE8B7",
INIT_30 => X"A10002E9754D000000000000000000000000000000000000000000000AAA4954",
INIT_31 => X"7400F780001FFAA84000AAFFD1401E7FFAA97555A2AEA8A10AAD568A00555168",
INIT_32 => X"7DFF7007BD5555AAD57DF55AAAEBDFEF007BE8A10AAAE8215D557BFDF55F7801",
INIT_33 => X"FEAA105D2EAAA005D2AAAA18AAAA975FF5D7BC21EFF7FBD7400F7FBC00BA5555",
INIT_34 => X"7FC01EF55043FEAAFF80021EFA2D1420BAAA8428AA2007FE8BFF080028BFFAAF",
INIT_35 => X"F84020AA0800154B2FF8402145A2AA954AA00043DE0000516AA10F7FBD740855",
INIT_36 => X"FFD140145007FE8BEF557BEAB55087FC215D555568A00AAFFEAA105D5155410F",
INIT_37 => X"0000000000AA80174AA082ABDF555D2A821EFAAFBC01FFF780155F7005140000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000000FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(0),               -- Port A write enable input
DIA(0)   => data_write_a(7),        -- Port A data input
DOA(0)   => data_read_a_lo_512(7),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(0),               -- Port B write enable input
DIB(0)   => data_write_b(7),        -- Port B data input
DOB(0)   => data_read_b_lo_512(7),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_8_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00000648E2840112C00000418000002700500030B3132000400812086",
INIT_01 => X"214009C21838284D042100000212026840000000180800080200080040510204",
INIT_02 => X"1021004000900110000006100088503000240800014400004808000000122160",
INIT_03 => X"0002004019110214044A82000121400C86000000000000860188008448400002",
INIT_04 => X"000402800031200A0000090214100889A5000000490090104800000224000400",
INIT_05 => X"10C025204289981000A820500344010428008500010080080909304040202004",
INIT_06 => X"8000440003280000340010208C04003420600000C6180810000C490703200010",
INIT_07 => X"130002000028000890240980A809012001020050000009F08004082640000082",
INIT_08 => X"20100402C4201041310041010008801201480200051023090024811008090A1A",
INIT_09 => X"0100001001248100308214528148A48008000008100004590711C04034000083",
INIT_0A => X"10804000801210140001C0103001088845010482004000008420041020008900",
INIT_0B => X"0004404002004400448000480004800048000480004800048000440022400200",
INIT_0C => X"880420000880204909004502D100A10C04205424010216010C26800805000004",
INIT_0D => X"8000801100509802082010400400018000488428800004082014000200010000",
INIT_0E => X"8000800A00000207A8BE7B00000200082040808000F07F80008000808000F07F",
INIT_0F => X"0002000402100000404CB1F8FC0000040000808000F07F80008000808000F07F",
INIT_10 => X"3E07800000004004080A000002072C3FCF0000020040804800040007687E3F00",
INIT_11 => X"10800018639EC00020100002C2F9B0000801016001008100000040120CB3067F",
INIT_12 => X"000200020000585EB6000100800030C73D8000402000001FC07FF80001000080",
INIT_13 => X"002EAE1FEC0000040200408000003C547E7B00000100801004000803551F8FC0",
INIT_14 => X"00000000440610C8000A808040000208901B86E568FE0C000000020080100400",
INIT_15 => X"0040100401004090240902449028D0230249850101349A98BAC0481000888810",
INIT_16 => X"0401004010040100401004010240902409024090240902409004010040100401",
INIT_17 => X"4010040100409024090240902409004010040100401004090240902409024090",
INIT_18 => X"543EBC57A10A1E75D6440A889050000000000000000040902409024010040100",
INIT_19 => X"79E79E79E79E79E79E79E79E79E79E79E79E79E7BF3CCD8DF5B2DB2CA4028A0A",
INIT_1A => X"4F87D3E1F4F87D3E1F4F87D3E1F4F87C3E1F0F87C3E1F0F87C3E79E79E79E79E",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000000D3E94F87D3E1F4F87D3E1F4F87D3E1F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"000000087BEAA10F7803DE00FFAEBFFFF0800155FF0000000000000000000000",
INIT_22 => X"7FC2145005155555F780155EFAAAEA8ABAAAFBFDE0055556AA005D0415555080",
INIT_23 => X"7AA974AAAAAA97555F784174BAF7D5555FF552AA8AAA557FC0010F780154105D",
INIT_24 => X"FFAE95555AAFFE8A00552EBFE00F7D17FF45F7FFFFF55AA80155FF087BFDF45F",
INIT_25 => X"5F7D140010552E821EFAAAABDF555555555EFAAFFFDFEFAAAAAAB455D556AA00",
INIT_26 => X"00AAAE955450055421FFFFFBC0010AAD5574BA557FFDFFF5504000AAAAAAA8B5",
INIT_27 => X"A00002EAAAAA082EA8A00002AA8A10F78402155AA8028A00A2D57FF45557BE8A",
INIT_28 => X"0000000000000000000000000000000000000000557BFDFFF55003DFFFF7FBEA",
INIT_29 => X"6AA10410E17555080E000280071E8A00EB8E3FE10F7AEBAFFF080A175D700000",
INIT_2A => X"1C2000FF8A17400557FC015514555757DFF8E175C7A2AAAAA82A2F1FAE105D55",
INIT_2B => X"8A105D71C7BFFF55FFA095482B6A49256DEB84104BAFFD1525FF492EA8AAA557",
INIT_2C => X"AAAAFB7D495F6AA10E3AE90555A2FBE8A38492ABDE10EBDF7AF6DE3FFF8F7DB6",
INIT_2D => X"550E00082B6A0AFB55F7D1420104124821D7AAA0BDF6D415B575D7AAF1FFFD7A",
INIT_2E => X"0B6D578F6D557FFDA00A2AE9756D145B401FFFFFFC7010BEDF524AA5571FDFEF",
INIT_2F => X"FF49003AFEFEBFBEAA001C2EA8A821C2EAAA001C2EA8A00F7800017DA2842FA0",
INIT_30 => X"BEF082E95545000000000000000000000000000000000000000000000497BFAF",
INIT_31 => X"8A10AAD568A00555168A10002E9754D082E820BA08556AA00AAAABFE00F7AEAA",
INIT_32 => X"401E7082EAAABA5D5140010F7AE974105D7BC21555D51575EFFFAA97555A2AEA",
INIT_33 => X"BEABFFAAFBEABFFF7AA80145557BFDF55F78017400F780001FFAA84000AAFFD1",
INIT_34 => X"7BD5555AAD57DF55AAAEBDFEF007BE8A10AAAE8215DA2FFE8ABA082ABFE00AAF",
INIT_35 => X"7FBC00BA55557DFF75D2E82010F7843DF45FFD540000000402145AA843FFFF00",
INIT_36 => X"F780021FFA2803DE10FFD16ABFF5D7BFDE10AAAA975FF5D7BC21EFF7FBD7400F",
INIT_37 => X"0000000000007FE8BFF080028BFFAAFFEAA105D2EAAA005D2AAAA185D2AAAA10",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000400000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(1),               -- Port A write enable input
DIA(0)   => data_write_a(8),        -- Port A data input
DOA(0)   => data_read_a_lo_512(8),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(1),               -- Port B write enable input
DIB(0)   => data_write_b(8),        -- Port B data input
DOB(0)   => data_read_b_lo_512(8),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_9_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000B0001800002840002C0000281800000030000000033022000000000002",
INIT_01 => X"8000098218302849180060000C004240413C0A61590001D90213C90008510200",
INIT_02 => X"000008700CB089100002061031200074810448800104008048080080001210E2",
INIT_03 => X"000200140C1822000A028010408100000628000140402080041A100040024840",
INIT_04 => X"41040000000400080002040200080800040000000B08D1055842080604600700",
INIT_05 => X"10002024000020102400010000026104200004000400800C8B0024E4E0010C40",
INIT_06 => X"8000440802280002700800008A840004A0610000C0000810000C590103600810",
INIT_07 => X"538600220028001890240980A80800200102025000000BF08200002440000883",
INIT_08 => X"00000402C220104131102101040810028528820005100003900E884000010007",
INIT_09 => X"00000005E000000600BCA284140200800C834948100004590111824404012080",
INIT_0A => X"04080000901012100A1141005922000245410002008880000032005080000800",
INIT_0B => X"2000020040044010440104401004010440100401044010040104400802008208",
INIT_0C => X"D1A1344420D2E100000808000000000481000000202002400006800825908402",
INIT_0D => X"0500000000109000000000000580008000080000C852240100068D0B4685A342",
INIT_0E => X"0500000A00000000000000000000028000408020000000050000208020000000",
INIT_0F => X"0000304002100020000000000000000900208004000000050000208004000000",
INIT_10 => X"0000000001200000000A00000000000000000000050000480008000000000000",
INIT_11 => X"009F0080000000004807C0200000000012000020000081000000040000000000",
INIT_12 => X"00000048F8000400000002403E0004000000009067E000000000000000000900",
INIT_13 => X"0000000000000000140000CEE001000000000000000A000036AC008000000000",
INIT_14 => X"03210000000400CA81000000619480D4000400000000000000004100000036E8",
INIT_15 => X"A368DA368DA3685A1685A1685A121A11A1419001512490040024001000008019",
INIT_16 => X"1685A1685A1685A1685A1685A368DA368DA368DA368DA368DA368DA368DA368D",
INIT_17 => X"685A1685A168DA368DA368DA368DA368DA368DA368DA3685A1685A1685A1685A",
INIT_18 => X"CCF48DE68A895C38E250080000000000000000000000685A1685A1685A1685A1",
INIT_19 => X"514514514514514514514514514D34D34D34D34D28E10040392482090157344C",
INIT_1A => X"4D268341A0D069349A0D069349A0D068341A0D068341A0D06834514514514514",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000001654D0D069349A0D068341A4D268341A",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"BE8B45002A974AAAA803DFFFAA843DF45FFFFEAABA0000000000000000000000",
INIT_22 => X"AEBDE00AAFBEAABA080000000087BEAA10F7803DE00FFAEBFFFF0800155FFAAF",
INIT_23 => X"AAEA8ABAAAFBFDE0055556AA005D0415555087BFDE00A2FBD7400F7FBFDFFFA2",
INIT_24 => X"005155555557BE8BEF007FFDEAAAAD1555EF0055401FFF7AEAAA10F780155EFA",
INIT_25 => X"0F7AA974AA082E80010A2AAAAA10552AA8AAA557FC0010F780154105D7FC2145",
INIT_26 => X"BA087BFDF45F7AA974AAAAAA97555F784174BAF7D5555FFF780154AA5D2AA8A1",
INIT_27 => X"F45F7FFFFF55AA80155FF080400145FFFBEAABAF7D17FEBAA2AEBDF45002EAAA",
INIT_28 => X"0000000000000000000000000000000000000000AAFFE8A00552EBFE00F7D17F",
INIT_29 => X"BAFFF080A175D7BEF1E8B6D002090482B68E38FC7BE8A3DF7DF7F5E8A9200000",
INIT_2A => X"BD0400FFF5FDFC7B6A0BDE38B6F5E8A92080E000280071E8A00EB8E3FE10F7AE",
INIT_2B => X"AAA8A38FF8E175C7A2AAAAA82A2F1FAE105D556AA10410E175550871FFE00A2F",
INIT_2C => X"F8A17400557FC015514555757D5D71E8BEF147BFAE82A2DB555C71C5B451D7FF",
INIT_2D => X"FF84174BA5D20AAA00E3AA904BA142A87010A2AEADA38492EA8AAA5571C2000F",
INIT_2E => X"AAAA0BFF7D0024ADA921C7BFFF55FFA095482B6A49256DEB84104BAFFD1525FF",
INIT_2F => X"38492ABDE10EBDF7AF6DE3FFF8F7DB68A105D7000400155FFFBEDA82FFD57DEB",
INIT_30 => X"FEFF7D16AA00000000000000000000000000000000000000000000000A2FBE8A",
INIT_31 => X"AA00AAAABFE00F7AEAABEF082E95545F7D568BEF080402000F7AAA8B55FFAABD",
INIT_32 => X"9754D00517DE00A2FFC2000F7D17FF55FF803FEAAFFD16AA00082E820BA08556",
INIT_33 => X"FD55555D7FD5555FFAAA8AAAFFAA97555A2AEA8A10AAD568A00555168A10002E",
INIT_34 => X"2EAAABA5D5140010F7AE974105D7BC21555D51575EF555568BEF5D7FE8A10AAF",
INIT_35 => X"A84000AAFFD1401E7FF80174AA5D0028A00AAAE800AA552A97400A2AEBDEAA08",
INIT_36 => X"F7FBFFE00FFD17FEAAA2803DFEF08043FE00557BFDF55F78017400F780001FFA",
INIT_37 => X"0000000000A2FFE8ABA082ABFE00AAFBEABFFAAFBEABFFF7AA80145080002145",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000800000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(1),               -- Port A write enable input
DIA(0)   => data_write_a(9),        -- Port A data input
DOA(0)   => data_read_a_lo_512(9),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(1),               -- Port B write enable input
DIB(0)   => data_write_b(9),        -- Port B data input
DOB(0)   => data_read_b_lo_512(9),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_10_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000B0001800002840002C0000281800020030000000033022000000180006",
INIT_01 => X"000008000000004C002000000010026840000000080000080200000000110200",
INIT_02 => X"0000004000800110000006100000003000040800010400004808000000120060",
INIT_03 => X"000200000810020000020000400100000600000000400000001A000040004800",
INIT_04 => X"0004000000000008000200020000000004000000080010004000000200000000",
INIT_05 => X"1000202000011010000000000000010520000400000080000000200000200004",
INIT_06 => X"80004408022800023000000088040004A061000040000810000C490103600000",
INIT_07 => X"120420020028000890240980A808002001020050000009F08000002440000082",
INIT_08 => X"00000402C0201051311001000000020201080200440400000000800000000000",
INIT_09 => X"0000105808000000000000000000008000008088100004590111800004000000",
INIT_0A => X"00804000801210440003C1411008800045000002000014000040009002800000",
INIT_0B => X"0400200000000000000004000040000000000000040000400000000000000221",
INIT_0C => X"0100802000000000000002802000000400100000000002000026000840011400",
INIT_0D => X"0500000000409002082010400400008000400008002044082000081004080204",
INIT_0E => X"0500000200000000000000000000028000400000000000050000200000000000",
INIT_0F => X"0000304002000000000000000000000900200000000000050000200000000000",
INIT_10 => X"0000000001200000000200000000000000000000050000400000000000000000",
INIT_11 => X"0082000000000000480080000000000012000101000080000000000000000000",
INIT_12 => X"0000004810000000000002400400000000000090400000000000000000000940",
INIT_13 => X"0000000000000000150000C00000000000000000000A40001400000000000000",
INIT_14 => X"02000000002400C2810000006000000000000000000000000000410040001400",
INIT_15 => X"020080200802008020080200800800220200840001309A08A848001000008000",
INIT_16 => X"0000000000000000000000000200802008020080200802008020080200802008",
INIT_17 => X"0080200802000000000000000000000000000000000000000000000000000000",
INIT_18 => X"940FE0D397124355520542821010000000000000000000802008020080200802",
INIT_19 => X"28A28A28A28A28A28A28A28A28A28A28A28A28A29554199854514514F546890A",
INIT_1A => X"32994CA6532995CAE572B94CA6532994CA6532994CA6532994CA28A28A28A28A",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000001867172B94CA6532994CA6572B95CAE5",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FC2155F7D155545AA80001EFAAFBEAB45557FFDE100000000000000000000000",
INIT_22 => X"FBE8BFFF78402155AAFBE8B45002A974AAAA803DFFFAA843DF45FFFFEAABA007",
INIT_23 => X"87BEAA10F7803DE00FFAEBFFFF0800155FF00042AB55FFD168B55AA8000010FF",
INIT_24 => X"AAFBEAABAA2FFD741055003DFEFF7AA801FFAAD16AABA002ABDE100800000000",
INIT_25 => X"FF7FBC0145F78028A00A2D142155087BFDE00A2FBD7400F7FBFDFFFA2AEBDE00",
INIT_26 => X"BAF780155EFAAAEA8ABAAAFBFDE0055556AA005D0415555007FD74105555555E",
INIT_27 => X"5EF0055401FFF7AEAAA105D042ABFF5D556AB55AAD168ABA002A975FFF7AEBDE",
INIT_28 => X"0000000000000000000000000000000000000000557BE8BEF007FFDEAAAAD155",
INIT_29 => X"3DF7DF7F5E8A92007BC217DEBDB55555AA8E071D7AAFBEFB455D71F8E0000000",
INIT_2A => X"B6DB55BE8E05000EBFFE8BC7E38E07145BEF1E8B6D002090482B68E38FC7BE8A",
INIT_2B => X"2EB8E00080E000280071E8A00EB8E3FE10F7AEBAFFF080A175D700042AB7DEBD",
INIT_2C => X"FF5FDFC7B6A0BDE38B6F5E8A92B6FBD5410490A3DFD7F7A4821D7A2D16FA8214",
INIT_2D => X"0071D54104951555D7EBF5C5155E3842AA00BED1421450871FFE00A2FBD0400F",
INIT_2E => X"20820955EFE3AEBDEAAFF8E175C7A2AAAAA82A2F1FAE105D556AA10410E17555",
INIT_2F => X"EF147BFAE82A2DB555C71C5B451D7FFAAA8A38410E2ABD749516FB55BED16FA8",
INIT_30 => X"F455D556AA000000000000000000000000000000000000000000000005D71E8B",
INIT_31 => X"2000F7AAA8B55FFAABDFEFF7D16AA00087FC01EFA2FFD7545AAAE97555A2FBFD",
INIT_32 => X"9554500042ABFFA2FFFFF45F7AE97400AAFFE8B45AAAA95545F7D568BEF08040",
INIT_33 => X"400155A2D57FE00552EA8A00082E820BA08556AA00AAAABFE00F7AEAABEF082E",
INIT_34 => X"517DE00A2FFC2000F7D17FF55FF803FEAAFFD16AA00FFFBD5400082EBFF45F78",
INIT_35 => X"55168A10002E9754D085155410085557555AAD557555A2802AA10FFD54214500",
INIT_36 => X"08557DF55F7D17FE000804155FFAAAABDEAAFFAA97555A2AEA8A10AAD568A005",
INIT_37 => X"0000000000555568BEF5D7FE8A10AAFFD55555D7FD5555FFAAA8AAA002AAAB45",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000008FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(1),               -- Port A write enable input
DIA(0)   => data_write_a(10),        -- Port A data input
DOA(0)   => data_read_a_lo_512(10),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(1),               -- Port B write enable input
DIB(0)   => data_write_b(10),        -- Port B data input
DOB(0)   => data_read_b_lo_512(10),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_11_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10180B05A0010402840602C2D001019000000300000000330A20080EC180002",
INIT_01 => X"AB400986B830284D1820E0000C3642484000000008000008820009080A512220",
INIT_02 => X"102A68440080011000000618062AD03502640800010410424908136019920868",
INIT_03 => X"004A0846191B22120642000442C110044600000101E9225CDC9A10844A9A4842",
INIT_04 => X"0094024000250808800216021138000B848000000800100040000102A0600200",
INIT_05 => X"7E4024242008A8102CA88A44010401042200444000888000000028000002A002",
INIT_06 => X"8088445712280000B18812288E0400253855200045C86810000C5B0503286A28",
INIT_07 => X"10008822A028004880200A80880208200122006C000015F0C20408264902C840",
INIT_08 => X"9390040280241041D1754100000018108728820024002B3A01A89540080824C8",
INIT_09 => X"A1001C41A1348498B080801010000080D00301081000045B0511D28D94012339",
INIT_0A => X"44080000901012428003414158230CBA4576708241C010908040341322008000",
INIT_0B => X"040464D280144050C72A0872A0C72A0872A0C72A0C72A0872A0C595043950421",
INIT_0C => X"0804001400000820110A42822204880CD81040442900021704E6000800001D54",
INIT_0D => X"80C62D0500409002082010404580018000404012004004192C10000000000000",
INIT_0E => X"80C62D5803161C526DB40506C120A806ABB0D808CC334A80A54B70D408CC32D2",
INIT_0F => X"2B5144D0DD903C54916D15458C0513005570D408CC334A80A54B70D808CC32D2",
INIT_10 => X"52148C4DB05621E363F813961C20EDA944016558C2347A080B10D8DD6422AA10",
INIT_11 => X"1880144D3345C65593800319C18BD1ECA1C9010112566F10AC4183C340DAE02D",
INIT_12 => X"5810503000633830DE3C2C9C00289A66AA8DE50E0800360614AC281430890600",
INIT_13 => X"0CD2A9CEA8199B6B082B55900314140365320485C4F00AD544407241C175C402",
INIT_14 => X"0000074044C4801832701A89D20A38093631425969020855A281844E00540404",
INIT_15 => X"0000000000000000000000000020C00200088101513492101280401000400200",
INIT_16 => X"2008020080200802008020080000000000000000000000000000000000000000",
INIT_17 => X"0080200802008020080200802008020080200802008020080200802008020080",
INIT_18 => X"804180C0B10A4210420140028400000000000000000000802008020080200802",
INIT_19 => X"000000000000000000000000000820820820820801C414947000000055062608",
INIT_1A => X"0000000004020000000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000001F87E000000000000010080000000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"ABDF5508557DF45002ABDFFFF7803DE10AA80000AA0000000000000000000000",
INIT_22 => X"FFE8A10A28000000007FC2155F7D155545AA80001EFAAFBEAB45557FFDE10082",
INIT_23 => X"02A974AAAA803DFFFAA843DF45FFFFEAABAA2AEBFF45FFAEBFEAA002A801FFF7",
INIT_24 => X"F78402155AAD155555A28428BFF002ABDE00A2AABFE10082ABFFEFAAFBE8B450",
INIT_25 => X"0002A80010A2842AAAA007BFFF4500042AB55FFD168B55AA8000010FFFBE8BFF",
INIT_26 => X"00080000000087BEAA10F7803DE00FFAEBFFFF0800155FF00557FF45557FC201",
INIT_27 => X"1FFAAD16AABA002ABDE10A2D168A10A284021FF5D00154BAF7FBE8BEFFFD5400",
INIT_28 => X"0000000000000000000000000000000000000000A2FFD741055003DFEFF7AA80",
INIT_29 => X"EFB455D71F8E00002EBDF6D005B78F7D142ABDFC7F78E3FE28B684070AA00000",
INIT_2A => X"0BDEAA1C2A801C7E3FFEFA10B68407038007BC217DEBDB55555AA8E071D7AAFB",
INIT_2B => X"20B8FEFBEF1E8B6D002090482B68E38FC7BE8A3DF7DF7F5E8A92BEAEBFF7DEBA",
INIT_2C => X"E8E05000EBFFE8BC7E38E07145B6D15756DA28A28BFF082ABAE10B6AAB8E2808",
INIT_2D => X"08517DF7D497BC5028142A87000A28A2AA92007FF8F7D00042AB7DEBDB6DB55B",
INIT_2E => X"2FFFFEFBC7E3DF42028080E000280071E8A00EB8E3FE10F7AEBAFFF080A175D7",
INIT_2F => X"10490A3DFD7F7A4821D7A2D16FA82142EB8E00B6DB6AA28A280001FF5D0A1048",
INIT_30 => X"EAAF784154BA000000000000000000000000000000000000000000000B6FBD54",
INIT_31 => X"7545AAAE97555A2FBFDF455D556AA00082EBFFEF007BE8BFF5D2ABDF55F7AABD",
INIT_32 => X"6AA00FFAEBFFEFAA803DEBA5D2E82155A2FBFDE00FF84154BA087FC01EFA2FFD",
INIT_33 => X"AAAA00FFAAA8AAA080028BFFF7D568BEF080402000F7AAA8B55FFAABDFEFF7D1",
INIT_34 => X"042ABFFA2FFFFF45F7AE97400AAFFE8B45AAAA95545F7D5555FFAAAAA8BFF002",
INIT_35 => X"7AEAABEF082E9554508557DFFF007BD54BA5D2E95400A2AEA8A00007FEABFF00",
INIT_36 => X"AA80001FF5D2E82000F7FFFFF45AAFFC20BA082E820BA08556AA00AAAABFE00F",
INIT_37 => X"0000000000FFFBD5400082EBFF45F78400155A2D57FE00552EA8A00FFFFE8AAA",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000800000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(1),               -- Port A write enable input
DIA(0)   => data_write_a(11),        -- Port A data input
DOA(0)   => data_read_a_lo_512(11),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(1),               -- Port B write enable input
DIB(0)   => data_write_b(11),        -- Port B data input
DOB(0)   => data_read_b_lo_512(11),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_12_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A500C4B01BC0268A6940312C0DE045196A831A300500032B333287E4FC812006",
INIT_01 => X"AF400D869830E84D5823E0000C1742484000000008000008820009280A553235",
INIT_02 => X"502A7144008001100000171C022BD13412762A000586235ECC09C8423B960866",
INIT_03 => X"31863846191BA218064204000281200406A10843010022DEDF0852944A9C014A",
INIT_04 => X"0014030000250409000014821038080B840000400800102040000302F0600233",
INIT_05 => X"7FC034348008A8102CA88F48010601042400048000188000000938000002E088",
INIT_06 => X"9CC96CC6F63A5001F12B56A0AC8601F47AC06400D1F80C10020C493F03343A38",
INIT_07 => X"1020002030280098A12048908A16BA311177124C000003F08A94282E5C262861",
INIT_08 => X"827A0602902A10491165E10000049010C52882008600A73A01E8974008092CF8",
INIT_09 => X"47000001A1248008F000000000000080000F010C100204593F11A6CDF48023BF",
INIT_0A => X"040000208010120ACA01400058010CBA4D277C86CCE802B380003C1360008000",
INIT_0B => X"011C46D3C7BC1EF083AF0C3AF083AF083AF0C3AF083AF083AF0C1D7861D78400",
INIT_0C => X"08040014C9001AE91D17E50AD79FEFC87C2154745F82131FFCCE00080000095E",
INIT_0D => X"807BF7118180984004000803D40001880001001400C005031010000000000000",
INIT_0E => X"807BF76A109C944B5891BF06C5EEB14FCBF0D90076D61C807BF7D0D80876D49C",
INIT_0F => X"6DE38EB9FB10350C00A99F7CA80757365E50D80876D61C807BF7D0D90076D49C",
INIT_10 => X"841BCC69A0D8C6F7F0AA001C943A65756A0976EB5A7E7FC8951018186334F311",
INIT_11 => X"D5A014481991C6A737D80211912970CDCDD1864116D6C7080651CB4661F33615",
INIT_12 => X"349E929300423224AE19B9BEC0289033238D4E6EA805892946A9B011A7B152CF",
INIT_13 => X"6244CD7AC01CAAA56B3E6D9001068715D64006D2A961CF9B44512A2504532182",
INIT_14 => X"00000439FDC25C58067A9FAB46095A0B5289A0282D2E1444ACB12A17CF9B4414",
INIT_15 => X"0000000000000000000000040026C00000288401513492909280401000F70A00",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"088881360A95090CB05442029010000000000000000000000000000000000000",
INIT_19 => X"1041041041041041041041041049249249249249200100002D4514510051B946",
INIT_1A => X"592C964B2592C964B2592C964B2592C86432190C86432190C864104104104104",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000002007F592C964B2592C964B2592C964B2",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"43FE0008557DFFF0800020105D557FEAA00557DE100000000000000000000000",
INIT_22 => X"557DFFFF7AA80000082ABDF5508557DF45002ABDFFFF7803DE10AA80000AAAA8",
INIT_23 => X"7D155545AA80001EFAAFBEAB45557FFDE10AAD5420000051555FFA2AA8200000",
INIT_24 => X"A28000000A2D155410F7FFFFEBA08003FE00082AA8AAAAAFFC00BA007FC2155F",
INIT_25 => X"0A2AABFE1055516ABEF5D517DEAAA2AEBFF45FFAEBFEAA002A801FFF7FFE8A10",
INIT_26 => X"55AAFBE8B45002A974AAAA803DFFFAA843DF45FFFFEAABA000028A105D2ABFE1",
INIT_27 => X"E00A2AABFE10082ABFFEF085542000000417555002A820AA08557DFFFF7AA821",
INIT_28 => X"0000000000000000000000000000000000000000AAD155555A28428BFF002ABD",
INIT_29 => X"3FE28B684070AABE803AE38145B78FD7000005010495B7AE921C517DE1000000",
INIT_2A => X"B505FFB6A487000005F7AFD7F7A482038002EBDF6D005B78F7D142ABDFC7F78E",
INIT_2B => X"F5C2082007BC217DEBDB55555AA8E071D7AAFBEFB455D71F8E00BED547038145",
INIT_2C => X"C2A801C7E3FFEFA10B68407038B6D550428FFF1FDE821C003FE001C2EAAAAAB6",
INIT_2D => X"00002FA285D20BDE28A2A4B8E10555B68BEF5D517DEAABEAEBFF7DEBA0BDEAA1",
INIT_2E => X"2005F7DFD7F7A482155BEF1E8B6D002090482B68E38FC7BE8A3DF7DF7F5E8A92",
INIT_2F => X"6DA28A28BFF082ABAE10B6AAB8E280820B8FEF085F4703814001055514208208",
INIT_30 => X"A0055517DE00000000000000000000000000000000000000000000000B6D1575",
INIT_31 => X"8BFF5D2ABDF55F7AABDEAAF784154BAF7802AABA5D7FEAB45080015410007FEA",
INIT_32 => X"6AA00F7D1554BA5D7BC01FFFF8015410007FEAB45F780020BA082EBFFEF007BE",
INIT_33 => X"43FE10552EAAAAAFFD140000087FC01EFA2FFD7545AAAE97555A2FBFDF455D55",
INIT_34 => X"AEBFFEFAA803DEBA5D2E82155A2FBFDE00FF84154BAF7D1400BAFFD57FE005D0",
INIT_35 => X"FAABDFEFF7D16AA0008003FEBA55003DEBAA28428A105D7FEABEF55557DEBAFF",
INIT_36 => X"550402145550000010087FFFF45F78402145F7D568BEF080402000F7AAA8B55F",
INIT_37 => X"0000000000F7D5555FFAAAAA8BFF002AAAA00FFAAA8AAA080028BFF087BD54AA",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000000FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(1),               -- Port A write enable input
DIA(0)   => data_write_a(12),        -- Port A data input
DOA(0)   => data_read_a_lo_512(12),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(1),               -- Port B write enable input
DIB(0)   => data_write_b(12),        -- Port B data input
DOB(0)   => data_read_b_lo_512(12),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_13_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10110A0441812402840402822007818000E00700000000330A3000000008042",
INIT_01 => X"A1400984B830C848180260000C0042604001000008220008A200100802110200",
INIT_02 => X"10A00860009141100000C6180C285035000E0800010431004908135980120C60",
INIT_03 => X"004E20441910221B06420C85D5013804060000000040324C441A108468024842",
INIT_04 => X"0184034010250089C00EA8021938325B04800002091090014880080200000900",
INIT_05 => X"18002424B008881024A8004E01040104270004E0000080090500604840000481",
INIT_06 => X"80004414022A2490B00A142C8C840005794540015E006810001C4B01032C7E20",
INIT_07 => X"510200028028004880280A808816002101022468000011F082040A264006C000",
INIT_08 => X"D2B00402B220104B531001000008001041080200B660E30B200C8040080A9206",
INIT_09 => X"A1000809A93484D21000000000000080C90391881000145B0111A30404015000",
INIT_0A => X"000000008010102A82014100101118BA4510008241480290882400900000A000",
INIT_0B => X"0284484000000000400000000040000000000000040000000000000020000000",
INIT_0C => X"A944AA2000A02000212800020000000D80004084A0000390002E001843210400",
INIT_0D => X"859C1881A04090000000000021800180010341179065441356150A1285094284",
INIT_0E => X"859C188810C65A72A617520252781EA02520D589B9A260859C1840DD81B9A0E0",
INIT_0F => X"0E71F1052D942748C19484E39442D15961C0DD81B9A260859C1840D589B9A0E0",
INIT_10 => X"E60605C0C12CBD400B0810C65A61AA459D0047398500D5889D26907356533C00",
INIT_11 => X"8F60CA1562094650CA28398A42C051E0332181010109294C8E1160CB8C80A561",
INIT_12 => X"2645056D073148580A3C065141942AC4128CA199180C5232575138094450AD0A",
INIT_13 => X"84CA93A2FC008962142B17301A9A1A5196A80245208E0AC5C853C8028163B8C0",
INIT_14 => X"0240034000E4DC8A84000014982372011FC1E475F0F0084A3961F5A80AC5C816",
INIT_15 => X"4250942509425094250942509428D421420882020120981812C8403000088212",
INIT_16 => X"2509425094250942509425094250942509425094250942509425094250942509",
INIT_17 => X"5094250942509425094250942509425094250942509425094250942509425094",
INIT_18 => X"FF3F7DF7FF3E9F7DF7E24502A800000000000000000050942509425094250942",
INIT_19 => X"EBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBF7DFDFDDD555555F7EFBBEE",
INIT_1A => X"7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAEBAEBAEBAEBA",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000000007F7EBF5FAFD7EBF5FAFD7EBF5FAFD",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5554BA087FFFF55557BD54AAF7FBC01FFA2802ABEF0000000000000000000000",
INIT_22 => X"2E80155AA802AB45AA843FE0008557DFFF0800020105D557FEAA00557DE10AAD",
INIT_23 => X"8557DF45002ABDFFFF7803DE10AA80000AA087BD75EF087FFFFEF557BEAB4555",
INIT_24 => X"F7AA80000AAD1420AA087BD7555FFD168AAAFFAE820AA5D5557555082ABDF550",
INIT_25 => X"5FFD157555085140010F7AEAABFFAAD5420000051555FFA2AA8200000557DFFF",
INIT_26 => X"45007FC2155F7D155545AA80001EFAAFBEAB45557FFDE10AAAEA8BFFA2FBD754",
INIT_27 => X"E00082AA8AAAAAFFC00BA00002AAAAF7D5574BA557BE8A10A284154BAFFAAAAB",
INIT_28 => X"0000000000000000000000000000000000000000A2D155410F7FFFFEBA08003F",
INIT_29 => X"7AE921C517DE10A2DB50482147FFAF554971D0492E3F1C71C7BE8A2ABD700000",
INIT_2A => X"FFAFD7497BE8B5555208217DBE8A2AB45BE803AE38145B78FD7000005010495B",
INIT_2B => X"5F5056D002EBDF6D005B78F7D142ABDFC7F78E3FE28B684070AA1C71D25D7007",
INIT_2C => X"6A487000005F7AFD7F7A482038AADF47092147FD257DFFD568A82FFA4870BA55",
INIT_2D => X"A2A0ADBC7A2FFD257DE3DF52555085142000FFAAAFBFFBED547038145B505FFB",
INIT_2E => X"0B680124BAFFAAAFB45007BC217DEBDB55555AA8E071D7AAFBEFB455D71F8E00",
INIT_2F => X"28FFF1FDE821C003FE001C2EAAAAAB6F5C20821C002AA92FFDF574824171EAA1",
INIT_30 => X"545F7AEA8B55000000000000000000000000000000000000000000000B6D5504",
INIT_31 => X"AB45080015410007FEAA0055517DE00A2FFC00105D7BE8B55085142010AAD157",
INIT_32 => X"154BA5D5140145007BE8B55087BEAB555D04001EFF7AAA8B55F7802AABA5D7FE",
INIT_33 => X"16AA10FF80174AA557FC21EF082EBFFEF007BE8BFF5D2ABDF55F7AABDEAAF784",
INIT_34 => X"D1554BA5D7BC01FFFF8015410007FEAB45F780020BAA2FFD54105D7FC21EFFFD",
INIT_35 => X"2FBFDF455D556AA00A2803FF45AAFFC21EFAAFBC0155085540000FFAEBFFEFF7",
INIT_36 => X"F7FBD5410085568A10FF80020AAFFAABFF55087FC01EFA2FFD7545AAAE97555A",
INIT_37 => X"0000000000F7D1400BAFFD57FE005D043FE10552EAAAAAFFD1400005D042AA00",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000CFFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(1),               -- Port A write enable input
DIA(0)   => data_write_a(13),        -- Port A data input
DOA(0)   => data_read_a_lo_512(13),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(1),               -- Port B write enable input
DIB(0)   => data_write_b(13),        -- Port B data input
DOB(0)   => data_read_b_lo_512(13),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_14_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10020A000180000284008280000281800000030000000033022000000580002",
INIT_01 => X"A140098018300848184860000C20C24040000000084000084200000000110200",
INIT_02 => X"1020006000900110000006102028503400040800010400204908012018120E64",
INIT_03 => X"000200441910221006420000400100040600000000E9E401209A108448004842",
INIT_04 => X"0004020000250008000200021038000804000000090090004800080200000000",
INIT_05 => X"500024240008881024A800400104010420000400000080080100204040000000",
INIT_06 => X"8000440102282015B10A10288E0400042345400040006810000C5901033D7880",
INIT_07 => X"1100000200280048802008828812002001220064000005F1C2850A2649204070",
INIT_08 => X"00B00402802010411110010000080010010802000400230B000C804008080002",
INIT_09 => X"01000009A92480001000000000000080C8038188100004590111B68404010000",
INIT_0A => X"0000000080101000000141001001088A45000082400000008020009000008000",
INIT_0B => X"0004404000000000400004000000000000004000000000000004000000000000",
INIT_0C => X"8904A0200080200001080002000000088000400420000200002E000841010400",
INIT_0D => X"0500000C80409000000000000000018000000000806044010014081204090204",
INIT_0E => X"0500005813A0210D072E8D012001028402908004000587050000108004000707",
INIT_0F => X"9004300044900812386A280E5800088980108020000587050000108020000707",
INIT_10 => X"DE00482E19E30002007813A02096038AE200880405200308828062A68C0BC700",
INIT_11 => X"00000E5A08E6000048001292B83280001208A1011004011060049A1C59192055",
INIT_12 => X"492060480256530650000240001DB011CC00009000032C4C979E3806180C0900",
INIT_13 => X"5A3433EDE00154181400000007BCBD858F120120541A0000000033757465B2C0",
INIT_14 => X"02002C000024008A84001A0902000422E3E99681004802115652594000000001",
INIT_15 => X"0240902409024090240902409028D021020880000120901812C8401000000210",
INIT_16 => X"2409024090240902409024090240902409024090240902409024090240902409",
INIT_17 => X"4090240902409024090240902409024090240902409024090240902409024090",
INIT_18 => X"5C8FF0F7BE9D5F7DF65040028000000000000000000040902409024090240902",
INIT_19 => X"79E79E79E79E79E79E79E79E79E79E79E79E79E7BF7DDDDDFCF3CF3DF5579B4E",
INIT_1A => X"3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE79E79E79E79E",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000003FF803F9FCFE7F3F9FCFE7F3F9FCFE7F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"BE8B55A2AE80000F7D5555555D2AAAABAAAD1420BA0000000000000000000000",
INIT_22 => X"00155EF0804155EFAAD5554BA087FFFF55557BD54AAF7FBC01FFA2802ABEFA2F",
INIT_23 => X"8557DFFF0800020105D557FEAA00557DE10A2AA801FFA28402000AAAE9554555",
INIT_24 => X"AA802AB4500516AA00A2AE800BAFFFFC20BAF7AEA8B45080417400AA843FE000",
INIT_25 => X"0A2843FEBAFFFBD7410A2D168BFF087BD75EF087FFFFEF557BEAB45552E80155",
INIT_26 => X"AA082ABDF5508557DF45002ABDFFFF7803DE10AA80000AA005568ABAA2840201",
INIT_27 => X"AAAFFAE820AA5D5557555002E80155A280000005D7FFDF4555517DFEF00043FE",
INIT_28 => X"0000000000000000000000000000000000000000AAD1420AA087BD7555FFD168",
INIT_29 => X"C71C7BE8A2ABD7A2FFEDB55B6A080038E3DB50555412AA8ABAAADB4009200000",
INIT_2A => X"402038AAAA955554900105FF0800175D7A2DB50482147FFAF554971D0492E3F1",
INIT_2B => X"0A12410BE803AE38145B78FD7000005010495B7AE921C517DE10A2AE851FFB68",
INIT_2C => X"97BE8B5555208217DBE8A2AB451C556FA00A2A0800BAE3F1C0092EBAAADB6D08",
INIT_2D => X"00516DABAA28402038B6803DE82F7F5D5410A2D568BC71C71D25D7007FFAFD74",
INIT_2E => X"55D5F78FD7000E3FEAA002EBDF6D005B78F7D142ABDFC7F78E3FE28B684070AA",
INIT_2F => X"92147FD257DFFD568A82FFA4870BA555F5056D002A80155B680000105D7FF8F4",
INIT_30 => X"AAAAAFFC2000000000000000000000000000000000000000000000000AADF470",
INIT_31 => X"8B55085142010AAD157545F7AEA8B55A2FBFFF55FF84000AAAAFBC0145002AA8",
INIT_32 => X"7DE00A2AA955FFFF80020BAAAAA975450800001EF080417555A2FFC00105D7BE",
INIT_33 => X"140000A2AEBFFEF082A82010F7802AABA5D7FEAB45080015410007FEAA005551",
INIT_34 => X"5140145007BE8B55087BEAB555D04001EFF7AAA8B555D557FE00A280020BAAAD",
INIT_35 => X"7AABDEAAF784154BA08557FEAAA284000AAFF803DE00FFD557400AAD56AB455D",
INIT_36 => X"F780020105D7BEAB45557BE8B45082EBFEBA082EBFFEF007BE8BFF5D2ABDF55F",
INIT_37 => X"0000000000A2FFD54105D7FC21EFFFD16AA10FF80174AA557FC21EF082A80145",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000000FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(1),               -- Port A write enable input
DIA(0)   => data_write_a(14),        -- Port A data input
DOA(0)   => data_read_a_lo_512(14),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(1),               -- Port B write enable input
DIB(0)   => data_write_b(14),        -- Port B data input
DOB(0)   => data_read_b_lo_512(14),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_15_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000A000000000284000280000001800020030000000033022000000180002",
INIT_01 => X"A140098018300848180060000C00424040000000080000080200000000110200",
INIT_02 => X"102100400C8011100000061000A8503401044880010430004808000180122378",
INIT_03 => X"000200541D102210064200000045000546080000400020000008108448400042",
INIT_04 => X"8094020000254C880000028A1018000844000000880013504000002600000000",
INIT_05 => X"10002424000AA81024A82040010C61062001440002988000000024808001004B",
INIT_06 => X"80004400022A00003C8912248E0400042854400040006810000C4901032B1800",
INIT_07 => X"50200000B0280048A0280A828801002101020040000005F38204082640000000",
INIT_08 => X"01F00402802610411100110000000010010802000400230A0008884008080004",
INIT_09 => X"01000001A12481041000000000000080C0030108100004590111820404000000",
INIT_0A => X"0000000080101000004140001001088A45000082000000008000001080008000",
INIT_0B => X"0004404000000000400004000040000400000000000000000004000020000200",
INIT_0C => X"0804000020024100012808020000000981004004A0200310000C000800000000",
INIT_0D => X"0000001180009000000000002100018000000000004004010010000000000000",
INIT_0E => X"00000008000002000000000000000000000080A40000000000000080A4000000",
INIT_0F => X"00000000001000204800000000000000000080A40000000000000080A4000000",
INIT_10 => X"000000000000000000080000020000000000000000000008000C020000000000",
INIT_11 => X"000000824000000000000020220000000001800100020300000004003420480A",
INIT_12 => X"0000000000040440000000000001048000000000000000100800400000000000",
INIT_13 => X"000800000000000000000000000100C220050000000000000000008220884400",
INIT_14 => X"000000000000000830000000000000000016101C5C1400000000000000000000",
INIT_15 => X"0000000000000000000000000020C00000088000012090101280401000000200",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000040028000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"000010082A954BA00003DFEF085155400F78428BEF0000000000000000000000",
INIT_22 => X"8015400FF84001EFA2FBE8B55A2AE80000F7D5555555D2AAAABAAAD1420BAFF8",
INIT_23 => X"87FFFF55557BD54AAF7FBC01FFA2802ABEFF7AE95555A2FBE8BEFA2843DE00AA",
INIT_24 => X"0804155EFFFFBE8BFF0800174AA557BFDE10A2FBEAB45F7D56AABAAAD5554BA0",
INIT_25 => X"5FFD568BEF087FE8A1055003FE00A2AA801FFA28402000AAAE955455500155EF",
INIT_26 => X"45AA843FE0008557DFFF0800020105D557FEAA00557DE10F7D1574AAA2D16AB5",
INIT_27 => X"0BAF7AEA8B45080417400FFFFC2145080015400AA802AA00AAAE800BA5D00155",
INIT_28 => X"000000000000000000000000000000000000000000516AA00A2AE800BAFFFFC2",
INIT_29 => X"A8ABAAADB40092E38E070280024904AA1C0438FD7005150438F78A2DBFF00000",
INIT_2A => X"FE8BC7BE8E38E10A28017400E38A051FFA2FFEDB55B6A080038E3DB50555412A",
INIT_2B => X"D16AABAA2DB50482147FFAF554971D0492E3F1C71C7BE8A2ABD7E3AA9257DA2F",
INIT_2C => X"AAA955554900105FF0800175D7E3FFEFBD70000124AA557FFDE10A2FBEDB6DF7",
INIT_2D => X"FFDF50482A2DB6AB45FFD56DBD7087BEAA38410038E38A2AE851FFB68402038A",
INIT_2E => X"0AAA085082550A1057DBE803AE38145B78FD7000005010495B7AE921C517DE10",
INIT_2F => X"00A2A0800BAE3F1C0092EBAAADB6D080A12410FFF1C017D140410400BE8E28A1",
INIT_30 => X"0AAF7AEBDFEF0000000000000000000000000000000000000000000001C556FA",
INIT_31 => X"00AAAAFBC0145002AA8AAAAAFFC2000AAAA974AA0800020BA550028B55085540",
INIT_32 => X"A8B55AAAE821EFAAFBEAB55F7AAA8A00AA8417400AAAE975EFA2FBFFF55FF840",
INIT_33 => X"BFFE10A2FFFFFEFF7D568ABAA2FFC00105D7BE8B55085142010AAD157545F7AE",
INIT_34 => X"AA955FFFF80020BAAAAA975450800001EF080417555AAFFFDF450804020AA557",
INIT_35 => X"07FEAA0055517DE00FFFBC2000AAFBE8B55F7D17DF45007FE8AAA08002AAAAA2",
INIT_36 => X"5D0000010F7AAA8A10AA8017400552A801EFF7802AABA5D7FEAB450800154100",
INIT_37 => X"00000000005D557FE00A280020BAAAD140000A2AEBFFEF082A82010FFD5421EF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000C00000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(1),               -- Port A write enable input
DIA(0)   => data_write_a(15),        -- Port A data input
DOA(0)   => data_read_a_lo_512(15),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(1),               -- Port B write enable input
DIB(0)   => data_write_b(15),        -- Port B data input
DOB(0)   => data_read_b_lo_512(15),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_16_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"DA22C618B1000482B688B186588884862A400438255FC38381441205BA803003",
INIT_01 => X"264AC80028404C211203A952A90341080B173340412000E1005D628000820484",
INIT_02 => X"400034C206C405000001A48202084004003008255040826EE008B440200E2042",
INIT_03 => X"A459C1240181AB20AD27315B7F1983CA1C900040422A005762010010000C0400",
INIT_04 => X"296E542B6E3A825C15FB385321B4ADFE16AB45FD2C400002E205231201290A28",
INIT_05 => X"B9E5815006028179808C00A0D2152B90707A1E0BD423CAC0000D610000000710",
INIT_06 => X"81F104A1415C292164280081C6AB88742086ACACDE240000A80090CE82A803B9",
INIT_07 => X"400800000ACCAA280940580400A37B8896CA4D000A80C1102A00001C14028009",
INIT_08 => X"0015452880C8D90409A02D965965200100104F2B00822512000000231520A024",
INIT_09 => X"A5AA80018120E00066000000000012C9000A0000D0A80000BF8028E87C1B9927",
INIT_0A => X"00520228080108039501200848002912300208092B940192D1000000000000A8",
INIT_0B => X"03561180063DB4F6110001100011000110001100011000110001080008800080",
INIT_0C => X"080200854409418B02ED0000502A02972000040BB401100010012B4C90000100",
INIT_0D => X"6D061A1F8D60D80820500101244AA8A2AA242E80000009200120000000000000",
INIT_0E => X"6D066210E5001DB4A5B400C7D553847165A99000C6564CDD051DC99000C65555",
INIT_0F => X"21D0C48F254946148107354292673D1F72C99000C6564CDD0565C99000C65555",
INIT_10 => X"952D2058F33225787810F5001D6121A9559224D1FF97D0272F04D89441A56D8A",
INIT_11 => X"6C1C74485B81E31306C71D1093AB8A64811BADC00992180D58033B1172F2A025",
INIT_12 => X"7B86DED8E3A212748F0E0CA638E890B7A8546120C0AFF5B548AC431FB1C7DB07",
INIT_13 => X"EFCE9B26DECA1AD36A2E4F40DF6AAAF260AF88899E8B8B93D12A877178DD0032",
INIT_14 => X"A8009F8B108C80A1021B9A8BB8056662CA1951596800FC01A38D4D4B072B922F",
INIT_15 => X"00000000000000000000000000044000102A0001148442A1108103595580A840",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"4C690DA64C1C4F68A36040000000000000000000000000000000000000000000",
INIT_19 => X"D14D14D14D14D14D14D14D14D14514514514514529E5F87869E79E78558D1154",
INIT_1A => X"3D1E8F47A7D3E9F4FA7D3E9F4FA7D3E9F47A7D1E9F47A7D1E9F4D14D14D14D14",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE000000000000000007D3E9F4FA7D3E8F47A3D1E8F47A",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFEFF7D168B55AAD17FFFF552EBFE00007FC00AA0000000000000000000000",
INIT_22 => X"04000BA552A821FFFF8000010082A954BA00003DFEF085155400F78428BEF087",
INIT_23 => X"2AE80000F7D5555555D2AAAABAAAD1420BA5D2E975EFF7D568BFFFF80175EF00",
INIT_24 => X"FF84001EF0000020AA5D00154005D043FF45555540000082EAABFFA2FBE8B55A",
INIT_25 => X"0087FD74BAAAAEBFFEF557FC00AAF7AE95555A2FBE8BEFA2843DE00AA8015400",
INIT_26 => X"FFAAD5554BA087FFFF55557BD54AAF7FBC01FFA2802ABEF557BEABEF5D041541",
INIT_27 => X"E10A2FBEAB45F7D56AABA082A97545F7D16ABFFFFAABFEAAFF84001FF002A821",
INIT_28 => X"0000000000000000000000000000000000000000FFFBE8BFF0800174AA557BFD",
INIT_29 => X"50438F78A2DBFF0871F8FC7E3D56AB6DBEDB7FFEF552AB8E38087FC209200000",
INIT_2A => X"16ABFFE38E175EF1400000BA412E871FFE38E070280024904AA1C0438FD70051",
INIT_2B => X"2EAFBD7A2FFEDB55B6A080038E3DB50555412AA8ABAAADB400924920925EFF7D",
INIT_2C => X"E8E38E10A28017400E38A051FF0804050BA410A1240055003FF6D5551420101C",
INIT_2D => X"4975EDBC7550E12410087FD74AAB6AABFFC7557FC00BAE3AA9257DA2FFE8BC7B",
INIT_2E => X"AF780051C70824851D7A2DB50482147FFAF554971D0492E3F1C71C7BE8A2ABD7",
INIT_2F => X"D70000124AA557FFDE10A2FBEDB6DF7D16AABA08249756DF7D168BC7F7AABAEA",
INIT_30 => X"AAA007BC0000000000000000000000000000000000000000000000000E3FFEFB",
INIT_31 => X"20BA550028B550855400AAF7AEBDFEF08516AB55A2D16ABEFFFFBFDFFF552AAA",
INIT_32 => X"C20000000021EFF7D568BFFA2AA955FF5D04020AA002A955EFAAAA974AA08000",
INIT_33 => X"03DFEF5D51420005D2ABFF45A2FBFFF55FF84000AAAAFBC0145002AA8AAAAAFF",
INIT_34 => X"AE821EFAAFBEAB55F7AAA8A00AA8417400AAAE975EF0800174BA002E820105D0",
INIT_35 => X"AD157545F7AEA8B5500557DF45552A82000007BD74AAF7AEBDF455D7BC20BAAA",
INIT_36 => X"F7D568B55FFAAAAABAFF8415545000015555A2FFC00105D7BE8B55085142010A",
INIT_37 => X"0000000000AAFFFDF450804020AA557BFFE10A2FFFFFEFF7D568ABA0804155FF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000400000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(2),               -- Port A write enable input
DIA(0)   => data_write_a(16),        -- Port A data input
DOA(0)   => data_read_a_lo_512(16),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(2),               -- Port B write enable input
DIB(0)   => data_write_b(16),        -- Port B data input
DOB(0)   => data_read_b_lo_512(16),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_17_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"5284CE4FB7BD2C8994A13392DBD02E14006B82AC7E800D44D3DD2FD5F9B961C0",
INIT_01 => X"F9BA301F7E03FC6793F2199B39FC233C11D93AE6F3BB92B32091DBC339B24542",
INIT_02 => X"1D5FC0C08F040404446965C0607FB8A217C400C33A908078551BD04222186338",
INIT_03 => X"8504930A37F65820CB24111B7F08014A0AB84A52B6D2AFF97C1B5AC757F06D6B",
INIT_04 => X"250834336D1E81500FDB38302292ADFE103B6DBD204037F202042075E2B1D00A",
INIT_05 => X"8F039786062C6CE092F5FE005236781C402A0807B4070670083DC68206D7E6D0",
INIT_06 => X"0CD26803C3582408962C58B183F8AEF42045919B30E085DD2ED57D4EED08CA6A",
INIT_07 => X"700000B30380670B8142500448E3E01E94EF1340A28AC1AC8156044D1400AA00",
INIT_08 => X"009F3A1B0120A1C51DFFC40C30E5F0182D0950190C0810BE00E9A76E4C6FFBE4",
INIT_09 => X"8FCCC200A59BDD2FFE3F3EC7C7DEF207000F00059D2ED56D7EED2ED3C9A867DC",
INIT_0A => X"0617112E46F05D02DD814102F800633F1D0A7CC9AE7A08BFF0001D35682AC0CE",
INIT_0B => X"8A3F06ABD73DBCF4FBCF4FBCF4FBCF4FBCF4FBCF4FBCF4FBCF4FBE7A7DE7A780",
INIT_0C => X"001000974F08518F5AFFC94B533FADA7FDE97D6BFF329E1B50FF99F086000D9E",
INIT_0D => X"F50B018F95EA3DED1652EC0B27E67F419E2E1E8000C0036340B8000000000000",
INIT_0E => X"F50B01C8DF7F96197DB4AFC8C8886AF672A1537F759299F50B03C1537F759199",
INIT_0F => X"6068331C5103E7EF0FBEED6BB6A9412007C1537F759299F50B03C1537F759199",
INIT_10 => X"21F2CD7F252CDABB3CE8CF7F963AB9FD6AD434201AA68B837FFD1F7B7125B68C",
INIT_11 => X"BD055EB6D555CB2949C15BA7270FF256526BBFD55BBE71D79F73C7AC6DB9BF37",
INIT_12 => X"94080BF82B74E4E1FE4ACA4E0ABD6DAAAB965293036FF6B652A99A6026027FBE",
INIT_13 => X"EF5CBA7A43482800FEFAFD06B8CFCCAB7550D0C2022EAEBD438697AD2EBA9168",
INIT_14 => X"AC00A8BBFC8B501CF7A0FED9A548FA19752C4A4EADAE42FCBC38C3B7BEBF42CF",
INIT_15 => X"0000000000000000000000000026E100002F382DBD9ECFE117805F20CFDAAB00",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"09EDCC4052E917114F981800C000000000000000000000000000000000000000",
INIT_19 => X"EBA69AEBA69A69AEBA69AEBA69A69A69A69A69A68698686981D75D7443720030",
INIT_1A => X"46A351A8D068341A0D068341A0D068341A0D46A341A0D46A341A69AEBA69A69A",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000000000046A351A8D46A351A8D46A351A8D",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFEFF7FBEAB450804001EFAAD57FEAA0000000000000000000000",
INIT_22 => X"51401EF087FD74AA087FFFFEFF7D168B55AAD17FFFF552EBFE00007FC00AA087",
INIT_23 => X"82A954BA00003DFEF085155400F78428BEFAAD168A000004020AA5D7BE8B4500",
INIT_24 => X"552A821FF5D00020BA552A82000552A821555D7FEAB55FF80175EFFF80000100",
INIT_25 => X"FAAFBC01EF5D0015555557BFDEBA5D2E975EFF7D568BFFFF80175EF0004000BA",
INIT_26 => X"BAA2FBE8B55A2AE80000F7D5555555D2AAAABAAAD1420BAFFFFFDF45AAD17FFF",
INIT_27 => X"F45555540000082EAABFF00516AA10552E820BA007FEABEF005555555A2D1554",
INIT_28 => X"00000000000000000000000000000000000000000000020AA5D00154005D043F",
INIT_29 => X"B8E38087FC2092147FFFFFFFFFBFDFC7EBF5E8B550000071EFB6DF7AE9200000",
INIT_2A => X"A07082497FEFB6D1451471EF007BD04920871F8FC7E3D56AB6DBEDB7FFEF552A",
INIT_2B => X"8E175FFE38E070280024904AA1C0438FD7005150438F78A2DBFFBED16AA381C0",
INIT_2C => X"38E175EF1400000BA412E871FF550A00092492A850105D2A80155417BEFB6DEB",
INIT_2D => X"FFF5FFF6DAADF7FFD7B6F1C71EF55001756D5D7BFAEBA4920925EFF7D16ABFFE",
INIT_2E => X"700515556DA2DF50492A2FFEDB55B6A080038E3DB50555412AA8ABAAADB40092",
INIT_2F => X"BA410A1240055003FF6D5551420101C2EAFBD7145B6AA28492487082007FEDBD",
INIT_30 => X"5EFFFFBEAA000000000000000000000000000000000000000000000000804050",
INIT_31 => X"ABEFFFFBFDFFF552AAAAAA007BC0000557FFDFEFF7FBFFF55A2D16AB55000017",
INIT_32 => X"BDFEFF7D568AAA5D2A97410007BFFFFF5551555EF087FC200008516AB55A2D16",
INIT_33 => X"A82155087FFFFEFAAAA975EFAAAA974AA0800020BA550028B550855400AAF7AE",
INIT_34 => X"00021EFF7D568BFFA2AA955FF5D04020AA002A955EF5D2E80010002A954005D2",
INIT_35 => X"02AA8AAAAAFFC2000FFD57DFFFAAFFFDF55FFD1575FF5504175EF5D7FEAAAA00",
INIT_36 => X"000415410007BFFF450051555EFA2FBC0000A2FBFFF55FF84000AAAAFBC01450",
INIT_37 => X"00000000000800174BA002E820105D003DFEF5D51420005D2ABFF45557FE8AAA",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000CFFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(2),               -- Port A write enable input
DIA(0)   => data_write_a(17),        -- Port A data input
DOA(0)   => data_read_a_lo_512(17),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(2),               -- Port B write enable input
DIB(0)   => data_write_b(17),        -- Port B data input
DOB(0)   => data_read_b_lo_512(17),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_18_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"69844019080000A21A611406840014122A641074155FC28A2024001001801003",
INIT_01 => X"01067920034004180005E9E3C90360C0041C0181002001602025800008440084",
INIT_02 => X"40AC3CAA22D605200000856E2481902400344A20F802C22054001000021E2379",
INIT_03 => X"A54C23B34C81EB2076471000800981140C010101750D1007E58040102B0E0100",
INIT_04 => X"22660C1C0065003C04040013236E105016A028402D618803EB092B9201490B2A",
INIT_05 => X"B8E080000000005889AC41E04508A99070200E010001C1CA11803850C8000100",
INIT_06 => X"800A4CE301545001F40050216C09950004C2047BCF1C8090C02800C0120886B3",
INIT_07 => X"814A0080064C1F300020080182001A9E02C03400082002700000217294007101",
INIT_08 => X"000117088080990419002D86184A01018030430700802541420440022030041A",
INIT_09 => X"7030C30B885200D274004008080003C32A10A19090C02010E102294406168800",
INIT_0A => X"00602A01880980037109700C04C44C92A88DCC2211E44174112840880000060D",
INIT_0B => X"11C0D95C20C2030A003080030800308003080030800308003080018400184004",
INIT_0C => X"8304E02809832E6021002020404042000F00008400811824AD4007ECD9436261",
INIT_0D => X"0AFCE5D22A82B20000520100C801F8A07E103000A1285C84000418360C1B060D",
INIT_0E => X"0AFCFD8CB17E5B4F045557575E6EFBE3942C1040A41D660AFCE1CC1040A41E66",
INIT_0F => X"8E7FFBB385661C08D1455ABA91E6FF5FDFCC1040A41D660AFCF9CC1040A41E66",
INIT_10 => X"015F82C006C3AF31E64CB17E5A9655017F1FC73FAF1D61B1040294C58AD1FF5F",
INIT_11 => X"B95454005BAA36DCF8E519001BF80DEB3EE2020EA678189C6EC32881F7F75648",
INIT_12 => X"67D7EDFCA320037E81BD77D728A800B7546DBDFF12904747A351145FC53ABF8D",
INIT_13 => X"92B764225C57C97EBE76E1254F0C0D4514A84F5573FE9DBA4A38E247C522CC0E",
INIT_14 => X"BE84370001B6922070440556B15F7FABBC40151D7C747D8220673C3B9DB84B20",
INIT_15 => X"06C1B06C1B06C1B06C1B06C1B0491069068000004060300A005A01183F240014",
INIT_16 => X"6C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B",
INIT_17 => X"C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B0",
INIT_18 => X"B80EE173C2300F7DF16000000000000000000000000041B06C1B06C1B06C1B06",
INIT_19 => X"AAAAAA28A28A28AAAAAAA28A28A28A28A28A28A2910591505C104104B28BBECE",
INIT_1A => X"128944A25128944A25128944A25128944A2552A954AA5128944AAAA28A28A28A",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000128944A25128944A25128944A25",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFDFEF5D2A974BA082E954000000000000000000000000",
INIT_22 => X"0028B55002E82000087FFFFFFFFFFFFFEFF7FBEAB450804001EFAAD57FEAA087",
INIT_23 => X"7D168B55AAD17FFFF552EBFE00007FC00AA087FFFFFFFFFBFDF45AAD568B5508",
INIT_24 => X"087FD74AAAAFFFDF45A2D16AB55F7FFFFFFF00043DE10AA843DE00087FFFFEFF",
INIT_25 => X"A55042ABEF5D7FD75FFAAD540145AAD168A000004020AA5D7BE8B450051401EF",
INIT_26 => X"45FF8000010082A954BA00003DFEF085155400F78428BEFAA80000000804154B",
INIT_27 => X"1555D7FEAB55FF80175EF5D00020105D2A97400082E95555085168A10557FD75",
INIT_28 => X"00000000000000000000000000000000000000005D00020BA552A82000552A82",
INIT_29 => X"071EFB6DF7AE921C7FFFFFFFFFFFFFFFF7FBFDFFF5D2A954AA082A9242800000",
INIT_2A => X"1FAF55A2DF6DB7D1C002AB7D002A82028147FFFFFFFFFBFDFC7EBF5E8B550000",
INIT_2B => X"8E38E280871F8FC7E3D56AB6DBEDB7FFEF552AB8E38087FC2092087FFDFC7E3F",
INIT_2C => X"97FEFB6D1451471EF007BD0492B6F1F8F55AADF6DB7DE3F5FAFC708003DE28B6",
INIT_2D => X"A28407038140410492550A2ABC7497BD25FFAADF4516DBED16AA381C0A070824",
INIT_2E => X"D1C516FA28417BD5545E38E070280024904AA1C0438FD7005150438F78A2DBFF",
INIT_2F => X"92492A850105D2A80155417BEFB6DEB8E175FF5D0E05000492097428002E9557",
INIT_30 => X"4AA082A820AA000000000000000000000000000000000000000000000550A000",
INIT_31 => X"FF55A2D16AB550000175EFFFFBEAA00557FFFFFFFFFFFDFEFF7FBFFFEF552E97",
INIT_32 => X"C0000087BFDF45AAD568B55AAFBFDFEF55042ABEF002A800AA557FFDFEFF7FBF",
INIT_33 => X"16AB4500043DEAAFFAEAAAAA08516AB55A2D16ABEFFFFBFDFFF552AAAAAA007B",
INIT_34 => X"D568AAA5D2A97410007BFFFFF5551555EF087FC2000FFD56AB45A2FFFDFFFAAD",
INIT_35 => X"855400AAF7AEBDFEFA280154BA550400000552AA8B45087FC01EFA2FFD55EFF7",
INIT_36 => X"0804154BA082A975EF5D517DEAA007BD5545AAAA974AA0800020BA550028B550",
INIT_37 => X"00000000005D2E80010002A954005D2A82155087FFFFEFAAAA975EF5D2E97400",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000400000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(2),               -- Port A write enable input
DIA(0)   => data_write_a(18),        -- Port A data input
DOA(0)   => data_read_a_lo_512(18),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(2),               -- Port B write enable input
DIB(0)   => data_write_b(18),        -- Port B data input
DOB(0)   => data_read_b_lo_512(18),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_19_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"042200000000000041088001001AA00000000000000000000000500802000003",
INIT_01 => X"074018000024000000000404000000000A22000800000800004A200000000001",
INIT_02 => X"0000048002C405000000000006A84000000000200893C246A20000000020031A",
INIT_03 => X"082A58E411004B2000071000000981000C000000002045000200000000000000",
INIT_04 => X"200604000000001C0400001320000000162000002C4000026201201200090800",
INIT_05 => X"1020800000000058840200204000099070200E010001C0400000000000000000",
INIT_06 => X"0012048037805421402850001402498820022802400480405008901100A00102",
INIT_07 => X"00000000020C0130481204919200010C82000000000006002A548902A0020109",
INIT_08 => X"0001150800009900000005861840000000004301000B000000000001C1C00000",
INIT_09 => X"001F00002024B20002000000000002C300000000405000103010204000000000",
INIT_0A => X"00000000000000000000000000000040002000044000000000000000000002F0",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000420003B00000000000000000040012C80000000",
INIT_0D => X"45001A03C0825A0D20800000000018A006001000000000000000000000000000",
INIT_0E => X"450002131E01A1F6EA0A0020211146E069C2ACC01AE80045001D82ACC01AE800",
INIT_0F => X"1188340C3E1CFAD27CC2E004481020892282ACC01AE80045000582ACC01AE800",
INIT_10 => X"DEA03228D810007019931E01A1E5BA02802008C06F029D4C7B76639CEC0A0020",
INIT_11 => X"428AA3592000000206C2A4DAC00000008113C246A181C03FE4662A84575768DF",
INIT_12 => X"08201090549B5800000000261546B24000000000C53807E7CC06618018C51210",
INIT_13 => X"13F6A185A0A0168128411ACB800C0E108A0720288C011046B5986247C5452291",
INIT_14 => X"0000C220010808C10D9A92A74CD7CF4A080031B1515B212143D841431046B58A",
INIT_15 => X"00000000000000000000000000000000000000000000000000000118030004E0",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"3F0C7010C660C744192000000000000000000000000000000000000000000000",
INIT_19 => X"1861861861869A61861861861861861861861861A8208C4C1534D34C07208BBA",
INIT_1A => X"0984C26130984C26130984C26130984D26930984C26130984C261861861869A6",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE000000000000000000984C26130984C26130984C2613",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF552A974AA0004174BA0000000000000000000000",
INIT_22 => X"2E974BAA2FFFFE10087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974BA082E95400F7F",
INIT_23 => X"FFFFFFEFF7FBEAB450804001EFAAD57FEAAF7FFFFFFFFFFFFFFFFF7FBFDFFF55",
INIT_24 => X"002E82000F7FFFFFFFFFFFFDFEFA2D568B550004001EFAAAEA8ABA087FFFFFFF",
INIT_25 => X"5AAD16ABEF5D2ABFF55080402010087FFFFFFFFFBFDF45AAD568B55080028B55",
INIT_26 => X"BA087FFFFEFF7D168B55AAD17FFFF552EBFE00007FC00AAF7FFFFFFFF7FBE8B5",
INIT_27 => X"FFF00043DE10AA843DE00557FFDFEFA2D16AB55A2FFFDFEF5D2EBFE00AAFFFFE",
INIT_28 => X"0000000000000000000000000000000000000000AAFFFDF45A2D16AB55F7FFFF",
INIT_29 => X"954AA082A92428E3FFFFFFFFFFFFFFFFFFFFFFFEF552A974AA0000104AA00000",
INIT_2A => X"FFDFEFF7F5FAFC7492A974AAB6F5F8E101C7FFFFFFFFFFFFFFFF7FBFDFFF5D2A",
INIT_2B => X"A4A8AAA147FFFFFFFFFBFDFC7EBF5E8B550000071EFB6DF7AE92EBFFFFFFFFFF",
INIT_2C => X"2DF6DB7D1C002AB7D002A82028FFFFFFFEFF7F1F8FD7AAD16AB450000001FFBE",
INIT_2D => X"F7FBF8FC7E3F5EAB45B6DF6FBEF5D2AB8F7D000000010087FFDFC7E3F1FAF55A",
INIT_2E => X"7412ABFE28B6F5F8E820871F8FC7E3D56AB6DBEDB7FFEF552AB8E38087FC2092",
INIT_2F => X"55AADF6DB7DE3F5FAFC708003DE28B68E38E284971F8FC7AAD56DB6DBEF5F8FD",
INIT_30 => X"4AA0004000AA000000000000000000000000000000000000000000000B6F1F8F",
INIT_31 => X"DFEFF7FBFFFEF552E974AA082A820AAA2FFFFFFFFFFFFFFFFFFFFFDFEF552E95",
INIT_32 => X"EAA00A2FFFFFFFF7FBFDFFFFFD568B55002A954AAF7D568A00557FFFFFFFFFFF",
INIT_33 => X"56AB450004001EFFF842AAAA557FFDFEFF7FBFFF55A2D16AB550000175EFFFFB",
INIT_34 => X"7BFDF45AAD568B55AAFBFDFEF55042ABEF002A800AAF7FBFDFEFF7D56AB45AAD",
INIT_35 => X"52AAAAAA007BC0000FFFBE8B55AAD168B55F7FFFFFFF552AA8BEF08040200008",
INIT_36 => X"A2D57FFFFF7D568B45002ABDEAAFFD16AA0008516AB55A2D16ABEFFFFBFDFFF5",
INIT_37 => X"0000000000FFD56AB45A2FFFDFFFAAD16AB4500043DEAAFFAEAAAAA08556AB55",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000800000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(2),               -- Port A write enable input
DIA(0)   => data_write_a(19),        -- Port A data input
DOA(0)   => data_read_a_lo_512(19),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(2),               -- Port B write enable input
DIB(0)   => data_write_b(19),        -- Port B data input
DOB(0)   => data_read_b_lo_512(19),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_20_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000003",
INIT_01 => X"A65FF80000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000048002CC070000000000000000000000002FF86100200000000220002362",
INIT_03 => X"0000000000080F6000977060009B87A03C000000000000000000000000000000",
INIT_04 => X"3F2EFC040388137C3E20C477600142019E6000003CC0000A6601601A000B0000",
INIT_05 => X"102F91D10802ABFB80000021C8010FB0F0F43E1FE867DFC04400390210000220",
INIT_06 => X"90492261000080003400000010008000004203FE400580000000803000200006",
INIT_07 => X"401000004FFDFF28C4300C0010200100004000002AA001F00000000014000000",
INIT_08 => X"0801F5780259FB00000007BEFBC010002008FF7F00000000010018A81000041C",
INIT_09 => X"00000000020000000000000000000ADF00000020000000800000802830011023",
INIT_0A => X"0000000000000200020000000000000000000000000000000200200290000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"08120000B9090A700000200000004000000400000080002000407FED80000000",
INIT_0D => X"000079804000F00000000000C01FF8A7FE003000000004008100000000000000",
INIT_0E => X"0000798201000000100000000135386000401000010000000079801000010000",
INIT_0F => X"0185C300020004000010000000000252C7801000010000000079801000010000",
INIT_10 => X"00000010C1F30F300002010000080000000000CD8A0000400400000010000000",
INIT_11 => X"008040000000000292C0080000000000A5604000000284000818505200080000",
INIT_12 => X"0015E1B00100000000001496008000000000052B000048080000000000FC3600",
INIT_13 => X"80000000000002BA280000800830300000000000B8B400000401881010000000",
INIT_14 => X"00000000020020020001000040283024E6FB8604020080000383383B00000400",
INIT_15 => X"000000000000000000000004010201001003020200000000000127DBFF004000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"038200010089120104D204002000000000000000000000000000000000000000",
INIT_19 => X"B2CB2CB2CB2CB2CB2CB2CB2CB2C30C30C30C30C306982121A1E79E79A0700030",
INIT_1A => X"432190C86432190C86432190C86432190C86432190C86432190CB2CB2CB2CB2C",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000432190C86432190C86432190C86",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA0804020100000000000000000000000",
INIT_22 => X"2E954AA000400000F7FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0004174BAFFF",
INIT_23 => X"FFFFFFFFFFFFFDFEF5D2A974BA082E95400007FFFFFFFFFFFFFFFFFFFFFFEF55",
INIT_24 => X"A2FFFFE10FFFFFFFFFFFFFFFFFFFFFBFDFFF5D2E954BA007FC00BA087FFFFFFF",
INIT_25 => X"FF7FBFFF550800020BAAAD56AAAAF7FFFFFFFFFFFFFFFFF7FBFDFFF552E974BA",
INIT_26 => X"10087FFFFFFFFFFFFFEFF7FBEAB450804001EFAAD57FEAA007FFFFFFFFFFFFFE",
INIT_27 => X"B550004001EFAAAEA8ABA5D7FFFFFFFFFFFDFEFF7D56AB450000021EFA2D57DE",
INIT_28 => X"0000000000000000000000000000000000000000F7FFFFFFFFFFFFDFEFA2D568",
INIT_29 => X"974AA0000104AAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA08000500000000",
INIT_2A => X"FFFFFFFFFBFDFEF5D2E974AA000A07000E3FFFFFFFFFFFFFFFFFFFFFFFEF552A",
INIT_2B => X"71C50BA1C7FFFFFFFFFFFFFFFF7FBFDFFF5D2A954AA082A92428087FFFFFFFFF",
INIT_2C => X"7F5FAFC7492A974AAB6F5F8E10E3FFFFFFFFFFFFFFEFF7FBFFFFF552E974AA00",
INIT_2D => X"1C7FFFFFFFFFBFDFEFE3F5F8F450004050AABEDF6FABAEBFFFFFFFFFFFFDFEFF",
INIT_2E => X"50804021FFB6D57DE28147FFFFFFFFFBFDFC7EBF5E8B550000071EFB6DF7AE92",
INIT_2F => X"EFF7F1F8FD7AAD16AB450000001FFBEA4A8AAA497FFFFFFF7FBF8FC7EBD168B4",
INIT_30 => X"4AA080017410000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFDFEF552E954AA0004000AAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A95",
INIT_32 => X"820AA087FFFFFFFFFFFFFEFF7FBFDFFF5D2A974AA002E95410A2FFFFFFFFFFFF",
INIT_33 => X"FFDFEF5D2E954AA0051554BA557FFFFFFFFFFFDFEFF7FBFFFEF552E974AA082A",
INIT_34 => X"FFFFFFFF7FBFDFFFFFD568B55002A954AAF7D568A00AAFFFFFFFFFFBFDFEFFFF",
INIT_35 => X"000175EFFFFBEAA005D7FFFFEFF7FBFDFFFAAD16AB450804174AAFFFFFFEBAA2",
INIT_36 => X"F7FFEAB45A2D568B550804001EFF7D57DEBA557FFDFEFF7FBFFF55A2D16AB550",
INIT_37 => X"0000000000F7FBFDFEFF7D56AB45AAD56AB450004001EFFF842AAAA087BFDFEF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000000FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(2),               -- Port A write enable input
DIA(0)   => data_write_a(20),        -- Port A data input
DOA(0)   => data_read_a_lo_512(20),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(2),               -- Port B write enable input
DIB(0)   => data_write_b(20),        -- Port B data input
DOB(0)   => data_read_b_lo_512(20),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_21_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"4A302428B824900A128C090A5C1800261500213C005FE812D10420054085A202",
INIT_01 => X"081FFE3440B609703B0427F801A40B8115BC4F655300340288A40D30040E4DD8",
INIT_02 => X"04CA478082CC1740002019824E0203100640303FF8C0B31061096E21A1840814",
INIT_03 => X"8C329E9204020FE002577800405B87047D5042129D8D0248903200013290C800",
INIT_04 => X"3E7FFE02482553FC3C020277E128080A1E6000003CC0000A6601E03A8B0F0008",
INIT_05 => X"F43F8140000203FFC806C8A1C1048FF0F0E07E1F00F7FFC00024010000468310",
INIT_06 => X"08710C10015E083D01A24404786BE0014114C3FE4187A009A663A680100B3096",
INIT_07 => X"200800008FDFFF00290000100211019812E210488228000000900260026C6058",
INIT_08 => X"0EF1F5FA0041FF080AC707FEFBC110008420F7FF388B70A20389346FE8000580",
INIT_09 => X"917FC30010107688862A28C54518DBFF00020004C0A6044901112A0908AA0A30",
INIT_0A => X"006309044081A001B188300E20806520398C6021569249C4B3007127080806FF",
INIT_0B => X"904595123203040D9228D9228D9228D9228D9228D9228D9228D99146C9146C84",
INIT_0C => X"88042090068008003120000806001402504110C48002403601887FEF80022A51",
INIT_0D => X"26C0AC404E43032CA0C205880A7FFAB7FE01409400400C0594A4002200110008",
INIT_0E => X"26C0AC086A170250454004C6012280129B034A080C0B0016A0D20346080C0A80",
INIT_0F => X"0B064092D85938C0112144050224120C500346080C0B0016A0D2034A080C0A80",
INIT_10 => X"40702E058355458967E86A170220D1800093414B0414782E4B5000D81480809A",
INIT_11 => X"081B1545104135443306C35901024F88A88049062A747512B76783C5D040E080",
INIT_12 => X"40160040D86B202049B22198362A8A208279854400A036801480031401900800",
INIT_13 => X"0DD001C002D38334000914028354008301008C0CF1480245108C7640A0604032",
INIT_14 => X"AC0496022300233104662848808E191526205018030060540284FA0C0044022C",
INIT_15 => X"004010040100401004010040102090010008000001C0E010020007DFFFC06E60",
INIT_16 => X"0401004010040100401004010040100401004010040100401004010040100401",
INIT_17 => X"4010040100401004010040100401004010040100401004010040100401004010",
INIT_18 => X"FF7FFDF7FF3E3DFDF7E000000000000000000000000040100401004010040100",
INIT_19 => X"FBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBFFDFDFFFCF3CF3FFFEF9FEE",
INIT_1A => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFEFF7FBFDFEFF7FBFDFEFBEFBEFBEFBE",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0004000100000000000000000000000",
INIT_22 => X"2A954BA0004154BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080402010FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF552A974AA0004174BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"000400000007FFFFFFFFFFFFFFFFFFFFFFEF552E974BA0804000AAF7FFFFFFFF",
INIT_25 => X"FFFFFFDFEF5D2E974BA002E97400007FFFFFFFFFFFFFFFFFFFFFFEF552E954AA",
INIT_26 => X"BA087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974BA082E95400007FFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2E954BA007FC00BA5D7FFFFFFFFFFFFFFFFFFBFDFEF5D2A954AA002E974",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFBFD",
INIT_29 => X"954AA080005000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA00000200000000",
INIT_2A => X"FFFFFFFFFFFFFFF552A974BA0000174AAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0A000AAE3FFFFFFFFFFFFFFFFFFFFFFFEF552A974AA0000104AAF7FFFFFFFFFF",
INIT_2C => X"FFBFDFEF5D2E974AA000A07000007FFFFFFFFFFFFFFFFFFFFDFEF552E954BA08",
INIT_2D => X"1C7FFFFFFFFFFFFFFFFFFBFDFEF5D2A974BA002A95400087FFFFFFFFFFFFFFFF",
INIT_2E => X"F552E974BA0020924BA1C7FFFFFFFFFFFFFFFF7FBFDFFF5D2A954AA082A92428",
INIT_2F => X"FFFFFFFFFEFF7FBFFFFF552E974AA0071C50BA557FFFFFFFFFFFFFFFF7FBFDFF",
INIT_30 => X"4BA000002000000000000000000000000000000000000000000000000E3FFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2A954AA080017410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"000AAF7FFFFFFFFFFFFFFFFFFFFFFFEF552A974BA0000174BAFFFFFFFFFFFFFF",
INIT_33 => X"BFDFEF5D2A954BA082E800AAA2FFFFFFFFFFFFFFFFFFFFFDFEF552E954AA0004",
INIT_34 => X"7FFFFFFFFFFFFFEFF7FBFDFFF5D2A974AA002E95410087FFFFFFFFFFFFFFFF7F",
INIT_35 => X"52E974AA082A820AA557FFFFFFFFFFFFFEFF7FBFFFFF552E954BA002E9741008",
INIT_36 => X"FFFBFDFEFF7FFFFFEF5D2A974BA0000020AA557FFFFFFFFFFFDFEFF7FBFFFEF5",
INIT_37 => X"0000000000AAFFFFFFFFFFBFDFEFFFFFFDFEF5D2E954AA0051554BA5D7FFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(2),               -- Port A write enable input
DIA(0)   => data_write_a(21),        -- Port A data input
DOA(0)   => data_read_a_lo_512(21),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(2),               -- Port B write enable input
DIB(0)   => data_write_b(21),        -- Port B data input
DOB(0)   => data_read_b_lo_512(21),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_22_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"5290F4CDE914905A14A43D33F488243E17122300F55FEB189B343A1140548380",
INIT_01 => X"A94007B259F6A975386262000C344BA9573C6FF57B18A5FB0ABFCD3C2C5F4F0C",
INIT_02 => X"D56B4302AC01005111011BD506AA5205274056900596A539584E2E6DFE4B2418",
INIT_03 => X"6B03F2F6151A2081F24001E8400008F401CB10C6594423C8923AD6B55AD0EB5A",
INIT_04 => X"8001023D37E50880436200808BC8492A0089249600101100008087248B64426E",
INIT_05 => X"A51035B41C0A88046CAEE8C23C08E040011C0020F8882001102D620A06D68301",
INIT_06 => X"B93FF975CF7889D085E997A2144E8FC2060B880081A26DCD4047EFF9EF018980",
INIT_07 => X"283800AA500200E8024AD03546A3262FB5AA5542A882040C7A64CBD64065F028",
INIT_08 => X"141008801018040E48D500400015805060040080A2A0F4A82381B4000A0905A0",
INIT_09 => X"4D0000002126F30C902A29C54539C020E11810098D4067EFF9FF284D483E2AB4",
INIT_0A => X"1400006100003202D040050220103D2A512C6A8C4F0008AA800470370000A000",
INIT_0B => X"013456520CA09281C2A81C2A81C2A81C2A81C2A81C2A81C2A81C9540E1540E00",
INIT_0C => X"A1402A13C0A10A893165281A1C2A7283516344C594A85536B1AD800214202C50",
INIT_0D => X"3C70FC20515808A0100820112300011000287B071105034406950A0285014280",
INIT_0E => X"3C70FC48E11CFC48400184CE0D6783139B0959A41606003C70FA0958AC160480",
INIT_0F => X"0D87E8B3B811B52048B10E0402AE1606D80958AC1606003C70FA0959A4160480",
INIT_10 => X"80F84E0185594581E088E11CFC38414020DD42CF909D7E0A551C02180300C0DD",
INIT_11 => X"441154C258012D86F3044A3133004A99BD8455300654458A1D588C4061403000",
INIT_12 => X"A096A240894626600953379822A984B0025B0DEC0345C9200680027181B44887",
INIT_13 => X"E2404160035482BE521C2C04A90783C18000D610B9D8070B12B1A2A62040202A",
INIT_14 => X"304244A91102C93A2D608D2A258DF8034284200C050070E40C80620C870B02C4",
INIT_15 => X"4411044110441104411044110466C440446CA06951D4EA801000980400646002",
INIT_16 => X"0100441104411044110441104411044110441104411044110441104411044110",
INIT_17 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_18 => X"FE8FF1F7DEBDDF7DF7D05122890000000003FFFFFFFF90040100401004010040",
INIT_19 => X"79E79E79E79E79E79E79E79E79E79E79E79E79E7BFFDFD7DDDF7DF7DF7DFBFDE",
INIT_1A => X"3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE79E79E79E79E",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE000000000000000003F9FCFE7F3F9FCFE7F3F9FCFE7F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0800000000000000000000000000000",
INIT_22 => X"2E974AA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000400010FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E954AA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"0004154BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA000015400FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF552A974AA0800154AAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA",
INIT_26 => X"BAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0004174BAFFFFFFFFFFFFFFFFF",
INIT_27 => X"FEF552E974BA0804000AAA2FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0000174",
INIT_28 => X"0000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040001000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E954AA000402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0417410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080005000FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF552A974BA0000174AAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA00",
INIT_2D => X"E3FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0804154BAF7FFFFFFFFFFFFFFFFF",
INIT_2E => X"F552E954BA000E124BAE3FFFFFFFFFFFFFFFFFFFFFFFEF552A974AA0000104AA",
INIT_2F => X"FFFFFFFFFFFFFFFFDFEF552E954BA080A000AAA2FFFFFFFFFFFFFFFFFFFFFFFE",
INIT_30 => X"4BA080400010000000000000000000000000000000000000000000000007FFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"17410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000400010FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF552A954BA000415400FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954AA0800",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFEF552A974BA0000174BAF7FFFFFFFFFFFFFFFFFFF",
INIT_35 => X"52E954AA0004000AAA2FFFFFFFFFFFFFFFFFFFFFDFEF552E974AA0804174AAF7",
INIT_36 => X"FFFFFFFFFFFFBFDFEF5D2E954BA002A820BAA2FFFFFFFFFFFFFFFFFFFFFDFEF5",
INIT_37 => X"0000000000087FFFFFFFFFFFFFFFF7FBFDFEF5D2A954BA082E800AAAAFFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000000FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(2),               -- Port A write enable input
DIA(0)   => data_write_a(22),        -- Port A data input
DOA(0)   => data_read_a_lo_512(22),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(2),               -- Port B write enable input
DIB(0)   => data_write_b(22),        -- Port B data input
DOB(0)   => data_read_b_lo_512(22),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_23_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"EF20906D902424807BC8241BC81801B97D38AD3C0800103362A6741C80A12A02",
INIT_01 => X"001FFF8409F089003B4422000D80C80106804A7951C5B9D1C828043EA28838F9",
INIT_02 => X"028406A002DC176444683862400003111001303FFC00F240D50146013B300500",
INIT_03 => X"001B243004080FE000177003145F87017D584B10D804034800200200A1008008",
INIT_04 => X"BEFFFC0248005FFC3C18A2FFE12222425E600000BDC0800AEE01E81A100F0A00",
INIT_05 => X"D03F8000000003FF810640A1C0008FF2F0E17E1F02FFFFC80100004044800080",
INIT_06 => X"800264B4854650040123428C204BF40F439647FF4807E189A477EF81DF0AF116",
INIT_07 => X"01000000FFDFFFE800401005C0A0008F86C60840AAAA100C68D1810C9F4A0020",
INIT_08 => X"1BE1F5F80003FF0002021FFEFBC80000000077FF184B03010004002FE1F29002",
INIT_09 => X"907FC308181204800600000000001BFFA800808189A657EF81DD0C00079CC800",
INIT_0A => X"0063090442A18001B188300C48907120AC810033149249C433200180082A06FF",
INIT_0B => X"9A41C1443243050C1010C1010C1010C1010C1010C1010C1010C1008608086084",
INIT_0C => X"000082A00600200080000500C000400800601200000254A000007FEFC1030221",
INIT_0D => X"0A9080400E0BF30C20CA858E087FFABFFE01409780214EE49620001000080004",
INIT_0E => X"0A908044294700701641005218521210150E5789F90A000A90800E5F81F90880",
INIT_0F => X"0E0220036864A7DCA190440301E2105C000E5F81F90A000A90800E5789F90880",
INIT_10 => X"C1400500C6CE5400032429470068924010164302048156305D66F8701681000E",
INIT_11 => X"2E0CCB0500013440600339C800004D8018000857A82920CE8CB220C81400A180",
INIT_12 => X"220344406739000009B0030019960A00026880C0422C52B01700044901488822",
INIT_13 => X"85C811A010428104128996465ADA020180804A040108A2658217C4008060300C",
INIT_14 => X"BE0692020328CA0028042054A92771C50FC070109000C1C819078280A265920E",
INIT_15 => X"020080200802008020080200800800200200000000000008004807DFFF000470",
INIT_16 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_17 => X"0080200802008020080200802008020080200802008020080200802008020080",
INIT_18 => X"0000000000000000000000000000000000000000000000802008020080200802",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000",
INIT_22 => X"2E974BA080002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E974BA000400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000400000FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF5D2E954AA080000010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA",
INIT_26 => X"10FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080402010FFFFFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2A954BA000015400FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA0804000",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E974BA080002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF5D2E954AA000402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA00",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080002010FFFFFFFFFFFFFFFFFFF",
INIT_2E => X"F5D2A954BA080407000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080005000",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF5D2A954BA000417410FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA080402000000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"02000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000010FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF5D2E974AA000402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0000",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000400010FFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"D2A954AA080017410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954AA080002000FF",
INIT_36 => X"FFFFFFFFFFFFFFFFFF552A954BA080015410FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_37 => X"0000000000F7FFFFFFFFFFFFFFFFFFFFFFFFF552A954BA000415400F7FFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000000FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(2),               -- Port A write enable input
DIA(0)   => data_write_a(23),        -- Port A data input
DOA(0)   => data_read_a_lo_512(23),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(2),               -- Port B write enable input
DIB(0)   => data_write_b(23),        -- Port B data input
DOB(0)   => data_read_b_lo_512(23),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_24_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100600007FFF000080108004000800020000840041000080808",
INIT_02 => X"0000068002CC07400000090C080002000000103FF811F150231000520ABE4404",
INIT_03 => X"8428180000080FE000177000001B87003D4000000E8B84010020000000008000",
INIT_04 => X"3E2FFC024800137C3C000077E00000001E6000003CC0000A6601E01A000F0200",
INIT_05 => X"103F8000000003FF80000021C0000FF0F0E03E1F0067FFC00000000000000000",
INIT_06 => X"00132412079001AD00810005E8000001401643FE4007E5501AA00000DC8C3006",
INIT_07 => X"000000000FDFFF62695A5685C094831D966000008002100C2040A178B600C240",
INIT_08 => X"08E1F5F80001FF00000007FEFBC00000000077FF000B00000000002FE0000000",
INIT_09 => X"107FC300000000000600000000001BFFA0000005501AA00000CE200000940000",
INIT_0A => X"00630104408180012188300C00814080008000010012414433000100080806FD",
INIT_0B => X"904181003003000C1000C1000C1000C1000C1000C1000C1000C1000608006084",
INIT_0C => X"00000080060000000000000012002C00000000000000000000007FEF80020201",
INIT_0D => X"440082404E0B332CA2C20188087FFAB7FE000082000000008220000000000000",
INIT_0E => X"4400824903210308074084210002460402009280010D80440084009280010F00",
INIT_0F => X"800A2400401A0C82183248060010280C20009280010D80440084009280010F00",
INIT_10 => X"C0A078160000404A0469032102981380202080026420020D06C002A08481C020",
INIT_11 => X"00164F400860000824059AD01802000208104817B00011306B2D9B0DD5082080",
INIT_12 => X"41021800B35A0300400041202C9E8010C0001040C5836CC01780018601030088",
INIT_13 => X"DB1011E000A140058220004AEFFC8101810021084301880030A8B77400603011",
INIT_14 => X"8C063C0220002201490418082010A57263E010000201033016085A40880030A1",
INIT_15 => X"000000000000000000000000000000000000000000000000000007DFFF0006E0",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"F6E7CC1132CDB444199000000000000000000000000000000000000000000000",
INIT_19 => X"79E79E79E79EFBEFBEFBEFBEFBEF9EF9EF9EF9EFA69861219575D75FF2D0AEEA",
INIT_1A => X"0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1EFBEFBEFBE79E",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE000000000000000000783C1E0F0783C1E0F0783C1E0F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020100000000000000000000000",
INIT_22 => X"2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"080002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_26 => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000400010FFFFFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2E974AA000400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0004000",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040201000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF5D2E974BA080002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFF",
INIT_2E => X"F5D2E974AA000400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF5D2E974AA000400000FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA080402010000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"00010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000010FFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002010FF",
INIT_36 => X"FFFFFFFFFFFFFFFFFF5D2E974AA000002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_37 => X"0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000402010FFFFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(3),               -- Port A write enable input
DIA(0)   => data_write_a(24),        -- Port A data input
DOA(0)   => data_read_a_lo_512(24),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(3),               -- Port B write enable input
DIB(0)   => data_write_b(24),        -- Port B data input
DOB(0)   => data_read_b_lo_512(24),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_25_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100200002000000080100004000000020000800041000080808",
INIT_02 => X"0000068002CC474000000800000002000000103FFCE302008000000880844A04",
INIT_03 => X"00000101C0200FF004177800081B87003D400000080000000020000000008000",
INIT_04 => X"3E2FFE024820137C3C004077F01000001E7249213CC1264A660DF05A000F9000",
INIT_05 => X"103F81C1002203FF80000021C1140FF8F0E03E1F0067FFE04800258280010052",
INIT_06 => X"80480AE20000000100000001C8608001401643FE4007C00000000000CC083006",
INIT_07 => X"280800000FDFFFEA4050140540B00100840000080002A00C2040810000000010",
INIT_08 => X"C8E1F5FA21C9FF80040007FEFBE031018C31F7FFBAEBC0020008086FE0000100",
INIT_09 => X"107FC301800000000600000000001BFFE00301000000000000CC020000140000",
INIT_0A => X"0077330C4889CC292588300C0080400000800001001243443B000100880806FD",
INIT_0B => X"904189003003000C1000C1000C1000C1000C1000C1000C1000C1000608006084",
INIT_0C => X"8B04228026824100000000000000000000000000000004A000007FEF80020201",
INIT_0D => X"400000400E03C30C20C2818C087FFAB7FE01409700C10007962418220C110608",
INIT_0E => X"4000000001010000004000000000400400001200000800400000001200000800",
INIT_0F => X"0008000000000480000040000000200000001200000800400000001200000800",
INIT_10 => X"0000001001000002000001010000100000000000202000000440000000800000",
INIT_11 => X"0000410000000008000008400000000200000806300400000820000020004880",
INIT_12 => X"0000080001080000000040000082000000001000000040800800000000020008",
INIT_13 => X"8100000000000000802000000840000200040000020008000000840000804000",
INIT_14 => X"8C04100200000200000610000000210000000018140000000008000008000000",
INIT_15 => X"04411044110441104411044510629041040D180400000010028047DFFF800C60",
INIT_16 => X"4411044110441104411044110441104411044110441104411044110441104411",
INIT_17 => X"4110441104411044110441104411044110441104411044110441104411044110",
INIT_18 => X"196A8C5A2932EC15DA080800002FFFFFFFFFFFFFFFFFC1104411044110441104",
INIT_19 => X"92492492492410410410410410410492410492412000531215A69A6BFBA2894A",
INIT_1A => X"B158AC562B158AC562B158AC562B1588C46231188C46231188C4924924924924",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000B158AC562B158AC562B158AC562",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000",
INIT_22 => X"2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF5D2E974BA080400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_26 => X"10FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0800000",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400000FFFFFFFFFFFFFFFFFFF",
INIT_2E => X"F5D2E974BA080000010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA080402000000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"02000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400000FF",
INIT_36 => X"FFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_37 => X"0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000000FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(3),               -- Port A write enable input
DIA(0)   => data_write_a(25),        -- Port A data input
DOA(0)   => data_read_a_lo_512(25),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(3),               -- Port B write enable input
DIB(0)   => data_write_b(25),        -- Port B data input
DOB(0)   => data_read_b_lo_512(25),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_26_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"E9264EAB20190CA3BA4997AA9002AE9C001006B0778015CFA17E0811039879C7",
INIT_01 => X"F1FFF9BB1F773C7F9BB07DFFFDD863FC5FFF3FEFFBBF9FFB22FFFBC7B9F30686",
INIT_02 => X"9B3184F8AFDEAF300029E4E300FC78A6258548EFFA71C00172082400003A2161",
INIT_03 => X"0213C3FDFFFC7F74FFBF737A603B87FEBE1A5294F65628A0001B9CE6CC606E73",
INIT_04 => X"7E2EFEBF6FFEB37C3FF3017776FFCDA43E7B6DFD7DEBFD8E6F5F78DF0BFBD644",
INIT_05 => X"902F87C74E8CCFFBB6FF70E1FE61FFBDF0FEBE1FFD67DFFEFFBDA7F7FED50870",
INIT_06 => X"213246200BCC8920360C1831CD7DF60A244B9BFEE00589DDBCEFEDC1DFA08957",
INIT_07 => X"B1D4223B4FFDFF21CC721C85DCE1458E8782484020A2C1FCA3468D77E0000300",
INIT_08 => X"2C05FD7BC471FBD13D980FBEFBEBF30B8D79FF7F451F33CFD60FE8FFFDF54003",
INIT_09 => X"19FFC71FEFED7B251E35768E8ED6BFDF3EB3EBF9DDBCE7FDC1DF8A760F3EACC0",
INIT_0A => X"56F7730ECCDBDF152199F51EDDCDEBCFF589807B7096CD4CF73AC1FC98884FFF",
INIT_0B => X"B867D3683A03A40F78C0D78C0D78C0D78C0D78C0D78C0D78C0D7A606BC606B8C",
INIT_0C => X"DFBFF5EB36DFE51FC3A80D73D840303983EE7F0EA03BDA680137FFFDFFD7E681",
INIT_0D => X"3F0080425E6BFF8DB0DAE19C09FFFFE7FE3EBEA8EB7AFEE5C9AEBD7F5EBFAF5F",
INIT_0E => X"3F00800DEC010280004000F808020290100FA2F60008003F00800FA2F6000800",
INIT_0F => X"00023002007BC0A14E00400003B8000D000FA2F60008003F00800FA2F6000800",
INIT_10 => X"01E0320007204008040DEC010300100000F600020581003F604D0700008000EE",
INIT_11 => X"201F21A2C40039006807C46426040E101A0259DFE82011A311AA042016040080",
INIT_12 => X"80020048F88C84C101C203403E434588007200D047F00090200007E0010009B0",
INIT_13 => X"0109000003E2000416C0804FE04140E80000F808010AB02033AC048A2A00003D",
INIT_14 => X"FFAFD082003B032FB987E04021D481D4000419060201E1A000044300B02033E8",
INIT_15 => X"AFEBFAFEBFAFEBFAFEBFAFEFFBFBFBFBBFCFBB0FFDFEFFEF2DFFFFFBFF802FFD",
INIT_16 => X"FEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBF",
INIT_17 => X"EBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFA",
INIT_18 => X"F491E166CC8553F86EDB5C88646FFFFFFFFFFFFFFFFFEBFAFEBFAFEBFAFEBFAF",
INIT_19 => X"1861861861861861861861861861869A69A61861AFBD54D5F871C71D475B15BC",
INIT_1A => X"0984C26130984C26130984C26130984C26130984C26130984C26186186186186",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE000000000000000000984C26130984C26130984C2613",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000",
INIT_22 => X"2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_26 => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFF",
INIT_2E => X"F5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA080402000000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"02010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_36 => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_37 => X"0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(3),               -- Port A write enable input
DIA(0)   => data_write_a(26),        -- Port A data input
DOA(0)   => data_read_a_lo_512(26),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(3),               -- Port B write enable input
DIB(0)   => data_write_b(26),        -- Port B data input
DOB(0)   => data_read_b_lo_512(26),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_27_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"00080A40000A41248002029000050A088000008242A0004404480002000A1155",
INIT_01 => X"F1FFF1C11F781C129C107DFFFE0860941E81258CA2B71C2220EC1B86E1A00002",
INIT_02 => X"183080988B2EAE00002BE001117C78C6848140CFFA0000800042008000011081",
INIT_03 => X"000003FDF3E47C74F7BCF36A203A47F6B8184210B6160820001318C60C204C63",
INIT_04 => X"7E28FEBF6FEEB3723F71017476DFC524397B6DF572EB6C8E175E70D90F539600",
INIT_05 => X"000F86064C8DDFE3B6FF50D1FC61DE39C8FCB91FF9671FE6B68984B5BCE40834",
INIT_06 => X"0000000800000042020C18300520620A80231BFE200181092CE7ED80DFC00147",
INIT_07 => X"8AC4AA3B0FD1FF201044110560884000840200520002080C23468D0300000282",
INIT_08 => X"2005F0784411E390A4880E3DF7E2FB0B8E717C7F411F3BC6D60B60FFDDE44001",
INIT_09 => X"18FFD757E7ED7A211E81C09818109E1F16B16B71092CE7ED81CF403601228C40",
INIT_0A => X"46FF730E5CCBCD55219AB55F0DEFABC7054880693016DD4C755AC16C1A884FFE",
INIT_0B => X"BC63F1683803C00E3440C3440C3440C3440C3440C3440C3440C3C2061A2061AD",
INIT_0C => X"56BF55CB165EC51D41880FA3F040202883B475062033186801137FF1BAD6F281",
INIT_0D => X"3B0000421E2B0F2E2AE215C808FFFA47FE62BAA86B1AB268E92AB56D5AB6AD5B",
INIT_0E => X"3B000025EC010080004000F808000098100F22520008003B00002F2252000800",
INIT_0F => X"00001042006BC0810600400003B80001002F22520008003B00002F2252000800",
INIT_10 => X"01E032000620000C0405EC010100100000F6000001C1003760410500008000EE",
INIT_11 => X"201D2120840039000817444404040E10020218DE282010A311AA002002040080",
INIT_12 => X"8000000AE888808101C20040BA4241080072001027F00080200007E0000001F0",
INIT_13 => X"0101000003E2000007C0800FE04040280000F8080002F02023AC04080A00003D",
INIT_14 => X"DDAFD082001B03249887E04001D481D4000009020201E1A000040100F02023E8",
INIT_15 => X"ADAB6ADAB6ADAB6ADAB6ADAB6BF1EBDABD8E270BF84A25C6ACB777E3FF800C6D",
INIT_16 => X"DAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6",
INIT_17 => X"AB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6A",
INIT_18 => X"100481CA860402104A471688747FFFFFFFFFFFFFFFFFAB6ADAB6ADAB6ADAB6AD",
INIT_19 => X"0000000000000000000000000008200000000000200072F210000001490E2168",
INIT_1A => X"A05028140A05028140A05028140A050080402010080402010080000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000A05028140A05028140A05028140",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000",
INIT_22 => X"2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_26 => X"10FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFF",
INIT_2E => X"F5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA080402000000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"02000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FF",
INIT_36 => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_37 => X"0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000000FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(3),               -- Port A write enable input
DIA(0)   => data_write_a(27),        -- Port A data input
DOA(0)   => data_read_a_lo_512(27),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(3),               -- Port B write enable input
DIB(0)   => data_write_b(27),        -- Port B data input
DOB(0)   => data_read_b_lo_512(27),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_28_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"02200AA400180030808802A900002A08001280A08A801044104A1000001818C3",
INIT_01 => X"50A00011460214428114180000882214413D0A71592A01D92213D28005210202",
INIT_02 => X"8A54800A210200111100C2110054289220810440030404010844000444410001",
INIT_03 => X"4200040822D4500001E0000028000002000211842010092000018C6295200631",
INIT_04 => X"00400000000B8000000140000005840C00000040002008808100048100100044",
INIT_05 => X"0000222200244400135110000135100000000000000000024CA0A01018000320",
INIT_06 => X"A004912008208040024489121144080400081000200008104000000020000041",
INIT_07 => X"A85800994000000A0200802004204420210001022AA8A0001122448142491008",
INIT_08 => X"0414000201800004080A000000124058200408000880004440004080160C4100",
INIT_09 => X"0080000206CB0821082B694D4D29400002002038104000000020003204000440",
INIT_0A => X"12000843066021001400040024440245400082D022040000400800081022C000",
INIT_0B => X"0002002C004001036050160501605016050160501605016050160280B0280B00",
INIT_0C => X"0012400810080414C0A800310840102182C62302A0194C08001680100E4040A0",
INIT_0D => X"05000002003004208208841401800040000A0000200814004198000400020001",
INIT_0E => X"0500000004000080000000000000028000002052000000050000002052000000",
INIT_0F => X"0000300000004001060000000000000900002052000000050000002052000000",
INIT_10 => X"0000000001200000000004000100000000000000050000002001050000000000",
INIT_11 => X"00002020840000004800040404040000120200A9000000010000002002040000",
INIT_12 => X"0000004800808081000002400040410800000090001000002000000000000910",
INIT_13 => X"0001000000000000144000010000402800000000000A1000010000080A000000",
INIT_14 => X"0080000000110006B08140000040000000000902000000000000410010000100",
INIT_15 => X"0080200802008020080200802101210810C39A66A90A85420413A82000000204",
INIT_16 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_17 => X"8020080200802008020080200802008020080200802008020080200802008020",
INIT_18 => X"110A00246972BD89A40A0C22E100000000000000000000200802008020080200",
INIT_19 => X"82082082082082082082082082082082082082080D35050758C30C31DE21102C",
INIT_1A => X"B0582C160B0582C160B0582C160B0580C06030180C06030180C0820820820820",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000B0582C160B0582C160B0582C160",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000",
INIT_22 => X"2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_26 => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFF",
INIT_2E => X"F5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA080402000000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"02000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_36 => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_37 => X"0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000000FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(3),               -- Port A write enable input
DIA(0)   => data_write_a(28),        -- Port A data input
DOA(0)   => data_read_a_lo_512(28),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(3),               -- Port B write enable input
DIB(0)   => data_write_b(28),        -- Port B data input
DOB(0)   => data_read_b_lo_512(28),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_29_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"79964E4BA01DACAB9E659792D00AAE160002829C7FDFEFCEE97C2815039D70C3",
INIT_01 => X"50BFF9AB0775343F9AB01DF80D5821FC0FFF3FEFD1AF9FF1207FFBC7B9720586",
INIT_02 => X"0D15846807D207200021C4E200D428A2018408600271C000720A0000003A2161",
INIT_03 => X"0002C009EEFC5F10F9B70178681B80FA3E000100765029A00019084345606421",
INIT_04 => X"3E6E023D27DA937C03E3407712E5CDA41E0924DC3D20B98AE905189F0BF8C000",
INIT_05 => X"902003C30E0447F877F930203E213F8CF01E3E00FC67C03A4D9C87525E510160",
INIT_06 => X"0012460003CC002036040811D919F402244293FEE00400CCB46BA4C164A08857",
INIT_07 => X"914800110FFC0001CC320C81D841418E82800100000041FCA1428575A0001108",
INIT_08 => X"0805FD0180E1F8C1111A0782082B50080508FF00048B124D4005C8AFF4154102",
INIT_09 => X"0180000ABFEF89250815568A8AD6ABC02A02A0B0CCB463B4C0748A720B1EA4C0",
INIT_0A => X"021410028450530014014002D445624DB481806A62840800C22800B8900042FF",
INIT_0B => X"0806522C0A40A50268D0068D0068D0068D0068D0068D0068D006A68034680300",
INIT_0C => X"8912E0A83289641F42A80561D040203182AC3D0AA0118A080036FFFC4F4164A0",
INIT_0D => X"050080424069F5A51250648801BFFFE0003E3E00A0685A85410C0816040B0205",
INIT_0E => X"050080080400028000000000000202900000A0F600000005008000A0F6000000",
INIT_0F => X"00023000001040214E0000000000000D0000A0F600000005008000A0F6000000",
INIT_10 => X"000000000120400800080400030000000000000205800008200D070000000000",
INIT_11 => X"000220A2C400000068008424260400001A0241DAC80001010000042016040000",
INIT_12 => X"00020048108484C10000034004414588000000D04010001020000000010009B0",
INIT_13 => X"000900000000000416C00041000140E800000000010AB0001100008A2A000000",
INIT_14 => X"A282C0000033010FB181E00020400000000419060000000000004300B0001100",
INIT_15 => X"02C0B02C0B02C0B02C0B02C4B12B312912831A27FCFE7FFB175B6FF800802594",
INIT_16 => X"2C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B",
INIT_17 => X"C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B0",
INIT_18 => X"EE7FFDF7FE783FFDFFEA0C00602FFFFFFFFFFFFFFFFFC0B02C0B02C0B02C0B02",
INIT_19 => X"BEFBEFBEFBEFBEFBEFBEFBEFBEEBAEBAEBAEBAEBBFFDF9FBEFFFFFFEBBCF9F96",
INIT_1A => X"FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFBEFBEFBEFBEF",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000FBFDFEFF7FBFDFEFF7FBFDFEFF7",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000",
INIT_22 => X"2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_26 => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFF",
INIT_2E => X"F5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA080402000000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"02000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_36 => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_37 => X"0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(3),               -- Port A write enable input
DIA(0)   => data_write_a(29),        -- Port A data input
DOA(0)   => data_read_a_lo_512(29),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(3),               -- Port B write enable input
DIB(0)   => data_write_b(29),        -- Port B data input
DOB(0)   => data_read_b_lo_512(29),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_30_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"FF9FE1F7FFBFFFFDFFD000000000000000000000000000000000000000000000",
INIT_19 => X"79E79E79E79E79E79E79E79E79E79E79E79E79E7AFBD75F5FDF7DF7FF7FFBFFE",
INIT_1A => X"3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE79E79E79E79E",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE000000000000000003F9FCFE7F3F9FCFE7F3F9FCFE7F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000",
INIT_22 => X"2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_26 => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFF",
INIT_2E => X"F5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA080402000000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"02000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_36 => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_37 => X"0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(3),               -- Port A write enable input
DIA(0)   => data_write_a(30),        -- Port A data input
DOA(0)   => data_read_a_lo_512(30),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(3),               -- Port B write enable input
DIB(0)   => data_write_b(30),        -- Port B data input
DOB(0)   => data_read_b_lo_512(30),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_31_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"129000008004A00804A40000400800020000000C005FEA005800200400050100",
INIT_01 => X"A15FF18019700810180065FFFC0040801E80258CA2951C2200EC0906A0804140",
INIT_02 => X"146000808A0C060444692000402850040400408FF80000000010000000004000",
INIT_03 => X"000003F5D1202C70F654716A001A07F438184210960600000012108518004842",
INIT_04 => X"3E28FE3F6FE513703F70007472DA4128187B6DB530C1240A060C70580B439200",
INIT_05 => X"000F84040C088BE3E4AE40C1FD04CE38C0FC381FF8671FE01009048084C40010",
INIT_06 => X"0000000000000008000810200420620E00030BFE000181092CE7ED80DF800106",
INIT_07 => X"000000220FD1FF200040100540800000840200408002000C2244890200000200",
INIT_08 => X"0011F0780011E38004800E3CF3E0B1118C31747F000B33820209206FC9E80000",
INIT_09 => X"187FC301B124F2001600000000001A1F00110101092CE7ED81CF000401228800",
INIT_0A => X"0477330C4889CC012188310E08812982050800A91012494C31004124080886FE",
INIT_0B => X"9861D1403803800C1000C1000C1000C1000C1000C1000C1000C1800608006084",
INIT_0C => X"020400830602410901000D02D0002008012054040022102001017FE190022201",
INIT_0D => X"3A0000401E030B0C20C20188087FFA07FE203A80010002608030102008100408",
INIT_0E => X"3A000005E8010000004000F808000010100F02000008003A00000F0200000800",
INIT_0F => X"00000002006B80800000400003B80000000F02000008003A00000F0200000800",
INIT_10 => X"01E03200060000080405E8010000100000F600000081003740400000008000EE",
INIT_11 => X"201D0100000039000007404000000E1000001846282010A211AA000000000080",
INIT_12 => X"80000000E808000001C200003A0200000072000007E00080000007E0000000A0",
INIT_13 => X"0100000003E200000280800EE04000000000F8080000A02022AC04000000003D",
INIT_14 => X"9C06D082000A03200806A040019481D4000000000201E1A000040000A02022E8",
INIT_15 => X"0401004010040100401004010060C040040C200950402090128057C3FF800C60",
INIT_16 => X"4010040100401004010040100401004010040100401004010040100401004010",
INIT_17 => X"0100401004010040100401004010040100401004010040100401004010040100",
INIT_18 => X"000000000000000000001000802FFFFFFFFFFFFFFFFF81004010040100401004",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000",
INIT_22 => X"2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_26 => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFF",
INIT_2E => X"F5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA080402000000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"02000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_36 => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_37 => X"0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512,               -- Port A enable input
WEA      => wbe_a_lo_512(3),               -- Port A write enable input
DIA(0)   => data_write_a(31),        -- Port A data input
DOA(0)   => data_read_a_lo_512(31),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512,               -- Port B enable input
WEB      => wbe_b_lo_512(3),               -- Port B write enable input
DIB(0)   => data_write_b(31),        -- Port B data input
DOB(0)   => data_read_b_lo_512(31),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_0_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"ED39BA795990D275FB4A6E96ACC4731DEA4598B0AFB54867F6EE4618C3749803",
INIT_01 => X"58A0047C8607844847CA180001E4A2404042106208408208C2002069161734B3",
INIT_02 => X"8B1EC9562121F8051500147A0E5629A302CF28400615F5787B09FBF999BB1EFD",
INIT_03 => X"404EFC0A2AD6100F01A88E851CE47803C280110521898F6996088862C7B22221",
INIT_04 => X"C0D001C0100AEC83C008E7880D01A64661800002C21A52C590D2012194804844",
INIT_05 => X"650002C3F08754001B51981E007910070F01C1E003980015A204C22F32328BAF",
INIT_06 => X"BCDA4677CAEE7CF5BB870E1DDB9889C5FBFC440129A0604442180238203F70C1",
INIT_07 => X"7AAE0088B02000C2EC3A0E829836E0AF3325372E2AA8FDF3C18306758B24197A",
INIT_08 => X"D7E40002F7AE005FFB4730010411400A61080000F7F4C464B58294901606D5A5",
INIT_09 => X"C4801C40469B0CA9881A28C141118000C5A85A60444210123820B43B40804274",
INIT_0A => X"400800219010107ED453C041B13216656074EA560F0092A24856B05312226900",
INIT_0B => X"27122C3E04E03383E2781EA781E2781EA781E2781EA781E2781C33C0613C0E29",
INIT_0C => X"74EB1F50D0758A9650E520610A6A57A5529E2B439499CF96B086000000B09870",
INIT_0D => X"04F07E024108F4E28638EC57250004480155C1375A97A9121F8BA749D3A4E9D2",
INIT_0E => X"04F07E42177EFDF8570184071575970F8FC07D5BFF078004F07E007D5BFF0780",
INIT_0F => X"8F85ECB1FE047F5FB7B30E0700461E5AF8007D5BFF078004F07E007D5BFF0780",
INIT_10 => X"C0184D07C1DF15C7E3E2177EFDF8C3C03009C3CDD47C7F403FB3FDF89701C011",
INIT_11 => X"4F80FE659C6104C6D7103F9D1D064189B5924418D65FE45DEE55BBEDE34CF900",
INIT_12 => X"6395F64207F3A3A1483136B881FCCB38C2098DACA01FFF603F80001F80FDC81F",
INIT_13 => X"FED151E01015C3BB507D3F811FBEC32B81840714F8D91F4FC513F37C8AE07002",
INIT_14 => X"61692F293185D8D724E15D3FCC6B7C236FE0691A9500125C1F83F8CC1F4FC507",
INIT_15 => X"E93A4E93A4E93A4E93A4E93A4F942F90E9628540052090650525A0000066A00B",
INIT_16 => X"93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4",
INIT_17 => X"3A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E",
INIT_18 => X"09B56C74DAB15D1CF13501AA495000000000000000003A4E93A4E93A4E93A4E9",
INIT_19 => X"2082082082082082082082082082082082082082082084E41DC71C7155F3898E",
INIT_1A => X"3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F8208208208208",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE5294A5294A52800003E1F0F87C3E1F0F87C3E1F0F87C",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000030FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"A975EFFFAABDE00FFAEBDFFF5D2EAAAAAF7AEBDEBA0000000000000000000000",
INIT_22 => X"8000155087FC0155F7D168B55007BFDF45085168ABA002E82145085155545F7A",
INIT_23 => X"FFFD7545AA8028A00A2802AABAFF8028BEF5D7FFFE10005542145557FD5545FF",
INIT_24 => X"F7AEAAAAAA2FFFDF4500043FE105D2E954BAF7FFC0010080017555555568AAAF",
INIT_25 => X"A5D5168A00A2D142155005142010FFAE820AAFF842AABAA2AE95545FFD168ABA",
INIT_26 => X"FF5D2A821550000000BA007FD55FF5D7FC0145007FD7400550415410002E974B",
INIT_27 => X"F455D5142000082E82145FFD17DFEFFFD168BFFF780000BA007FE8AAAFF803FF",
INIT_28 => X"0000000000000000000000000000000000000000AAFBEAA00007BFDFFF082EBD",
INIT_29 => X"AABEA495FC716F002A975FFE3AA95E00EBAEBDFD75D2AA8A80EA8E2FE3F00000",
INIT_2A => X"56A16D557BC257D415E0216FA3F1E8FC0145B68B551475FAF6D1C556F0AA1C24",
INIT_2B => X"7FD24AFE3D02DAAAE12BD5545A2803AA0000542A0070071C50BAFEF1FAE0016D",
INIT_2C => X"A8B50F55A2F150005A3A438BD04AFAB8F550A8010E004924874825D7FEAA8548",
INIT_2D => X"A2A5504001C74BA42A1571E8028E3DB7816D0120155EA568E870BAEB8A05A2AE",
INIT_2E => X"2FFAFD2A82485FD2415A105C21451ED42A002545E055FFBE81D0BE8EA8A3AA05",
INIT_2F => X"100AA1D0F6F480B6A555A2A57A002A3D5FDB6A5C7E3DFFFE90B45B47ABA497A8",
INIT_30 => X"A0AFE80A8B0A000000000000000000000000000000000000000000000B55EAAA",
INIT_31 => X"ABEF5D557FEBA55022A3F70C6B405F4D2AE975EFAAAAB5E1AF3AABFF45592E88",
INIT_32 => X"411A8DED57CE1055555E5F58EFFC01FE2CACB65F520EBE9EF67D7BEA1FD5D556",
INIT_33 => X"A4AD0079C75D6070CC5CBB0280C029ABAA3EBC114728007521170821CE0FDE69",
INIT_34 => X"2A95E02A2AAB5EB0F280800EFAEE9F5D18F3142341D5DEEBEF55080034E0A592",
INIT_35 => X"B69C30E02116220415A9540AA854140A0A2047F353AAF6C77F7F20D968BF5781",
INIT_36 => X"ABEBE1B4D792A4AD1183454180DD3FDCAAAB7C91565455C141E41887D58AC448",
INIT_37 => X"F0000001FF01EABC4B8014174FF7DA80F52FEDE6BE93172D7D625B556EEAB157",
INIT_38 => X"FF0000001FF0000001FF0000001FF0000001FF0000001FF0000001FF0000001F",
INIT_39 => X"0000000000000000000000000001FF0000001FF0000001FF0000001FF0000001",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000100000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(0),               -- Port A write enable input
DIA(0)   => data_write_a(0),        -- Port A data input
DOA(0)   => data_read_a_hi_512(0),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(0),               -- Port B write enable input
DIB(0)   => data_write_b(0),        -- Port B data input
DOB(0)   => data_read_b_hi_512(0),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_1_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"212C001411984004084D000508C53810A03D1450E839B003342114428A000803",
INIT_01 => X"08000011400A100A81160000008C005400400002000000000000028001340000",
INIT_02 => X"C084484000002014400205851002007030450E0000A606C8C44CB4C6666C00E0",
INIT_03 => X"33DF380008164004000002000C80400002031943000101091608463061120118",
INIT_04 => X"4140008000000002000064000400004201000000000210458010070080100433",
INIT_05 => X"8500101040200000010009100000000508000100000000002010600100208D04",
INIT_06 => X"B5EDFDE24618AD433060C182BA860044204C000008A004100008000820280020",
INIT_07 => X"581E02100020000A81244890AA20263030517F122AA801F0983060AC564BF808",
INIT_08 => X"00820800C7A00045B103200000140A02234808000584000004808400020011A4",
INIT_09 => X"0000104000020082800808111008400000200204100000100820800144000414",
INIT_0A => X"12804062945211441E13C051156E800008402802060C94000040901102800000",
INIT_0B => X"24002006406401918C191AC191A4191A4191AC191AC191A4191A00C8560C8D29",
INIT_0C => X"0408010040050880383820080F105F05800302E0E08842422006000000041032",
INIT_0D => X"05000600000090C1841808172580000000008008020084082080204010200810",
INIT_0E => X"0500066210000178470184000000878402C000001E07800500062000001E0780",
INIT_0F => X"00003C404600000011A30E0700000009382000001E07800500062000001E0780",
INIT_10 => X"C0180000012010C20022100000F0C3C03000000055200340000000F88701C000",
INIT_11 => X"05800241186100004D100098190240001290002050068000001010486140F900",
INIT_12 => X"0000164A001303204800026880048230C2000094A0000F601F8000000001C908",
INIT_13 => X"12D051E01000000154200580003C030381840000004B08014401025480E07000",
INIT_14 => X"40082300218450C2800010094000482142E0601895001000000041C408014400",
INIT_15 => X"0802008020080200802008020080008208600500A82A15008000000000468000",
INIT_16 => X"8020080200802008020080200802008020080200802008020080200802008020",
INIT_17 => X"0200802008020080200802008020080200802008020080200802008020080200",
INIT_18 => X"BABEFC54A0810C7452B5420A1000000000000000000002008020080200802008",
INIT_19 => X"AAAAAAAAAAAAAAAAAAAAAAAAAAA28A28A28A28A2A8218D2C0C92492581328A46",
INIT_1A => X"2E974BA5D2E974BA5D2E974BA5D2E975BADD6EB75BADD6EB75BAAAAAAAAAAAAA",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFF6318C6318C63000002E974BA5D2E974BA5D2E974BA5D",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"00000000000000000000000C0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"002155557FFFFFF007FC21EFA2FFD74AAAAD5555550000000000000000000000",
INIT_22 => X"7FD75FFAAAA800AAF7AA974BAFFFBE8B45F7AEBDF455D2EAABEFF7FFE8BFF5D0",
INIT_23 => X"0557DF45AAD1400BAA2AE801550051555EFF7AA95400552AAAABAFFD1574105D",
INIT_24 => X"FFFBEAB55F780020AAAA80020AA082EAAB5500517DF555D2EAAA105500001550",
INIT_25 => X"AF7AE820AA0851574BAA2D1574AA5D7BFDEBAFFD540155557FD5400F78028BFF",
INIT_26 => X"FFFFD56AAAAFFFFD7555AAD168B45AAAEAAABAFF842ABEF5D517DF55552A974A",
INIT_27 => X"4BAF7AE80010082A97410557FEABFFAAFBE8BEFAAD1575EF557FFFE10557FFFF",
INIT_28 => X"00000000000000000000000000000000000000005D7FFDF4500043FE105D2E95",
INIT_29 => X"A8BC2EBDFEAF7F1F840017D4975D2FEF147FC51C7A2FBD5490BFD1C056A00000",
INIT_2A => X"AA8AAAE3D145410F7F1D55D71C002DABAEBAA974BAF7FFEFB45FFAABDF55492A",
INIT_2B => X"0E2AE85028B40155145F7AF6DBED5450AA1C2080BEF495FC71D54124924385FA",
INIT_2C => X"571D2E28E38E0216FA2D1E8E80140F45082B4002D082082AB8B6DBEDB7DF7F54",
INIT_2D => X"A97F7AF6D417E92482BF84020BA495557E3FF78E021FF1471FDEAAFFD56F16D5",
INIT_2E => X"7002FD74951D71EDFFABFD16FAAAE92BD5545A2DA3FB7DAAD4AAAAF487BC70BF",
INIT_2F => X"550A8010E00492487482FFFE82A85EBAE2FFC55554ADBD7A2FFC7BEFF6FFD7FC",
INIT_30 => X"400FBF9424F7000000000000000000000000000000000000000000000547AB8F",
INIT_31 => X"DF55F7AABFF55082CA8B4DF6C1E8F5E5400021EF005162BEF047FD5545AAFBF7",
INIT_32 => X"404547184164AA5D2EBEEB0A2D555410D3555714F8338AAAA1D0AE974AAF7FFF",
INIT_33 => X"AEABFFDF79DCBF755962010BDCBBC21455D7FEABEF75550ACBB7582225FF5843",
INIT_34 => X"D57D412F7D55F5E50C7F401BAAE8403CF5A3FFEAAEB083BC1000FF8409000512",
INIT_35 => X"2AA9FEAFDF7F431A9F7FFE81FF013A8001AFF801F8BA0C57740BDAA0688E5405",
INIT_36 => X"A2FBF7FED2C7F955445079E280A00C56145EF5D16BABAA3EBC3157ABD5FFE55F",
INIT_37 => X"0000000000596EBEF55080034E0A592A4AD00FB863550229BCABEB7DA403FFFD",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000100000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(0),               -- Port A write enable input
DIA(0)   => data_write_a(1),        -- Port A data input
DOA(0)   => data_read_a_hi_512(1),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(0),               -- Port B write enable input
DIB(0)   => data_write_b(1),        -- Port B data input
DOB(0)   => data_read_b_hi_512(1),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_2_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10E006600180111284380310006289800480032283E000A34301002001A0817",
INIT_01 => X"A14AC00A1079284D04A044A54E504368404000720885800802000006ECD10200",
INIT_02 => X"92250052A0348C310102048800A8507000040C8550200000480E0080001321E0",
INIT_03 => X"020204E4593C0824400C2220483042809292430400440180000890A4C9400242",
INIT_04 => X"486854B141002252142241502460480031B94420634850069A42241009610A04",
INIT_05 => X"800504244080892105AA6010A44882144840910A21220A8C820025E4A0000B00",
INIT_06 => X"A000442802280000340810209C444804206000AC800088096A0EA8C022208012",
INIT_07 => X"309820A848E0AA09826489A5CC49002001020112028201F8A20488260000108A",
INIT_08 => X"2400582881E0C1419D12041455509341A539C42A0D8208099002801700D10103",
INIT_09 => X"110D525861263100009200151409130A3C80C8C8096A06B8C12088400A9C2080",
INIT_0A => X"0451394CD0391A441583C04B580040089581001342801044877200D002A00DE0",
INIT_0B => X"144423040240450114901149013C9011C9013C9011C90134901144801A4808A5",
INIT_0C => X"D8A5345206D2C10082080A90C00000188150100C202A4640000E2B4081969420",
INIT_0D => X"050080400A0391A51240C480000AA902AA009028C83220008086952B4285A54A",
INIT_0E => X"05008021C00000000040000000020288000500000008000500802A0000000800",
INIT_0F => X"0002300000428000000040000000000D002A0000000800050080250000000800",
INIT_10 => X"0000000001204004000508000000100000000002054000130000000000800000",
INIT_11 => X"000C00000000000068144000000000001A000106200010021002000000000080",
INIT_12 => X"0002004A880000000000034098000000000000D024A000000000000001000900",
INIT_13 => X"00000000000000041400000A8000000000000000010A00000284000000000000",
INIT_14 => X"012100000002000280000000011080C000000000000000000000430000000260",
INIT_15 => X"A769DA769DA769DA368DA36CDA3A9A13A14801404134DA84A024024155000399",
INIT_16 => X"168DA769DA769DA769DA368DA368DA368DA769DA769DA769DA368DA368DA368D",
INIT_17 => X"68DA168DA169DA569DA569DA568DA168DA168DA169DA569DA569DA568DA168DA",
INIT_18 => X"138D70C030B51C50C7D000A2012F81F81F83F03F03F069DA569DA569DA568DA1",
INIT_19 => X"1041041041041041041041041041041041041041024860208165965975960040",
INIT_1A => X"25128944A25128944A25128944A25128944A25128944A2512894104104104104",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFF8421084210840703F25128944A25128944A25128944A",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"00000000000000000000000F0FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"415555087BFFF55A2AA800BAFFAE9540008002AA000000000000000000000000",
INIT_22 => X"7FE8B555551421455D0002145552EBFEBA007FC21EFA2FFD75EFAA8415410AA8",
INIT_23 => X"FFFE8B45552EBDF45FFAEAABFFF7FFE8B55F784155EFA2AEBDEAAA2FBEAABA5D",
INIT_24 => X"5D2AAAAAA5D2E820BAA2FBEAB5555557DF55A2AEBDF555D2E954BAA2AA974BAF",
INIT_25 => X"A5D04021EF557FC21FFAA8428BFFAAAA954AAAAAAAAAAAFFD1574105D7FFFF55",
INIT_26 => X"EFF7800215500557DF55AA80001FFAA80001550055575EFFF84021555D043DEA",
INIT_27 => X"B5500517DF555D042AA10A284154005D0015410085568A00FF80175FFA2D17DF",
INIT_28 => X"00000000000000000000000000000000000000005D00020AAAA80020AA082EAA",
INIT_29 => X"D55D2BE800042AFE8E1557D0075D2F45BEAA800AAFFAA9543A080038A2A00000",
INIT_2A => X"0BDEAAA2FBF8AAA557BE8B6D5D5FFABEF49040017D5D20B8EAA007FC51C7A2FB",
INIT_2B => X"0E174BFA02A974BAF7F5EFB455D2ABDF55492AA8BC7EBDFEAFEFFD00105FFBC2",
INIT_2C => X"3D155E105571D55D71C002DABA5524820BAB6FFEFB6D555578F7DB6A0BDF7D48",
INIT_2D => X"092A071555D5E3AE821D00001FF0871C016DBED1FDE90E3A497492B6AAADAAAE",
INIT_2E => X"0E3DA3DFD5E3DFFFBD5A38A021551C5F7AF6DBE8F401D7B6A0001470155C51D0",
INIT_2F => X"82B4002D082082AB8B6D1C5B7DF7FF78E075C5BE8555400550A38428007FED00",
INIT_30 => X"4AA00042AAA2000000000000000000000000000000000000000000000410F450",
INIT_31 => X"AAAA007FD5555AAFBD7545FBB8020A3F7AE975EF005560B55F7AA800AAF7AA95",
INIT_32 => X"E8F5EFF84165EFF7802BAB0A2FFEAABA557BEABEF057D68F5F5A00021EF55042",
INIT_33 => X"52ABFFFF841FFE75CA882108202E974AAF7D57DF55D7AABFF5428ACA8F45A6C1",
INIT_34 => X"84174A8FFAEBFEB0A2D55541051555694F002CA8AA80800020AAF7FBFFFEF045",
INIT_35 => X"7AAA155F595542455512A975455D3AA8A005500151FF0C57401E5F3D1E00A1A8",
INIT_36 => X"5D2A8A0B882FFFFE10AAAAAB755A66B6AF56A2AA801455D7FE8BFFF680800FFF",
INIT_37 => X"00000000000C3BC1000FF8409000512AEABFF5D79FCAF774AE005BE789555400",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000200000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(0),               -- Port A write enable input
DIA(0)   => data_write_a(2),        -- Port A data input
DOA(0)   => data_read_a_hi_512(2),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(0),               -- Port B write enable input
DIB(0)   => data_write_b(2),        -- Port B data input
DOB(0)   => data_read_b_hi_512(2),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_3_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"210C44A20020248B08431120001604B8156023104C4077133420400A02380202",
INIT_01 => X"015A2A424080216D3C2462C99E104B49404040028804A0080A000C16A0D90A0C",
INIT_02 => X"C0A4065000F0A95011000D1501005270B4045AB330860281CC08008222170060",
INIT_03 => X"AD22014098340394A4021320080841C40B411B4298042180002846B06900811A",
INIT_04 => X"244B32A86D20014A0D20403194904900071A24110F0BF400F85F92420E0C946E",
INIT_05 => X"80331030442898B4812840D0500008C528280B063006A64CA30004E5A4E40304",
INIT_06 => X"90016CA00E380042302040A0BC47160424428198C0038C89904E640023600816",
INIT_07 => X"1288020843A66620816049908AA0061011CA0142000009F0A810292E7402F088",
INIT_08 => X"20003C9984A0AC411102014D34EC2200214D5099048823019603A01A49410103",
INIT_09 => X"001CD74C4826220010A8891451284B661CA24A4C899046740121824004100080",
INIT_0A => X"44C9516DC0135C45159BE45F112B48804DC10203021290400772C0F402820D4C",
INIT_0B => X"B400624402404501A49018490184901A4901A4901849018C901A648056480C2D",
INIT_0C => X"D7A9B54000D7C10820680D08C420180381211081A022160000266723E1909021",
INIT_0D => X"400080200E199A4A2CA2994C0399981666409800CA52E4890806BD6B56BDAB52",
INIT_0E => X"40008008E00000000000000000024008000C8000000000400080028000000000",
INIT_0F => X"000A000000588000000000000000200400088000000000400080078000000000",
INIT_10 => X"0000001000004004000D800000000000000000022040000B4000000000000000",
INIT_11 => X"001A0000000000082006C000000000020804087220000122000A000000000000",
INIT_12 => X"00020800B8000000000041002E00000000001040466000000000000001020080",
INIT_13 => X"00000000000000048200004A600000000000000003008000320C000000000000",
INIT_14 => X"432900000222200871028000210400C4000000000000000000080200800030E0",
INIT_15 => X"AF6A5AF6A5AF6A5AF6A5AF6E5AFADA91AB68000101B4D20C08EC461733804A19",
INIT_16 => X"B6B5AF6A5AF6A5AF6A5AF6A5AF6A5AF6A5AB6B5AB6B5AB6B5AB6B5AB6B5AB6B5",
INIT_17 => X"6BDAB6B5A96ADAF6A5AD6ADAF6A5AD6ADAF6A5AD6BDAB6B5A96BDAB6B5A96BDA",
INIT_18 => X"C78C706428A14C586290008A044D54AAB556AA9556AAEBDAB6B5A96BDAB6B5A9",
INIT_19 => X"92492492492492492492492492410410410410412821600001249249015303C0",
INIT_1A => X"351A8D46A351A8D46A351A8D46A351A9D4EA753A9D4EA753A9D4924924924924",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000001543B351A8D46A351A8D46A351A8D46A",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"43DF55FFAA955EFA2D168B55557BEAA000055420000000000000000000000000",
INIT_22 => X"7BE8BFFA2D155410AA8415555087BFFF55A2AA800BAFFAE9554508002AA00AA8",
INIT_23 => X"52ABFEBA007FC21EF007FD75FFAA841541008002AB55AAAA955EF005568A0008",
INIT_24 => X"005168B455D042AB45F7FFD741000042AA10AAAABFF5508003FF555D00021455",
INIT_25 => X"0A2D1575FFF7AA975555D2E80145F78415545082EBDEAAA2FBEAABA5D7FC0155",
INIT_26 => X"55552A954BAFFFFE8B55552EBDE00F7AEAABFFF7FBEAB55F7AABDEBA5D7FC201",
INIT_27 => X"F55A2AEBDF555D2E954BA002EAAABA002A821EF5555554AA087BC01FFFFAAAAB",
INIT_28 => X"0000000000000000000000000000000000000000082E820BAA2FBEAB5555557D",
INIT_29 => X"95578080038A2AA28E3AF55E3A0BA5D7AADB6FB7D5D7FEAA3808554203A00000",
INIT_2A => X"0925D7085F6AA10087FEABD7AAD57AEBAB68E1557D1475FAF45BEAA800AAFFAA",
INIT_2B => X"04AAFFA41040017D5D20B8EAA007FC51C7A2FBD55D7BE80004AA1E8E2AB55B6A",
INIT_2C => X"2FBE80AA557BE8B6D5D5FFABEF49002FB55FFF5D0438140E2FA38B6AEBFF6D1D",
INIT_2D => X"AB8ABAE925D21C7010EADB525D7FFAE975C75D0A901FFFF801557D1C20B8EAAA",
INIT_2E => X"20875C21D5EB8AA8FFF012A954BAFFF5EFB455D20BDE00EBAAA8BC7EBDFEAFEF",
INIT_2F => X"BAB6FFEFB6D555578F7DB6A0BDF7DEB8E125FF002EADA921420871D74971D248",
INIT_30 => X"ABA0051400A20000000000000000000000000000000000000000000001C24820",
INIT_31 => X"8B55F7AA800BAF7AA955EF00042AAA2A2AEAAB55A28408145AAFFFFFFF5D7FEA",
INIT_32 => X"020A35D2ABEF55F7800015F087FEAA00007FEAB55FAD568AA2AFAE975EF55516",
INIT_33 => X"ABFEAAF7AE9DFF759A82AEF70800021EF55042AAAA007FD55558A7BD7145FBB8",
INIT_34 => X"84175EF55002AAB0A2FFEAABA557BEA3EF057968F575D003FF55F7D5420BA5D2",
INIT_35 => X"A8429F45A7D5EAF5FFBAEAAA10554155400AAFFD5145FBAC9755F05040255FFD",
INIT_36 => X"550415557085540000005156155FE90A8F5C082E974AAF7D57DF45552A3FF10A",
INIT_37 => X"00000000005500020AAF7FBFFFEF04552ABFFFF843FFE77C80825BC052ABFE10",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000100000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(0),               -- Port A write enable input
DIA(0)   => data_write_a(3),        -- Port A data input
DOA(0)   => data_read_a_hi_512(3),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(0),               -- Port B write enable input
DIB(0)   => data_write_b(3),        -- Port B data input
DOB(0)   => data_read_b_hi_512(3),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_4_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A108400020612C80284210081034849800A000303100048B3432C82904204002",
INIT_01 => X"21066802000820491C00650E1E004360403008418984014902030906A8D10200",
INIT_02 => X"120404E00E4C0600000206100008402005040C00F104008040080080001310E0",
INIT_03 => X"DCA201514D1C0D706C5CF010083A0708BA0841945004010000080084C1000002",
INIT_04 => X"5C4CF21C48B133483C80417570D000083A62488074C1350EA60D785C0A6B0619",
INIT_05 => X"000F0400028083B381A60001E5546EB5C0E2B81E4166DE000139200004E50940",
INIT_06 => X"80004408020800023000102098000204A040038600018019004B800123208806",
INIT_07 => X"120C20204665E1008024188488800000001A01520000A1F08044892400001088",
INIT_08 => X"0801007AC0A1EB413102063CF3E0B3028D29F407059B0B000205A801C2200102",
INIT_09 => X"106052400922D00406BE1002C6150F41200280001900439001FD8A0004142000",
INIT_0A => X"047F2201D899BA503583504B58AB80804540001202805544314041B48A888EC5",
INIT_0B => X"1441E3443043410C5010C3010C1010C3010C1010C1010C3010C14086980861A5",
INIT_0C => X"020000A02600000805400502C0A0004A00625015000A12000026E1E180011220",
INIT_0D => X"400000000E43930C20C20188120782861E4004A800600401A030001008080400",
INIT_0E => X"40000021A8800000000000000000400800170024000000400000310024000000",
INIT_0F => X"0008000000AA80200800000000002000003400240000004000003B0024000000",
INIT_10 => X"00000010000000040004A080000000000000000020400006C008020000000000",
INIT_11 => X"002C008200000008001B4020200000020000090760000200110A040010000000",
INIT_12 => X"00000803E004040000004000E801040000001000086000000000000000020040",
INIT_13 => X"0000000000000000810000164001008000000000020040002240008020000000",
INIT_14 => X"04001040026026004000000002940040000410000000000000080000400000B8",
INIT_15 => X"040080201004008060000001806AC000004890015124D880100886D8F0014420",
INIT_16 => X"4010000180600000018020100400802010000080601000008020000401802000",
INIT_17 => X"0100000004008020180600000000000180600802010000000401802018020000",
INIT_18 => X"3807E05000140634504048820064B261934D964C326980004010000080600806",
INIT_19 => X"AAAAAAAAAAAAAAAAAAAAAAAAAAA28A28A28A28A2934C8D0CCD145144C0A28A06",
INIT_1A => X"068341A0D068341A0D068341A0D068351A8D46A351A8D46A351AAAAAAAAAAAAA",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000000173F068341A0D068341A0D068341A0D",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"57FE10FFFBEAA10007FD7410FFAA97555082A800AA0000000000000000000000",
INIT_22 => X"7FEAA00007BE8AAAAA843DF55FFAA955EFA2D168B55557BEAB45005542000005",
INIT_23 => X"87BFFF55A2AA800BAFFAE9555508002AA000055574105D2A800AA00043FEBA5D",
INIT_24 => X"A2D17DE1000517FE10AAAAA8AAA002E97545557BC00AAA2FFEAAAAAA84155550",
INIT_25 => X"0A2D157400AAAE974AAAAAA974BA08002AB55A2AA955EF005568A00087BE8BFF",
INIT_26 => X"BA080002145552ABFEAA007FC21EF007FD75FFAA8417410A2D140000F7FBC201",
INIT_27 => X"A10AAAABFF5508003FF55F7D568A00552EA8BEFA2AABDEAA087BEAAAAA2FBD54",
INIT_28 => X"000000000000000000000000000000000000000055042AB45F7FFD741000042A",
INIT_29 => X"EAB7808554203A145178E00FFFBE8A101475D5400F7A49057D0824850B800000",
INIT_2A => X"E8008200043FE925571EFA380871C7028A28E3AF55F7A0925D7AADB6FB7D5D7F",
INIT_2B => X"F5FDA38BE8E1557D1475FAF45BEAA800AAFFAA9557D080038AAA145157428492",
INIT_2C => X"85F6AA10087FEABD7AAD57AEBA08517DE00AAAEA8A9200249056D4175C5092AA",
INIT_2D => X"FEDB42028EBFBC2028BED152438AAA092492AAA4954281C0E2FB55B6A0925D70",
INIT_2E => X"A0875EDA80BEF1C743840040017D5520B8EAA007FC51C7007BD55D7BE80004AA",
INIT_2F => X"55FFF5D0438140E2FA38B6AEBFF6DBE84AAEBAF7DF6AA00412EAABFFAA803DEB",
INIT_30 => X"1EF0800154B200000000000000000000000000000000000000000000041002FB",
INIT_31 => X"0145AAFFFFFEF5D7FEABFF0051400A25D5568A00FFFFEAA105D5155410FF8402",
INIT_32 => X"2AAA25555410BA082E8201000043FE005D517DEBA0851574B2AAAEAAB55F7840",
INIT_33 => X"4001FF005575408AA557FEB2FFAE975EF555168B55F7AA800BAF7AA955EF0004",
INIT_34 => X"2ABFF55F7800015F087FEAA00007FEAB55FAD568AA200557DE00AAAAAAA00080",
INIT_35 => X"87BD6145FAAC000A2A6FBC00BAAAFBC00BAF7D1550AAAA8002010F2AC154B25F",
INIT_36 => X"082EA8BFFAA843FEBA08517DE00F3F9574B30800021EF55042AAAA007FD55550",
INIT_37 => X"000000000008003FF55F7D5420BA5D2ABFEAAF7AEBDFF779A82AA43F7FBE8A00",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000200000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(0),               -- Port A write enable input
DIA(0)   => data_write_a(4),        -- Port A data input
DOA(0)   => data_read_a_hi_512(4),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(0),               -- Port B write enable input
DIB(0)   => data_write_b(4),        -- Port B data input
DOB(0)   => data_read_b_hi_512(4),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_5_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50DF4A0791B3FCB694379283C81FD996A091832102004A337A20E07C0C1E006",
INIT_01 => X"294014468000A04D5C6A60000C34C24841280A00084000C8C212892EEAD53235",
INIT_02 => X"50AE41540CA1D9100002171C1F0A5171134E2A200D8633F8CD09DBFBBB970E7C",
INIT_03 => X"214E3C521D16021B64430CC51C45B8154689094241898749920842946B90010A",
INIT_04 => X"A2F20F7D7A314CB5C208E28A1BF0224A448920028A185340D0C20B2690000C22",
INIT_05 => X"7520B430B20B984809A8886E230C6106371146E1829941C58310402C600381CF",
INIT_06 => X"9CC96CD7C63A7495B9A356ACBC4601C57FD44F8549A46490261C4B39203F7080",
INIT_07 => X"12A88800B029E0C0A12C4B92AA36A2111167357C220095F3C8952A2E5D26F078",
INIT_08 => X"F3F00503B4AE105B534711820C0C0A1043080300F7E0E728B1829C2FEA0A95A1",
INIT_09 => X"C5184F084136848C9298A8560688F480C58858449026145B3830F40944906234",
INIT_0A => X"50EB4124D2B3902BF5C9700C1199DCA84DF46A974F92C7E28F1630D38088A438",
INIT_0B => X"B3144E5636E3178C86B8CC6B8CA6B8CE6B8C86B8CE6B8CA6B8CC15C6435C670C",
INIT_0C => X"79E51E70E070AA8132252008360A7E91504104C8948047D6B0AE1FE440B28A71",
INIT_0D => X"05F0FE40014090400400080329FF8089FF49611F589765923E139F09C78CE7C6",
INIT_0E => X"05F0FE64037FFD7857418407157797878F005F0DFF0F8005F0FE205F0DFF0F80",
INIT_0F => X"8F87FCB1F8053FDEB9B34E0700461E5FF8205F29FF0F8005F0FE205F29FF0F80",
INIT_10 => X"C0184D07C1FF55C3E3E0037FFCF8D3C03009C3CFD53C7E001FF2FAF89781C011",
INIT_11 => X"4E0CDF47186104C6FF177BD939024189BF900401165D645CEEF5BBCDF148F980",
INIT_12 => X"6397F64AEF7F2320483137F8A9BF8A30C2098DFCA06FFFE01F80001F81FDC94F",
INIT_13 => X"FFD051E01015C3BF553D3E0E5FFE838381840714F9DB4F4FA213F774A0E07002",
INIT_14 => X"8B652E2B3120C81284641D3E8DBF7D636FE070189500125C1F83FBCC4F4F80EF",
INIT_15 => X"E7394E339CE138CE5394E33D4E1E0E30E1208C251134921C12A44103F064014B",
INIT_16 => X"7384E3394E338CE538CE1394E3384E738CE139CE1394E7384E339CE139CE5384",
INIT_17 => X"38CE139CE1384E7384E7394E3384E738CE539CE139CE538CE5384E3394E7384E",
INIT_18 => X"7F7B9DB7FF3A1B6DB7ED438A9C3124B2DA6924965B4D384E7384E339CE138CE5",
INIT_19 => X"FBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEF9F7CFDFDDCF3CF3DF5E5BB4E",
INIT_1A => X"7BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEFBEFBEFBEFBE",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE000000000000118D27BBDDEEF77BBDDEEF77BBDDEEF7",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"E955450055421FFFFFBC0010AAD5574BA557FFDFFF0000000000000000000000",
INIT_22 => X"D5575EF55517FF5500557FE10FFFBEAA10007FD7410FFAA97410082A800AAAAA",
INIT_23 => X"FAA955EFA2D168B55557BEAB55005542000007FD74000055574BA5D7FD7555A2",
INIT_24 => X"007BC00AAAAAEBDF45A28428B45FFD168BFF00002AABA5D2ABFFFFAA843DF55F",
INIT_25 => X"AFF80174BAAAD1555EF5555555550055574105D2A800AA00043FEBA5D7FEAA00",
INIT_26 => X"FFAA8415555087BFFF55A2AA800BAFFAE95555080028A00A2FFFDE00F7D57FEB",
INIT_27 => X"545557BC00AAA2FFEAAAA082A97545F7D5420BA5D2E821FFA2D5554BA557BD75",
INIT_28 => X"000000000000000000000000000000000000000000517FE10AAAAA8AAA002E97",
INIT_29 => X"9043D0824850B8A2AE9756D145B401FFFFFFC7010BEDF524AA5571FDFEF00000",
INIT_2A => X"1524BA5571D757DB6D5525EF555178F6D145178E00EBFBE8A101475D5400F7A4",
INIT_2B => X"24BFFFFA28E3AF55F7A0925D7AADB6FB7D5D7FEAB7D0855420BA1471D7438085",
INIT_2C => X"0043FE925571EFA380871C7028B6AEBDF45B68A28B6DEBDF6DBEF1C0A28AAA55",
INIT_2D => X"A2FBF8E10EBD578EAAFF8415482BED1555EF55555057D145152428492E800820",
INIT_2E => X"FB6DF574A85575C55EFBE8E1557D1475FAF45BEAA800AAFFAA9557D080038AAA",
INIT_2F => X"00AAAEA8A9200249056D4175C50920875FDA381C209256DFFDF420BA552A821F",
INIT_30 => X"0BA55557DFF700000000000000000000000000000000000000000000008517DE",
INIT_31 => X"AA105D5155410FF84020AA0800154B2AAAA975FF5D7BC21EFF7FBD7400F7FBC0",
INIT_32 => X"400A25551554BA0051400BA5551575EFF7D1401FF5D5568BE7555568A00AAFFE",
INIT_33 => X"FFDFFF552EA8AAA55043DFF7AAAEAAB55F78400145AAFFFFFEF5D7FEABFF0051",
INIT_34 => X"55400BA082E8201000043FE005D517DEBA0851574B2FFAABFF45FFAAAABFFAAF",
INIT_35 => X"7AA955EF00002AAA2A2FBE8A00A2D16AAAAFF8002410FFD5575EF5555421E755",
INIT_36 => X"FFFFC00BA552A821EFFFFFD74BA5D51575F7FFAE975EF555168B55F7AA800BAF",
INIT_37 => X"000000000000557DE00AAAAAAA000804001FF0055554088A557FEB25D00021FF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000C00000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(0),               -- Port A write enable input
DIA(0)   => data_write_a(5),        -- Port A data input
DOA(0)   => data_read_a_hi_512(5),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(0),               -- Port B write enable input
DIB(0)   => data_write_b(5),        -- Port B data input
DOB(0)   => data_read_b_hi_512(5),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_6_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10800B0061A01002840002C03002818000402322520070B313301C4389B2082",
INIT_01 => X"274008482009404C18A160000C52424841000000090800090210000008510200",
INIT_02 => X"102430600C800110000006100009D070012408000000000648080000001210E0",
INIT_03 => X"000200501D1D02140C420200480140040608010040400104681A0084490C4802",
INIT_04 => X"404402820021000A00824002141000980500000808001114C000080624600600",
INIT_05 => X"120024204209981001A806500304610528000500000080000000300000012940",
INIT_06 => X"2000440832280002300010209C4400142061207A024008900008000220600220",
INIT_07 => X"130C8A220FF41F00902008808800182001020150000001F0800408264000100A",
INIT_08 => X"001BF002C4A01041B1120101000010128568837F04842B080020890008080342",
INIT_09 => X"011847140126805432A62A1596C8B5DF10000008900000100220C00084000008",
INIT_0A => X"44EB4104D09392053589F11C59898888454010830212C54081000410A0088C00",
INIT_0B => X"B0044245B25B456C0096C0096C4096C4096C2096C2096C6096C444B6004B600C",
INIT_0C => X"09040020280010000B3002820110101D0012402CC00802410C26800860070621",
INIT_0D => X"0500819D0000900208201040C4007920004884080000448C281018100C000200",
INIT_0E => X"05008182100000000000000000022AE800C00004000000050081A00004000000",
INIT_0F => X"0002330006000000080000000000000D07A00020000000050081A00020000000",
INIT_10 => X"0000000001204A340002100000000000000000020F4001400000020000000000",
INIT_11 => X"019300020000000068D08000200000001A692121000280000000000010000000",
INIT_12 => X"000201FA100400000000034696010000000000D3478000000000000001003F00",
INIT_13 => X"00000000000000043C0001C0A000008000000000012E000054AC000020000000",
INIT_14 => X"0200000040A410C2810800016000809400001000000000000000433300007600",
INIT_15 => X"060180400000008060180404002AC0200208940041309210B28048180F028000",
INIT_16 => X"2008000100601802000000100601800000000180600800000020180600000000",
INIT_17 => X"0180600000008040100200800000060100000802010040180200002018040100",
INIT_18 => X"7F8FF0F4FA955F7CF7F40A80907638C31C71C718638E00006018040080200004",
INIT_19 => X"38E38E38E38E38E38E38E38E38E38E38E38E38E39B6CEDECDDF7DF7DF5F78BCE",
INIT_1A => X"3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE38E38E38E38E",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFF000000000000196A03F9FCFE7F3F9FCFE7F3F9FCFE7F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"00000000000000000000000C0FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"BFDF45F7AA974AAAAAA97555F784174BAF7D5555FF0000000000000000000000",
INIT_22 => X"FBD7410AA8428AAAAAAE955450055421FFFFFBC0010AAD5574BA557FFDFFF087",
INIT_23 => X"FFBEAA10007FD7410FFAA97400082A800AA08515555508043FE00F7AA97555A2",
INIT_24 => X"55517FF55A2AA97400552AAAB45082E80155F7D1575EFFFAA9555500557FE10F",
INIT_25 => X"FF7AAA8A10082EAAB45A2FFC2000007FD74000055574BA5D7FD7555A2D5575EF",
INIT_26 => X"FFAA843DF55FFAA955EFA2D168B55557BEAB5500554200000003DE10FFD5401F",
INIT_27 => X"BFF00002AABA5D2ABFFFF087BD5545007BFDE10AA803FE105D516AABAFF843FF",
INIT_28 => X"0000000000000000000000000000000000000000AAAEBDF45A28428B45FFD168",
INIT_29 => X"524AA5571FDFEF1C7BFFF55FFA095482B6A49256DEB84104BAFFD1525FF00000",
INIT_2A => X"03DE28F7A49057DAAF5D2428A2842AAAAA2AE9756D145B401FFFFFFC7010BEDF",
INIT_2B => X"A49756D145178E00EBFBE8A101475D5400F7A4904380824850381C5B5057D1C0",
INIT_2C => X"571D757DB6D5525EF555178F6DAAA495428412AAFB451C2A8017DE3DF525FFFF",
INIT_2D => X"1C0E3FE00E3DB471EFE3AAAAA00082EA8B6DA2F1C50381471D74380851524BA5",
INIT_2E => X"049516AAB8FF8428FEFA28E3AF55F7A0925D7AADB6FB7D5D7FEAB7D0855420BA",
INIT_2F => X"45B68A28B6DEBDF6DBEF1C0A28AAA5524BFFFF1C7BD057D1C71FFE10A28038E1",
INIT_30 => X"0AAFFD1401E7000000000000000000000000000000000000000000000B6AEBDF",
INIT_31 => X"21EFF7FBD7400F7FBC00BA55557DFF7557BFDF55F78017400F780001FFAA8400",
INIT_32 => X"154B2557FC01EF55043FEAAFF80021EFA2D1420BAAA8428AA2AAAA975FF5D7BC",
INIT_33 => X"A821EFAAFBC01FFF780155F7555568A00AAFFEAA105D5155410FF84020AA0800",
INIT_34 => X"51554BA0051400BA5551575EFF7D1401FF5D5568BE7AA80174AA082ABDF555D2",
INIT_35 => X"D7FEABFF0051400A25D2EBFE10AAFFD55EFA2AEA8A10082EA8BEFAAD5554B255",
INIT_36 => X"55557DE00AA842AA0000516AABAFF8428BE7AAAEAAB55F78400145AAFFFFFEF5",
INIT_37 => X"0000000000FFAABFF45FFAAAABFFAAFFFDFFF552EA8AAA55043DFF7557BC01EF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000900000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(0),               -- Port A write enable input
DIA(0)   => data_write_a(6),        -- Port A data input
DOA(0)   => data_read_a_hi_512(6),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(0),               -- Port B write enable input
DIB(0)   => data_write_b(6),        -- Port B data input
DOB(0)   => data_read_b_hi_512(6),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_7_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10844B00482258A2842112C02450418800002300500030B313300C418992002",
INIT_01 => X"234008422008604D1C20E0000E11426840000000080000080200090000110204",
INIT_02 => X"1025207000B08910000206101188D03080144880010400044808000000122160",
INIT_03 => X"000200401914821004420000CA01000C0600010000605114291A008449484802",
INIT_04 => X"40440200002100080006500210101019040000000B085024D842080244000000",
INIT_05 => X"1A8024200009981001A8224001040104200204000000800CC2092CE4A0004900",
INIT_06 => X"A000440822280002340010209C040014A061200052500810000C490323208E28",
INIT_07 => X"128802020028000890240980A809102001020140000009F0800408264000100A",
INIT_08 => X"001A0602C4A01051B13281010408881203480200448423199046821008082351",
INIT_09 => X"336784144126811054809C1040140A001C8648481000045903318B80A400310A",
INIT_0A => X"000800009010100014114110312388984502148282A08415B032095048008100",
INIT_0B => X"20CDC1C483484D201192011920119201192051920519205192074C9018C90188",
INIT_0C => X"D8A5B44001D2C12901228F82F005310D293054048A2212004466000DA1908528",
INIT_0D => X"800F8108A0D09802082010408580008000000008C85264010816851B428DA146",
INIT_0E => X"800F81321000020000261900E28A204040E000A0000007800F814000A0000007",
INIT_0F => X"7072024807000020400000581C01C1A406400084000007800F81400084000007",
INIT_10 => X"060180E83800E820101210000200000CC3003C32080201C0000C000000160700",
INIT_11 => X"81DD00804086423120B74020023090644840A34000828800000004000420020B",
INIT_12 => X"1C6A0186E8000446120C8905BA0004810C84624237E00010001878007F0030C0",
INIT_13 => X"00080208E4083C44230201AEE0010040261900E30520C0806EAC0082000984C0",
INIT_14 => X"0121011088A600C032128201519480D40005802448160403E0700622C0806EE8",
INIT_15 => X"A1685A1685A168DA368DA36CDA30DA13A108810111349A943AA4401000928A19",
INIT_16 => X"368DA768DA1685A1685A5685A368DA368DA7685A1685A1685A768DA368DA368D",
INIT_17 => X"685A1685A169DA368DA1685A1695A368DA3685A1685A168DA368DA1685A1685A",
INIT_18 => X"00000000000000000000400A8448410400020820800069DA1685A168DA369DA3",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000003667B000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"0155EFAAAEA8ABAAAFBFDE0055556AA005D04155550000000000000000000000",
INIT_22 => X"556AA00FFAE95555087BFDF45F7AA974AAAAAA97555F784174BAF7D5555FFF78",
INIT_23 => X"055421FFFFFBC0010AAD5574BA557FFDFFF5555555EFAAFFFDFEFAAAAAAB455D",
INIT_24 => X"AA8428AAA557BFDFFF55003DFFFF7FBEAA00002EAAAAA082EA8A00AAAE955450",
INIT_25 => X"0552EBDE00007BEAAAAA2D14000008515555508043FE00F7AA97555A2FBD7410",
INIT_26 => X"FF00557FE10FFFBEAA10007FD7410FFAA97400082A800AAF7AE975FFA2800001",
INIT_27 => X"155F7D1575EFFFAA955555D51574AAAAFFD5545087FEAB455D516AB55557BD55",
INIT_28 => X"0000000000000000000000000000000000000000A2AA97400552AAAB45082E80",
INIT_29 => X"104BAFFD1525FFFF8E175C7A2AAAAA82A2F1FAE105D556AA10410E1755500000",
INIT_2A => X"1FFFD7AAAAAFB7D495F6AA10E3AE905551C7BFFF55FFA095482B6A49256DEB84",
INIT_2B => X"2EAAA00A2AE9756D145B401FFFFFFC7010BEDF524AA5571FDFEF415B575D7AAF",
INIT_2C => X"7A49057DAAF5D2428A2842AAAA497BFAFFF49003AFEFEBFBEAA001C2EA8A821C",
INIT_2D => X"F7A4905C7A28A070384120BDE100075EAA82BEDB470101C5B5057D1C003DE28F",
INIT_2E => X"D555F6AB57417BC05D7145178E00EBFBE8A101475D5400F7A490438082485038",
INIT_2F => X"28412AAFB451C2A8017DE3DF525FFFFA49756D495150492BEF1D2555087BE8B7",
INIT_30 => X"A10002E9754D000000000000000000000000000000000000000000000AAA4954",
INIT_31 => X"7400F780001FFAA84000AAFFD1401E7FFAA97555A2AEA8A10AAD568A00555168",
INIT_32 => X"7DFF7007BD5555AAD57DF55AAAEBDFEF007BE8A10AAAE8215D557BFDF55F7801",
INIT_33 => X"FEAA105D2EAAA005D2AAAA18AAAA975FF5D7BC21EFF7FBD7400F7FBC00BA5555",
INIT_34 => X"7FC01EF55043FEAAFF80021EFA2D1420BAAA8428AA2007FE8BFF080028BFFAAF",
INIT_35 => X"F84020AA0800154B2FF8402145A2AA954AA00043DE0000516AA10F7FBD740855",
INIT_36 => X"FFD140145007FE8BEF557BEAB55087FC215D555568A00AAFFEAA105D5155410F",
INIT_37 => X"0000000000AA80174AA082ABDF555D2A821EFAAFBC01FFF780155F7005140000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000000FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(0),               -- Port A write enable input
DIA(0)   => data_write_a(7),        -- Port A data input
DOA(0)   => data_read_a_hi_512(7),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(0),               -- Port B write enable input
DIB(0)   => data_write_b(7),        -- Port B data input
DOB(0)   => data_read_b_hi_512(7),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_8_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00000648E2840112C00000418000002700500030B3132000400812086",
INIT_01 => X"214009C21838284D042100000212026840000000180800080200080040510204",
INIT_02 => X"1021004000900110000006100088503000240800014400004808000000122160",
INIT_03 => X"0002004019110214044A82000121400C86000000000000860188008448400002",
INIT_04 => X"000402800031200A0000090214100889A5000000490090104800000224000400",
INIT_05 => X"10C025204289981000A820500344010428008500010080080909304040202004",
INIT_06 => X"8000440003280000340010208C04003420600000C6180810000C490703200010",
INIT_07 => X"130002000028000890240980A809012001020050000009F08004082640000082",
INIT_08 => X"20100402C4201041310041010008801201480200051023090024811008090A1A",
INIT_09 => X"0100001001248100308214528148A48008000008100004590711C04034000083",
INIT_0A => X"10804000801210140001C0103001088845010482004000008420041020008900",
INIT_0B => X"0004404002004400448000480004800048000480004800048000440022400200",
INIT_0C => X"880420000880204909004502D100A10C04205424010216010C26800805000004",
INIT_0D => X"8000801100509802082010400400018000488428800004082014000200010000",
INIT_0E => X"8000800A00000207A8BE7B00000200082040808000F07F80008000808000F07F",
INIT_0F => X"0002000402100000404CB1F8FC0000040000808000F07F80008000808000F07F",
INIT_10 => X"3E07800000004004080A000002072C3FCF0000020040804800040007687E3F00",
INIT_11 => X"10800018639EC00020100002C2F9B0000801016001008100000040120CB3067F",
INIT_12 => X"000200020000585EB6000100800030C73D8000402000001FC07FF80001000080",
INIT_13 => X"002EAE1FEC0000040200408000003C547E7B00000100801004000803551F8FC0",
INIT_14 => X"00000000440610C8000A808040000208901B86E568FE0C000000020080100400",
INIT_15 => X"0040100401004090240902449028D0230249850101349A98BAC0481000888810",
INIT_16 => X"0401004010040100401004010240902409024090240902409004010040100401",
INIT_17 => X"4010040100409024090240902409004010040100401004090240902409024090",
INIT_18 => X"543EBC57A10A1E75D6440A889050000000000000000040902409024010040100",
INIT_19 => X"79E79E79E79E79E79E79E79E79E79E79E79E79E7BF3CCD8DF5B2DB2CA4028A0A",
INIT_1A => X"4F87D3E1F4F87D3E1F4F87D3E1F4F87C3E1F0F87C3E1F0F87C3E79E79E79E79E",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000000D3E94F87D3E1F4F87D3E1F4F87D3E1F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"000000087BEAA10F7803DE00FFAEBFFFF0800155FF0000000000000000000000",
INIT_22 => X"7FC2145005155555F780155EFAAAEA8ABAAAFBFDE0055556AA005D0415555080",
INIT_23 => X"7AA974AAAAAA97555F784174BAF7D5555FF552AA8AAA557FC0010F780154105D",
INIT_24 => X"FFAE95555AAFFE8A00552EBFE00F7D17FF45F7FFFFF55AA80155FF087BFDF45F",
INIT_25 => X"5F7D140010552E821EFAAAABDF555555555EFAAFFFDFEFAAAAAAB455D556AA00",
INIT_26 => X"00AAAE955450055421FFFFFBC0010AAD5574BA557FFDFFF5504000AAAAAAA8B5",
INIT_27 => X"A00002EAAAAA082EA8A00002AA8A10F78402155AA8028A00A2D57FF45557BE8A",
INIT_28 => X"0000000000000000000000000000000000000000557BFDFFF55003DFFFF7FBEA",
INIT_29 => X"6AA10410E17555080E000280071E8A00EB8E3FE10F7AEBAFFF080A175D700000",
INIT_2A => X"1C2000FF8A17400557FC015514555757DFF8E175C7A2AAAAA82A2F1FAE105D55",
INIT_2B => X"8A105D71C7BFFF55FFA095482B6A49256DEB84104BAFFD1525FF492EA8AAA557",
INIT_2C => X"AAAAFB7D495F6AA10E3AE90555A2FBE8A38492ABDE10EBDF7AF6DE3FFF8F7DB6",
INIT_2D => X"550E00082B6A0AFB55F7D1420104124821D7AAA0BDF6D415B575D7AAF1FFFD7A",
INIT_2E => X"0B6D578F6D557FFDA00A2AE9756D145B401FFFFFFC7010BEDF524AA5571FDFEF",
INIT_2F => X"FF49003AFEFEBFBEAA001C2EA8A821C2EAAA001C2EA8A00F7800017DA2842FA0",
INIT_30 => X"BEF082E95545000000000000000000000000000000000000000000000497BFAF",
INIT_31 => X"8A10AAD568A00555168A10002E9754D082E820BA08556AA00AAAABFE00F7AEAA",
INIT_32 => X"401E7082EAAABA5D5140010F7AE974105D7BC21555D51575EFFFAA97555A2AEA",
INIT_33 => X"BEABFFAAFBEABFFF7AA80145557BFDF55F78017400F780001FFAA84000AAFFD1",
INIT_34 => X"7BD5555AAD57DF55AAAEBDFEF007BE8A10AAAE8215DA2FFE8ABA082ABFE00AAF",
INIT_35 => X"7FBC00BA55557DFF75D2E82010F7843DF45FFD540000000402145AA843FFFF00",
INIT_36 => X"F780021FFA2803DE10FFD16ABFF5D7BFDE10AAAA975FF5D7BC21EFF7FBD7400F",
INIT_37 => X"0000000000007FE8BFF080028BFFAAFFEAA105D2EAAA005D2AAAA185D2AAAA10",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000400000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(1),               -- Port A write enable input
DIA(0)   => data_write_a(8),        -- Port A data input
DOA(0)   => data_read_a_hi_512(8),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(1),               -- Port B write enable input
DIB(0)   => data_write_b(8),        -- Port B data input
DOB(0)   => data_read_b_hi_512(8),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_9_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000B0001800002840002C0000281800000030000000033022000000000002",
INIT_01 => X"8000098218302849180060000C004240413C0A61590001D90213C90008510200",
INIT_02 => X"000008700CB089100002061031200074810448800104008048080080001210E2",
INIT_03 => X"000200140C1822000A028010408100000628000140402080041A100040024840",
INIT_04 => X"41040000000400080002040200080800040000000B08D1055842080604600700",
INIT_05 => X"10002024000020102400010000026104200004000400800C8B0024E4E0010C40",
INIT_06 => X"8000440802280002700800008A840004A0610000C0000810000C590103600810",
INIT_07 => X"538600220028001890240980A80800200102025000000BF08200002440000883",
INIT_08 => X"00000402C220104131102101040810028528820005100003900E884000010007",
INIT_09 => X"00000005E000000600BCA284140200800C834948100004590111824404012080",
INIT_0A => X"04080000901012100A1141005922000245410002008880000032005080000800",
INIT_0B => X"2000020040044010440104401004010440100401044010040104400802008208",
INIT_0C => X"D1A1344420D2E100000808000000000481000000202002400006800825908402",
INIT_0D => X"0500000000109000000000000580008000080000C852240100068D0B4685A342",
INIT_0E => X"0500000A00000000000000000000028000408020000000050000208020000000",
INIT_0F => X"0000304002100020000000000000000900208004000000050000208004000000",
INIT_10 => X"0000000001200000000A00000000000000000000050000480008000000000000",
INIT_11 => X"009F0080000000004807C0200000000012000020000081000000040000000000",
INIT_12 => X"00000048F8000400000002403E0004000000009067E000000000000000000900",
INIT_13 => X"0000000000000000140000CEE001000000000000000A000036AC008000000000",
INIT_14 => X"03210000000400CA81000000619480D4000400000000000000004100000036E8",
INIT_15 => X"A368DA368DA3685A1685A1685A121A11A1419001512490040024001000008019",
INIT_16 => X"1685A1685A1685A1685A1685A368DA368DA368DA368DA368DA368DA368DA368D",
INIT_17 => X"685A1685A168DA368DA368DA368DA368DA368DA368DA3685A1685A1685A1685A",
INIT_18 => X"CCF48DE68A895C38E250080000000000000000000000685A1685A1685A1685A1",
INIT_19 => X"514514514514514514514514514D34D34D34D34D28E10040392482090157344C",
INIT_1A => X"4D268341A0D069349A0D069349A0D068341A0D068341A0D06834514514514514",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000001654D0D069349A0D068341A4D268341A",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"BE8B45002A974AAAA803DFFFAA843DF45FFFFEAABA0000000000000000000000",
INIT_22 => X"AEBDE00AAFBEAABA080000000087BEAA10F7803DE00FFAEBFFFF0800155FFAAF",
INIT_23 => X"AAEA8ABAAAFBFDE0055556AA005D0415555087BFDE00A2FBD7400F7FBFDFFFA2",
INIT_24 => X"005155555557BE8BEF007FFDEAAAAD1555EF0055401FFF7AEAAA10F780155EFA",
INIT_25 => X"0F7AA974AA082E80010A2AAAAA10552AA8AAA557FC0010F780154105D7FC2145",
INIT_26 => X"BA087BFDF45F7AA974AAAAAA97555F784174BAF7D5555FFF780154AA5D2AA8A1",
INIT_27 => X"F45F7FFFFF55AA80155FF080400145FFFBEAABAF7D17FEBAA2AEBDF45002EAAA",
INIT_28 => X"0000000000000000000000000000000000000000AAFFE8A00552EBFE00F7D17F",
INIT_29 => X"BAFFF080A175D7BEF1E8B6D002090482B68E38FC7BE8A3DF7DF7F5E8A9200000",
INIT_2A => X"BD0400FFF5FDFC7B6A0BDE38B6F5E8A92080E000280071E8A00EB8E3FE10F7AE",
INIT_2B => X"AAA8A38FF8E175C7A2AAAAA82A2F1FAE105D556AA10410E175550871FFE00A2F",
INIT_2C => X"F8A17400557FC015514555757D5D71E8BEF147BFAE82A2DB555C71C5B451D7FF",
INIT_2D => X"FF84174BA5D20AAA00E3AA904BA142A87010A2AEADA38492EA8AAA5571C2000F",
INIT_2E => X"AAAA0BFF7D0024ADA921C7BFFF55FFA095482B6A49256DEB84104BAFFD1525FF",
INIT_2F => X"38492ABDE10EBDF7AF6DE3FFF8F7DB68A105D7000400155FFFBEDA82FFD57DEB",
INIT_30 => X"FEFF7D16AA00000000000000000000000000000000000000000000000A2FBE8A",
INIT_31 => X"AA00AAAABFE00F7AEAABEF082E95545F7D568BEF080402000F7AAA8B55FFAABD",
INIT_32 => X"9754D00517DE00A2FFC2000F7D17FF55FF803FEAAFFD16AA00082E820BA08556",
INIT_33 => X"FD55555D7FD5555FFAAA8AAAFFAA97555A2AEA8A10AAD568A00555168A10002E",
INIT_34 => X"2EAAABA5D5140010F7AE974105D7BC21555D51575EF555568BEF5D7FE8A10AAF",
INIT_35 => X"A84000AAFFD1401E7FF80174AA5D0028A00AAAE800AA552A97400A2AEBDEAA08",
INIT_36 => X"F7FBFFE00FFD17FEAAA2803DFEF08043FE00557BFDF55F78017400F780001FFA",
INIT_37 => X"0000000000A2FFE8ABA082ABFE00AAFBEABFFAAFBEABFFF7AA80145080002145",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000800000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(1),               -- Port A write enable input
DIA(0)   => data_write_a(9),        -- Port A data input
DOA(0)   => data_read_a_hi_512(9),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(1),               -- Port B write enable input
DIB(0)   => data_write_b(9),        -- Port B data input
DOB(0)   => data_read_b_hi_512(9),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_10_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000B0001800002840002C0000281800020030000000033022000000180006",
INIT_01 => X"000008000000004C002000000010026840000000080000080200000000110200",
INIT_02 => X"0000004000800110000006100000003000040800010400004808000000120060",
INIT_03 => X"000200000810020000020000400100000600000000400000001A000040004800",
INIT_04 => X"0004000000000008000200020000000004000000080010004000000200000000",
INIT_05 => X"1000202000011010000000000000010520000400000080000000200000200004",
INIT_06 => X"80004408022800023000000088040004A061000040000810000C490103600000",
INIT_07 => X"120420020028000890240980A808002001020050000009F08000002440000082",
INIT_08 => X"00000402C0201051311001000000020201080200440400000000800000000000",
INIT_09 => X"0000105808000000000000000000008000008088100004590111800004000000",
INIT_0A => X"00804000801210440003C1411008800045000002000014000040009002800000",
INIT_0B => X"0400200000000000000004000040000000000000040000400000000000000221",
INIT_0C => X"0100802000000000000002802000000400100000000002000026000840011400",
INIT_0D => X"0500000000409002082010400400008000400008002044082000081004080204",
INIT_0E => X"0500000200000000000000000000028000400000000000050000200000000000",
INIT_0F => X"0000304002000000000000000000000900200000000000050000200000000000",
INIT_10 => X"0000000001200000000200000000000000000000050000400000000000000000",
INIT_11 => X"0082000000000000480080000000000012000101000080000000000000000000",
INIT_12 => X"0000004810000000000002400400000000000090400000000000000000000940",
INIT_13 => X"0000000000000000150000C00000000000000000000A40001400000000000000",
INIT_14 => X"02000000002400C2810000006000000000000000000000000000410040001400",
INIT_15 => X"020080200802008020080200800800220200840001309A08A848001000008000",
INIT_16 => X"0000000000000000000000000200802008020080200802008020080200802008",
INIT_17 => X"0080200802000000000000000000000000000000000000000000000000000000",
INIT_18 => X"940FE0D397124355520542821010000000000000000000802008020080200802",
INIT_19 => X"28A28A28A28A28A28A28A28A28A28A28A28A28A29554199854514514F546890A",
INIT_1A => X"32994CA6532995CAE572B94CA6532994CA6532994CA6532994CA28A28A28A28A",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000001867172B94CA6532994CA6572B95CAE5",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FC2155F7D155545AA80001EFAAFBEAB45557FFDE100000000000000000000000",
INIT_22 => X"FBE8BFFF78402155AAFBE8B45002A974AAAA803DFFFAA843DF45FFFFEAABA007",
INIT_23 => X"87BEAA10F7803DE00FFAEBFFFF0800155FF00042AB55FFD168B55AA8000010FF",
INIT_24 => X"AAFBEAABAA2FFD741055003DFEFF7AA801FFAAD16AABA002ABDE100800000000",
INIT_25 => X"FF7FBC0145F78028A00A2D142155087BFDE00A2FBD7400F7FBFDFFFA2AEBDE00",
INIT_26 => X"BAF780155EFAAAEA8ABAAAFBFDE0055556AA005D0415555007FD74105555555E",
INIT_27 => X"5EF0055401FFF7AEAAA105D042ABFF5D556AB55AAD168ABA002A975FFF7AEBDE",
INIT_28 => X"0000000000000000000000000000000000000000557BE8BEF007FFDEAAAAD155",
INIT_29 => X"3DF7DF7F5E8A92007BC217DEBDB55555AA8E071D7AAFBEFB455D71F8E0000000",
INIT_2A => X"B6DB55BE8E05000EBFFE8BC7E38E07145BEF1E8B6D002090482B68E38FC7BE8A",
INIT_2B => X"2EB8E00080E000280071E8A00EB8E3FE10F7AEBAFFF080A175D700042AB7DEBD",
INIT_2C => X"FF5FDFC7B6A0BDE38B6F5E8A92B6FBD5410490A3DFD7F7A4821D7A2D16FA8214",
INIT_2D => X"0071D54104951555D7EBF5C5155E3842AA00BED1421450871FFE00A2FBD0400F",
INIT_2E => X"20820955EFE3AEBDEAAFF8E175C7A2AAAAA82A2F1FAE105D556AA10410E17555",
INIT_2F => X"EF147BFAE82A2DB555C71C5B451D7FFAAA8A38410E2ABD749516FB55BED16FA8",
INIT_30 => X"F455D556AA000000000000000000000000000000000000000000000005D71E8B",
INIT_31 => X"2000F7AAA8B55FFAABDFEFF7D16AA00087FC01EFA2FFD7545AAAE97555A2FBFD",
INIT_32 => X"9554500042ABFFA2FFFFF45F7AE97400AAFFE8B45AAAA95545F7D568BEF08040",
INIT_33 => X"400155A2D57FE00552EA8A00082E820BA08556AA00AAAABFE00F7AEAABEF082E",
INIT_34 => X"517DE00A2FFC2000F7D17FF55FF803FEAAFFD16AA00FFFBD5400082EBFF45F78",
INIT_35 => X"55168A10002E9754D085155410085557555AAD557555A2802AA10FFD54214500",
INIT_36 => X"08557DF55F7D17FE000804155FFAAAABDEAAFFAA97555A2AEA8A10AAD568A005",
INIT_37 => X"0000000000555568BEF5D7FE8A10AAFFD55555D7FD5555FFAAA8AAA002AAAB45",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000008FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(1),               -- Port A write enable input
DIA(0)   => data_write_a(10),        -- Port A data input
DOA(0)   => data_read_a_hi_512(10),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(1),               -- Port B write enable input
DIB(0)   => data_write_b(10),        -- Port B data input
DOB(0)   => data_read_b_hi_512(10),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_11_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10180B05A0010402840602C2D001019000000300000000330A20080EC180002",
INIT_01 => X"AB400986B830284D1820E0000C3642484000000008000008820009080A512220",
INIT_02 => X"102A68440080011000000618062AD03502640800010410424908136019920868",
INIT_03 => X"004A0846191B22120642000442C110044600000101E9225CDC9A10844A9A4842",
INIT_04 => X"0094024000250808800216021138000B848000000800100040000102A0600200",
INIT_05 => X"7E4024242008A8102CA88A44010401042200444000888000000028000002A002",
INIT_06 => X"8088445712280000B18812288E0400253855200045C86810000C5B0503286A28",
INIT_07 => X"10008822A028004880200A80880208200122006C000015F0C20408264902C840",
INIT_08 => X"9390040280241041D1754100000018108728820024002B3A01A89540080824C8",
INIT_09 => X"A1001C41A1348498B080801010000080D00301081000045B0511D28D94012339",
INIT_0A => X"44080000901012428003414158230CBA4576708241C010908040341322008000",
INIT_0B => X"040464D280144050C72A0872A0C72A0872A0C72A0C72A0872A0C595043950421",
INIT_0C => X"0804001400000820110A42822204880CD81040442900021704E6000800001D54",
INIT_0D => X"80C62D0500409002082010404580018000404012004004192C10000000000000",
INIT_0E => X"80C62D5803161C526DB40506C120A806ABB0D808CC334A80A54B70D408CC32D2",
INIT_0F => X"2B5144D0DD903C54916D15458C0513005570D408CC334A80A54B70D808CC32D2",
INIT_10 => X"52148C4DB05621E363F813961C20EDA944016558C2347A080B10D8DD6422AA10",
INIT_11 => X"1880144D3345C65593800319C18BD1ECA1C9010112566F10AC4183C340DAE02D",
INIT_12 => X"5810503000633830DE3C2C9C00289A66AA8DE50E0800360614AC281430890600",
INIT_13 => X"0CD2A9CEA8199B6B082B55900314140365320485C4F00AD544407241C175C402",
INIT_14 => X"0000074044C4801832701A89D20A38093631425969020855A281844E00540404",
INIT_15 => X"0000000000000000000000000020C00200088101513492101280401000400200",
INIT_16 => X"2008020080200802008020080000000000000000000000000000000000000000",
INIT_17 => X"0080200802008020080200802008020080200802008020080200802008020080",
INIT_18 => X"804180C0B10A4210420140028400000000000000000000802008020080200802",
INIT_19 => X"000000000000000000000000000820820820820801C414947000000055062608",
INIT_1A => X"0000000004020000000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000001F87E000000000000010080000000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"ABDF5508557DF45002ABDFFFF7803DE10AA80000AA0000000000000000000000",
INIT_22 => X"FFE8A10A28000000007FC2155F7D155545AA80001EFAAFBEAB45557FFDE10082",
INIT_23 => X"02A974AAAA803DFFFAA843DF45FFFFEAABAA2AEBFF45FFAEBFEAA002A801FFF7",
INIT_24 => X"F78402155AAD155555A28428BFF002ABDE00A2AABFE10082ABFFEFAAFBE8B450",
INIT_25 => X"0002A80010A2842AAAA007BFFF4500042AB55FFD168B55AA8000010FFFBE8BFF",
INIT_26 => X"00080000000087BEAA10F7803DE00FFAEBFFFF0800155FF00557FF45557FC201",
INIT_27 => X"1FFAAD16AABA002ABDE10A2D168A10A284021FF5D00154BAF7FBE8BEFFFD5400",
INIT_28 => X"0000000000000000000000000000000000000000A2FFD741055003DFEFF7AA80",
INIT_29 => X"EFB455D71F8E00002EBDF6D005B78F7D142ABDFC7F78E3FE28B684070AA00000",
INIT_2A => X"0BDEAA1C2A801C7E3FFEFA10B68407038007BC217DEBDB55555AA8E071D7AAFB",
INIT_2B => X"20B8FEFBEF1E8B6D002090482B68E38FC7BE8A3DF7DF7F5E8A92BEAEBFF7DEBA",
INIT_2C => X"E8E05000EBFFE8BC7E38E07145B6D15756DA28A28BFF082ABAE10B6AAB8E2808",
INIT_2D => X"08517DF7D497BC5028142A87000A28A2AA92007FF8F7D00042AB7DEBDB6DB55B",
INIT_2E => X"2FFFFEFBC7E3DF42028080E000280071E8A00EB8E3FE10F7AEBAFFF080A175D7",
INIT_2F => X"10490A3DFD7F7A4821D7A2D16FA82142EB8E00B6DB6AA28A280001FF5D0A1048",
INIT_30 => X"EAAF784154BA000000000000000000000000000000000000000000000B6FBD54",
INIT_31 => X"7545AAAE97555A2FBFDF455D556AA00082EBFFEF007BE8BFF5D2ABDF55F7AABD",
INIT_32 => X"6AA00FFAEBFFEFAA803DEBA5D2E82155A2FBFDE00FF84154BA087FC01EFA2FFD",
INIT_33 => X"AAAA00FFAAA8AAA080028BFFF7D568BEF080402000F7AAA8B55FFAABDFEFF7D1",
INIT_34 => X"042ABFFA2FFFFF45F7AE97400AAFFE8B45AAAA95545F7D5555FFAAAAA8BFF002",
INIT_35 => X"7AEAABEF082E9554508557DFFF007BD54BA5D2E95400A2AEA8A00007FEABFF00",
INIT_36 => X"AA80001FF5D2E82000F7FFFFF45AAFFC20BA082E820BA08556AA00AAAABFE00F",
INIT_37 => X"0000000000FFFBD5400082EBFF45F78400155A2D57FE00552EA8A00FFFFE8AAA",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000800000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(1),               -- Port A write enable input
DIA(0)   => data_write_a(11),        -- Port A data input
DOA(0)   => data_read_a_hi_512(11),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(1),               -- Port B write enable input
DIB(0)   => data_write_b(11),        -- Port B data input
DOB(0)   => data_read_b_hi_512(11),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_12_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A500C4B01BC0268A6940312C0DE045196A831A300500032B333287E4FC812006",
INIT_01 => X"AF400D869830E84D5823E0000C1742484000000008000008820009280A553235",
INIT_02 => X"502A7144008001100000171C022BD13412762A000586235ECC09C8423B960866",
INIT_03 => X"31863846191BA218064204000281200406A10843010022DEDF0852944A9C014A",
INIT_04 => X"0014030000250409000014821038080B840000400800102040000302F0600233",
INIT_05 => X"7FC034348008A8102CA88F48010601042400048000188000000938000002E088",
INIT_06 => X"9CC96CC6F63A5001F12B56A0AC8601F47AC06400D1F80C10020C493F03343A38",
INIT_07 => X"1020002030280098A12048908A16BA311177124C000003F08A94282E5C262861",
INIT_08 => X"827A0602902A10491165E10000049010C52882008600A73A01E8974008092CF8",
INIT_09 => X"47000001A1248008F000000000000080000F010C100204593F11A6CDF48023BF",
INIT_0A => X"040000208010120ACA01400058010CBA4D277C86CCE802B380003C1360008000",
INIT_0B => X"011C46D3C7BC1EF083AF0C3AF083AF083AF0C3AF083AF083AF0C1D7861D78400",
INIT_0C => X"08040014C9001AE91D17E50AD79FEFC87C2154745F82131FFCCE00080000095E",
INIT_0D => X"807BF7118180984004000803D40001880001001400C005031010000000000000",
INIT_0E => X"807BF76A109C944B5891BF06C5EEB14FCBF0D90076D61C807BF7D0D80876D49C",
INIT_0F => X"6DE38EB9FB10350C00A99F7CA80757365E50D80876D61C807BF7D0D90076D49C",
INIT_10 => X"841BCC69A0D8C6F7F0AA001C943A65756A0976EB5A7E7FC8951018186334F311",
INIT_11 => X"D5A014481991C6A737D80211912970CDCDD1864116D6C7080651CB4661F33615",
INIT_12 => X"349E929300423224AE19B9BEC0289033238D4E6EA805892946A9B011A7B152CF",
INIT_13 => X"6244CD7AC01CAAA56B3E6D9001068715D64006D2A961CF9B44512A2504532182",
INIT_14 => X"00000439FDC25C58067A9FAB46095A0B5289A0282D2E1444ACB12A17CF9B4414",
INIT_15 => X"0000000000000000000000040026C00000288401513492909280401000F70A00",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"088881360A95090CB05442029010000000000000000000000000000000000000",
INIT_19 => X"1041041041041041041041041049249249249249200100002D4514510051B946",
INIT_1A => X"592C964B2592C964B2592C964B2592C86432190C86432190C864104104104104",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000002007F592C964B2592C964B2592C964B2",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"43FE0008557DFFF0800020105D557FEAA00557DE100000000000000000000000",
INIT_22 => X"557DFFFF7AA80000082ABDF5508557DF45002ABDFFFF7803DE10AA80000AAAA8",
INIT_23 => X"7D155545AA80001EFAAFBEAB45557FFDE10AAD5420000051555FFA2AA8200000",
INIT_24 => X"A28000000A2D155410F7FFFFEBA08003FE00082AA8AAAAAFFC00BA007FC2155F",
INIT_25 => X"0A2AABFE1055516ABEF5D517DEAAA2AEBFF45FFAEBFEAA002A801FFF7FFE8A10",
INIT_26 => X"55AAFBE8B45002A974AAAA803DFFFAA843DF45FFFFEAABA000028A105D2ABFE1",
INIT_27 => X"E00A2AABFE10082ABFFEF085542000000417555002A820AA08557DFFFF7AA821",
INIT_28 => X"0000000000000000000000000000000000000000AAD155555A28428BFF002ABD",
INIT_29 => X"3FE28B684070AABE803AE38145B78FD7000005010495B7AE921C517DE1000000",
INIT_2A => X"B505FFB6A487000005F7AFD7F7A482038002EBDF6D005B78F7D142ABDFC7F78E",
INIT_2B => X"F5C2082007BC217DEBDB55555AA8E071D7AAFBEFB455D71F8E00BED547038145",
INIT_2C => X"C2A801C7E3FFEFA10B68407038B6D550428FFF1FDE821C003FE001C2EAAAAAB6",
INIT_2D => X"00002FA285D20BDE28A2A4B8E10555B68BEF5D517DEAABEAEBFF7DEBA0BDEAA1",
INIT_2E => X"2005F7DFD7F7A482155BEF1E8B6D002090482B68E38FC7BE8A3DF7DF7F5E8A92",
INIT_2F => X"6DA28A28BFF082ABAE10B6AAB8E280820B8FEF085F4703814001055514208208",
INIT_30 => X"A0055517DE00000000000000000000000000000000000000000000000B6D1575",
INIT_31 => X"8BFF5D2ABDF55F7AABDEAAF784154BAF7802AABA5D7FEAB45080015410007FEA",
INIT_32 => X"6AA00F7D1554BA5D7BC01FFFF8015410007FEAB45F780020BA082EBFFEF007BE",
INIT_33 => X"43FE10552EAAAAAFFD140000087FC01EFA2FFD7545AAAE97555A2FBFDF455D55",
INIT_34 => X"AEBFFEFAA803DEBA5D2E82155A2FBFDE00FF84154BAF7D1400BAFFD57FE005D0",
INIT_35 => X"FAABDFEFF7D16AA0008003FEBA55003DEBAA28428A105D7FEABEF55557DEBAFF",
INIT_36 => X"550402145550000010087FFFF45F78402145F7D568BEF080402000F7AAA8B55F",
INIT_37 => X"0000000000F7D5555FFAAAAA8BFF002AAAA00FFAAA8AAA080028BFF087BD54AA",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000000FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(1),               -- Port A write enable input
DIA(0)   => data_write_a(12),        -- Port A data input
DOA(0)   => data_read_a_hi_512(12),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(1),               -- Port B write enable input
DIB(0)   => data_write_b(12),        -- Port B data input
DOB(0)   => data_read_b_hi_512(12),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_13_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10110A0441812402840402822007818000E00700000000330A3000000008042",
INIT_01 => X"A1400984B830C848180260000C0042604001000008220008A200100802110200",
INIT_02 => X"10A00860009141100000C6180C285035000E0800010431004908135980120C60",
INIT_03 => X"004E20441910221B06420C85D5013804060000000040324C441A108468024842",
INIT_04 => X"0184034010250089C00EA8021938325B04800002091090014880080200000900",
INIT_05 => X"18002424B008881024A8004E01040104270004E0000080090500604840000481",
INIT_06 => X"80004414022A2490B00A142C8C840005794540015E006810001C4B01032C7E20",
INIT_07 => X"510200028028004880280A808816002101022468000011F082040A264006C000",
INIT_08 => X"D2B00402B220104B531001000008001041080200B660E30B200C8040080A9206",
INIT_09 => X"A1000809A93484D21000000000000080C90391881000145B0111A30404015000",
INIT_0A => X"000000008010102A82014100101118BA4510008241480290882400900000A000",
INIT_0B => X"0284484000000000400000000040000000000000040000000000000020000000",
INIT_0C => X"A944AA2000A02000212800020000000D80004084A0000390002E001843210400",
INIT_0D => X"859C1881A04090000000000021800180010341179065441356150A1285094284",
INIT_0E => X"859C188810C65A72A617520252781EA02520D589B9A260859C1840DD81B9A0E0",
INIT_0F => X"0E71F1052D942748C19484E39442D15961C0DD81B9A260859C1840D589B9A0E0",
INIT_10 => X"E60605C0C12CBD400B0810C65A61AA459D0047398500D5889D26907356533C00",
INIT_11 => X"8F60CA1562094650CA28398A42C051E0332181010109294C8E1160CB8C80A561",
INIT_12 => X"2645056D073148580A3C065141942AC4128CA199180C5232575138094450AD0A",
INIT_13 => X"84CA93A2FC008962142B17301A9A1A5196A80245208E0AC5C853C8028163B8C0",
INIT_14 => X"0240034000E4DC8A84000014982372011FC1E475F0F0084A3961F5A80AC5C816",
INIT_15 => X"4250942509425094250942509428D421420882020120981812C8403000088212",
INIT_16 => X"2509425094250942509425094250942509425094250942509425094250942509",
INIT_17 => X"5094250942509425094250942509425094250942509425094250942509425094",
INIT_18 => X"FF3F7DF7FF3E9F7DF7E24502A800000000000000000050942509425094250942",
INIT_19 => X"EBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBF7DFDFDDD555555F7EFBBEE",
INIT_1A => X"7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAEBAEBAEBAEBA",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000000007F7EBF5FAFD7EBF5FAFD7EBF5FAFD",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5554BA087FFFF55557BD54AAF7FBC01FFA2802ABEF0000000000000000000000",
INIT_22 => X"2E80155AA802AB45AA843FE0008557DFFF0800020105D557FEAA00557DE10AAD",
INIT_23 => X"8557DF45002ABDFFFF7803DE10AA80000AA087BD75EF087FFFFEF557BEAB4555",
INIT_24 => X"F7AA80000AAD1420AA087BD7555FFD168AAAFFAE820AA5D5557555082ABDF550",
INIT_25 => X"5FFD157555085140010F7AEAABFFAAD5420000051555FFA2AA8200000557DFFF",
INIT_26 => X"45007FC2155F7D155545AA80001EFAAFBEAB45557FFDE10AAAEA8BFFA2FBD754",
INIT_27 => X"E00082AA8AAAAAFFC00BA00002AAAAF7D5574BA557BE8A10A284154BAFFAAAAB",
INIT_28 => X"0000000000000000000000000000000000000000A2D155410F7FFFFEBA08003F",
INIT_29 => X"7AE921C517DE10A2DB50482147FFAF554971D0492E3F1C71C7BE8A2ABD700000",
INIT_2A => X"FFAFD7497BE8B5555208217DBE8A2AB45BE803AE38145B78FD7000005010495B",
INIT_2B => X"5F5056D002EBDF6D005B78F7D142ABDFC7F78E3FE28B684070AA1C71D25D7007",
INIT_2C => X"6A487000005F7AFD7F7A482038AADF47092147FD257DFFD568A82FFA4870BA55",
INIT_2D => X"A2A0ADBC7A2FFD257DE3DF52555085142000FFAAAFBFFBED547038145B505FFB",
INIT_2E => X"0B680124BAFFAAAFB45007BC217DEBDB55555AA8E071D7AAFBEFB455D71F8E00",
INIT_2F => X"28FFF1FDE821C003FE001C2EAAAAAB6F5C20821C002AA92FFDF574824171EAA1",
INIT_30 => X"545F7AEA8B55000000000000000000000000000000000000000000000B6D5504",
INIT_31 => X"AB45080015410007FEAA0055517DE00A2FFC00105D7BE8B55085142010AAD157",
INIT_32 => X"154BA5D5140145007BE8B55087BEAB555D04001EFF7AAA8B55F7802AABA5D7FE",
INIT_33 => X"16AA10FF80174AA557FC21EF082EBFFEF007BE8BFF5D2ABDF55F7AABDEAAF784",
INIT_34 => X"D1554BA5D7BC01FFFF8015410007FEAB45F780020BAA2FFD54105D7FC21EFFFD",
INIT_35 => X"2FBFDF455D556AA00A2803FF45AAFFC21EFAAFBC0155085540000FFAEBFFEFF7",
INIT_36 => X"F7FBD5410085568A10FF80020AAFFAABFF55087FC01EFA2FFD7545AAAE97555A",
INIT_37 => X"0000000000F7D1400BAFFD57FE005D043FE10552EAAAAAFFD1400005D042AA00",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000CFFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(1),               -- Port A write enable input
DIA(0)   => data_write_a(13),        -- Port A data input
DOA(0)   => data_read_a_hi_512(13),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(1),               -- Port B write enable input
DIB(0)   => data_write_b(13),        -- Port B data input
DOB(0)   => data_read_b_hi_512(13),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_14_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10020A000180000284008280000281800000030000000033022000000580002",
INIT_01 => X"A140098018300848184860000C20C24040000000084000084200000000110200",
INIT_02 => X"1020006000900110000006102028503400040800010400204908012018120E64",
INIT_03 => X"000200441910221006420000400100040600000000E9E401209A108448004842",
INIT_04 => X"0004020000250008000200021038000804000000090090004800080200000000",
INIT_05 => X"500024240008881024A800400104010420000400000080080100204040000000",
INIT_06 => X"8000440102282015B10A10288E0400042345400040006810000C5901033D7880",
INIT_07 => X"1100000200280048802008828812002001220064000005F1C2850A2649204070",
INIT_08 => X"00B00402802010411110010000080010010802000400230B000C804008080002",
INIT_09 => X"01000009A92480001000000000000080C8038188100004590111B68404010000",
INIT_0A => X"0000000080101000000141001001088A45000082400000008020009000008000",
INIT_0B => X"0004404000000000400004000000000000004000000000000004000000000000",
INIT_0C => X"8904A0200080200001080002000000088000400420000200002E000841010400",
INIT_0D => X"0500000C80409000000000000000018000000000806044010014081204090204",
INIT_0E => X"0500005813A0210D072E8D012001028402908004000587050000108004000707",
INIT_0F => X"9004300044900812386A280E5800088980108020000587050000108020000707",
INIT_10 => X"DE00482E19E30002007813A02096038AE200880405200308828062A68C0BC700",
INIT_11 => X"00000E5A08E6000048001292B83280001208A1011004011060049A1C59192055",
INIT_12 => X"492060480256530650000240001DB011CC00009000032C4C979E3806180C0900",
INIT_13 => X"5A3433EDE00154181400000007BCBD858F120120541A0000000033757465B2C0",
INIT_14 => X"02002C000024008A84001A0902000422E3E99681004802115652594000000001",
INIT_15 => X"0240902409024090240902409028D021020880000120901812C8401000000210",
INIT_16 => X"2409024090240902409024090240902409024090240902409024090240902409",
INIT_17 => X"4090240902409024090240902409024090240902409024090240902409024090",
INIT_18 => X"5C8FF0F7BE9D5F7DF65040028000000000000000000040902409024090240902",
INIT_19 => X"79E79E79E79E79E79E79E79E79E79E79E79E79E7BF7DDDDDFCF3CF3DF5579B4E",
INIT_1A => X"3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE79E79E79E79E",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000003FF803F9FCFE7F3F9FCFE7F3F9FCFE7F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"BE8B55A2AE80000F7D5555555D2AAAABAAAD1420BA0000000000000000000000",
INIT_22 => X"00155EF0804155EFAAD5554BA087FFFF55557BD54AAF7FBC01FFA2802ABEFA2F",
INIT_23 => X"8557DFFF0800020105D557FEAA00557DE10A2AA801FFA28402000AAAE9554555",
INIT_24 => X"AA802AB4500516AA00A2AE800BAFFFFC20BAF7AEA8B45080417400AA843FE000",
INIT_25 => X"0A2843FEBAFFFBD7410A2D168BFF087BD75EF087FFFFEF557BEAB45552E80155",
INIT_26 => X"AA082ABDF5508557DF45002ABDFFFF7803DE10AA80000AA005568ABAA2840201",
INIT_27 => X"AAAFFAE820AA5D5557555002E80155A280000005D7FFDF4555517DFEF00043FE",
INIT_28 => X"0000000000000000000000000000000000000000AAD1420AA087BD7555FFD168",
INIT_29 => X"C71C7BE8A2ABD7A2FFEDB55B6A080038E3DB50555412AA8ABAAADB4009200000",
INIT_2A => X"402038AAAA955554900105FF0800175D7A2DB50482147FFAF554971D0492E3F1",
INIT_2B => X"0A12410BE803AE38145B78FD7000005010495B7AE921C517DE10A2AE851FFB68",
INIT_2C => X"97BE8B5555208217DBE8A2AB451C556FA00A2A0800BAE3F1C0092EBAAADB6D08",
INIT_2D => X"00516DABAA28402038B6803DE82F7F5D5410A2D568BC71C71D25D7007FFAFD74",
INIT_2E => X"55D5F78FD7000E3FEAA002EBDF6D005B78F7D142ABDFC7F78E3FE28B684070AA",
INIT_2F => X"92147FD257DFFD568A82FFA4870BA555F5056D002A80155B680000105D7FF8F4",
INIT_30 => X"AAAAAFFC2000000000000000000000000000000000000000000000000AADF470",
INIT_31 => X"8B55085142010AAD157545F7AEA8B55A2FBFFF55FF84000AAAAFBC0145002AA8",
INIT_32 => X"7DE00A2AA955FFFF80020BAAAAA975450800001EF080417555A2FFC00105D7BE",
INIT_33 => X"140000A2AEBFFEF082A82010F7802AABA5D7FEAB45080015410007FEAA005551",
INIT_34 => X"5140145007BE8B55087BEAB555D04001EFF7AAA8B555D557FE00A280020BAAAD",
INIT_35 => X"7AABDEAAF784154BA08557FEAAA284000AAFF803DE00FFD557400AAD56AB455D",
INIT_36 => X"F780020105D7BEAB45557BE8B45082EBFEBA082EBFFEF007BE8BFF5D2ABDF55F",
INIT_37 => X"0000000000A2FFD54105D7FC21EFFFD16AA10FF80174AA557FC21EF082A80145",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000000FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(1),               -- Port A write enable input
DIA(0)   => data_write_a(14),        -- Port A data input
DOA(0)   => data_read_a_hi_512(14),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(1),               -- Port B write enable input
DIB(0)   => data_write_b(14),        -- Port B data input
DOB(0)   => data_read_b_hi_512(14),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_15_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000A000000000284000280000001800020030000000033022000000180002",
INIT_01 => X"A140098018300848180060000C00424040000000080000080200000000110200",
INIT_02 => X"102100400C8011100000061000A8503401044880010430004808000180122378",
INIT_03 => X"000200541D102210064200000045000546080000400020000008108448400042",
INIT_04 => X"8094020000254C880000028A1018000844000000880013504000002600000000",
INIT_05 => X"10002424000AA81024A82040010C61062001440002988000000024808001004B",
INIT_06 => X"80004400022A00003C8912248E0400042854400040006810000C4901032B1800",
INIT_07 => X"50200000B0280048A0280A828801002101020040000005F38204082640000000",
INIT_08 => X"01F00402802610411100110000000010010802000400230A0008884008080004",
INIT_09 => X"01000001A12481041000000000000080C0030108100004590111820404000000",
INIT_0A => X"0000000080101000004140001001088A45000082000000008000001080008000",
INIT_0B => X"0004404000000000400004000040000400000000000000000004000020000200",
INIT_0C => X"0804000020024100012808020000000981004004A0200310000C000800000000",
INIT_0D => X"0000001180009000000000002100018000000000004004010010000000000000",
INIT_0E => X"00000008000002000000000000000000000080A40000000000000080A4000000",
INIT_0F => X"00000000001000204800000000000000000080A40000000000000080A4000000",
INIT_10 => X"000000000000000000080000020000000000000000000008000C020000000000",
INIT_11 => X"000000824000000000000020220000000001800100020300000004003420480A",
INIT_12 => X"0000000000040440000000000001048000000000000000100800400000000000",
INIT_13 => X"000800000000000000000000000100C220050000000000000000008220884400",
INIT_14 => X"000000000000000830000000000000000016101C5C1400000000000000000000",
INIT_15 => X"0000000000000000000000000020C00000088000012090101280401000000200",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000040028000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"000010082A954BA00003DFEF085155400F78428BEF0000000000000000000000",
INIT_22 => X"8015400FF84001EFA2FBE8B55A2AE80000F7D5555555D2AAAABAAAD1420BAFF8",
INIT_23 => X"87FFFF55557BD54AAF7FBC01FFA2802ABEFF7AE95555A2FBE8BEFA2843DE00AA",
INIT_24 => X"0804155EFFFFBE8BFF0800174AA557BFDE10A2FBEAB45F7D56AABAAAD5554BA0",
INIT_25 => X"5FFD568BEF087FE8A1055003FE00A2AA801FFA28402000AAAE955455500155EF",
INIT_26 => X"45AA843FE0008557DFFF0800020105D557FEAA00557DE10F7D1574AAA2D16AB5",
INIT_27 => X"0BAF7AEA8B45080417400FFFFC2145080015400AA802AA00AAAE800BA5D00155",
INIT_28 => X"000000000000000000000000000000000000000000516AA00A2AE800BAFFFFC2",
INIT_29 => X"A8ABAAADB40092E38E070280024904AA1C0438FD7005150438F78A2DBFF00000",
INIT_2A => X"FE8BC7BE8E38E10A28017400E38A051FFA2FFEDB55B6A080038E3DB50555412A",
INIT_2B => X"D16AABAA2DB50482147FFAF554971D0492E3F1C71C7BE8A2ABD7E3AA9257DA2F",
INIT_2C => X"AAA955554900105FF0800175D7E3FFEFBD70000124AA557FFDE10A2FBEDB6DF7",
INIT_2D => X"FFDF50482A2DB6AB45FFD56DBD7087BEAA38410038E38A2AE851FFB68402038A",
INIT_2E => X"0AAA085082550A1057DBE803AE38145B78FD7000005010495B7AE921C517DE10",
INIT_2F => X"00A2A0800BAE3F1C0092EBAAADB6D080A12410FFF1C017D140410400BE8E28A1",
INIT_30 => X"0AAF7AEBDFEF0000000000000000000000000000000000000000000001C556FA",
INIT_31 => X"00AAAAFBC0145002AA8AAAAAFFC2000AAAA974AA0800020BA550028B55085540",
INIT_32 => X"A8B55AAAE821EFAAFBEAB55F7AAA8A00AA8417400AAAE975EFA2FBFFF55FF840",
INIT_33 => X"BFFE10A2FFFFFEFF7D568ABAA2FFC00105D7BE8B55085142010AAD157545F7AE",
INIT_34 => X"AA955FFFF80020BAAAAA975450800001EF080417555AAFFFDF450804020AA557",
INIT_35 => X"07FEAA0055517DE00FFFBC2000AAFBE8B55F7D17DF45007FE8AAA08002AAAAA2",
INIT_36 => X"5D0000010F7AAA8A10AA8017400552A801EFF7802AABA5D7FEAB450800154100",
INIT_37 => X"00000000005D557FE00A280020BAAAD140000A2AEBFFEF082A82010FFD5421EF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000C00000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(1),               -- Port A write enable input
DIA(0)   => data_write_a(15),        -- Port A data input
DOA(0)   => data_read_a_hi_512(15),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(1),               -- Port B write enable input
DIB(0)   => data_write_b(15),        -- Port B data input
DOB(0)   => data_read_b_hi_512(15),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_16_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"DA22C618B1000482B688B186588884862A400438255FC38381441205BA803003",
INIT_01 => X"264AC80028404C211203A952A90341080B173340412000E1005D628000820484",
INIT_02 => X"400034C206C405000001A48202084004003008255040826EE008B440200E2042",
INIT_03 => X"A459C1240181AB20AD27315B7F1983CA1C900040422A005762010010000C0400",
INIT_04 => X"296E542B6E3A825C15FB385321B4ADFE16AB45FD2C400002E205231201290A28",
INIT_05 => X"B9E5815006028179808C00A0D2152B90707A1E0BD423CAC0000D610000000710",
INIT_06 => X"81F104A1415C292164280081C6AB88742086ACACDE240000A80090CE82A803B9",
INIT_07 => X"400800000ACCAA280940580400A37B8896CA4D000A80C1102A00001C14028009",
INIT_08 => X"0015452880C8D90409A02D965965200100104F2B00822512000000231520A024",
INIT_09 => X"A5AA80018120E00066000000000012C9000A0000D0A80000BF8028E87C1B9927",
INIT_0A => X"00520228080108039501200848002912300208092B940192D1000000000000A8",
INIT_0B => X"03561180063DB4F6110001100011000110001100011000110001080008800080",
INIT_0C => X"080200854409418B02ED0000502A02972000040BB401100010012B4C90000100",
INIT_0D => X"6D061A1F8D60D80820500101244AA8A2AA242E80000009200120000000000000",
INIT_0E => X"6D066210E5001DB4A5B400C7D553847165A99000C6564CDD051DC99000C65555",
INIT_0F => X"21D0C48F254946148107354292673D1F72C99000C6564CDD0565C99000C65555",
INIT_10 => X"952D2058F33225787810F5001D6121A9559224D1FF97D0272F04D89441A56D8A",
INIT_11 => X"6C1C74485B81E31306C71D1093AB8A64811BADC00992180D58033B1172F2A025",
INIT_12 => X"7B86DED8E3A212748F0E0CA638E890B7A8546120C0AFF5B548AC431FB1C7DB07",
INIT_13 => X"EFCE9B26DECA1AD36A2E4F40DF6AAAF260AF88899E8B8B93D12A877178DD0032",
INIT_14 => X"A8009F8B108C80A1021B9A8BB8056662CA1951596800FC01A38D4D4B072B922F",
INIT_15 => X"00000000000000000000000000044000102A0001148442A1108103595580A840",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"4C690DA64C1C4F68A36040000000000000000000000000000000000000000000",
INIT_19 => X"D14D14D14D14D14D14D14D14D14514514514514529E5F87869E79E78558D1154",
INIT_1A => X"3D1E8F47A7D3E9F4FA7D3E9F4FA7D3E9F47A7D1E9F47A7D1E9F4D14D14D14D14",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE000000000000000007D3E9F4FA7D3E8F47A3D1E8F47A",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFEFF7D168B55AAD17FFFF552EBFE00007FC00AA0000000000000000000000",
INIT_22 => X"04000BA552A821FFFF8000010082A954BA00003DFEF085155400F78428BEF087",
INIT_23 => X"2AE80000F7D5555555D2AAAABAAAD1420BA5D2E975EFF7D568BFFFF80175EF00",
INIT_24 => X"FF84001EF0000020AA5D00154005D043FF45555540000082EAABFFA2FBE8B55A",
INIT_25 => X"0087FD74BAAAAEBFFEF557FC00AAF7AE95555A2FBE8BEFA2843DE00AA8015400",
INIT_26 => X"FFAAD5554BA087FFFF55557BD54AAF7FBC01FFA2802ABEF557BEABEF5D041541",
INIT_27 => X"E10A2FBEAB45F7D56AABA082A97545F7D16ABFFFFAABFEAAFF84001FF002A821",
INIT_28 => X"0000000000000000000000000000000000000000FFFBE8BFF0800174AA557BFD",
INIT_29 => X"50438F78A2DBFF0871F8FC7E3D56AB6DBEDB7FFEF552AB8E38087FC209200000",
INIT_2A => X"16ABFFE38E175EF1400000BA412E871FFE38E070280024904AA1C0438FD70051",
INIT_2B => X"2EAFBD7A2FFEDB55B6A080038E3DB50555412AA8ABAAADB400924920925EFF7D",
INIT_2C => X"E8E38E10A28017400E38A051FF0804050BA410A1240055003FF6D5551420101C",
INIT_2D => X"4975EDBC7550E12410087FD74AAB6AABFFC7557FC00BAE3AA9257DA2FFE8BC7B",
INIT_2E => X"AF780051C70824851D7A2DB50482147FFAF554971D0492E3F1C71C7BE8A2ABD7",
INIT_2F => X"D70000124AA557FFDE10A2FBEDB6DF7D16AABA08249756DF7D168BC7F7AABAEA",
INIT_30 => X"AAA007BC0000000000000000000000000000000000000000000000000E3FFEFB",
INIT_31 => X"20BA550028B550855400AAF7AEBDFEF08516AB55A2D16ABEFFFFBFDFFF552AAA",
INIT_32 => X"C20000000021EFF7D568BFFA2AA955FF5D04020AA002A955EFAAAA974AA08000",
INIT_33 => X"03DFEF5D51420005D2ABFF45A2FBFFF55FF84000AAAAFBC0145002AA8AAAAAFF",
INIT_34 => X"AE821EFAAFBEAB55F7AAA8A00AA8417400AAAE975EF0800174BA002E820105D0",
INIT_35 => X"AD157545F7AEA8B5500557DF45552A82000007BD74AAF7AEBDF455D7BC20BAAA",
INIT_36 => X"F7D568B55FFAAAAABAFF8415545000015555A2FFC00105D7BE8B55085142010A",
INIT_37 => X"0000000000AAFFFDF450804020AA557BFFE10A2FFFFFEFF7D568ABA0804155FF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000400000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(2),               -- Port A write enable input
DIA(0)   => data_write_a(16),        -- Port A data input
DOA(0)   => data_read_a_hi_512(16),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(2),               -- Port B write enable input
DIB(0)   => data_write_b(16),        -- Port B data input
DOB(0)   => data_read_b_hi_512(16),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_17_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"5284CE4FB7BD2C8994A13392DBD02E14006B82AC7E800D44D3DD2FD5F9B961C0",
INIT_01 => X"F9BA301F7E03FC6793F2199B39FC233C11D93AE6F3BB92B32091DBC339B24542",
INIT_02 => X"1D5FC0C08F040404446965C0607FB8A217C400C33A908078551BD04222186338",
INIT_03 => X"8504930A37F65820CB24111B7F08014A0AB84A52B6D2AFF97C1B5AC757F06D6B",
INIT_04 => X"250834336D1E81500FDB38302292ADFE103B6DBD204037F202042075E2B1D00A",
INIT_05 => X"8F039786062C6CE092F5FE005236781C402A0807B4070670083DC68206D7E6D0",
INIT_06 => X"0CD26803C3582408962C58B183F8AEF42045919B30E085DD2ED57D4EED08CA6A",
INIT_07 => X"700000B30380670B8142500448E3E01E94EF1340A28AC1AC8156044D1400AA00",
INIT_08 => X"009F3A1B0120A1C51DFFC40C30E5F0182D0950190C0810BE00E9A76E4C6FFBE4",
INIT_09 => X"8FCCC200A59BDD2FFE3F3EC7C7DEF207000F00059D2ED56D7EED2ED3C9A867DC",
INIT_0A => X"0617112E46F05D02DD814102F800633F1D0A7CC9AE7A08BFF0001D35682AC0CE",
INIT_0B => X"8A3F06ABD73DBCF4FBCF4FBCF4FBCF4FBCF4FBCF4FBCF4FBCF4FBE7A7DE7A780",
INIT_0C => X"001000974F08518F5AFFC94B533FADA7FDE97D6BFF329E1B50FF99F086000D9E",
INIT_0D => X"F50B018F95EA3DED1652EC0B27E67F419E2E1E8000C0036340B8000000000000",
INIT_0E => X"F50B01C8DF7F96197DB4AFC8C8886AF672A1537F759299F50B03C1537F759199",
INIT_0F => X"6068331C5103E7EF0FBEED6BB6A9412007C1537F759299F50B03C1537F759199",
INIT_10 => X"21F2CD7F252CDABB3CE8CF7F963AB9FD6AD434201AA68B837FFD1F7B7125B68C",
INIT_11 => X"BD055EB6D555CB2949C15BA7270FF256526BBFD55BBE71D79F73C7AC6DB9BF37",
INIT_12 => X"94080BF82B74E4E1FE4ACA4E0ABD6DAAAB965293036FF6B652A99A6026027FBE",
INIT_13 => X"EF5CBA7A43482800FEFAFD06B8CFCCAB7550D0C2022EAEBD438697AD2EBA9168",
INIT_14 => X"AC00A8BBFC8B501CF7A0FED9A548FA19752C4A4EADAE42FCBC38C3B7BEBF42CF",
INIT_15 => X"0000000000000000000000000026E100002F382DBD9ECFE117805F20CFDAAB00",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"09EDCC4052E917114F981800C000000000000000000000000000000000000000",
INIT_19 => X"EBA69AEBA69A69AEBA69AEBA69A69A69A69A69A68698686981D75D7443720030",
INIT_1A => X"46A351A8D068341A0D068341A0D068341A0D46A341A0D46A341A69AEBA69A69A",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000000000046A351A8D46A351A8D46A351A8D",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFEFF7FBEAB450804001EFAAD57FEAA0000000000000000000000",
INIT_22 => X"51401EF087FD74AA087FFFFEFF7D168B55AAD17FFFF552EBFE00007FC00AA087",
INIT_23 => X"82A954BA00003DFEF085155400F78428BEFAAD168A000004020AA5D7BE8B4500",
INIT_24 => X"552A821FF5D00020BA552A82000552A821555D7FEAB55FF80175EFFF80000100",
INIT_25 => X"FAAFBC01EF5D0015555557BFDEBA5D2E975EFF7D568BFFFF80175EF0004000BA",
INIT_26 => X"BAA2FBE8B55A2AE80000F7D5555555D2AAAABAAAD1420BAFFFFFDF45AAD17FFF",
INIT_27 => X"F45555540000082EAABFF00516AA10552E820BA007FEABEF005555555A2D1554",
INIT_28 => X"00000000000000000000000000000000000000000000020AA5D00154005D043F",
INIT_29 => X"B8E38087FC2092147FFFFFFFFFBFDFC7EBF5E8B550000071EFB6DF7AE9200000",
INIT_2A => X"A07082497FEFB6D1451471EF007BD04920871F8FC7E3D56AB6DBEDB7FFEF552A",
INIT_2B => X"8E175FFE38E070280024904AA1C0438FD7005150438F78A2DBFFBED16AA381C0",
INIT_2C => X"38E175EF1400000BA412E871FF550A00092492A850105D2A80155417BEFB6DEB",
INIT_2D => X"FFF5FFF6DAADF7FFD7B6F1C71EF55001756D5D7BFAEBA4920925EFF7D16ABFFE",
INIT_2E => X"700515556DA2DF50492A2FFEDB55B6A080038E3DB50555412AA8ABAAADB40092",
INIT_2F => X"BA410A1240055003FF6D5551420101C2EAFBD7145B6AA28492487082007FEDBD",
INIT_30 => X"5EFFFFBEAA000000000000000000000000000000000000000000000000804050",
INIT_31 => X"ABEFFFFBFDFFF552AAAAAA007BC0000557FFDFEFF7FBFFF55A2D16AB55000017",
INIT_32 => X"BDFEFF7D568AAA5D2A97410007BFFFFF5551555EF087FC200008516AB55A2D16",
INIT_33 => X"A82155087FFFFEFAAAA975EFAAAA974AA0800020BA550028B550855400AAF7AE",
INIT_34 => X"00021EFF7D568BFFA2AA955FF5D04020AA002A955EF5D2E80010002A954005D2",
INIT_35 => X"02AA8AAAAAFFC2000FFD57DFFFAAFFFDF55FFD1575FF5504175EF5D7FEAAAA00",
INIT_36 => X"000415410007BFFF450051555EFA2FBC0000A2FBFFF55FF84000AAAAFBC01450",
INIT_37 => X"00000000000800174BA002E820105D003DFEF5D51420005D2ABFF45557FE8AAA",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000CFFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(2),               -- Port A write enable input
DIA(0)   => data_write_a(17),        -- Port A data input
DOA(0)   => data_read_a_hi_512(17),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(2),               -- Port B write enable input
DIB(0)   => data_write_b(17),        -- Port B data input
DOB(0)   => data_read_b_hi_512(17),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_18_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"69844019080000A21A611406840014122A641074155FC28A2024001001801003",
INIT_01 => X"01067920034004180005E9E3C90360C0041C0181002001602025800008440084",
INIT_02 => X"40AC3CAA22D605200000856E2481902400344A20F802C22054001000021E2379",
INIT_03 => X"A54C23B34C81EB2076471000800981140C010101750D1007E58040102B0E0100",
INIT_04 => X"22660C1C0065003C04040013236E105016A028402D618803EB092B9201490B2A",
INIT_05 => X"B8E080000000005889AC41E04508A99070200E010001C1CA11803850C8000100",
INIT_06 => X"800A4CE301545001F40050216C09950004C2047BCF1C8090C02800C0120886B3",
INIT_07 => X"814A0080064C1F300020080182001A9E02C03400082002700000217294007101",
INIT_08 => X"000117088080990419002D86184A01018030430700802541420440022030041A",
INIT_09 => X"7030C30B885200D274004008080003C32A10A19090C02010E102294406168800",
INIT_0A => X"00602A01880980037109700C04C44C92A88DCC2211E44174112840880000060D",
INIT_0B => X"11C0D95C20C2030A003080030800308003080030800308003080018400184004",
INIT_0C => X"8304E02809832E6021002020404042000F00008400811824AD4007ECD9436261",
INIT_0D => X"0AFCE5D22A82B20000520100C801F8A07E103000A1285C84000418360C1B060D",
INIT_0E => X"0AFCFD8CB17E5B4F045557575E6EFBE3942C1040A41D660AFCE1CC1040A41E66",
INIT_0F => X"8E7FFBB385661C08D1455ABA91E6FF5FDFCC1040A41D660AFCF9CC1040A41E66",
INIT_10 => X"015F82C006C3AF31E64CB17E5A9655017F1FC73FAF1D61B1040294C58AD1FF5F",
INIT_11 => X"B95454005BAA36DCF8E519001BF80DEB3EE2020EA678189C6EC32881F7F75648",
INIT_12 => X"67D7EDFCA320037E81BD77D728A800B7546DBDFF12904747A351145FC53ABF8D",
INIT_13 => X"92B764225C57C97EBE76E1254F0C0D4514A84F5573FE9DBA4A38E247C522CC0E",
INIT_14 => X"BE84370001B6922070440556B15F7FABBC40151D7C747D8220673C3B9DB84B20",
INIT_15 => X"06C1B06C1B06C1B06C1B06C1B0491069068000004060300A005A01183F240014",
INIT_16 => X"6C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B",
INIT_17 => X"C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B0",
INIT_18 => X"B80EE173C2300F7DF16000000000000000000000000041B06C1B06C1B06C1B06",
INIT_19 => X"AAAAAA28A28A28AAAAAAA28A28A28A28A28A28A2910591505C104104B28BBECE",
INIT_1A => X"128944A25128944A25128944A25128944A2552A954AA5128944AAAA28A28A28A",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000128944A25128944A25128944A25",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFDFEF5D2A974BA082E954000000000000000000000000",
INIT_22 => X"0028B55002E82000087FFFFFFFFFFFFFEFF7FBEAB450804001EFAAD57FEAA087",
INIT_23 => X"7D168B55AAD17FFFF552EBFE00007FC00AA087FFFFFFFFFBFDF45AAD568B5508",
INIT_24 => X"087FD74AAAAFFFDF45A2D16AB55F7FFFFFFF00043DE10AA843DE00087FFFFEFF",
INIT_25 => X"A55042ABEF5D7FD75FFAAD540145AAD168A000004020AA5D7BE8B450051401EF",
INIT_26 => X"45FF8000010082A954BA00003DFEF085155400F78428BEFAA80000000804154B",
INIT_27 => X"1555D7FEAB55FF80175EF5D00020105D2A97400082E95555085168A10557FD75",
INIT_28 => X"00000000000000000000000000000000000000005D00020BA552A82000552A82",
INIT_29 => X"071EFB6DF7AE921C7FFFFFFFFFFFFFFFF7FBFDFFF5D2A954AA082A9242800000",
INIT_2A => X"1FAF55A2DF6DB7D1C002AB7D002A82028147FFFFFFFFFBFDFC7EBF5E8B550000",
INIT_2B => X"8E38E280871F8FC7E3D56AB6DBEDB7FFEF552AB8E38087FC2092087FFDFC7E3F",
INIT_2C => X"97FEFB6D1451471EF007BD0492B6F1F8F55AADF6DB7DE3F5FAFC708003DE28B6",
INIT_2D => X"A28407038140410492550A2ABC7497BD25FFAADF4516DBED16AA381C0A070824",
INIT_2E => X"D1C516FA28417BD5545E38E070280024904AA1C0438FD7005150438F78A2DBFF",
INIT_2F => X"92492A850105D2A80155417BEFB6DEB8E175FF5D0E05000492097428002E9557",
INIT_30 => X"4AA082A820AA000000000000000000000000000000000000000000000550A000",
INIT_31 => X"FF55A2D16AB550000175EFFFFBEAA00557FFFFFFFFFFFDFEFF7FBFFFEF552E97",
INIT_32 => X"C0000087BFDF45AAD568B55AAFBFDFEF55042ABEF002A800AA557FFDFEFF7FBF",
INIT_33 => X"16AB4500043DEAAFFAEAAAAA08516AB55A2D16ABEFFFFBFDFFF552AAAAAA007B",
INIT_34 => X"D568AAA5D2A97410007BFFFFF5551555EF087FC2000FFD56AB45A2FFFDFFFAAD",
INIT_35 => X"855400AAF7AEBDFEFA280154BA550400000552AA8B45087FC01EFA2FFD55EFF7",
INIT_36 => X"0804154BA082A975EF5D517DEAA007BD5545AAAA974AA0800020BA550028B550",
INIT_37 => X"00000000005D2E80010002A954005D2A82155087FFFFEFAAAA975EF5D2E97400",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000400000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(2),               -- Port A write enable input
DIA(0)   => data_write_a(18),        -- Port A data input
DOA(0)   => data_read_a_hi_512(18),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(2),               -- Port B write enable input
DIB(0)   => data_write_b(18),        -- Port B data input
DOB(0)   => data_read_b_hi_512(18),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_19_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"042200000000000041088001001AA00000000000000000000000500802000003",
INIT_01 => X"074018000024000000000404000000000A22000800000800004A200000000001",
INIT_02 => X"0000048002C405000000000006A84000000000200893C246A20000000020031A",
INIT_03 => X"082A58E411004B2000071000000981000C000000002045000200000000000000",
INIT_04 => X"200604000000001C0400001320000000162000002C4000026201201200090800",
INIT_05 => X"1020800000000058840200204000099070200E010001C0400000000000000000",
INIT_06 => X"0012048037805421402850001402498820022802400480405008901100A00102",
INIT_07 => X"00000000020C0130481204919200010C82000000000006002A548902A0020109",
INIT_08 => X"0001150800009900000005861840000000004301000B000000000001C1C00000",
INIT_09 => X"001F00002024B20002000000000002C300000000405000103010204000000000",
INIT_0A => X"00000000000000000000000000000040002000044000000000000000000002F0",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000420003B00000000000000000040012C80000000",
INIT_0D => X"45001A03C0825A0D20800000000018A006001000000000000000000000000000",
INIT_0E => X"450002131E01A1F6EA0A0020211146E069C2ACC01AE80045001D82ACC01AE800",
INIT_0F => X"1188340C3E1CFAD27CC2E004481020892282ACC01AE80045000582ACC01AE800",
INIT_10 => X"DEA03228D810007019931E01A1E5BA02802008C06F029D4C7B76639CEC0A0020",
INIT_11 => X"428AA3592000000206C2A4DAC00000008113C246A181C03FE4662A84575768DF",
INIT_12 => X"08201090549B5800000000261546B24000000000C53807E7CC06618018C51210",
INIT_13 => X"13F6A185A0A0168128411ACB800C0E108A0720288C011046B5986247C5452291",
INIT_14 => X"0000C220010808C10D9A92A74CD7CF4A080031B1515B212143D841431046B58A",
INIT_15 => X"00000000000000000000000000000000000000000000000000000118030004E0",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"3F0C7010C660C744192000000000000000000000000000000000000000000000",
INIT_19 => X"1861861861869A61861861861861861861861861A8208C4C1534D34C07208BBA",
INIT_1A => X"0984C26130984C26130984C26130984D26930984C26130984C261861861869A6",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE000000000000000000984C26130984C26130984C2613",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF552A974AA0004174BA0000000000000000000000",
INIT_22 => X"2E974BAA2FFFFE10087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974BA082E95400F7F",
INIT_23 => X"FFFFFFEFF7FBEAB450804001EFAAD57FEAAF7FFFFFFFFFFFFFFFFF7FBFDFFF55",
INIT_24 => X"002E82000F7FFFFFFFFFFFFDFEFA2D568B550004001EFAAAEA8ABA087FFFFFFF",
INIT_25 => X"5AAD16ABEF5D2ABFF55080402010087FFFFFFFFFBFDF45AAD568B55080028B55",
INIT_26 => X"BA087FFFFEFF7D168B55AAD17FFFF552EBFE00007FC00AAF7FFFFFFFF7FBE8B5",
INIT_27 => X"FFF00043DE10AA843DE00557FFDFEFA2D16AB55A2FFFDFEF5D2EBFE00AAFFFFE",
INIT_28 => X"0000000000000000000000000000000000000000AAFFFDF45A2D16AB55F7FFFF",
INIT_29 => X"954AA082A92428E3FFFFFFFFFFFFFFFFFFFFFFFEF552A974AA0000104AA00000",
INIT_2A => X"FFDFEFF7F5FAFC7492A974AAB6F5F8E101C7FFFFFFFFFFFFFFFF7FBFDFFF5D2A",
INIT_2B => X"A4A8AAA147FFFFFFFFFBFDFC7EBF5E8B550000071EFB6DF7AE92EBFFFFFFFFFF",
INIT_2C => X"2DF6DB7D1C002AB7D002A82028FFFFFFFEFF7F1F8FD7AAD16AB450000001FFBE",
INIT_2D => X"F7FBF8FC7E3F5EAB45B6DF6FBEF5D2AB8F7D000000010087FFDFC7E3F1FAF55A",
INIT_2E => X"7412ABFE28B6F5F8E820871F8FC7E3D56AB6DBEDB7FFEF552AB8E38087FC2092",
INIT_2F => X"55AADF6DB7DE3F5FAFC708003DE28B68E38E284971F8FC7AAD56DB6DBEF5F8FD",
INIT_30 => X"4AA0004000AA000000000000000000000000000000000000000000000B6F1F8F",
INIT_31 => X"DFEFF7FBFFFEF552E974AA082A820AAA2FFFFFFFFFFFFFFFFFFFFFDFEF552E95",
INIT_32 => X"EAA00A2FFFFFFFF7FBFDFFFFFD568B55002A954AAF7D568A00557FFFFFFFFFFF",
INIT_33 => X"56AB450004001EFFF842AAAA557FFDFEFF7FBFFF55A2D16AB550000175EFFFFB",
INIT_34 => X"7BFDF45AAD568B55AAFBFDFEF55042ABEF002A800AAF7FBFDFEFF7D56AB45AAD",
INIT_35 => X"52AAAAAA007BC0000FFFBE8B55AAD168B55F7FFFFFFF552AA8BEF08040200008",
INIT_36 => X"A2D57FFFFF7D568B45002ABDEAAFFD16AA0008516AB55A2D16ABEFFFFBFDFFF5",
INIT_37 => X"0000000000FFD56AB45A2FFFDFFFAAD16AB4500043DEAAFFAEAAAAA08556AB55",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000800000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(2),               -- Port A write enable input
DIA(0)   => data_write_a(19),        -- Port A data input
DOA(0)   => data_read_a_hi_512(19),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(2),               -- Port B write enable input
DIB(0)   => data_write_b(19),        -- Port B data input
DOB(0)   => data_read_b_hi_512(19),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_20_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000003",
INIT_01 => X"A65FF80000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000048002CC070000000000000000000000002FF86100200000000220002362",
INIT_03 => X"0000000000080F6000977060009B87A03C000000000000000000000000000000",
INIT_04 => X"3F2EFC040388137C3E20C477600142019E6000003CC0000A6601601A000B0000",
INIT_05 => X"102F91D10802ABFB80000021C8010FB0F0F43E1FE867DFC04400390210000220",
INIT_06 => X"90492261000080003400000010008000004203FE400580000000803000200006",
INIT_07 => X"401000004FFDFF28C4300C0010200100004000002AA001F00000000014000000",
INIT_08 => X"0801F5780259FB00000007BEFBC010002008FF7F00000000010018A81000041C",
INIT_09 => X"00000000020000000000000000000ADF00000020000000800000802830011023",
INIT_0A => X"0000000000000200020000000000000000000000000000000200200290000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"08120000B9090A700000200000004000000400000080002000407FED80000000",
INIT_0D => X"000079804000F00000000000C01FF8A7FE003000000004008100000000000000",
INIT_0E => X"0000798201000000100000000135386000401000010000000079801000010000",
INIT_0F => X"0185C300020004000010000000000252C7801000010000000079801000010000",
INIT_10 => X"00000010C1F30F300002010000080000000000CD8A0000400400000010000000",
INIT_11 => X"008040000000000292C0080000000000A5604000000284000818505200080000",
INIT_12 => X"0015E1B00100000000001496008000000000052B000048080000000000FC3600",
INIT_13 => X"80000000000002BA280000800830300000000000B8B400000401881010000000",
INIT_14 => X"00000000020020020001000040283024E6FB8604020080000383383B00000400",
INIT_15 => X"000000000000000000000004010201001003020200000000000127DBFF004000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"038200010089120104D204002000000000000000000000000000000000000000",
INIT_19 => X"B2CB2CB2CB2CB2CB2CB2CB2CB2C30C30C30C30C306982121A1E79E79A0700030",
INIT_1A => X"432190C86432190C86432190C86432190C86432190C86432190CB2CB2CB2CB2C",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000432190C86432190C86432190C86",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA0804020100000000000000000000000",
INIT_22 => X"2E954AA000400000F7FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0004174BAFFF",
INIT_23 => X"FFFFFFFFFFFFFDFEF5D2A974BA082E95400007FFFFFFFFFFFFFFFFFFFFFFEF55",
INIT_24 => X"A2FFFFE10FFFFFFFFFFFFFFFFFFFFFBFDFFF5D2E954BA007FC00BA087FFFFFFF",
INIT_25 => X"FF7FBFFF550800020BAAAD56AAAAF7FFFFFFFFFFFFFFFFF7FBFDFFF552E974BA",
INIT_26 => X"10087FFFFFFFFFFFFFEFF7FBEAB450804001EFAAD57FEAA007FFFFFFFFFFFFFE",
INIT_27 => X"B550004001EFAAAEA8ABA5D7FFFFFFFFFFFDFEFF7D56AB450000021EFA2D57DE",
INIT_28 => X"0000000000000000000000000000000000000000F7FFFFFFFFFFFFDFEFA2D568",
INIT_29 => X"974AA0000104AAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA08000500000000",
INIT_2A => X"FFFFFFFFFBFDFEF5D2E974AA000A07000E3FFFFFFFFFFFFFFFFFFFFFFFEF552A",
INIT_2B => X"71C50BA1C7FFFFFFFFFFFFFFFF7FBFDFFF5D2A954AA082A92428087FFFFFFFFF",
INIT_2C => X"7F5FAFC7492A974AAB6F5F8E10E3FFFFFFFFFFFFFFEFF7FBFFFFF552E974AA00",
INIT_2D => X"1C7FFFFFFFFFBFDFEFE3F5F8F450004050AABEDF6FABAEBFFFFFFFFFFFFDFEFF",
INIT_2E => X"50804021FFB6D57DE28147FFFFFFFFFBFDFC7EBF5E8B550000071EFB6DF7AE92",
INIT_2F => X"EFF7F1F8FD7AAD16AB450000001FFBEA4A8AAA497FFFFFFF7FBF8FC7EBD168B4",
INIT_30 => X"4AA080017410000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFDFEF552E954AA0004000AAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A95",
INIT_32 => X"820AA087FFFFFFFFFFFFFEFF7FBFDFFF5D2A974AA002E95410A2FFFFFFFFFFFF",
INIT_33 => X"FFDFEF5D2E954AA0051554BA557FFFFFFFFFFFDFEFF7FBFFFEF552E974AA082A",
INIT_34 => X"FFFFFFFF7FBFDFFFFFD568B55002A954AAF7D568A00AAFFFFFFFFFFBFDFEFFFF",
INIT_35 => X"000175EFFFFBEAA005D7FFFFEFF7FBFDFFFAAD16AB450804174AAFFFFFFEBAA2",
INIT_36 => X"F7FFEAB45A2D568B550804001EFF7D57DEBA557FFDFEFF7FBFFF55A2D16AB550",
INIT_37 => X"0000000000F7FBFDFEFF7D56AB45AAD56AB450004001EFFF842AAAA087BFDFEF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000000FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(2),               -- Port A write enable input
DIA(0)   => data_write_a(20),        -- Port A data input
DOA(0)   => data_read_a_hi_512(20),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(2),               -- Port B write enable input
DIB(0)   => data_write_b(20),        -- Port B data input
DOB(0)   => data_read_b_hi_512(20),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_21_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"4A302428B824900A128C090A5C1800261500213C005FE812D10420054085A202",
INIT_01 => X"081FFE3440B609703B0427F801A40B8115BC4F655300340288A40D30040E4DD8",
INIT_02 => X"04CA478082CC1740002019824E0203100640303FF8C0B31061096E21A1840814",
INIT_03 => X"8C329E9204020FE002577800405B87047D5042129D8D0248903200013290C800",
INIT_04 => X"3E7FFE02482553FC3C020277E128080A1E6000003CC0000A6601E03A8B0F0008",
INIT_05 => X"F43F8140000203FFC806C8A1C1048FF0F0E07E1F00F7FFC00024010000468310",
INIT_06 => X"08710C10015E083D01A24404786BE0014114C3FE4187A009A663A680100B3096",
INIT_07 => X"200800008FDFFF00290000100211019812E210488228000000900260026C6058",
INIT_08 => X"0EF1F5FA0041FF080AC707FEFBC110008420F7FF388B70A20389346FE8000580",
INIT_09 => X"917FC30010107688862A28C54518DBFF00020004C0A6044901112A0908AA0A30",
INIT_0A => X"006309044081A001B188300E20806520398C6021569249C4B3007127080806FF",
INIT_0B => X"904595123203040D9228D9228D9228D9228D9228D9228D9228D99146C9146C84",
INIT_0C => X"88042090068008003120000806001402504110C48002403601887FEF80022A51",
INIT_0D => X"26C0AC404E43032CA0C205880A7FFAB7FE01409400400C0594A4002200110008",
INIT_0E => X"26C0AC086A170250454004C6012280129B034A080C0B0016A0D20346080C0A80",
INIT_0F => X"0B064092D85938C0112144050224120C500346080C0B0016A0D2034A080C0A80",
INIT_10 => X"40702E058355458967E86A170220D1800093414B0414782E4B5000D81480809A",
INIT_11 => X"081B1545104135443306C35901024F88A88049062A747512B76783C5D040E080",
INIT_12 => X"40160040D86B202049B22198362A8A208279854400A036801480031401900800",
INIT_13 => X"0DD001C002D38334000914028354008301008C0CF1480245108C7640A0604032",
INIT_14 => X"AC0496022300233104662848808E191526205018030060540284FA0C0044022C",
INIT_15 => X"004010040100401004010040102090010008000001C0E010020007DFFFC06E60",
INIT_16 => X"0401004010040100401004010040100401004010040100401004010040100401",
INIT_17 => X"4010040100401004010040100401004010040100401004010040100401004010",
INIT_18 => X"FF7FFDF7FF3E3DFDF7E000000000000000000000000040100401004010040100",
INIT_19 => X"FBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBFFDFDFFFCF3CF3FFFEF9FEE",
INIT_1A => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFEFF7FBFDFEFF7FBFDFEFBEFBEFBEFBE",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0004000100000000000000000000000",
INIT_22 => X"2A954BA0004154BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080402010FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF552A974AA0004174BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"000400000007FFFFFFFFFFFFFFFFFFFFFFEF552E974BA0804000AAF7FFFFFFFF",
INIT_25 => X"FFFFFFDFEF5D2E974BA002E97400007FFFFFFFFFFFFFFFFFFFFFFEF552E954AA",
INIT_26 => X"BA087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974BA082E95400007FFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2E954BA007FC00BA5D7FFFFFFFFFFFFFFFFFFBFDFEF5D2A954AA002E974",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFBFD",
INIT_29 => X"954AA080005000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA00000200000000",
INIT_2A => X"FFFFFFFFFFFFFFF552A974BA0000174AAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0A000AAE3FFFFFFFFFFFFFFFFFFFFFFFEF552A974AA0000104AAF7FFFFFFFFFF",
INIT_2C => X"FFBFDFEF5D2E974AA000A07000007FFFFFFFFFFFFFFFFFFFFDFEF552E954BA08",
INIT_2D => X"1C7FFFFFFFFFFFFFFFFFFBFDFEF5D2A974BA002A95400087FFFFFFFFFFFFFFFF",
INIT_2E => X"F552E974BA0020924BA1C7FFFFFFFFFFFFFFFF7FBFDFFF5D2A954AA082A92428",
INIT_2F => X"FFFFFFFFFEFF7FBFFFFF552E974AA0071C50BA557FFFFFFFFFFFFFFFF7FBFDFF",
INIT_30 => X"4BA000002000000000000000000000000000000000000000000000000E3FFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2A954AA080017410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"000AAF7FFFFFFFFFFFFFFFFFFFFFFFEF552A974BA0000174BAFFFFFFFFFFFFFF",
INIT_33 => X"BFDFEF5D2A954BA082E800AAA2FFFFFFFFFFFFFFFFFFFFFDFEF552E954AA0004",
INIT_34 => X"7FFFFFFFFFFFFFEFF7FBFDFFF5D2A974AA002E95410087FFFFFFFFFFFFFFFF7F",
INIT_35 => X"52E974AA082A820AA557FFFFFFFFFFFFFEFF7FBFFFFF552E954BA002E9741008",
INIT_36 => X"FFFBFDFEFF7FFFFFEF5D2A974BA0000020AA557FFFFFFFFFFFDFEFF7FBFFFEF5",
INIT_37 => X"0000000000AAFFFFFFFFFFBFDFEFFFFFFDFEF5D2E954AA0051554BA5D7FFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(2),               -- Port A write enable input
DIA(0)   => data_write_a(21),        -- Port A data input
DOA(0)   => data_read_a_hi_512(21),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(2),               -- Port B write enable input
DIB(0)   => data_write_b(21),        -- Port B data input
DOB(0)   => data_read_b_hi_512(21),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_22_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"5290F4CDE914905A14A43D33F488243E17122300F55FEB189B343A1140548380",
INIT_01 => X"A94007B259F6A975386262000C344BA9573C6FF57B18A5FB0ABFCD3C2C5F4F0C",
INIT_02 => X"D56B4302AC01005111011BD506AA5205274056900596A539584E2E6DFE4B2418",
INIT_03 => X"6B03F2F6151A2081F24001E8400008F401CB10C6594423C8923AD6B55AD0EB5A",
INIT_04 => X"8001023D37E50880436200808BC8492A0089249600101100008087248B64426E",
INIT_05 => X"A51035B41C0A88046CAEE8C23C08E040011C0020F8882001102D620A06D68301",
INIT_06 => X"B93FF975CF7889D085E997A2144E8FC2060B880081A26DCD4047EFF9EF018980",
INIT_07 => X"283800AA500200E8024AD03546A3262FB5AA5542A882040C7A64CBD64065F028",
INIT_08 => X"141008801018040E48D500400015805060040080A2A0F4A82381B4000A0905A0",
INIT_09 => X"4D0000002126F30C902A29C54539C020E11810098D4067EFF9FF284D483E2AB4",
INIT_0A => X"1400006100003202D040050220103D2A512C6A8C4F0008AA800470370000A000",
INIT_0B => X"013456520CA09281C2A81C2A81C2A81C2A81C2A81C2A81C2A81C9540E1540E00",
INIT_0C => X"A1402A13C0A10A893165281A1C2A7283516344C594A85536B1AD800214202C50",
INIT_0D => X"3C70FC20515808A0100820112300011000287B071105034406950A0285014280",
INIT_0E => X"3C70FC48E11CFC48400184CE0D6783139B0959A41606003C70FA0958AC160480",
INIT_0F => X"0D87E8B3B811B52048B10E0402AE1606D80958AC1606003C70FA0959A4160480",
INIT_10 => X"80F84E0185594581E088E11CFC38414020DD42CF909D7E0A551C02180300C0DD",
INIT_11 => X"441154C258012D86F3044A3133004A99BD8455300654458A1D588C4061403000",
INIT_12 => X"A096A240894626600953379822A984B0025B0DEC0345C9200680027181B44887",
INIT_13 => X"E2404160035482BE521C2C04A90783C18000D610B9D8070B12B1A2A62040202A",
INIT_14 => X"304244A91102C93A2D608D2A258DF8034284200C050070E40C80620C870B02C4",
INIT_15 => X"4411044110441104411044110466C440446CA06951D4EA801000980400646002",
INIT_16 => X"0100441104411044110441104411044110441104411044110441104411044110",
INIT_17 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_18 => X"FE8FF1F7DEBDDF7DF7D05122890000000003FFFFFFFF90040100401004010040",
INIT_19 => X"79E79E79E79E79E79E79E79E79E79E79E79E79E7BFFDFD7DDDF7DF7DF7DFBFDE",
INIT_1A => X"3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE79E79E79E79E",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE000000000000000003F9FCFE7F3F9FCFE7F3F9FCFE7F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0800000000000000000000000000000",
INIT_22 => X"2E974AA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000400010FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E954AA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"0004154BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA000015400FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF552A974AA0800154AAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA",
INIT_26 => X"BAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0004174BAFFFFFFFFFFFFFFFFF",
INIT_27 => X"FEF552E974BA0804000AAA2FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0000174",
INIT_28 => X"0000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040001000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E954AA000402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0417410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080005000FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF552A974BA0000174AAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA00",
INIT_2D => X"E3FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0804154BAF7FFFFFFFFFFFFFFFFF",
INIT_2E => X"F552E954BA000E124BAE3FFFFFFFFFFFFFFFFFFFFFFFEF552A974AA0000104AA",
INIT_2F => X"FFFFFFFFFFFFFFFFDFEF552E954BA080A000AAA2FFFFFFFFFFFFFFFFFFFFFFFE",
INIT_30 => X"4BA080400010000000000000000000000000000000000000000000000007FFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"17410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000400010FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF552A954BA000415400FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954AA0800",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFEF552A974BA0000174BAF7FFFFFFFFFFFFFFFFFFF",
INIT_35 => X"52E954AA0004000AAA2FFFFFFFFFFFFFFFFFFFFFDFEF552E974AA0804174AAF7",
INIT_36 => X"FFFFFFFFFFFFBFDFEF5D2E954BA002A820BAA2FFFFFFFFFFFFFFFFFFFFFDFEF5",
INIT_37 => X"0000000000087FFFFFFFFFFFFFFFF7FBFDFEF5D2A954BA082E800AAAAFFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000000FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(2),               -- Port A write enable input
DIA(0)   => data_write_a(22),        -- Port A data input
DOA(0)   => data_read_a_hi_512(22),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(2),               -- Port B write enable input
DIB(0)   => data_write_b(22),        -- Port B data input
DOB(0)   => data_read_b_hi_512(22),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_23_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"EF20906D902424807BC8241BC81801B97D38AD3C0800103362A6741C80A12A02",
INIT_01 => X"001FFF8409F089003B4422000D80C80106804A7951C5B9D1C828043EA28838F9",
INIT_02 => X"028406A002DC176444683862400003111001303FFC00F240D50146013B300500",
INIT_03 => X"001B243004080FE000177003145F87017D584B10D804034800200200A1008008",
INIT_04 => X"BEFFFC0248005FFC3C18A2FFE12222425E600000BDC0800AEE01E81A100F0A00",
INIT_05 => X"D03F8000000003FF810640A1C0008FF2F0E17E1F02FFFFC80100004044800080",
INIT_06 => X"800264B4854650040123428C204BF40F439647FF4807E189A477EF81DF0AF116",
INIT_07 => X"01000000FFDFFFE800401005C0A0008F86C60840AAAA100C68D1810C9F4A0020",
INIT_08 => X"1BE1F5F80003FF0002021FFEFBC80000000077FF184B03010004002FE1F29002",
INIT_09 => X"907FC308181204800600000000001BFFA800808189A657EF81DD0C00079CC800",
INIT_0A => X"0063090442A18001B188300C48907120AC810033149249C433200180082A06FF",
INIT_0B => X"9A41C1443243050C1010C1010C1010C1010C1010C1010C1010C1008608086084",
INIT_0C => X"000082A00600200080000500C000400800601200000254A000007FEFC1030221",
INIT_0D => X"0A9080400E0BF30C20CA858E087FFABFFE01409780214EE49620001000080004",
INIT_0E => X"0A908044294700701641005218521210150E5789F90A000A90800E5F81F90880",
INIT_0F => X"0E0220036864A7DCA190440301E2105C000E5F81F90A000A90800E5789F90880",
INIT_10 => X"C1400500C6CE5400032429470068924010164302048156305D66F8701681000E",
INIT_11 => X"2E0CCB0500013440600339C800004D8018000857A82920CE8CB220C81400A180",
INIT_12 => X"220344406739000009B0030019960A00026880C0422C52B01700044901488822",
INIT_13 => X"85C811A010428104128996465ADA020180804A040108A2658217C4008060300C",
INIT_14 => X"BE0692020328CA0028042054A92771C50FC070109000C1C819078280A265920E",
INIT_15 => X"020080200802008020080200800800200200000000000008004807DFFF000470",
INIT_16 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_17 => X"0080200802008020080200802008020080200802008020080200802008020080",
INIT_18 => X"0000000000000000000000000000000000000000000000802008020080200802",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000",
INIT_22 => X"2E974BA080002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E974BA000400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000400000FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF5D2E954AA080000010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA",
INIT_26 => X"10FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080402010FFFFFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2A954BA000015400FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA0804000",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E974BA080002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF5D2E954AA000402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA00",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080002010FFFFFFFFFFFFFFFFFFF",
INIT_2E => X"F5D2A954BA080407000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080005000",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF5D2A954BA000417410FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA080402000000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"02000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000010FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF5D2E974AA000402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0000",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000400010FFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"D2A954AA080017410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954AA080002000FF",
INIT_36 => X"FFFFFFFFFFFFFFFFFF552A954BA080015410FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_37 => X"0000000000F7FFFFFFFFFFFFFFFFFFFFFFFFF552A954BA000415400F7FFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000000FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(2),               -- Port A write enable input
DIA(0)   => data_write_a(23),        -- Port A data input
DOA(0)   => data_read_a_hi_512(23),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(2),               -- Port B write enable input
DIB(0)   => data_write_b(23),        -- Port B data input
DOB(0)   => data_read_b_hi_512(23),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_24_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100600007FFF000080108004000800020000840041000080808",
INIT_02 => X"0000068002CC07400000090C080002000000103FF811F150231000520ABE4404",
INIT_03 => X"8428180000080FE000177000001B87003D4000000E8B84010020000000008000",
INIT_04 => X"3E2FFC024800137C3C000077E00000001E6000003CC0000A6601E01A000F0200",
INIT_05 => X"103F8000000003FF80000021C0000FF0F0E03E1F0067FFC00000000000000000",
INIT_06 => X"00132412079001AD00810005E8000001401643FE4007E5501AA00000DC8C3006",
INIT_07 => X"000000000FDFFF62695A5685C094831D966000008002100C2040A178B600C240",
INIT_08 => X"08E1F5F80001FF00000007FEFBC00000000077FF000B00000000002FE0000000",
INIT_09 => X"107FC300000000000600000000001BFFA0000005501AA00000CE200000940000",
INIT_0A => X"00630104408180012188300C00814080008000010012414433000100080806FD",
INIT_0B => X"904181003003000C1000C1000C1000C1000C1000C1000C1000C1000608006084",
INIT_0C => X"00000080060000000000000012002C00000000000000000000007FEF80020201",
INIT_0D => X"440082404E0B332CA2C20188087FFAB7FE000082000000008220000000000000",
INIT_0E => X"4400824903210308074084210002460402009280010D80440084009280010F00",
INIT_0F => X"800A2400401A0C82183248060010280C20009280010D80440084009280010F00",
INIT_10 => X"C0A078160000404A0469032102981380202080026420020D06C002A08481C020",
INIT_11 => X"00164F400860000824059AD01802000208104817B00011306B2D9B0DD5082080",
INIT_12 => X"41021800B35A0300400041202C9E8010C0001040C5836CC01780018601030088",
INIT_13 => X"DB1011E000A140058220004AEFFC8101810021084301880030A8B77400603011",
INIT_14 => X"8C063C0220002201490418082010A57263E010000201033016085A40880030A1",
INIT_15 => X"000000000000000000000000000000000000000000000000000007DFFF0006E0",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"F6E7CC1132CDB444199000000000000000000000000000000000000000000000",
INIT_19 => X"79E79E79E79EFBEFBEFBEFBEFBEF9EF9EF9EF9EFA69861219575D75FF2D0AEEA",
INIT_1A => X"0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1EFBEFBEFBE79E",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE000000000000000000783C1E0F0783C1E0F0783C1E0F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020100000000000000000000000",
INIT_22 => X"2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"080002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_26 => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000400010FFFFFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2E974AA000400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0004000",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040201000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF5D2E974BA080002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFF",
INIT_2E => X"F5D2E974AA000400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF5D2E974AA000400000FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA080402010000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"00010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000010FFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002010FF",
INIT_36 => X"FFFFFFFFFFFFFFFFFF5D2E974AA000002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_37 => X"0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000402010FFFFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(3),               -- Port A write enable input
DIA(0)   => data_write_a(24),        -- Port A data input
DOA(0)   => data_read_a_hi_512(24),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(3),               -- Port B write enable input
DIB(0)   => data_write_b(24),        -- Port B data input
DOB(0)   => data_read_b_hi_512(24),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_25_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100200002000000080100004000000020000800041000080808",
INIT_02 => X"0000068002CC474000000800000002000000103FFCE302008000000880844A04",
INIT_03 => X"00000101C0200FF004177800081B87003D400000080000000020000000008000",
INIT_04 => X"3E2FFE024820137C3C004077F01000001E7249213CC1264A660DF05A000F9000",
INIT_05 => X"103F81C1002203FF80000021C1140FF8F0E03E1F0067FFE04800258280010052",
INIT_06 => X"80480AE20000000100000001C8608001401643FE4007C00000000000CC083006",
INIT_07 => X"280800000FDFFFEA4050140540B00100840000080002A00C2040810000000010",
INIT_08 => X"C8E1F5FA21C9FF80040007FEFBE031018C31F7FFBAEBC0020008086FE0000100",
INIT_09 => X"107FC301800000000600000000001BFFE00301000000000000CC020000140000",
INIT_0A => X"0077330C4889CC292588300C0080400000800001001243443B000100880806FD",
INIT_0B => X"904189003003000C1000C1000C1000C1000C1000C1000C1000C1000608006084",
INIT_0C => X"8B04228026824100000000000000000000000000000004A000007FEF80020201",
INIT_0D => X"400000400E03C30C20C2818C087FFAB7FE01409700C10007962418220C110608",
INIT_0E => X"4000000001010000004000000000400400001200000800400000001200000800",
INIT_0F => X"0008000000000480000040000000200000001200000800400000001200000800",
INIT_10 => X"0000001001000002000001010000100000000000202000000440000000800000",
INIT_11 => X"0000410000000008000008400000000200000806300400000820000020004880",
INIT_12 => X"0000080001080000000040000082000000001000000040800800000000020008",
INIT_13 => X"8100000000000000802000000840000200040000020008000000840000804000",
INIT_14 => X"8C04100200000200000610000000210000000018140000000008000008000000",
INIT_15 => X"04411044110441104411044510629041040D180400000010028047DFFF800C60",
INIT_16 => X"4411044110441104411044110441104411044110441104411044110441104411",
INIT_17 => X"4110441104411044110441104411044110441104411044110441104411044110",
INIT_18 => X"196A8C5A2932EC15DA080800002FFFFFFFFFFFFFFFFFC1104411044110441104",
INIT_19 => X"92492492492410410410410410410492410492412000531215A69A6BFBA2894A",
INIT_1A => X"B158AC562B158AC562B158AC562B1588C46231188C46231188C4924924924924",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000B158AC562B158AC562B158AC562",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000",
INIT_22 => X"2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF5D2E974BA080400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_26 => X"10FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0800000",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400000FFFFFFFFFFFFFFFFFFF",
INIT_2E => X"F5D2E974BA080000010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA080402000000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"02000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400000FF",
INIT_36 => X"FFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_37 => X"0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000000FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(3),               -- Port A write enable input
DIA(0)   => data_write_a(25),        -- Port A data input
DOA(0)   => data_read_a_hi_512(25),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(3),               -- Port B write enable input
DIB(0)   => data_write_b(25),        -- Port B data input
DOB(0)   => data_read_b_hi_512(25),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_26_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"E9264EAB20190CA3BA4997AA9002AE9C001006B0778015CFA17E0811039879C7",
INIT_01 => X"F1FFF9BB1F773C7F9BB07DFFFDD863FC5FFF3FEFFBBF9FFB22FFFBC7B9F30686",
INIT_02 => X"9B3184F8AFDEAF300029E4E300FC78A6258548EFFA71C00172082400003A2161",
INIT_03 => X"0213C3FDFFFC7F74FFBF737A603B87FEBE1A5294F65628A0001B9CE6CC606E73",
INIT_04 => X"7E2EFEBF6FFEB37C3FF3017776FFCDA43E7B6DFD7DEBFD8E6F5F78DF0BFBD644",
INIT_05 => X"902F87C74E8CCFFBB6FF70E1FE61FFBDF0FEBE1FFD67DFFEFFBDA7F7FED50870",
INIT_06 => X"213246200BCC8920360C1831CD7DF60A244B9BFEE00589DDBCEFEDC1DFA08957",
INIT_07 => X"B1D4223B4FFDFF21CC721C85DCE1458E8782484020A2C1FCA3468D77E0000300",
INIT_08 => X"2C05FD7BC471FBD13D980FBEFBEBF30B8D79FF7F451F33CFD60FE8FFFDF54003",
INIT_09 => X"19FFC71FEFED7B251E35768E8ED6BFDF3EB3EBF9DDBCE7FDC1DF8A760F3EACC0",
INIT_0A => X"56F7730ECCDBDF152199F51EDDCDEBCFF589807B7096CD4CF73AC1FC98884FFF",
INIT_0B => X"B867D3683A03A40F78C0D78C0D78C0D78C0D78C0D78C0D78C0D7A606BC606B8C",
INIT_0C => X"DFBFF5EB36DFE51FC3A80D73D840303983EE7F0EA03BDA680137FFFDFFD7E681",
INIT_0D => X"3F0080425E6BFF8DB0DAE19C09FFFFE7FE3EBEA8EB7AFEE5C9AEBD7F5EBFAF5F",
INIT_0E => X"3F00800DEC010280004000F808020290100FA2F60008003F00800FA2F6000800",
INIT_0F => X"00023002007BC0A14E00400003B8000D000FA2F60008003F00800FA2F6000800",
INIT_10 => X"01E0320007204008040DEC010300100000F600020581003F604D0700008000EE",
INIT_11 => X"201F21A2C40039006807C46426040E101A0259DFE82011A311AA042016040080",
INIT_12 => X"80020048F88C84C101C203403E434588007200D047F00090200007E0010009B0",
INIT_13 => X"0109000003E2000416C0804FE04140E80000F808010AB02033AC048A2A00003D",
INIT_14 => X"FFAFD082003B032FB987E04021D481D4000419060201E1A000044300B02033E8",
INIT_15 => X"AFEBFAFEBFAFEBFAFEBFAFEFFBFBFBFBBFCFBB0FFDFEFFEF2DFFFFFBFF802FFD",
INIT_16 => X"FEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBF",
INIT_17 => X"EBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFA",
INIT_18 => X"F491E166CC8553F86EDB5C88646FFFFFFFFFFFFFFFFFEBFAFEBFAFEBFAFEBFAF",
INIT_19 => X"1861861861861861861861861861869A69A61861AFBD54D5F871C71D475B15BC",
INIT_1A => X"0984C26130984C26130984C26130984C26130984C26130984C26186186186186",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE000000000000000000984C26130984C26130984C2613",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000",
INIT_22 => X"2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_26 => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFF",
INIT_2E => X"F5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA080402000000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"02010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_36 => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_37 => X"0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(3),               -- Port A write enable input
DIA(0)   => data_write_a(26),        -- Port A data input
DOA(0)   => data_read_a_hi_512(26),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(3),               -- Port B write enable input
DIB(0)   => data_write_b(26),        -- Port B data input
DOB(0)   => data_read_b_hi_512(26),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_27_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"00080A40000A41248002029000050A088000008242A0004404480002000A1155",
INIT_01 => X"F1FFF1C11F781C129C107DFFFE0860941E81258CA2B71C2220EC1B86E1A00002",
INIT_02 => X"183080988B2EAE00002BE001117C78C6848140CFFA0000800042008000011081",
INIT_03 => X"000003FDF3E47C74F7BCF36A203A47F6B8184210B6160820001318C60C204C63",
INIT_04 => X"7E28FEBF6FEEB3723F71017476DFC524397B6DF572EB6C8E175E70D90F539600",
INIT_05 => X"000F86064C8DDFE3B6FF50D1FC61DE39C8FCB91FF9671FE6B68984B5BCE40834",
INIT_06 => X"0000000800000042020C18300520620A80231BFE200181092CE7ED80DFC00147",
INIT_07 => X"8AC4AA3B0FD1FF201044110560884000840200520002080C23468D0300000282",
INIT_08 => X"2005F0784411E390A4880E3DF7E2FB0B8E717C7F411F3BC6D60B60FFDDE44001",
INIT_09 => X"18FFD757E7ED7A211E81C09818109E1F16B16B71092CE7ED81CF403601228C40",
INIT_0A => X"46FF730E5CCBCD55219AB55F0DEFABC7054880693016DD4C755AC16C1A884FFE",
INIT_0B => X"BC63F1683803C00E3440C3440C3440C3440C3440C3440C3440C3C2061A2061AD",
INIT_0C => X"56BF55CB165EC51D41880FA3F040202883B475062033186801137FF1BAD6F281",
INIT_0D => X"3B0000421E2B0F2E2AE215C808FFFA47FE62BAA86B1AB268E92AB56D5AB6AD5B",
INIT_0E => X"3B000025EC010080004000F808000098100F22520008003B00002F2252000800",
INIT_0F => X"00001042006BC0810600400003B80001002F22520008003B00002F2252000800",
INIT_10 => X"01E032000620000C0405EC010100100000F6000001C1003760410500008000EE",
INIT_11 => X"201D2120840039000817444404040E10020218DE282010A311AA002002040080",
INIT_12 => X"8000000AE888808101C20040BA4241080072001027F00080200007E0000001F0",
INIT_13 => X"0101000003E2000007C0800FE04040280000F8080002F02023AC04080A00003D",
INIT_14 => X"DDAFD082001B03249887E04001D481D4000009020201E1A000040100F02023E8",
INIT_15 => X"ADAB6ADAB6ADAB6ADAB6ADAB6BF1EBDABD8E270BF84A25C6ACB777E3FF800C6D",
INIT_16 => X"DAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6",
INIT_17 => X"AB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6A",
INIT_18 => X"100481CA860402104A471688747FFFFFFFFFFFFFFFFFAB6ADAB6ADAB6ADAB6AD",
INIT_19 => X"0000000000000000000000000008200000000000200072F210000001490E2168",
INIT_1A => X"A05028140A05028140A05028140A050080402010080402010080000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000A05028140A05028140A05028140",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000",
INIT_22 => X"2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_26 => X"10FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFF",
INIT_2E => X"F5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA080402000000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"02000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FF",
INIT_36 => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_37 => X"0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000000FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(3),               -- Port A write enable input
DIA(0)   => data_write_a(27),        -- Port A data input
DOA(0)   => data_read_a_hi_512(27),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(3),               -- Port B write enable input
DIB(0)   => data_write_b(27),        -- Port B data input
DOB(0)   => data_read_b_hi_512(27),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_28_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"02200AA400180030808802A900002A08001280A08A801044104A1000001818C3",
INIT_01 => X"50A00011460214428114180000882214413D0A71592A01D92213D28005210202",
INIT_02 => X"8A54800A210200111100C2110054289220810440030404010844000444410001",
INIT_03 => X"4200040822D4500001E0000028000002000211842010092000018C6295200631",
INIT_04 => X"00400000000B8000000140000005840C00000040002008808100048100100044",
INIT_05 => X"0000222200244400135110000135100000000000000000024CA0A01018000320",
INIT_06 => X"A004912008208040024489121144080400081000200008104000000020000041",
INIT_07 => X"A85800994000000A0200802004204420210001022AA8A0001122448142491008",
INIT_08 => X"0414000201800004080A000000124058200408000880004440004080160C4100",
INIT_09 => X"0080000206CB0821082B694D4D29400002002038104000000020003204000440",
INIT_0A => X"12000843066021001400040024440245400082D022040000400800081022C000",
INIT_0B => X"0002002C004001036050160501605016050160501605016050160280B0280B00",
INIT_0C => X"0012400810080414C0A800310840102182C62302A0194C08001680100E4040A0",
INIT_0D => X"05000002003004208208841401800040000A0000200814004198000400020001",
INIT_0E => X"0500000004000080000000000000028000002052000000050000002052000000",
INIT_0F => X"0000300000004001060000000000000900002052000000050000002052000000",
INIT_10 => X"0000000001200000000004000100000000000000050000002001050000000000",
INIT_11 => X"00002020840000004800040404040000120200A9000000010000002002040000",
INIT_12 => X"0000004800808081000002400040410800000090001000002000000000000910",
INIT_13 => X"0001000000000000144000010000402800000000000A1000010000080A000000",
INIT_14 => X"0080000000110006B08140000040000000000902000000000000410010000100",
INIT_15 => X"0080200802008020080200802101210810C39A66A90A85420413A82000000204",
INIT_16 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_17 => X"8020080200802008020080200802008020080200802008020080200802008020",
INIT_18 => X"110A00246972BD89A40A0C22E100000000000000000000200802008020080200",
INIT_19 => X"82082082082082082082082082082082082082080D35050758C30C31DE21102C",
INIT_1A => X"B0582C160B0582C160B0582C160B0580C06030180C06030180C0820820820820",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000B0582C160B0582C160B0582C160",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000",
INIT_22 => X"2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_26 => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFF",
INIT_2E => X"F5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA080402000000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"02000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_36 => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_37 => X"0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000000FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(3),               -- Port A write enable input
DIA(0)   => data_write_a(28),        -- Port A data input
DOA(0)   => data_read_a_hi_512(28),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(3),               -- Port B write enable input
DIB(0)   => data_write_b(28),        -- Port B data input
DOB(0)   => data_read_b_hi_512(28),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_29_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"79964E4BA01DACAB9E659792D00AAE160002829C7FDFEFCEE97C2815039D70C3",
INIT_01 => X"50BFF9AB0775343F9AB01DF80D5821FC0FFF3FEFD1AF9FF1207FFBC7B9720586",
INIT_02 => X"0D15846807D207200021C4E200D428A2018408600271C000720A0000003A2161",
INIT_03 => X"0002C009EEFC5F10F9B70178681B80FA3E000100765029A00019084345606421",
INIT_04 => X"3E6E023D27DA937C03E3407712E5CDA41E0924DC3D20B98AE905189F0BF8C000",
INIT_05 => X"902003C30E0447F877F930203E213F8CF01E3E00FC67C03A4D9C87525E510160",
INIT_06 => X"0012460003CC002036040811D919F402244293FEE00400CCB46BA4C164A08857",
INIT_07 => X"914800110FFC0001CC320C81D841418E82800100000041FCA1428575A0001108",
INIT_08 => X"0805FD0180E1F8C1111A0782082B50080508FF00048B124D4005C8AFF4154102",
INIT_09 => X"0180000ABFEF89250815568A8AD6ABC02A02A0B0CCB463B4C0748A720B1EA4C0",
INIT_0A => X"021410028450530014014002D445624DB481806A62840800C22800B8900042FF",
INIT_0B => X"0806522C0A40A50268D0068D0068D0068D0068D0068D0068D006A68034680300",
INIT_0C => X"8912E0A83289641F42A80561D040203182AC3D0AA0118A080036FFFC4F4164A0",
INIT_0D => X"050080424069F5A51250648801BFFFE0003E3E00A0685A85410C0816040B0205",
INIT_0E => X"050080080400028000000000000202900000A0F600000005008000A0F6000000",
INIT_0F => X"00023000001040214E0000000000000D0000A0F600000005008000A0F6000000",
INIT_10 => X"000000000120400800080400030000000000000205800008200D070000000000",
INIT_11 => X"000220A2C400000068008424260400001A0241DAC80001010000042016040000",
INIT_12 => X"00020048108484C10000034004414588000000D04010001020000000010009B0",
INIT_13 => X"000900000000000416C00041000140E800000000010AB0001100008A2A000000",
INIT_14 => X"A282C0000033010FB181E00020400000000419060000000000004300B0001100",
INIT_15 => X"02C0B02C0B02C0B02C0B02C4B12B312912831A27FCFE7FFB175B6FF800802594",
INIT_16 => X"2C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B",
INIT_17 => X"C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B0",
INIT_18 => X"EE7FFDF7FE783FFDFFEA0C00602FFFFFFFFFFFFFFFFFC0B02C0B02C0B02C0B02",
INIT_19 => X"BEFBEFBEFBEFBEFBEFBEFBEFBEEBAEBAEBAEBAEBBFFDF9FBEFFFFFFEBBCF9F96",
INIT_1A => X"FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFBEFBEFBEFBEF",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000FBFDFEFF7FBFDFEFF7FBFDFEFF7",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000",
INIT_22 => X"2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_26 => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFF",
INIT_2E => X"F5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA080402000000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"02000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_36 => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_37 => X"0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(3),               -- Port A write enable input
DIA(0)   => data_write_a(29),        -- Port A data input
DOA(0)   => data_read_a_hi_512(29),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(3),               -- Port B write enable input
DIB(0)   => data_write_b(29),        -- Port B data input
DOB(0)   => data_read_b_hi_512(29),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_30_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"FF9FE1F7FFBFFFFDFFD000000000000000000000000000000000000000000000",
INIT_19 => X"79E79E79E79E79E79E79E79E79E79E79E79E79E7AFBD75F5FDF7DF7FF7FFBFFE",
INIT_1A => X"3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE79E79E79E79E",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE000000000000000003F9FCFE7F3F9FCFE7F3F9FCFE7F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000",
INIT_22 => X"2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_26 => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFF",
INIT_2E => X"F5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA080402000000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"02000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_36 => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_37 => X"0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(3),               -- Port A write enable input
DIA(0)   => data_write_a(30),        -- Port A data input
DOA(0)   => data_read_a_hi_512(30),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(3),               -- Port B write enable input
DIB(0)   => data_write_b(30),        -- Port B data input
DOB(0)   => data_read_b_hi_512(30),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_31_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"129000008004A00804A40000400800020000000C005FEA005800200400050100",
INIT_01 => X"A15FF18019700810180065FFFC0040801E80258CA2951C2200EC0906A0804140",
INIT_02 => X"146000808A0C060444692000402850040400408FF80000000010000000004000",
INIT_03 => X"000003F5D1202C70F654716A001A07F438184210960600000012108518004842",
INIT_04 => X"3E28FE3F6FE513703F70007472DA4128187B6DB530C1240A060C70580B439200",
INIT_05 => X"000F84040C088BE3E4AE40C1FD04CE38C0FC381FF8671FE01009048084C40010",
INIT_06 => X"0000000000000008000810200420620E00030BFE000181092CE7ED80DF800106",
INIT_07 => X"000000220FD1FF200040100540800000840200408002000C2244890200000200",
INIT_08 => X"0011F0780011E38004800E3CF3E0B1118C31747F000B33820209206FC9E80000",
INIT_09 => X"187FC301B124F2001600000000001A1F00110101092CE7ED81CF000401228800",
INIT_0A => X"0477330C4889CC012188310E08812982050800A91012494C31004124080886FE",
INIT_0B => X"9861D1403803800C1000C1000C1000C1000C1000C1000C1000C1800608006084",
INIT_0C => X"020400830602410901000D02D0002008012054040022102001017FE190022201",
INIT_0D => X"3A0000401E030B0C20C20188087FFA07FE203A80010002608030102008100408",
INIT_0E => X"3A000005E8010000004000F808000010100F02000008003A00000F0200000800",
INIT_0F => X"00000002006B80800000400003B80000000F02000008003A00000F0200000800",
INIT_10 => X"01E03200060000080405E8010000100000F600000081003740400000008000EE",
INIT_11 => X"201D0100000039000007404000000E1000001846282010A211AA000000000080",
INIT_12 => X"80000000E808000001C200003A0200000072000007E00080000007E0000000A0",
INIT_13 => X"0100000003E200000280800EE04000000000F8080000A02022AC04000000003D",
INIT_14 => X"9C06D082000A03200806A040019481D4000000000201E1A000040000A02022E8",
INIT_15 => X"0401004010040100401004010060C040040C200950402090128057C3FF800C60",
INIT_16 => X"4010040100401004010040100401004010040100401004010040100401004010",
INIT_17 => X"0100401004010040100401004010040100401004010040100401004010040100",
INIT_18 => X"000000000000000000001000802FFFFFFFFFFFFFFFFF81004010040100401004",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000",
INIT_22 => X"2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_26 => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFF",
INIT_2E => X"F5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA080402000000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"02000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_36 => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_37 => X"0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512,               -- Port A enable input
WEA      => wbe_a_hi_512(3),               -- Port A write enable input
DIA(0)   => data_write_a(31),        -- Port A data input
DOA(0)   => data_read_a_hi_512(31),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512,               -- Port B enable input
WEB      => wbe_b_hi_512(3),               -- Port B write enable input
DIB(0)   => data_write_b(31),        -- Port B data input
DOB(0)   => data_read_b_hi_512(31),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_0_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"ED39BA795990D275FB4A6E96ACC4731DEA4598B0AFB54867F6EE4618C3749803",
INIT_01 => X"58A0047C8607844847CA180001E4A2404042106208408208C2002069161734B3",
INIT_02 => X"8B1EC9562121F8051500147A0E5629A302CF28400615F5787B09FBF999BB1EFD",
INIT_03 => X"404EFC0A2AD6100F01A88E851CE47803C280110521898F6996088862C7B22221",
INIT_04 => X"C0D001C0100AEC83C008E7880D01A64661800002C21A52C590D2012194804844",
INIT_05 => X"650002C3F08754001B51981E007910070F01C1E003980015A204C22F32328BAF",
INIT_06 => X"BCDA4677CAEE7CF5BB870E1DDB9889C5FBFC440129A0604442180238203F70C1",
INIT_07 => X"7AAE0088B02000C2EC3A0E829836E0AF3325372E2AA8FDF3C18306758B24197A",
INIT_08 => X"D7E40002F7AE005FFB4730010411400A61080000F7F4C464B58294901606D5A5",
INIT_09 => X"C4801C40469B0CA9881A28C141118000C5A85A60444210123820B43B40804274",
INIT_0A => X"400800219010107ED453C041B13216656074EA560F0092A24856B05312226900",
INIT_0B => X"27122C3E04E03383E2781EA781E2781EA781E2781EA781E2781C33C0613C0E29",
INIT_0C => X"74EB1F50D0758A9650E520610A6A57A5529E2B439499CF96B086000000B09870",
INIT_0D => X"04F07E024108F4E28638EC57250004480155C1375A97A9121F8BA749D3A4E9D2",
INIT_0E => X"04F07E42177EFDF8570184071575970F8FC07D5BFF078004F07E007D5BFF0780",
INIT_0F => X"8F85ECB1FE047F5FB7B30E0700461E5AF8007D5BFF078004F07E007D5BFF0780",
INIT_10 => X"C0184D07C1DF15C7E3E2177EFDF8C3C03009C3CDD47C7F403FB3FDF89701C011",
INIT_11 => X"4F80FE659C6104C6D7103F9D1D064189B5924418D65FE45DEE55BBEDE34CF900",
INIT_12 => X"6395F64207F3A3A1483136B881FCCB38C2098DACA01FFF603F80001F80FDC81F",
INIT_13 => X"FED151E01015C3BB507D3F811FBEC32B81840714F8D91F4FC513F37C8AE07002",
INIT_14 => X"61692F293185D8D724E15D3FCC6B7C236FE0691A9500125C1F83F8CC1F4FC507",
INIT_15 => X"E93A4E93A4E93A4E93A4E93A4F942F90E9628540052090650525A0000066A00B",
INIT_16 => X"93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4",
INIT_17 => X"3A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E",
INIT_18 => X"09B56C74DAB15D1CF13501AA495000000000000000003A4E93A4E93A4E93A4E9",
INIT_19 => X"2082082082082082082082082082082082082082082084E41DC71C7155F3898E",
INIT_1A => X"3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F8208208208208",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE5294A5294A52800003E1F0F87C3E1F0F87C3E1F0F87C",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000030FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"A975EFFFAABDE00FFAEBDFFF5D2EAAAAAF7AEBDEBA0000000000000000000000",
INIT_22 => X"8000155087FC0155F7D168B55007BFDF45085168ABA002E82145085155545F7A",
INIT_23 => X"FFFD7545AA8028A00A2802AABAFF8028BEF5D7FFFE10005542145557FD5545FF",
INIT_24 => X"F7AEAAAAAA2FFFDF4500043FE105D2E954BAF7FFC0010080017555555568AAAF",
INIT_25 => X"A5D5168A00A2D142155005142010FFAE820AAFF842AABAA2AE95545FFD168ABA",
INIT_26 => X"FF5D2A821550000000BA007FD55FF5D7FC0145007FD7400550415410002E974B",
INIT_27 => X"F455D5142000082E82145FFD17DFEFFFD168BFFF780000BA007FE8AAAFF803FF",
INIT_28 => X"0000000000000000000000000000000000000000AAFBEAA00007BFDFFF082EBD",
INIT_29 => X"AABEA495FC716F002A975FFE3AA95E00EBAEBDFD75D2AA8A80EA8E2FE3F00000",
INIT_2A => X"56A16D557BC257D415E0216FA3F1E8FC0145B68B551475FAF6D1C556F0AA1C24",
INIT_2B => X"7FD24AFE3D02DAAAE12BD5545A2803AA0000542A0070071C50BAFEF1FAE0016D",
INIT_2C => X"A8B50F55A2F150005A3A438BD04AFAB8F550A8010E004924874825D7FEAA8548",
INIT_2D => X"A2A5504001C74BA42A1571E8028E3DB7816D0120155EA568E870BAEB8A05A2AE",
INIT_2E => X"2FFAFD2A82485FD2415A105C21451ED42A002545E055FFBE81D0BE8EA8A3AA05",
INIT_2F => X"100AA1D0F6F480B6A555A2A57A002A3D5FDB6A5C7E3DFFFE90B45B47ABA497A8",
INIT_30 => X"A0AFE80A8B0A000000000000000000000000000000000000000000000B55EAAA",
INIT_31 => X"ABEF5D557FEBA55022A3F70C6B405F4D2AE975EFAAAAB5E1AF3AABFF45592E88",
INIT_32 => X"411A8DED57CE1055555E5F58EFFC01FE2CACB65F520EBE9EF67D7BEA1FD5D556",
INIT_33 => X"A4AD0079C75D6070CC5CBB0280C029ABAA3EBC114728007521170821CE0FDE69",
INIT_34 => X"2A95E02A2AAB5EB0F280800EFAEE9F5D18F3142341D5DEEBEF55080034E0A592",
INIT_35 => X"B69C30E02116220415A9540AA854140A0A2047F353AAF6C77F7F20D968BF5781",
INIT_36 => X"ABEBE1B4D792A4AD1183454180DD3FDCAAAB7C91565455C141E41887D58AC448",
INIT_37 => X"F0000001FF01EABC4B8014174FF7DA80F52FEDE6BE93172D7D625B556EEAB157",
INIT_38 => X"FF0000001FF0000001FF0000001FF0000001FF0000001FF0000001FF0000001F",
INIT_39 => X"0000000000000000000000000001FF0000001FF0000001FF0000001FF0000001",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000100000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(0),               -- Port A write enable input
DIA(0)   => data_write_a(0),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(0),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(0),               -- Port B write enable input
DIB(0)   => data_write_b(0),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(0),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_1_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"212C001411984004084D000508C53810A03D1450E839B003342114428A000803",
INIT_01 => X"08000011400A100A81160000008C005400400002000000000000028001340000",
INIT_02 => X"C084484000002014400205851002007030450E0000A606C8C44CB4C6666C00E0",
INIT_03 => X"33DF380008164004000002000C80400002031943000101091608463061120118",
INIT_04 => X"4140008000000002000064000400004201000000000210458010070080100433",
INIT_05 => X"8500101040200000010009100000000508000100000000002010600100208D04",
INIT_06 => X"B5EDFDE24618AD433060C182BA860044204C000008A004100008000820280020",
INIT_07 => X"581E02100020000A81244890AA20263030517F122AA801F0983060AC564BF808",
INIT_08 => X"00820800C7A00045B103200000140A02234808000584000004808400020011A4",
INIT_09 => X"0000104000020082800808111008400000200204100000100820800144000414",
INIT_0A => X"12804062945211441E13C051156E800008402802060C94000040901102800000",
INIT_0B => X"24002006406401918C191AC191A4191A4191AC191AC191A4191A00C8560C8D29",
INIT_0C => X"0408010040050880383820080F105F05800302E0E08842422006000000041032",
INIT_0D => X"05000600000090C1841808172580000000008008020084082080204010200810",
INIT_0E => X"0500066210000178470184000000878402C000001E07800500062000001E0780",
INIT_0F => X"00003C404600000011A30E0700000009382000001E07800500062000001E0780",
INIT_10 => X"C0180000012010C20022100000F0C3C03000000055200340000000F88701C000",
INIT_11 => X"05800241186100004D100098190240001290002050068000001010486140F900",
INIT_12 => X"0000164A001303204800026880048230C2000094A0000F601F8000000001C908",
INIT_13 => X"12D051E01000000154200580003C030381840000004B08014401025480E07000",
INIT_14 => X"40082300218450C2800010094000482142E0601895001000000041C408014400",
INIT_15 => X"0802008020080200802008020080008208600500A82A15008000000000468000",
INIT_16 => X"8020080200802008020080200802008020080200802008020080200802008020",
INIT_17 => X"0200802008020080200802008020080200802008020080200802008020080200",
INIT_18 => X"BABEFC54A0810C7452B5420A1000000000000000000002008020080200802008",
INIT_19 => X"AAAAAAAAAAAAAAAAAAAAAAAAAAA28A28A28A28A2A8218D2C0C92492581328A46",
INIT_1A => X"2E974BA5D2E974BA5D2E974BA5D2E975BADD6EB75BADD6EB75BAAAAAAAAAAAAA",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFF6318C6318C63000002E974BA5D2E974BA5D2E974BA5D",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"00000000000000000000000C0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"002155557FFFFFF007FC21EFA2FFD74AAAAD5555550000000000000000000000",
INIT_22 => X"7FD75FFAAAA800AAF7AA974BAFFFBE8B45F7AEBDF455D2EAABEFF7FFE8BFF5D0",
INIT_23 => X"0557DF45AAD1400BAA2AE801550051555EFF7AA95400552AAAABAFFD1574105D",
INIT_24 => X"FFFBEAB55F780020AAAA80020AA082EAAB5500517DF555D2EAAA105500001550",
INIT_25 => X"AF7AE820AA0851574BAA2D1574AA5D7BFDEBAFFD540155557FD5400F78028BFF",
INIT_26 => X"FFFFD56AAAAFFFFD7555AAD168B45AAAEAAABAFF842ABEF5D517DF55552A974A",
INIT_27 => X"4BAF7AE80010082A97410557FEABFFAAFBE8BEFAAD1575EF557FFFE10557FFFF",
INIT_28 => X"00000000000000000000000000000000000000005D7FFDF4500043FE105D2E95",
INIT_29 => X"A8BC2EBDFEAF7F1F840017D4975D2FEF147FC51C7A2FBD5490BFD1C056A00000",
INIT_2A => X"AA8AAAE3D145410F7F1D55D71C002DABAEBAA974BAF7FFEFB45FFAABDF55492A",
INIT_2B => X"0E2AE85028B40155145F7AF6DBED5450AA1C2080BEF495FC71D54124924385FA",
INIT_2C => X"571D2E28E38E0216FA2D1E8E80140F45082B4002D082082AB8B6DBEDB7DF7F54",
INIT_2D => X"A97F7AF6D417E92482BF84020BA495557E3FF78E021FF1471FDEAAFFD56F16D5",
INIT_2E => X"7002FD74951D71EDFFABFD16FAAAE92BD5545A2DA3FB7DAAD4AAAAF487BC70BF",
INIT_2F => X"550A8010E00492487482FFFE82A85EBAE2FFC55554ADBD7A2FFC7BEFF6FFD7FC",
INIT_30 => X"400FBF9424F7000000000000000000000000000000000000000000000547AB8F",
INIT_31 => X"DF55F7AABFF55082CA8B4DF6C1E8F5E5400021EF005162BEF047FD5545AAFBF7",
INIT_32 => X"404547184164AA5D2EBEEB0A2D555410D3555714F8338AAAA1D0AE974AAF7FFF",
INIT_33 => X"AEABFFDF79DCBF755962010BDCBBC21455D7FEABEF75550ACBB7582225FF5843",
INIT_34 => X"D57D412F7D55F5E50C7F401BAAE8403CF5A3FFEAAEB083BC1000FF8409000512",
INIT_35 => X"2AA9FEAFDF7F431A9F7FFE81FF013A8001AFF801F8BA0C57740BDAA0688E5405",
INIT_36 => X"A2FBF7FED2C7F955445079E280A00C56145EF5D16BABAA3EBC3157ABD5FFE55F",
INIT_37 => X"0000000000596EBEF55080034E0A592A4AD00FB863550229BCABEB7DA403FFFD",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000100000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(0),               -- Port A write enable input
DIA(0)   => data_write_a(1),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(1),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(0),               -- Port B write enable input
DIB(0)   => data_write_b(1),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(1),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_2_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10E006600180111284380310006289800480032283E000A34301002001A0817",
INIT_01 => X"A14AC00A1079284D04A044A54E504368404000720885800802000006ECD10200",
INIT_02 => X"92250052A0348C310102048800A8507000040C8550200000480E0080001321E0",
INIT_03 => X"020204E4593C0824400C2220483042809292430400440180000890A4C9400242",
INIT_04 => X"486854B141002252142241502460480031B94420634850069A42241009610A04",
INIT_05 => X"800504244080892105AA6010A44882144840910A21220A8C820025E4A0000B00",
INIT_06 => X"A000442802280000340810209C444804206000AC800088096A0EA8C022208012",
INIT_07 => X"309820A848E0AA09826489A5CC49002001020112028201F8A20488260000108A",
INIT_08 => X"2400582881E0C1419D12041455509341A539C42A0D8208099002801700D10103",
INIT_09 => X"110D525861263100009200151409130A3C80C8C8096A06B8C12088400A9C2080",
INIT_0A => X"0451394CD0391A441583C04B580040089581001342801044877200D002A00DE0",
INIT_0B => X"144423040240450114901149013C9011C9013C9011C90134901144801A4808A5",
INIT_0C => X"D8A5345206D2C10082080A90C00000188150100C202A4640000E2B4081969420",
INIT_0D => X"050080400A0391A51240C480000AA902AA009028C83220008086952B4285A54A",
INIT_0E => X"05008021C00000000040000000020288000500000008000500802A0000000800",
INIT_0F => X"0002300000428000000040000000000D002A0000000800050080250000000800",
INIT_10 => X"0000000001204004000508000000100000000002054000130000000000800000",
INIT_11 => X"000C00000000000068144000000000001A000106200010021002000000000080",
INIT_12 => X"0002004A880000000000034098000000000000D024A000000000000001000900",
INIT_13 => X"00000000000000041400000A8000000000000000010A00000284000000000000",
INIT_14 => X"012100000002000280000000011080C000000000000000000000430000000260",
INIT_15 => X"A769DA769DA769DA368DA36CDA3A9A13A14801404134DA84A024024155000399",
INIT_16 => X"168DA769DA769DA769DA368DA368DA368DA769DA769DA769DA368DA368DA368D",
INIT_17 => X"68DA168DA169DA569DA569DA568DA168DA168DA169DA569DA569DA568DA168DA",
INIT_18 => X"138D70C030B51C50C7D000A2012F81F81F83F03F03F069DA569DA569DA568DA1",
INIT_19 => X"1041041041041041041041041041041041041041024860208165965975960040",
INIT_1A => X"25128944A25128944A25128944A25128944A25128944A2512894104104104104",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFF8421084210840703F25128944A25128944A25128944A",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"00000000000000000000000F0FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"415555087BFFF55A2AA800BAFFAE9540008002AA000000000000000000000000",
INIT_22 => X"7FE8B555551421455D0002145552EBFEBA007FC21EFA2FFD75EFAA8415410AA8",
INIT_23 => X"FFFE8B45552EBDF45FFAEAABFFF7FFE8B55F784155EFA2AEBDEAAA2FBEAABA5D",
INIT_24 => X"5D2AAAAAA5D2E820BAA2FBEAB5555557DF55A2AEBDF555D2E954BAA2AA974BAF",
INIT_25 => X"A5D04021EF557FC21FFAA8428BFFAAAA954AAAAAAAAAAAFFD1574105D7FFFF55",
INIT_26 => X"EFF7800215500557DF55AA80001FFAA80001550055575EFFF84021555D043DEA",
INIT_27 => X"B5500517DF555D042AA10A284154005D0015410085568A00FF80175FFA2D17DF",
INIT_28 => X"00000000000000000000000000000000000000005D00020AAAA80020AA082EAA",
INIT_29 => X"D55D2BE800042AFE8E1557D0075D2F45BEAA800AAFFAA9543A080038A2A00000",
INIT_2A => X"0BDEAAA2FBF8AAA557BE8B6D5D5FFABEF49040017D5D20B8EAA007FC51C7A2FB",
INIT_2B => X"0E174BFA02A974BAF7F5EFB455D2ABDF55492AA8BC7EBDFEAFEFFD00105FFBC2",
INIT_2C => X"3D155E105571D55D71C002DABA5524820BAB6FFEFB6D555578F7DB6A0BDF7D48",
INIT_2D => X"092A071555D5E3AE821D00001FF0871C016DBED1FDE90E3A497492B6AAADAAAE",
INIT_2E => X"0E3DA3DFD5E3DFFFBD5A38A021551C5F7AF6DBE8F401D7B6A0001470155C51D0",
INIT_2F => X"82B4002D082082AB8B6D1C5B7DF7FF78E075C5BE8555400550A38428007FED00",
INIT_30 => X"4AA00042AAA2000000000000000000000000000000000000000000000410F450",
INIT_31 => X"AAAA007FD5555AAFBD7545FBB8020A3F7AE975EF005560B55F7AA800AAF7AA95",
INIT_32 => X"E8F5EFF84165EFF7802BAB0A2FFEAABA557BEABEF057D68F5F5A00021EF55042",
INIT_33 => X"52ABFFFF841FFE75CA882108202E974AAF7D57DF55D7AABFF5428ACA8F45A6C1",
INIT_34 => X"84174A8FFAEBFEB0A2D55541051555694F002CA8AA80800020AAF7FBFFFEF045",
INIT_35 => X"7AAA155F595542455512A975455D3AA8A005500151FF0C57401E5F3D1E00A1A8",
INIT_36 => X"5D2A8A0B882FFFFE10AAAAAB755A66B6AF56A2AA801455D7FE8BFFF680800FFF",
INIT_37 => X"00000000000C3BC1000FF8409000512AEABFF5D79FCAF774AE005BE789555400",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000200000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(0),               -- Port A write enable input
DIA(0)   => data_write_a(2),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(2),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(0),               -- Port B write enable input
DIB(0)   => data_write_b(2),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(2),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_3_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"210C44A20020248B08431120001604B8156023104C4077133420400A02380202",
INIT_01 => X"015A2A424080216D3C2462C99E104B49404040028804A0080A000C16A0D90A0C",
INIT_02 => X"C0A4065000F0A95011000D1501005270B4045AB330860281CC08008222170060",
INIT_03 => X"AD22014098340394A4021320080841C40B411B4298042180002846B06900811A",
INIT_04 => X"244B32A86D20014A0D20403194904900071A24110F0BF400F85F92420E0C946E",
INIT_05 => X"80331030442898B4812840D0500008C528280B063006A64CA30004E5A4E40304",
INIT_06 => X"90016CA00E380042302040A0BC47160424428198C0038C89904E640023600816",
INIT_07 => X"1288020843A66620816049908AA0061011CA0142000009F0A810292E7402F088",
INIT_08 => X"20003C9984A0AC411102014D34EC2200214D5099048823019603A01A49410103",
INIT_09 => X"001CD74C4826220010A8891451284B661CA24A4C899046740121824004100080",
INIT_0A => X"44C9516DC0135C45159BE45F112B48804DC10203021290400772C0F402820D4C",
INIT_0B => X"B400624402404501A49018490184901A4901A4901849018C901A648056480C2D",
INIT_0C => X"D7A9B54000D7C10820680D08C420180381211081A022160000266723E1909021",
INIT_0D => X"400080200E199A4A2CA2994C0399981666409800CA52E4890806BD6B56BDAB52",
INIT_0E => X"40008008E00000000000000000024008000C8000000000400080028000000000",
INIT_0F => X"000A000000588000000000000000200400088000000000400080078000000000",
INIT_10 => X"0000001000004004000D800000000000000000022040000B4000000000000000",
INIT_11 => X"001A0000000000082006C000000000020804087220000122000A000000000000",
INIT_12 => X"00020800B8000000000041002E00000000001040466000000000000001020080",
INIT_13 => X"00000000000000048200004A600000000000000003008000320C000000000000",
INIT_14 => X"432900000222200871028000210400C4000000000000000000080200800030E0",
INIT_15 => X"AF6A5AF6A5AF6A5AF6A5AF6E5AFADA91AB68000101B4D20C08EC461733804A19",
INIT_16 => X"B6B5AF6A5AF6A5AF6A5AF6A5AF6A5AF6A5AB6B5AB6B5AB6B5AB6B5AB6B5AB6B5",
INIT_17 => X"6BDAB6B5A96ADAF6A5AD6ADAF6A5AD6ADAF6A5AD6BDAB6B5A96BDAB6B5A96BDA",
INIT_18 => X"C78C706428A14C586290008A044D54AAB556AA9556AAEBDAB6B5A96BDAB6B5A9",
INIT_19 => X"92492492492492492492492492410410410410412821600001249249015303C0",
INIT_1A => X"351A8D46A351A8D46A351A8D46A351A9D4EA753A9D4EA753A9D4924924924924",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000001543B351A8D46A351A8D46A351A8D46A",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"43DF55FFAA955EFA2D168B55557BEAA000055420000000000000000000000000",
INIT_22 => X"7BE8BFFA2D155410AA8415555087BFFF55A2AA800BAFFAE9554508002AA00AA8",
INIT_23 => X"52ABFEBA007FC21EF007FD75FFAA841541008002AB55AAAA955EF005568A0008",
INIT_24 => X"005168B455D042AB45F7FFD741000042AA10AAAABFF5508003FF555D00021455",
INIT_25 => X"0A2D1575FFF7AA975555D2E80145F78415545082EBDEAAA2FBEAABA5D7FC0155",
INIT_26 => X"55552A954BAFFFFE8B55552EBDE00F7AEAABFFF7FBEAB55F7AABDEBA5D7FC201",
INIT_27 => X"F55A2AEBDF555D2E954BA002EAAABA002A821EF5555554AA087BC01FFFFAAAAB",
INIT_28 => X"0000000000000000000000000000000000000000082E820BAA2FBEAB5555557D",
INIT_29 => X"95578080038A2AA28E3AF55E3A0BA5D7AADB6FB7D5D7FEAA3808554203A00000",
INIT_2A => X"0925D7085F6AA10087FEABD7AAD57AEBAB68E1557D1475FAF45BEAA800AAFFAA",
INIT_2B => X"04AAFFA41040017D5D20B8EAA007FC51C7A2FBD55D7BE80004AA1E8E2AB55B6A",
INIT_2C => X"2FBE80AA557BE8B6D5D5FFABEF49002FB55FFF5D0438140E2FA38B6AEBFF6D1D",
INIT_2D => X"AB8ABAE925D21C7010EADB525D7FFAE975C75D0A901FFFF801557D1C20B8EAAA",
INIT_2E => X"20875C21D5EB8AA8FFF012A954BAFFF5EFB455D20BDE00EBAAA8BC7EBDFEAFEF",
INIT_2F => X"BAB6FFEFB6D555578F7DB6A0BDF7DEB8E125FF002EADA921420871D74971D248",
INIT_30 => X"ABA0051400A20000000000000000000000000000000000000000000001C24820",
INIT_31 => X"8B55F7AA800BAF7AA955EF00042AAA2A2AEAAB55A28408145AAFFFFFFF5D7FEA",
INIT_32 => X"020A35D2ABEF55F7800015F087FEAA00007FEAB55FAD568AA2AFAE975EF55516",
INIT_33 => X"ABFEAAF7AE9DFF759A82AEF70800021EF55042AAAA007FD55558A7BD7145FBB8",
INIT_34 => X"84175EF55002AAB0A2FFEAABA557BEA3EF057968F575D003FF55F7D5420BA5D2",
INIT_35 => X"A8429F45A7D5EAF5FFBAEAAA10554155400AAFFD5145FBAC9755F05040255FFD",
INIT_36 => X"550415557085540000005156155FE90A8F5C082E974AAF7D57DF45552A3FF10A",
INIT_37 => X"00000000005500020AAF7FBFFFEF04552ABFFFF843FFE77C80825BC052ABFE10",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000100000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(0),               -- Port A write enable input
DIA(0)   => data_write_a(3),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(3),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(0),               -- Port B write enable input
DIB(0)   => data_write_b(3),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(3),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_4_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A108400020612C80284210081034849800A000303100048B3432C82904204002",
INIT_01 => X"21066802000820491C00650E1E004360403008418984014902030906A8D10200",
INIT_02 => X"120404E00E4C0600000206100008402005040C00F104008040080080001310E0",
INIT_03 => X"DCA201514D1C0D706C5CF010083A0708BA0841945004010000080084C1000002",
INIT_04 => X"5C4CF21C48B133483C80417570D000083A62488074C1350EA60D785C0A6B0619",
INIT_05 => X"000F0400028083B381A60001E5546EB5C0E2B81E4166DE000139200004E50940",
INIT_06 => X"80004408020800023000102098000204A040038600018019004B800123208806",
INIT_07 => X"120C20204665E1008024188488800000001A01520000A1F08044892400001088",
INIT_08 => X"0801007AC0A1EB413102063CF3E0B3028D29F407059B0B000205A801C2200102",
INIT_09 => X"106052400922D00406BE1002C6150F41200280001900439001FD8A0004142000",
INIT_0A => X"047F2201D899BA503583504B58AB80804540001202805544314041B48A888EC5",
INIT_0B => X"1441E3443043410C5010C3010C1010C3010C1010C1010C3010C14086980861A5",
INIT_0C => X"020000A02600000805400502C0A0004A00625015000A12000026E1E180011220",
INIT_0D => X"400000000E43930C20C20188120782861E4004A800600401A030001008080400",
INIT_0E => X"40000021A8800000000000000000400800170024000000400000310024000000",
INIT_0F => X"0008000000AA80200800000000002000003400240000004000003B0024000000",
INIT_10 => X"00000010000000040004A080000000000000000020400006C008020000000000",
INIT_11 => X"002C008200000008001B4020200000020000090760000200110A040010000000",
INIT_12 => X"00000803E004040000004000E801040000001000086000000000000000020040",
INIT_13 => X"0000000000000000810000164001008000000000020040002240008020000000",
INIT_14 => X"04001040026026004000000002940040000410000000000000080000400000B8",
INIT_15 => X"040080201004008060000001806AC000004890015124D880100886D8F0014420",
INIT_16 => X"4010000180600000018020100400802010000080601000008020000401802000",
INIT_17 => X"0100000004008020180600000000000180600802010000000401802018020000",
INIT_18 => X"3807E05000140634504048820064B261934D964C326980004010000080600806",
INIT_19 => X"AAAAAAAAAAAAAAAAAAAAAAAAAAA28A28A28A28A2934C8D0CCD145144C0A28A06",
INIT_1A => X"068341A0D068341A0D068341A0D068351A8D46A351A8D46A351AAAAAAAAAAAAA",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000000173F068341A0D068341A0D068341A0D",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"57FE10FFFBEAA10007FD7410FFAA97555082A800AA0000000000000000000000",
INIT_22 => X"7FEAA00007BE8AAAAA843DF55FFAA955EFA2D168B55557BEAB45005542000005",
INIT_23 => X"87BFFF55A2AA800BAFFAE9555508002AA000055574105D2A800AA00043FEBA5D",
INIT_24 => X"A2D17DE1000517FE10AAAAA8AAA002E97545557BC00AAA2FFEAAAAAA84155550",
INIT_25 => X"0A2D157400AAAE974AAAAAA974BA08002AB55A2AA955EF005568A00087BE8BFF",
INIT_26 => X"BA080002145552ABFEAA007FC21EF007FD75FFAA8417410A2D140000F7FBC201",
INIT_27 => X"A10AAAABFF5508003FF55F7D568A00552EA8BEFA2AABDEAA087BEAAAAA2FBD54",
INIT_28 => X"000000000000000000000000000000000000000055042AB45F7FFD741000042A",
INIT_29 => X"EAB7808554203A145178E00FFFBE8A101475D5400F7A49057D0824850B800000",
INIT_2A => X"E8008200043FE925571EFA380871C7028A28E3AF55F7A0925D7AADB6FB7D5D7F",
INIT_2B => X"F5FDA38BE8E1557D1475FAF45BEAA800AAFFAA9557D080038AAA145157428492",
INIT_2C => X"85F6AA10087FEABD7AAD57AEBA08517DE00AAAEA8A9200249056D4175C5092AA",
INIT_2D => X"FEDB42028EBFBC2028BED152438AAA092492AAA4954281C0E2FB55B6A0925D70",
INIT_2E => X"A0875EDA80BEF1C743840040017D5520B8EAA007FC51C7007BD55D7BE80004AA",
INIT_2F => X"55FFF5D0438140E2FA38B6AEBFF6DBE84AAEBAF7DF6AA00412EAABFFAA803DEB",
INIT_30 => X"1EF0800154B200000000000000000000000000000000000000000000041002FB",
INIT_31 => X"0145AAFFFFFEF5D7FEABFF0051400A25D5568A00FFFFEAA105D5155410FF8402",
INIT_32 => X"2AAA25555410BA082E8201000043FE005D517DEBA0851574B2AAAEAAB55F7840",
INIT_33 => X"4001FF005575408AA557FEB2FFAE975EF555168B55F7AA800BAF7AA955EF0004",
INIT_34 => X"2ABFF55F7800015F087FEAA00007FEAB55FAD568AA200557DE00AAAAAAA00080",
INIT_35 => X"87BD6145FAAC000A2A6FBC00BAAAFBC00BAF7D1550AAAA8002010F2AC154B25F",
INIT_36 => X"082EA8BFFAA843FEBA08517DE00F3F9574B30800021EF55042AAAA007FD55550",
INIT_37 => X"000000000008003FF55F7D5420BA5D2ABFEAAF7AEBDFF779A82AA43F7FBE8A00",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000200000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(0),               -- Port A write enable input
DIA(0)   => data_write_a(4),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(4),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(0),               -- Port B write enable input
DIB(0)   => data_write_b(4),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(4),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_5_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50DF4A0791B3FCB694379283C81FD996A091832102004A337A20E07C0C1E006",
INIT_01 => X"294014468000A04D5C6A60000C34C24841280A00084000C8C212892EEAD53235",
INIT_02 => X"50AE41540CA1D9100002171C1F0A5171134E2A200D8633F8CD09DBFBBB970E7C",
INIT_03 => X"214E3C521D16021B64430CC51C45B8154689094241898749920842946B90010A",
INIT_04 => X"A2F20F7D7A314CB5C208E28A1BF0224A448920028A185340D0C20B2690000C22",
INIT_05 => X"7520B430B20B984809A8886E230C6106371146E1829941C58310402C600381CF",
INIT_06 => X"9CC96CD7C63A7495B9A356ACBC4601C57FD44F8549A46490261C4B39203F7080",
INIT_07 => X"12A88800B029E0C0A12C4B92AA36A2111167357C220095F3C8952A2E5D26F078",
INIT_08 => X"F3F00503B4AE105B534711820C0C0A1043080300F7E0E728B1829C2FEA0A95A1",
INIT_09 => X"C5184F084136848C9298A8560688F480C58858449026145B3830F40944906234",
INIT_0A => X"50EB4124D2B3902BF5C9700C1199DCA84DF46A974F92C7E28F1630D38088A438",
INIT_0B => X"B3144E5636E3178C86B8CC6B8CA6B8CE6B8C86B8CE6B8CA6B8CC15C6435C670C",
INIT_0C => X"79E51E70E070AA8132252008360A7E91504104C8948047D6B0AE1FE440B28A71",
INIT_0D => X"05F0FE40014090400400080329FF8089FF49611F589765923E139F09C78CE7C6",
INIT_0E => X"05F0FE64037FFD7857418407157797878F005F0DFF0F8005F0FE205F0DFF0F80",
INIT_0F => X"8F87FCB1F8053FDEB9B34E0700461E5FF8205F29FF0F8005F0FE205F29FF0F80",
INIT_10 => X"C0184D07C1FF55C3E3E0037FFCF8D3C03009C3CFD53C7E001FF2FAF89781C011",
INIT_11 => X"4E0CDF47186104C6FF177BD939024189BF900401165D645CEEF5BBCDF148F980",
INIT_12 => X"6397F64AEF7F2320483137F8A9BF8A30C2098DFCA06FFFE01F80001F81FDC94F",
INIT_13 => X"FFD051E01015C3BF553D3E0E5FFE838381840714F9DB4F4FA213F774A0E07002",
INIT_14 => X"8B652E2B3120C81284641D3E8DBF7D636FE070189500125C1F83FBCC4F4F80EF",
INIT_15 => X"E7394E339CE138CE5394E33D4E1E0E30E1208C251134921C12A44103F064014B",
INIT_16 => X"7384E3394E338CE538CE1394E3384E738CE139CE1394E7384E339CE139CE5384",
INIT_17 => X"38CE139CE1384E7384E7394E3384E738CE539CE139CE538CE5384E3394E7384E",
INIT_18 => X"7F7B9DB7FF3A1B6DB7ED438A9C3124B2DA6924965B4D384E7384E339CE138CE5",
INIT_19 => X"FBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEF9F7CFDFDDCF3CF3DF5E5BB4E",
INIT_1A => X"7BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEFBEFBEFBEFBE",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE000000000000118D27BBDDEEF77BBDDEEF77BBDDEEF7",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"E955450055421FFFFFBC0010AAD5574BA557FFDFFF0000000000000000000000",
INIT_22 => X"D5575EF55517FF5500557FE10FFFBEAA10007FD7410FFAA97410082A800AAAAA",
INIT_23 => X"FAA955EFA2D168B55557BEAB55005542000007FD74000055574BA5D7FD7555A2",
INIT_24 => X"007BC00AAAAAEBDF45A28428B45FFD168BFF00002AABA5D2ABFFFFAA843DF55F",
INIT_25 => X"AFF80174BAAAD1555EF5555555550055574105D2A800AA00043FEBA5D7FEAA00",
INIT_26 => X"FFAA8415555087BFFF55A2AA800BAFFAE95555080028A00A2FFFDE00F7D57FEB",
INIT_27 => X"545557BC00AAA2FFEAAAA082A97545F7D5420BA5D2E821FFA2D5554BA557BD75",
INIT_28 => X"000000000000000000000000000000000000000000517FE10AAAAA8AAA002E97",
INIT_29 => X"9043D0824850B8A2AE9756D145B401FFFFFFC7010BEDF524AA5571FDFEF00000",
INIT_2A => X"1524BA5571D757DB6D5525EF555178F6D145178E00EBFBE8A101475D5400F7A4",
INIT_2B => X"24BFFFFA28E3AF55F7A0925D7AADB6FB7D5D7FEAB7D0855420BA1471D7438085",
INIT_2C => X"0043FE925571EFA380871C7028B6AEBDF45B68A28B6DEBDF6DBEF1C0A28AAA55",
INIT_2D => X"A2FBF8E10EBD578EAAFF8415482BED1555EF55555057D145152428492E800820",
INIT_2E => X"FB6DF574A85575C55EFBE8E1557D1475FAF45BEAA800AAFFAA9557D080038AAA",
INIT_2F => X"00AAAEA8A9200249056D4175C50920875FDA381C209256DFFDF420BA552A821F",
INIT_30 => X"0BA55557DFF700000000000000000000000000000000000000000000008517DE",
INIT_31 => X"AA105D5155410FF84020AA0800154B2AAAA975FF5D7BC21EFF7FBD7400F7FBC0",
INIT_32 => X"400A25551554BA0051400BA5551575EFF7D1401FF5D5568BE7555568A00AAFFE",
INIT_33 => X"FFDFFF552EA8AAA55043DFF7AAAEAAB55F78400145AAFFFFFEF5D7FEABFF0051",
INIT_34 => X"55400BA082E8201000043FE005D517DEBA0851574B2FFAABFF45FFAAAABFFAAF",
INIT_35 => X"7AA955EF00002AAA2A2FBE8A00A2D16AAAAFF8002410FFD5575EF5555421E755",
INIT_36 => X"FFFFC00BA552A821EFFFFFD74BA5D51575F7FFAE975EF555168B55F7AA800BAF",
INIT_37 => X"000000000000557DE00AAAAAAA000804001FF0055554088A557FEB25D00021FF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000C00000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(0),               -- Port A write enable input
DIA(0)   => data_write_a(5),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(5),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(0),               -- Port B write enable input
DIB(0)   => data_write_b(5),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(5),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_6_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10800B0061A01002840002C03002818000402322520070B313301C4389B2082",
INIT_01 => X"274008482009404C18A160000C52424841000000090800090210000008510200",
INIT_02 => X"102430600C800110000006100009D070012408000000000648080000001210E0",
INIT_03 => X"000200501D1D02140C420200480140040608010040400104681A0084490C4802",
INIT_04 => X"404402820021000A00824002141000980500000808001114C000080624600600",
INIT_05 => X"120024204209981001A806500304610528000500000080000000300000012940",
INIT_06 => X"2000440832280002300010209C4400142061207A024008900008000220600220",
INIT_07 => X"130C8A220FF41F00902008808800182001020150000001F0800408264000100A",
INIT_08 => X"001BF002C4A01041B1120101000010128568837F04842B080020890008080342",
INIT_09 => X"011847140126805432A62A1596C8B5DF10000008900000100220C00084000008",
INIT_0A => X"44EB4104D09392053589F11C59898888454010830212C54081000410A0088C00",
INIT_0B => X"B0044245B25B456C0096C0096C4096C4096C2096C2096C6096C444B6004B600C",
INIT_0C => X"09040020280010000B3002820110101D0012402CC00802410C26800860070621",
INIT_0D => X"0500819D0000900208201040C4007920004884080000448C281018100C000200",
INIT_0E => X"05008182100000000000000000022AE800C00004000000050081A00004000000",
INIT_0F => X"0002330006000000080000000000000D07A00020000000050081A00020000000",
INIT_10 => X"0000000001204A340002100000000000000000020F4001400000020000000000",
INIT_11 => X"019300020000000068D08000200000001A692121000280000000000010000000",
INIT_12 => X"000201FA100400000000034696010000000000D3478000000000000001003F00",
INIT_13 => X"00000000000000043C0001C0A000008000000000012E000054AC000020000000",
INIT_14 => X"0200000040A410C2810800016000809400001000000000000000433300007600",
INIT_15 => X"060180400000008060180404002AC0200208940041309210B28048180F028000",
INIT_16 => X"2008000100601802000000100601800000000180600800000020180600000000",
INIT_17 => X"0180600000008040100200800000060100000802010040180200002018040100",
INIT_18 => X"7F8FF0F4FA955F7CF7F40A80907638C31C71C718638E00006018040080200004",
INIT_19 => X"38E38E38E38E38E38E38E38E38E38E38E38E38E39B6CEDECDDF7DF7DF5F78BCE",
INIT_1A => X"3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE38E38E38E38E",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFF000000000000196A03F9FCFE7F3F9FCFE7F3F9FCFE7F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"00000000000000000000000C0FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"BFDF45F7AA974AAAAAA97555F784174BAF7D5555FF0000000000000000000000",
INIT_22 => X"FBD7410AA8428AAAAAAE955450055421FFFFFBC0010AAD5574BA557FFDFFF087",
INIT_23 => X"FFBEAA10007FD7410FFAA97400082A800AA08515555508043FE00F7AA97555A2",
INIT_24 => X"55517FF55A2AA97400552AAAB45082E80155F7D1575EFFFAA9555500557FE10F",
INIT_25 => X"FF7AAA8A10082EAAB45A2FFC2000007FD74000055574BA5D7FD7555A2D5575EF",
INIT_26 => X"FFAA843DF55FFAA955EFA2D168B55557BEAB5500554200000003DE10FFD5401F",
INIT_27 => X"BFF00002AABA5D2ABFFFF087BD5545007BFDE10AA803FE105D516AABAFF843FF",
INIT_28 => X"0000000000000000000000000000000000000000AAAEBDF45A28428B45FFD168",
INIT_29 => X"524AA5571FDFEF1C7BFFF55FFA095482B6A49256DEB84104BAFFD1525FF00000",
INIT_2A => X"03DE28F7A49057DAAF5D2428A2842AAAAA2AE9756D145B401FFFFFFC7010BEDF",
INIT_2B => X"A49756D145178E00EBFBE8A101475D5400F7A4904380824850381C5B5057D1C0",
INIT_2C => X"571D757DB6D5525EF555178F6DAAA495428412AAFB451C2A8017DE3DF525FFFF",
INIT_2D => X"1C0E3FE00E3DB471EFE3AAAAA00082EA8B6DA2F1C50381471D74380851524BA5",
INIT_2E => X"049516AAB8FF8428FEFA28E3AF55F7A0925D7AADB6FB7D5D7FEAB7D0855420BA",
INIT_2F => X"45B68A28B6DEBDF6DBEF1C0A28AAA5524BFFFF1C7BD057D1C71FFE10A28038E1",
INIT_30 => X"0AAFFD1401E7000000000000000000000000000000000000000000000B6AEBDF",
INIT_31 => X"21EFF7FBD7400F7FBC00BA55557DFF7557BFDF55F78017400F780001FFAA8400",
INIT_32 => X"154B2557FC01EF55043FEAAFF80021EFA2D1420BAAA8428AA2AAAA975FF5D7BC",
INIT_33 => X"A821EFAAFBC01FFF780155F7555568A00AAFFEAA105D5155410FF84020AA0800",
INIT_34 => X"51554BA0051400BA5551575EFF7D1401FF5D5568BE7AA80174AA082ABDF555D2",
INIT_35 => X"D7FEABFF0051400A25D2EBFE10AAFFD55EFA2AEA8A10082EA8BEFAAD5554B255",
INIT_36 => X"55557DE00AA842AA0000516AABAFF8428BE7AAAEAAB55F78400145AAFFFFFEF5",
INIT_37 => X"0000000000FFAABFF45FFAAAABFFAAFFFDFFF552EA8AAA55043DFF7557BC01EF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000900000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(0),               -- Port A write enable input
DIA(0)   => data_write_a(6),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(6),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(0),               -- Port B write enable input
DIB(0)   => data_write_b(6),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(6),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_7_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10844B00482258A2842112C02450418800002300500030B313300C418992002",
INIT_01 => X"234008422008604D1C20E0000E11426840000000080000080200090000110204",
INIT_02 => X"1025207000B08910000206101188D03080144880010400044808000000122160",
INIT_03 => X"000200401914821004420000CA01000C0600010000605114291A008449484802",
INIT_04 => X"40440200002100080006500210101019040000000B085024D842080244000000",
INIT_05 => X"1A8024200009981001A8224001040104200204000000800CC2092CE4A0004900",
INIT_06 => X"A000440822280002340010209C040014A061200052500810000C490323208E28",
INIT_07 => X"128802020028000890240980A809102001020140000009F0800408264000100A",
INIT_08 => X"001A0602C4A01051B13281010408881203480200448423199046821008082351",
INIT_09 => X"336784144126811054809C1040140A001C8648481000045903318B80A400310A",
INIT_0A => X"000800009010100014114110312388984502148282A08415B032095048008100",
INIT_0B => X"20CDC1C483484D201192011920119201192051920519205192074C9018C90188",
INIT_0C => X"D8A5B44001D2C12901228F82F005310D293054048A2212004466000DA1908528",
INIT_0D => X"800F8108A0D09802082010408580008000000008C85264010816851B428DA146",
INIT_0E => X"800F81321000020000261900E28A204040E000A0000007800F814000A0000007",
INIT_0F => X"7072024807000020400000581C01C1A406400084000007800F81400084000007",
INIT_10 => X"060180E83800E820101210000200000CC3003C32080201C0000C000000160700",
INIT_11 => X"81DD00804086423120B74020023090644840A34000828800000004000420020B",
INIT_12 => X"1C6A0186E8000446120C8905BA0004810C84624237E00010001878007F0030C0",
INIT_13 => X"00080208E4083C44230201AEE0010040261900E30520C0806EAC0082000984C0",
INIT_14 => X"0121011088A600C032128201519480D40005802448160403E0700622C0806EE8",
INIT_15 => X"A1685A1685A168DA368DA36CDA30DA13A108810111349A943AA4401000928A19",
INIT_16 => X"368DA768DA1685A1685A5685A368DA368DA7685A1685A1685A768DA368DA368D",
INIT_17 => X"685A1685A169DA368DA1685A1695A368DA3685A1685A168DA368DA1685A1685A",
INIT_18 => X"00000000000000000000400A8448410400020820800069DA1685A168DA369DA3",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000003667B000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"0155EFAAAEA8ABAAAFBFDE0055556AA005D04155550000000000000000000000",
INIT_22 => X"556AA00FFAE95555087BFDF45F7AA974AAAAAA97555F784174BAF7D5555FFF78",
INIT_23 => X"055421FFFFFBC0010AAD5574BA557FFDFFF5555555EFAAFFFDFEFAAAAAAB455D",
INIT_24 => X"AA8428AAA557BFDFFF55003DFFFF7FBEAA00002EAAAAA082EA8A00AAAE955450",
INIT_25 => X"0552EBDE00007BEAAAAA2D14000008515555508043FE00F7AA97555A2FBD7410",
INIT_26 => X"FF00557FE10FFFBEAA10007FD7410FFAA97400082A800AAF7AE975FFA2800001",
INIT_27 => X"155F7D1575EFFFAA955555D51574AAAAFFD5545087FEAB455D516AB55557BD55",
INIT_28 => X"0000000000000000000000000000000000000000A2AA97400552AAAB45082E80",
INIT_29 => X"104BAFFD1525FFFF8E175C7A2AAAAA82A2F1FAE105D556AA10410E1755500000",
INIT_2A => X"1FFFD7AAAAAFB7D495F6AA10E3AE905551C7BFFF55FFA095482B6A49256DEB84",
INIT_2B => X"2EAAA00A2AE9756D145B401FFFFFFC7010BEDF524AA5571FDFEF415B575D7AAF",
INIT_2C => X"7A49057DAAF5D2428A2842AAAA497BFAFFF49003AFEFEBFBEAA001C2EA8A821C",
INIT_2D => X"F7A4905C7A28A070384120BDE100075EAA82BEDB470101C5B5057D1C003DE28F",
INIT_2E => X"D555F6AB57417BC05D7145178E00EBFBE8A101475D5400F7A490438082485038",
INIT_2F => X"28412AAFB451C2A8017DE3DF525FFFFA49756D495150492BEF1D2555087BE8B7",
INIT_30 => X"A10002E9754D000000000000000000000000000000000000000000000AAA4954",
INIT_31 => X"7400F780001FFAA84000AAFFD1401E7FFAA97555A2AEA8A10AAD568A00555168",
INIT_32 => X"7DFF7007BD5555AAD57DF55AAAEBDFEF007BE8A10AAAE8215D557BFDF55F7801",
INIT_33 => X"FEAA105D2EAAA005D2AAAA18AAAA975FF5D7BC21EFF7FBD7400F7FBC00BA5555",
INIT_34 => X"7FC01EF55043FEAAFF80021EFA2D1420BAAA8428AA2007FE8BFF080028BFFAAF",
INIT_35 => X"F84020AA0800154B2FF8402145A2AA954AA00043DE0000516AA10F7FBD740855",
INIT_36 => X"FFD140145007FE8BEF557BEAB55087FC215D555568A00AAFFEAA105D5155410F",
INIT_37 => X"0000000000AA80174AA082ABDF555D2A821EFAAFBC01FFF780155F7005140000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000000FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(0),               -- Port A write enable input
DIA(0)   => data_write_a(7),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(7),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(0),               -- Port B write enable input
DIB(0)   => data_write_b(7),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(7),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_8_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00000648E2840112C00000418000002700500030B3132000400812086",
INIT_01 => X"214009C21838284D042100000212026840000000180800080200080040510204",
INIT_02 => X"1021004000900110000006100088503000240800014400004808000000122160",
INIT_03 => X"0002004019110214044A82000121400C86000000000000860188008448400002",
INIT_04 => X"000402800031200A0000090214100889A5000000490090104800000224000400",
INIT_05 => X"10C025204289981000A820500344010428008500010080080909304040202004",
INIT_06 => X"8000440003280000340010208C04003420600000C6180810000C490703200010",
INIT_07 => X"130002000028000890240980A809012001020050000009F08004082640000082",
INIT_08 => X"20100402C4201041310041010008801201480200051023090024811008090A1A",
INIT_09 => X"0100001001248100308214528148A48008000008100004590711C04034000083",
INIT_0A => X"10804000801210140001C0103001088845010482004000008420041020008900",
INIT_0B => X"0004404002004400448000480004800048000480004800048000440022400200",
INIT_0C => X"880420000880204909004502D100A10C04205424010216010C26800805000004",
INIT_0D => X"8000801100509802082010400400018000488428800004082014000200010000",
INIT_0E => X"8000800A00000207A8BE7B00000200082040808000F07F80008000808000F07F",
INIT_0F => X"0002000402100000404CB1F8FC0000040000808000F07F80008000808000F07F",
INIT_10 => X"3E07800000004004080A000002072C3FCF0000020040804800040007687E3F00",
INIT_11 => X"10800018639EC00020100002C2F9B0000801016001008100000040120CB3067F",
INIT_12 => X"000200020000585EB6000100800030C73D8000402000001FC07FF80001000080",
INIT_13 => X"002EAE1FEC0000040200408000003C547E7B00000100801004000803551F8FC0",
INIT_14 => X"00000000440610C8000A808040000208901B86E568FE0C000000020080100400",
INIT_15 => X"0040100401004090240902449028D0230249850101349A98BAC0481000888810",
INIT_16 => X"0401004010040100401004010240902409024090240902409004010040100401",
INIT_17 => X"4010040100409024090240902409004010040100401004090240902409024090",
INIT_18 => X"543EBC57A10A1E75D6440A889050000000000000000040902409024010040100",
INIT_19 => X"79E79E79E79E79E79E79E79E79E79E79E79E79E7BF3CCD8DF5B2DB2CA4028A0A",
INIT_1A => X"4F87D3E1F4F87D3E1F4F87D3E1F4F87C3E1F0F87C3E1F0F87C3E79E79E79E79E",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000000D3E94F87D3E1F4F87D3E1F4F87D3E1F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"000000087BEAA10F7803DE00FFAEBFFFF0800155FF0000000000000000000000",
INIT_22 => X"7FC2145005155555F780155EFAAAEA8ABAAAFBFDE0055556AA005D0415555080",
INIT_23 => X"7AA974AAAAAA97555F784174BAF7D5555FF552AA8AAA557FC0010F780154105D",
INIT_24 => X"FFAE95555AAFFE8A00552EBFE00F7D17FF45F7FFFFF55AA80155FF087BFDF45F",
INIT_25 => X"5F7D140010552E821EFAAAABDF555555555EFAAFFFDFEFAAAAAAB455D556AA00",
INIT_26 => X"00AAAE955450055421FFFFFBC0010AAD5574BA557FFDFFF5504000AAAAAAA8B5",
INIT_27 => X"A00002EAAAAA082EA8A00002AA8A10F78402155AA8028A00A2D57FF45557BE8A",
INIT_28 => X"0000000000000000000000000000000000000000557BFDFFF55003DFFFF7FBEA",
INIT_29 => X"6AA10410E17555080E000280071E8A00EB8E3FE10F7AEBAFFF080A175D700000",
INIT_2A => X"1C2000FF8A17400557FC015514555757DFF8E175C7A2AAAAA82A2F1FAE105D55",
INIT_2B => X"8A105D71C7BFFF55FFA095482B6A49256DEB84104BAFFD1525FF492EA8AAA557",
INIT_2C => X"AAAAFB7D495F6AA10E3AE90555A2FBE8A38492ABDE10EBDF7AF6DE3FFF8F7DB6",
INIT_2D => X"550E00082B6A0AFB55F7D1420104124821D7AAA0BDF6D415B575D7AAF1FFFD7A",
INIT_2E => X"0B6D578F6D557FFDA00A2AE9756D145B401FFFFFFC7010BEDF524AA5571FDFEF",
INIT_2F => X"FF49003AFEFEBFBEAA001C2EA8A821C2EAAA001C2EA8A00F7800017DA2842FA0",
INIT_30 => X"BEF082E95545000000000000000000000000000000000000000000000497BFAF",
INIT_31 => X"8A10AAD568A00555168A10002E9754D082E820BA08556AA00AAAABFE00F7AEAA",
INIT_32 => X"401E7082EAAABA5D5140010F7AE974105D7BC21555D51575EFFFAA97555A2AEA",
INIT_33 => X"BEABFFAAFBEABFFF7AA80145557BFDF55F78017400F780001FFAA84000AAFFD1",
INIT_34 => X"7BD5555AAD57DF55AAAEBDFEF007BE8A10AAAE8215DA2FFE8ABA082ABFE00AAF",
INIT_35 => X"7FBC00BA55557DFF75D2E82010F7843DF45FFD540000000402145AA843FFFF00",
INIT_36 => X"F780021FFA2803DE10FFD16ABFF5D7BFDE10AAAA975FF5D7BC21EFF7FBD7400F",
INIT_37 => X"0000000000007FE8BFF080028BFFAAFFEAA105D2EAAA005D2AAAA185D2AAAA10",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000400000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(1),               -- Port A write enable input
DIA(0)   => data_write_a(8),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(8),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(1),               -- Port B write enable input
DIB(0)   => data_write_b(8),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(8),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_9_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000B0001800002840002C0000281800000030000000033022000000000002",
INIT_01 => X"8000098218302849180060000C004240413C0A61590001D90213C90008510200",
INIT_02 => X"000008700CB089100002061031200074810448800104008048080080001210E2",
INIT_03 => X"000200140C1822000A028010408100000628000140402080041A100040024840",
INIT_04 => X"41040000000400080002040200080800040000000B08D1055842080604600700",
INIT_05 => X"10002024000020102400010000026104200004000400800C8B0024E4E0010C40",
INIT_06 => X"8000440802280002700800008A840004A0610000C0000810000C590103600810",
INIT_07 => X"538600220028001890240980A80800200102025000000BF08200002440000883",
INIT_08 => X"00000402C220104131102101040810028528820005100003900E884000010007",
INIT_09 => X"00000005E000000600BCA284140200800C834948100004590111824404012080",
INIT_0A => X"04080000901012100A1141005922000245410002008880000032005080000800",
INIT_0B => X"2000020040044010440104401004010440100401044010040104400802008208",
INIT_0C => X"D1A1344420D2E100000808000000000481000000202002400006800825908402",
INIT_0D => X"0500000000109000000000000580008000080000C852240100068D0B4685A342",
INIT_0E => X"0500000A00000000000000000000028000408020000000050000208020000000",
INIT_0F => X"0000304002100020000000000000000900208004000000050000208004000000",
INIT_10 => X"0000000001200000000A00000000000000000000050000480008000000000000",
INIT_11 => X"009F0080000000004807C0200000000012000020000081000000040000000000",
INIT_12 => X"00000048F8000400000002403E0004000000009067E000000000000000000900",
INIT_13 => X"0000000000000000140000CEE001000000000000000A000036AC008000000000",
INIT_14 => X"03210000000400CA81000000619480D4000400000000000000004100000036E8",
INIT_15 => X"A368DA368DA3685A1685A1685A121A11A1419001512490040024001000008019",
INIT_16 => X"1685A1685A1685A1685A1685A368DA368DA368DA368DA368DA368DA368DA368D",
INIT_17 => X"685A1685A168DA368DA368DA368DA368DA368DA368DA3685A1685A1685A1685A",
INIT_18 => X"CCF48DE68A895C38E250080000000000000000000000685A1685A1685A1685A1",
INIT_19 => X"514514514514514514514514514D34D34D34D34D28E10040392482090157344C",
INIT_1A => X"4D268341A0D069349A0D069349A0D068341A0D068341A0D06834514514514514",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000001654D0D069349A0D068341A4D268341A",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"BE8B45002A974AAAA803DFFFAA843DF45FFFFEAABA0000000000000000000000",
INIT_22 => X"AEBDE00AAFBEAABA080000000087BEAA10F7803DE00FFAEBFFFF0800155FFAAF",
INIT_23 => X"AAEA8ABAAAFBFDE0055556AA005D0415555087BFDE00A2FBD7400F7FBFDFFFA2",
INIT_24 => X"005155555557BE8BEF007FFDEAAAAD1555EF0055401FFF7AEAAA10F780155EFA",
INIT_25 => X"0F7AA974AA082E80010A2AAAAA10552AA8AAA557FC0010F780154105D7FC2145",
INIT_26 => X"BA087BFDF45F7AA974AAAAAA97555F784174BAF7D5555FFF780154AA5D2AA8A1",
INIT_27 => X"F45F7FFFFF55AA80155FF080400145FFFBEAABAF7D17FEBAA2AEBDF45002EAAA",
INIT_28 => X"0000000000000000000000000000000000000000AAFFE8A00552EBFE00F7D17F",
INIT_29 => X"BAFFF080A175D7BEF1E8B6D002090482B68E38FC7BE8A3DF7DF7F5E8A9200000",
INIT_2A => X"BD0400FFF5FDFC7B6A0BDE38B6F5E8A92080E000280071E8A00EB8E3FE10F7AE",
INIT_2B => X"AAA8A38FF8E175C7A2AAAAA82A2F1FAE105D556AA10410E175550871FFE00A2F",
INIT_2C => X"F8A17400557FC015514555757D5D71E8BEF147BFAE82A2DB555C71C5B451D7FF",
INIT_2D => X"FF84174BA5D20AAA00E3AA904BA142A87010A2AEADA38492EA8AAA5571C2000F",
INIT_2E => X"AAAA0BFF7D0024ADA921C7BFFF55FFA095482B6A49256DEB84104BAFFD1525FF",
INIT_2F => X"38492ABDE10EBDF7AF6DE3FFF8F7DB68A105D7000400155FFFBEDA82FFD57DEB",
INIT_30 => X"FEFF7D16AA00000000000000000000000000000000000000000000000A2FBE8A",
INIT_31 => X"AA00AAAABFE00F7AEAABEF082E95545F7D568BEF080402000F7AAA8B55FFAABD",
INIT_32 => X"9754D00517DE00A2FFC2000F7D17FF55FF803FEAAFFD16AA00082E820BA08556",
INIT_33 => X"FD55555D7FD5555FFAAA8AAAFFAA97555A2AEA8A10AAD568A00555168A10002E",
INIT_34 => X"2EAAABA5D5140010F7AE974105D7BC21555D51575EF555568BEF5D7FE8A10AAF",
INIT_35 => X"A84000AAFFD1401E7FF80174AA5D0028A00AAAE800AA552A97400A2AEBDEAA08",
INIT_36 => X"F7FBFFE00FFD17FEAAA2803DFEF08043FE00557BFDF55F78017400F780001FFA",
INIT_37 => X"0000000000A2FFE8ABA082ABFE00AAFBEABFFAAFBEABFFF7AA80145080002145",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000800000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(1),               -- Port A write enable input
DIA(0)   => data_write_a(9),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(9),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(1),               -- Port B write enable input
DIB(0)   => data_write_b(9),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(9),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_10_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000B0001800002840002C0000281800020030000000033022000000180006",
INIT_01 => X"000008000000004C002000000010026840000000080000080200000000110200",
INIT_02 => X"0000004000800110000006100000003000040800010400004808000000120060",
INIT_03 => X"000200000810020000020000400100000600000000400000001A000040004800",
INIT_04 => X"0004000000000008000200020000000004000000080010004000000200000000",
INIT_05 => X"1000202000011010000000000000010520000400000080000000200000200004",
INIT_06 => X"80004408022800023000000088040004A061000040000810000C490103600000",
INIT_07 => X"120420020028000890240980A808002001020050000009F08000002440000082",
INIT_08 => X"00000402C0201051311001000000020201080200440400000000800000000000",
INIT_09 => X"0000105808000000000000000000008000008088100004590111800004000000",
INIT_0A => X"00804000801210440003C1411008800045000002000014000040009002800000",
INIT_0B => X"0400200000000000000004000040000000000000040000400000000000000221",
INIT_0C => X"0100802000000000000002802000000400100000000002000026000840011400",
INIT_0D => X"0500000000409002082010400400008000400008002044082000081004080204",
INIT_0E => X"0500000200000000000000000000028000400000000000050000200000000000",
INIT_0F => X"0000304002000000000000000000000900200000000000050000200000000000",
INIT_10 => X"0000000001200000000200000000000000000000050000400000000000000000",
INIT_11 => X"0082000000000000480080000000000012000101000080000000000000000000",
INIT_12 => X"0000004810000000000002400400000000000090400000000000000000000940",
INIT_13 => X"0000000000000000150000C00000000000000000000A40001400000000000000",
INIT_14 => X"02000000002400C2810000006000000000000000000000000000410040001400",
INIT_15 => X"020080200802008020080200800800220200840001309A08A848001000008000",
INIT_16 => X"0000000000000000000000000200802008020080200802008020080200802008",
INIT_17 => X"0080200802000000000000000000000000000000000000000000000000000000",
INIT_18 => X"940FE0D397124355520542821010000000000000000000802008020080200802",
INIT_19 => X"28A28A28A28A28A28A28A28A28A28A28A28A28A29554199854514514F546890A",
INIT_1A => X"32994CA6532995CAE572B94CA6532994CA6532994CA6532994CA28A28A28A28A",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000001867172B94CA6532994CA6572B95CAE5",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FC2155F7D155545AA80001EFAAFBEAB45557FFDE100000000000000000000000",
INIT_22 => X"FBE8BFFF78402155AAFBE8B45002A974AAAA803DFFFAA843DF45FFFFEAABA007",
INIT_23 => X"87BEAA10F7803DE00FFAEBFFFF0800155FF00042AB55FFD168B55AA8000010FF",
INIT_24 => X"AAFBEAABAA2FFD741055003DFEFF7AA801FFAAD16AABA002ABDE100800000000",
INIT_25 => X"FF7FBC0145F78028A00A2D142155087BFDE00A2FBD7400F7FBFDFFFA2AEBDE00",
INIT_26 => X"BAF780155EFAAAEA8ABAAAFBFDE0055556AA005D0415555007FD74105555555E",
INIT_27 => X"5EF0055401FFF7AEAAA105D042ABFF5D556AB55AAD168ABA002A975FFF7AEBDE",
INIT_28 => X"0000000000000000000000000000000000000000557BE8BEF007FFDEAAAAD155",
INIT_29 => X"3DF7DF7F5E8A92007BC217DEBDB55555AA8E071D7AAFBEFB455D71F8E0000000",
INIT_2A => X"B6DB55BE8E05000EBFFE8BC7E38E07145BEF1E8B6D002090482B68E38FC7BE8A",
INIT_2B => X"2EB8E00080E000280071E8A00EB8E3FE10F7AEBAFFF080A175D700042AB7DEBD",
INIT_2C => X"FF5FDFC7B6A0BDE38B6F5E8A92B6FBD5410490A3DFD7F7A4821D7A2D16FA8214",
INIT_2D => X"0071D54104951555D7EBF5C5155E3842AA00BED1421450871FFE00A2FBD0400F",
INIT_2E => X"20820955EFE3AEBDEAAFF8E175C7A2AAAAA82A2F1FAE105D556AA10410E17555",
INIT_2F => X"EF147BFAE82A2DB555C71C5B451D7FFAAA8A38410E2ABD749516FB55BED16FA8",
INIT_30 => X"F455D556AA000000000000000000000000000000000000000000000005D71E8B",
INIT_31 => X"2000F7AAA8B55FFAABDFEFF7D16AA00087FC01EFA2FFD7545AAAE97555A2FBFD",
INIT_32 => X"9554500042ABFFA2FFFFF45F7AE97400AAFFE8B45AAAA95545F7D568BEF08040",
INIT_33 => X"400155A2D57FE00552EA8A00082E820BA08556AA00AAAABFE00F7AEAABEF082E",
INIT_34 => X"517DE00A2FFC2000F7D17FF55FF803FEAAFFD16AA00FFFBD5400082EBFF45F78",
INIT_35 => X"55168A10002E9754D085155410085557555AAD557555A2802AA10FFD54214500",
INIT_36 => X"08557DF55F7D17FE000804155FFAAAABDEAAFFAA97555A2AEA8A10AAD568A005",
INIT_37 => X"0000000000555568BEF5D7FE8A10AAFFD55555D7FD5555FFAAA8AAA002AAAB45",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000008FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(1),               -- Port A write enable input
DIA(0)   => data_write_a(10),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(10),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(1),               -- Port B write enable input
DIB(0)   => data_write_b(10),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(10),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_11_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10180B05A0010402840602C2D001019000000300000000330A20080EC180002",
INIT_01 => X"AB400986B830284D1820E0000C3642484000000008000008820009080A512220",
INIT_02 => X"102A68440080011000000618062AD03502640800010410424908136019920868",
INIT_03 => X"004A0846191B22120642000442C110044600000101E9225CDC9A10844A9A4842",
INIT_04 => X"0094024000250808800216021138000B848000000800100040000102A0600200",
INIT_05 => X"7E4024242008A8102CA88A44010401042200444000888000000028000002A002",
INIT_06 => X"8088445712280000B18812288E0400253855200045C86810000C5B0503286A28",
INIT_07 => X"10008822A028004880200A80880208200122006C000015F0C20408264902C840",
INIT_08 => X"9390040280241041D1754100000018108728820024002B3A01A89540080824C8",
INIT_09 => X"A1001C41A1348498B080801010000080D00301081000045B0511D28D94012339",
INIT_0A => X"44080000901012428003414158230CBA4576708241C010908040341322008000",
INIT_0B => X"040464D280144050C72A0872A0C72A0872A0C72A0C72A0872A0C595043950421",
INIT_0C => X"0804001400000820110A42822204880CD81040442900021704E6000800001D54",
INIT_0D => X"80C62D0500409002082010404580018000404012004004192C10000000000000",
INIT_0E => X"80C62D5803161C526DB40506C120A806ABB0D808CC334A80A54B70D408CC32D2",
INIT_0F => X"2B5144D0DD903C54916D15458C0513005570D408CC334A80A54B70D808CC32D2",
INIT_10 => X"52148C4DB05621E363F813961C20EDA944016558C2347A080B10D8DD6422AA10",
INIT_11 => X"1880144D3345C65593800319C18BD1ECA1C9010112566F10AC4183C340DAE02D",
INIT_12 => X"5810503000633830DE3C2C9C00289A66AA8DE50E0800360614AC281430890600",
INIT_13 => X"0CD2A9CEA8199B6B082B55900314140365320485C4F00AD544407241C175C402",
INIT_14 => X"0000074044C4801832701A89D20A38093631425969020855A281844E00540404",
INIT_15 => X"0000000000000000000000000020C00200088101513492101280401000400200",
INIT_16 => X"2008020080200802008020080000000000000000000000000000000000000000",
INIT_17 => X"0080200802008020080200802008020080200802008020080200802008020080",
INIT_18 => X"804180C0B10A4210420140028400000000000000000000802008020080200802",
INIT_19 => X"000000000000000000000000000820820820820801C414947000000055062608",
INIT_1A => X"0000000004020000000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000001F87E000000000000010080000000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"ABDF5508557DF45002ABDFFFF7803DE10AA80000AA0000000000000000000000",
INIT_22 => X"FFE8A10A28000000007FC2155F7D155545AA80001EFAAFBEAB45557FFDE10082",
INIT_23 => X"02A974AAAA803DFFFAA843DF45FFFFEAABAA2AEBFF45FFAEBFEAA002A801FFF7",
INIT_24 => X"F78402155AAD155555A28428BFF002ABDE00A2AABFE10082ABFFEFAAFBE8B450",
INIT_25 => X"0002A80010A2842AAAA007BFFF4500042AB55FFD168B55AA8000010FFFBE8BFF",
INIT_26 => X"00080000000087BEAA10F7803DE00FFAEBFFFF0800155FF00557FF45557FC201",
INIT_27 => X"1FFAAD16AABA002ABDE10A2D168A10A284021FF5D00154BAF7FBE8BEFFFD5400",
INIT_28 => X"0000000000000000000000000000000000000000A2FFD741055003DFEFF7AA80",
INIT_29 => X"EFB455D71F8E00002EBDF6D005B78F7D142ABDFC7F78E3FE28B684070AA00000",
INIT_2A => X"0BDEAA1C2A801C7E3FFEFA10B68407038007BC217DEBDB55555AA8E071D7AAFB",
INIT_2B => X"20B8FEFBEF1E8B6D002090482B68E38FC7BE8A3DF7DF7F5E8A92BEAEBFF7DEBA",
INIT_2C => X"E8E05000EBFFE8BC7E38E07145B6D15756DA28A28BFF082ABAE10B6AAB8E2808",
INIT_2D => X"08517DF7D497BC5028142A87000A28A2AA92007FF8F7D00042AB7DEBDB6DB55B",
INIT_2E => X"2FFFFEFBC7E3DF42028080E000280071E8A00EB8E3FE10F7AEBAFFF080A175D7",
INIT_2F => X"10490A3DFD7F7A4821D7A2D16FA82142EB8E00B6DB6AA28A280001FF5D0A1048",
INIT_30 => X"EAAF784154BA000000000000000000000000000000000000000000000B6FBD54",
INIT_31 => X"7545AAAE97555A2FBFDF455D556AA00082EBFFEF007BE8BFF5D2ABDF55F7AABD",
INIT_32 => X"6AA00FFAEBFFEFAA803DEBA5D2E82155A2FBFDE00FF84154BA087FC01EFA2FFD",
INIT_33 => X"AAAA00FFAAA8AAA080028BFFF7D568BEF080402000F7AAA8B55FFAABDFEFF7D1",
INIT_34 => X"042ABFFA2FFFFF45F7AE97400AAFFE8B45AAAA95545F7D5555FFAAAAA8BFF002",
INIT_35 => X"7AEAABEF082E9554508557DFFF007BD54BA5D2E95400A2AEA8A00007FEABFF00",
INIT_36 => X"AA80001FF5D2E82000F7FFFFF45AAFFC20BA082E820BA08556AA00AAAABFE00F",
INIT_37 => X"0000000000FFFBD5400082EBFF45F78400155A2D57FE00552EA8A00FFFFE8AAA",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000800000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(1),               -- Port A write enable input
DIA(0)   => data_write_a(11),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(11),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(1),               -- Port B write enable input
DIB(0)   => data_write_b(11),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(11),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_12_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A500C4B01BC0268A6940312C0DE045196A831A300500032B333287E4FC812006",
INIT_01 => X"AF400D869830E84D5823E0000C1742484000000008000008820009280A553235",
INIT_02 => X"502A7144008001100000171C022BD13412762A000586235ECC09C8423B960866",
INIT_03 => X"31863846191BA218064204000281200406A10843010022DEDF0852944A9C014A",
INIT_04 => X"0014030000250409000014821038080B840000400800102040000302F0600233",
INIT_05 => X"7FC034348008A8102CA88F48010601042400048000188000000938000002E088",
INIT_06 => X"9CC96CC6F63A5001F12B56A0AC8601F47AC06400D1F80C10020C493F03343A38",
INIT_07 => X"1020002030280098A12048908A16BA311177124C000003F08A94282E5C262861",
INIT_08 => X"827A0602902A10491165E10000049010C52882008600A73A01E8974008092CF8",
INIT_09 => X"47000001A1248008F000000000000080000F010C100204593F11A6CDF48023BF",
INIT_0A => X"040000208010120ACA01400058010CBA4D277C86CCE802B380003C1360008000",
INIT_0B => X"011C46D3C7BC1EF083AF0C3AF083AF083AF0C3AF083AF083AF0C1D7861D78400",
INIT_0C => X"08040014C9001AE91D17E50AD79FEFC87C2154745F82131FFCCE00080000095E",
INIT_0D => X"807BF7118180984004000803D40001880001001400C005031010000000000000",
INIT_0E => X"807BF76A109C944B5891BF06C5EEB14FCBF0D90076D61C807BF7D0D80876D49C",
INIT_0F => X"6DE38EB9FB10350C00A99F7CA80757365E50D80876D61C807BF7D0D90076D49C",
INIT_10 => X"841BCC69A0D8C6F7F0AA001C943A65756A0976EB5A7E7FC8951018186334F311",
INIT_11 => X"D5A014481991C6A737D80211912970CDCDD1864116D6C7080651CB4661F33615",
INIT_12 => X"349E929300423224AE19B9BEC0289033238D4E6EA805892946A9B011A7B152CF",
INIT_13 => X"6244CD7AC01CAAA56B3E6D9001068715D64006D2A961CF9B44512A2504532182",
INIT_14 => X"00000439FDC25C58067A9FAB46095A0B5289A0282D2E1444ACB12A17CF9B4414",
INIT_15 => X"0000000000000000000000040026C00000288401513492909280401000F70A00",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"088881360A95090CB05442029010000000000000000000000000000000000000",
INIT_19 => X"1041041041041041041041041049249249249249200100002D4514510051B946",
INIT_1A => X"592C964B2592C964B2592C964B2592C86432190C86432190C864104104104104",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000002007F592C964B2592C964B2592C964B2",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"43FE0008557DFFF0800020105D557FEAA00557DE100000000000000000000000",
INIT_22 => X"557DFFFF7AA80000082ABDF5508557DF45002ABDFFFF7803DE10AA80000AAAA8",
INIT_23 => X"7D155545AA80001EFAAFBEAB45557FFDE10AAD5420000051555FFA2AA8200000",
INIT_24 => X"A28000000A2D155410F7FFFFEBA08003FE00082AA8AAAAAFFC00BA007FC2155F",
INIT_25 => X"0A2AABFE1055516ABEF5D517DEAAA2AEBFF45FFAEBFEAA002A801FFF7FFE8A10",
INIT_26 => X"55AAFBE8B45002A974AAAA803DFFFAA843DF45FFFFEAABA000028A105D2ABFE1",
INIT_27 => X"E00A2AABFE10082ABFFEF085542000000417555002A820AA08557DFFFF7AA821",
INIT_28 => X"0000000000000000000000000000000000000000AAD155555A28428BFF002ABD",
INIT_29 => X"3FE28B684070AABE803AE38145B78FD7000005010495B7AE921C517DE1000000",
INIT_2A => X"B505FFB6A487000005F7AFD7F7A482038002EBDF6D005B78F7D142ABDFC7F78E",
INIT_2B => X"F5C2082007BC217DEBDB55555AA8E071D7AAFBEFB455D71F8E00BED547038145",
INIT_2C => X"C2A801C7E3FFEFA10B68407038B6D550428FFF1FDE821C003FE001C2EAAAAAB6",
INIT_2D => X"00002FA285D20BDE28A2A4B8E10555B68BEF5D517DEAABEAEBFF7DEBA0BDEAA1",
INIT_2E => X"2005F7DFD7F7A482155BEF1E8B6D002090482B68E38FC7BE8A3DF7DF7F5E8A92",
INIT_2F => X"6DA28A28BFF082ABAE10B6AAB8E280820B8FEF085F4703814001055514208208",
INIT_30 => X"A0055517DE00000000000000000000000000000000000000000000000B6D1575",
INIT_31 => X"8BFF5D2ABDF55F7AABDEAAF784154BAF7802AABA5D7FEAB45080015410007FEA",
INIT_32 => X"6AA00F7D1554BA5D7BC01FFFF8015410007FEAB45F780020BA082EBFFEF007BE",
INIT_33 => X"43FE10552EAAAAAFFD140000087FC01EFA2FFD7545AAAE97555A2FBFDF455D55",
INIT_34 => X"AEBFFEFAA803DEBA5D2E82155A2FBFDE00FF84154BAF7D1400BAFFD57FE005D0",
INIT_35 => X"FAABDFEFF7D16AA0008003FEBA55003DEBAA28428A105D7FEABEF55557DEBAFF",
INIT_36 => X"550402145550000010087FFFF45F78402145F7D568BEF080402000F7AAA8B55F",
INIT_37 => X"0000000000F7D5555FFAAAAA8BFF002AAAA00FFAAA8AAA080028BFF087BD54AA",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000000FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(1),               -- Port A write enable input
DIA(0)   => data_write_a(12),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(12),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(1),               -- Port B write enable input
DIB(0)   => data_write_b(12),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(12),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_13_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10110A0441812402840402822007818000E00700000000330A3000000008042",
INIT_01 => X"A1400984B830C848180260000C0042604001000008220008A200100802110200",
INIT_02 => X"10A00860009141100000C6180C285035000E0800010431004908135980120C60",
INIT_03 => X"004E20441910221B06420C85D5013804060000000040324C441A108468024842",
INIT_04 => X"0184034010250089C00EA8021938325B04800002091090014880080200000900",
INIT_05 => X"18002424B008881024A8004E01040104270004E0000080090500604840000481",
INIT_06 => X"80004414022A2490B00A142C8C840005794540015E006810001C4B01032C7E20",
INIT_07 => X"510200028028004880280A808816002101022468000011F082040A264006C000",
INIT_08 => X"D2B00402B220104B531001000008001041080200B660E30B200C8040080A9206",
INIT_09 => X"A1000809A93484D21000000000000080C90391881000145B0111A30404015000",
INIT_0A => X"000000008010102A82014100101118BA4510008241480290882400900000A000",
INIT_0B => X"0284484000000000400000000040000000000000040000000000000020000000",
INIT_0C => X"A944AA2000A02000212800020000000D80004084A0000390002E001843210400",
INIT_0D => X"859C1881A04090000000000021800180010341179065441356150A1285094284",
INIT_0E => X"859C188810C65A72A617520252781EA02520D589B9A260859C1840DD81B9A0E0",
INIT_0F => X"0E71F1052D942748C19484E39442D15961C0DD81B9A260859C1840D589B9A0E0",
INIT_10 => X"E60605C0C12CBD400B0810C65A61AA459D0047398500D5889D26907356533C00",
INIT_11 => X"8F60CA1562094650CA28398A42C051E0332181010109294C8E1160CB8C80A561",
INIT_12 => X"2645056D073148580A3C065141942AC4128CA199180C5232575138094450AD0A",
INIT_13 => X"84CA93A2FC008962142B17301A9A1A5196A80245208E0AC5C853C8028163B8C0",
INIT_14 => X"0240034000E4DC8A84000014982372011FC1E475F0F0084A3961F5A80AC5C816",
INIT_15 => X"4250942509425094250942509428D421420882020120981812C8403000088212",
INIT_16 => X"2509425094250942509425094250942509425094250942509425094250942509",
INIT_17 => X"5094250942509425094250942509425094250942509425094250942509425094",
INIT_18 => X"FF3F7DF7FF3E9F7DF7E24502A800000000000000000050942509425094250942",
INIT_19 => X"EBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBF7DFDFDDD555555F7EFBBEE",
INIT_1A => X"7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAEBAEBAEBAEBA",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000000007F7EBF5FAFD7EBF5FAFD7EBF5FAFD",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5554BA087FFFF55557BD54AAF7FBC01FFA2802ABEF0000000000000000000000",
INIT_22 => X"2E80155AA802AB45AA843FE0008557DFFF0800020105D557FEAA00557DE10AAD",
INIT_23 => X"8557DF45002ABDFFFF7803DE10AA80000AA087BD75EF087FFFFEF557BEAB4555",
INIT_24 => X"F7AA80000AAD1420AA087BD7555FFD168AAAFFAE820AA5D5557555082ABDF550",
INIT_25 => X"5FFD157555085140010F7AEAABFFAAD5420000051555FFA2AA8200000557DFFF",
INIT_26 => X"45007FC2155F7D155545AA80001EFAAFBEAB45557FFDE10AAAEA8BFFA2FBD754",
INIT_27 => X"E00082AA8AAAAAFFC00BA00002AAAAF7D5574BA557BE8A10A284154BAFFAAAAB",
INIT_28 => X"0000000000000000000000000000000000000000A2D155410F7FFFFEBA08003F",
INIT_29 => X"7AE921C517DE10A2DB50482147FFAF554971D0492E3F1C71C7BE8A2ABD700000",
INIT_2A => X"FFAFD7497BE8B5555208217DBE8A2AB45BE803AE38145B78FD7000005010495B",
INIT_2B => X"5F5056D002EBDF6D005B78F7D142ABDFC7F78E3FE28B684070AA1C71D25D7007",
INIT_2C => X"6A487000005F7AFD7F7A482038AADF47092147FD257DFFD568A82FFA4870BA55",
INIT_2D => X"A2A0ADBC7A2FFD257DE3DF52555085142000FFAAAFBFFBED547038145B505FFB",
INIT_2E => X"0B680124BAFFAAAFB45007BC217DEBDB55555AA8E071D7AAFBEFB455D71F8E00",
INIT_2F => X"28FFF1FDE821C003FE001C2EAAAAAB6F5C20821C002AA92FFDF574824171EAA1",
INIT_30 => X"545F7AEA8B55000000000000000000000000000000000000000000000B6D5504",
INIT_31 => X"AB45080015410007FEAA0055517DE00A2FFC00105D7BE8B55085142010AAD157",
INIT_32 => X"154BA5D5140145007BE8B55087BEAB555D04001EFF7AAA8B55F7802AABA5D7FE",
INIT_33 => X"16AA10FF80174AA557FC21EF082EBFFEF007BE8BFF5D2ABDF55F7AABDEAAF784",
INIT_34 => X"D1554BA5D7BC01FFFF8015410007FEAB45F780020BAA2FFD54105D7FC21EFFFD",
INIT_35 => X"2FBFDF455D556AA00A2803FF45AAFFC21EFAAFBC0155085540000FFAEBFFEFF7",
INIT_36 => X"F7FBD5410085568A10FF80020AAFFAABFF55087FC01EFA2FFD7545AAAE97555A",
INIT_37 => X"0000000000F7D1400BAFFD57FE005D043FE10552EAAAAAFFD1400005D042AA00",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000CFFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(1),               -- Port A write enable input
DIA(0)   => data_write_a(13),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(13),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(1),               -- Port B write enable input
DIB(0)   => data_write_b(13),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(13),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_14_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10020A000180000284008280000281800000030000000033022000000580002",
INIT_01 => X"A140098018300848184860000C20C24040000000084000084200000000110200",
INIT_02 => X"1020006000900110000006102028503400040800010400204908012018120E64",
INIT_03 => X"000200441910221006420000400100040600000000E9E401209A108448004842",
INIT_04 => X"0004020000250008000200021038000804000000090090004800080200000000",
INIT_05 => X"500024240008881024A800400104010420000400000080080100204040000000",
INIT_06 => X"8000440102282015B10A10288E0400042345400040006810000C5901033D7880",
INIT_07 => X"1100000200280048802008828812002001220064000005F1C2850A2649204070",
INIT_08 => X"00B00402802010411110010000080010010802000400230B000C804008080002",
INIT_09 => X"01000009A92480001000000000000080C8038188100004590111B68404010000",
INIT_0A => X"0000000080101000000141001001088A45000082400000008020009000008000",
INIT_0B => X"0004404000000000400004000000000000004000000000000004000000000000",
INIT_0C => X"8904A0200080200001080002000000088000400420000200002E000841010400",
INIT_0D => X"0500000C80409000000000000000018000000000806044010014081204090204",
INIT_0E => X"0500005813A0210D072E8D012001028402908004000587050000108004000707",
INIT_0F => X"9004300044900812386A280E5800088980108020000587050000108020000707",
INIT_10 => X"DE00482E19E30002007813A02096038AE200880405200308828062A68C0BC700",
INIT_11 => X"00000E5A08E6000048001292B83280001208A1011004011060049A1C59192055",
INIT_12 => X"492060480256530650000240001DB011CC00009000032C4C979E3806180C0900",
INIT_13 => X"5A3433EDE00154181400000007BCBD858F120120541A0000000033757465B2C0",
INIT_14 => X"02002C000024008A84001A0902000422E3E99681004802115652594000000001",
INIT_15 => X"0240902409024090240902409028D021020880000120901812C8401000000210",
INIT_16 => X"2409024090240902409024090240902409024090240902409024090240902409",
INIT_17 => X"4090240902409024090240902409024090240902409024090240902409024090",
INIT_18 => X"5C8FF0F7BE9D5F7DF65040028000000000000000000040902409024090240902",
INIT_19 => X"79E79E79E79E79E79E79E79E79E79E79E79E79E7BF7DDDDDFCF3CF3DF5579B4E",
INIT_1A => X"3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE79E79E79E79E",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000003FF803F9FCFE7F3F9FCFE7F3F9FCFE7F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"BE8B55A2AE80000F7D5555555D2AAAABAAAD1420BA0000000000000000000000",
INIT_22 => X"00155EF0804155EFAAD5554BA087FFFF55557BD54AAF7FBC01FFA2802ABEFA2F",
INIT_23 => X"8557DFFF0800020105D557FEAA00557DE10A2AA801FFA28402000AAAE9554555",
INIT_24 => X"AA802AB4500516AA00A2AE800BAFFFFC20BAF7AEA8B45080417400AA843FE000",
INIT_25 => X"0A2843FEBAFFFBD7410A2D168BFF087BD75EF087FFFFEF557BEAB45552E80155",
INIT_26 => X"AA082ABDF5508557DF45002ABDFFFF7803DE10AA80000AA005568ABAA2840201",
INIT_27 => X"AAAFFAE820AA5D5557555002E80155A280000005D7FFDF4555517DFEF00043FE",
INIT_28 => X"0000000000000000000000000000000000000000AAD1420AA087BD7555FFD168",
INIT_29 => X"C71C7BE8A2ABD7A2FFEDB55B6A080038E3DB50555412AA8ABAAADB4009200000",
INIT_2A => X"402038AAAA955554900105FF0800175D7A2DB50482147FFAF554971D0492E3F1",
INIT_2B => X"0A12410BE803AE38145B78FD7000005010495B7AE921C517DE10A2AE851FFB68",
INIT_2C => X"97BE8B5555208217DBE8A2AB451C556FA00A2A0800BAE3F1C0092EBAAADB6D08",
INIT_2D => X"00516DABAA28402038B6803DE82F7F5D5410A2D568BC71C71D25D7007FFAFD74",
INIT_2E => X"55D5F78FD7000E3FEAA002EBDF6D005B78F7D142ABDFC7F78E3FE28B684070AA",
INIT_2F => X"92147FD257DFFD568A82FFA4870BA555F5056D002A80155B680000105D7FF8F4",
INIT_30 => X"AAAAAFFC2000000000000000000000000000000000000000000000000AADF470",
INIT_31 => X"8B55085142010AAD157545F7AEA8B55A2FBFFF55FF84000AAAAFBC0145002AA8",
INIT_32 => X"7DE00A2AA955FFFF80020BAAAAA975450800001EF080417555A2FFC00105D7BE",
INIT_33 => X"140000A2AEBFFEF082A82010F7802AABA5D7FEAB45080015410007FEAA005551",
INIT_34 => X"5140145007BE8B55087BEAB555D04001EFF7AAA8B555D557FE00A280020BAAAD",
INIT_35 => X"7AABDEAAF784154BA08557FEAAA284000AAFF803DE00FFD557400AAD56AB455D",
INIT_36 => X"F780020105D7BEAB45557BE8B45082EBFEBA082EBFFEF007BE8BFF5D2ABDF55F",
INIT_37 => X"0000000000A2FFD54105D7FC21EFFFD16AA10FF80174AA557FC21EF082A80145",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000000FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(1),               -- Port A write enable input
DIA(0)   => data_write_a(14),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(14),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(1),               -- Port B write enable input
DIB(0)   => data_write_b(14),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(14),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_15_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000A000000000284000280000001800020030000000033022000000180002",
INIT_01 => X"A140098018300848180060000C00424040000000080000080200000000110200",
INIT_02 => X"102100400C8011100000061000A8503401044880010430004808000180122378",
INIT_03 => X"000200541D102210064200000045000546080000400020000008108448400042",
INIT_04 => X"8094020000254C880000028A1018000844000000880013504000002600000000",
INIT_05 => X"10002424000AA81024A82040010C61062001440002988000000024808001004B",
INIT_06 => X"80004400022A00003C8912248E0400042854400040006810000C4901032B1800",
INIT_07 => X"50200000B0280048A0280A828801002101020040000005F38204082640000000",
INIT_08 => X"01F00402802610411100110000000010010802000400230A0008884008080004",
INIT_09 => X"01000001A12481041000000000000080C0030108100004590111820404000000",
INIT_0A => X"0000000080101000004140001001088A45000082000000008000001080008000",
INIT_0B => X"0004404000000000400004000040000400000000000000000004000020000200",
INIT_0C => X"0804000020024100012808020000000981004004A0200310000C000800000000",
INIT_0D => X"0000001180009000000000002100018000000000004004010010000000000000",
INIT_0E => X"00000008000002000000000000000000000080A40000000000000080A4000000",
INIT_0F => X"00000000001000204800000000000000000080A40000000000000080A4000000",
INIT_10 => X"000000000000000000080000020000000000000000000008000C020000000000",
INIT_11 => X"000000824000000000000020220000000001800100020300000004003420480A",
INIT_12 => X"0000000000040440000000000001048000000000000000100800400000000000",
INIT_13 => X"000800000000000000000000000100C220050000000000000000008220884400",
INIT_14 => X"000000000000000830000000000000000016101C5C1400000000000000000000",
INIT_15 => X"0000000000000000000000000020C00000088000012090101280401000000200",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000040028000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"000010082A954BA00003DFEF085155400F78428BEF0000000000000000000000",
INIT_22 => X"8015400FF84001EFA2FBE8B55A2AE80000F7D5555555D2AAAABAAAD1420BAFF8",
INIT_23 => X"87FFFF55557BD54AAF7FBC01FFA2802ABEFF7AE95555A2FBE8BEFA2843DE00AA",
INIT_24 => X"0804155EFFFFBE8BFF0800174AA557BFDE10A2FBEAB45F7D56AABAAAD5554BA0",
INIT_25 => X"5FFD568BEF087FE8A1055003FE00A2AA801FFA28402000AAAE955455500155EF",
INIT_26 => X"45AA843FE0008557DFFF0800020105D557FEAA00557DE10F7D1574AAA2D16AB5",
INIT_27 => X"0BAF7AEA8B45080417400FFFFC2145080015400AA802AA00AAAE800BA5D00155",
INIT_28 => X"000000000000000000000000000000000000000000516AA00A2AE800BAFFFFC2",
INIT_29 => X"A8ABAAADB40092E38E070280024904AA1C0438FD7005150438F78A2DBFF00000",
INIT_2A => X"FE8BC7BE8E38E10A28017400E38A051FFA2FFEDB55B6A080038E3DB50555412A",
INIT_2B => X"D16AABAA2DB50482147FFAF554971D0492E3F1C71C7BE8A2ABD7E3AA9257DA2F",
INIT_2C => X"AAA955554900105FF0800175D7E3FFEFBD70000124AA557FFDE10A2FBEDB6DF7",
INIT_2D => X"FFDF50482A2DB6AB45FFD56DBD7087BEAA38410038E38A2AE851FFB68402038A",
INIT_2E => X"0AAA085082550A1057DBE803AE38145B78FD7000005010495B7AE921C517DE10",
INIT_2F => X"00A2A0800BAE3F1C0092EBAAADB6D080A12410FFF1C017D140410400BE8E28A1",
INIT_30 => X"0AAF7AEBDFEF0000000000000000000000000000000000000000000001C556FA",
INIT_31 => X"00AAAAFBC0145002AA8AAAAAFFC2000AAAA974AA0800020BA550028B55085540",
INIT_32 => X"A8B55AAAE821EFAAFBEAB55F7AAA8A00AA8417400AAAE975EFA2FBFFF55FF840",
INIT_33 => X"BFFE10A2FFFFFEFF7D568ABAA2FFC00105D7BE8B55085142010AAD157545F7AE",
INIT_34 => X"AA955FFFF80020BAAAAA975450800001EF080417555AAFFFDF450804020AA557",
INIT_35 => X"07FEAA0055517DE00FFFBC2000AAFBE8B55F7D17DF45007FE8AAA08002AAAAA2",
INIT_36 => X"5D0000010F7AAA8A10AA8017400552A801EFF7802AABA5D7FEAB450800154100",
INIT_37 => X"00000000005D557FE00A280020BAAAD140000A2AEBFFEF082A82010FFD5421EF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000C00000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(1),               -- Port A write enable input
DIA(0)   => data_write_a(15),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(15),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(1),               -- Port B write enable input
DIB(0)   => data_write_b(15),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(15),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_16_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"DA22C618B1000482B688B186588884862A400438255FC38381441205BA803003",
INIT_01 => X"264AC80028404C211203A952A90341080B173340412000E1005D628000820484",
INIT_02 => X"400034C206C405000001A48202084004003008255040826EE008B440200E2042",
INIT_03 => X"A459C1240181AB20AD27315B7F1983CA1C900040422A005762010010000C0400",
INIT_04 => X"296E542B6E3A825C15FB385321B4ADFE16AB45FD2C400002E205231201290A28",
INIT_05 => X"B9E5815006028179808C00A0D2152B90707A1E0BD423CAC0000D610000000710",
INIT_06 => X"81F104A1415C292164280081C6AB88742086ACACDE240000A80090CE82A803B9",
INIT_07 => X"400800000ACCAA280940580400A37B8896CA4D000A80C1102A00001C14028009",
INIT_08 => X"0015452880C8D90409A02D965965200100104F2B00822512000000231520A024",
INIT_09 => X"A5AA80018120E00066000000000012C9000A0000D0A80000BF8028E87C1B9927",
INIT_0A => X"00520228080108039501200848002912300208092B940192D1000000000000A8",
INIT_0B => X"03561180063DB4F6110001100011000110001100011000110001080008800080",
INIT_0C => X"080200854409418B02ED0000502A02972000040BB401100010012B4C90000100",
INIT_0D => X"6D061A1F8D60D80820500101244AA8A2AA242E80000009200120000000000000",
INIT_0E => X"6D066210E5001DB4A5B400C7D553847165A99000C6564CDD051DC99000C65555",
INIT_0F => X"21D0C48F254946148107354292673D1F72C99000C6564CDD0565C99000C65555",
INIT_10 => X"952D2058F33225787810F5001D6121A9559224D1FF97D0272F04D89441A56D8A",
INIT_11 => X"6C1C74485B81E31306C71D1093AB8A64811BADC00992180D58033B1172F2A025",
INIT_12 => X"7B86DED8E3A212748F0E0CA638E890B7A8546120C0AFF5B548AC431FB1C7DB07",
INIT_13 => X"EFCE9B26DECA1AD36A2E4F40DF6AAAF260AF88899E8B8B93D12A877178DD0032",
INIT_14 => X"A8009F8B108C80A1021B9A8BB8056662CA1951596800FC01A38D4D4B072B922F",
INIT_15 => X"00000000000000000000000000044000102A0001148442A1108103595580A840",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"4C690DA64C1C4F68A36040000000000000000000000000000000000000000000",
INIT_19 => X"D14D14D14D14D14D14D14D14D14514514514514529E5F87869E79E78558D1154",
INIT_1A => X"3D1E8F47A7D3E9F4FA7D3E9F4FA7D3E9F47A7D1E9F47A7D1E9F4D14D14D14D14",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE000000000000000007D3E9F4FA7D3E8F47A3D1E8F47A",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFEFF7D168B55AAD17FFFF552EBFE00007FC00AA0000000000000000000000",
INIT_22 => X"04000BA552A821FFFF8000010082A954BA00003DFEF085155400F78428BEF087",
INIT_23 => X"2AE80000F7D5555555D2AAAABAAAD1420BA5D2E975EFF7D568BFFFF80175EF00",
INIT_24 => X"FF84001EF0000020AA5D00154005D043FF45555540000082EAABFFA2FBE8B55A",
INIT_25 => X"0087FD74BAAAAEBFFEF557FC00AAF7AE95555A2FBE8BEFA2843DE00AA8015400",
INIT_26 => X"FFAAD5554BA087FFFF55557BD54AAF7FBC01FFA2802ABEF557BEABEF5D041541",
INIT_27 => X"E10A2FBEAB45F7D56AABA082A97545F7D16ABFFFFAABFEAAFF84001FF002A821",
INIT_28 => X"0000000000000000000000000000000000000000FFFBE8BFF0800174AA557BFD",
INIT_29 => X"50438F78A2DBFF0871F8FC7E3D56AB6DBEDB7FFEF552AB8E38087FC209200000",
INIT_2A => X"16ABFFE38E175EF1400000BA412E871FFE38E070280024904AA1C0438FD70051",
INIT_2B => X"2EAFBD7A2FFEDB55B6A080038E3DB50555412AA8ABAAADB400924920925EFF7D",
INIT_2C => X"E8E38E10A28017400E38A051FF0804050BA410A1240055003FF6D5551420101C",
INIT_2D => X"4975EDBC7550E12410087FD74AAB6AABFFC7557FC00BAE3AA9257DA2FFE8BC7B",
INIT_2E => X"AF780051C70824851D7A2DB50482147FFAF554971D0492E3F1C71C7BE8A2ABD7",
INIT_2F => X"D70000124AA557FFDE10A2FBEDB6DF7D16AABA08249756DF7D168BC7F7AABAEA",
INIT_30 => X"AAA007BC0000000000000000000000000000000000000000000000000E3FFEFB",
INIT_31 => X"20BA550028B550855400AAF7AEBDFEF08516AB55A2D16ABEFFFFBFDFFF552AAA",
INIT_32 => X"C20000000021EFF7D568BFFA2AA955FF5D04020AA002A955EFAAAA974AA08000",
INIT_33 => X"03DFEF5D51420005D2ABFF45A2FBFFF55FF84000AAAAFBC0145002AA8AAAAAFF",
INIT_34 => X"AE821EFAAFBEAB55F7AAA8A00AA8417400AAAE975EF0800174BA002E820105D0",
INIT_35 => X"AD157545F7AEA8B5500557DF45552A82000007BD74AAF7AEBDF455D7BC20BAAA",
INIT_36 => X"F7D568B55FFAAAAABAFF8415545000015555A2FFC00105D7BE8B55085142010A",
INIT_37 => X"0000000000AAFFFDF450804020AA557BFFE10A2FFFFFEFF7D568ABA0804155FF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000400000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(2),               -- Port A write enable input
DIA(0)   => data_write_a(16),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(16),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(2),               -- Port B write enable input
DIB(0)   => data_write_b(16),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(16),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_17_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"5284CE4FB7BD2C8994A13392DBD02E14006B82AC7E800D44D3DD2FD5F9B961C0",
INIT_01 => X"F9BA301F7E03FC6793F2199B39FC233C11D93AE6F3BB92B32091DBC339B24542",
INIT_02 => X"1D5FC0C08F040404446965C0607FB8A217C400C33A908078551BD04222186338",
INIT_03 => X"8504930A37F65820CB24111B7F08014A0AB84A52B6D2AFF97C1B5AC757F06D6B",
INIT_04 => X"250834336D1E81500FDB38302292ADFE103B6DBD204037F202042075E2B1D00A",
INIT_05 => X"8F039786062C6CE092F5FE005236781C402A0807B4070670083DC68206D7E6D0",
INIT_06 => X"0CD26803C3582408962C58B183F8AEF42045919B30E085DD2ED57D4EED08CA6A",
INIT_07 => X"700000B30380670B8142500448E3E01E94EF1340A28AC1AC8156044D1400AA00",
INIT_08 => X"009F3A1B0120A1C51DFFC40C30E5F0182D0950190C0810BE00E9A76E4C6FFBE4",
INIT_09 => X"8FCCC200A59BDD2FFE3F3EC7C7DEF207000F00059D2ED56D7EED2ED3C9A867DC",
INIT_0A => X"0617112E46F05D02DD814102F800633F1D0A7CC9AE7A08BFF0001D35682AC0CE",
INIT_0B => X"8A3F06ABD73DBCF4FBCF4FBCF4FBCF4FBCF4FBCF4FBCF4FBCF4FBE7A7DE7A780",
INIT_0C => X"001000974F08518F5AFFC94B533FADA7FDE97D6BFF329E1B50FF99F086000D9E",
INIT_0D => X"F50B018F95EA3DED1652EC0B27E67F419E2E1E8000C0036340B8000000000000",
INIT_0E => X"F50B01C8DF7F96197DB4AFC8C8886AF672A1537F759299F50B03C1537F759199",
INIT_0F => X"6068331C5103E7EF0FBEED6BB6A9412007C1537F759299F50B03C1537F759199",
INIT_10 => X"21F2CD7F252CDABB3CE8CF7F963AB9FD6AD434201AA68B837FFD1F7B7125B68C",
INIT_11 => X"BD055EB6D555CB2949C15BA7270FF256526BBFD55BBE71D79F73C7AC6DB9BF37",
INIT_12 => X"94080BF82B74E4E1FE4ACA4E0ABD6DAAAB965293036FF6B652A99A6026027FBE",
INIT_13 => X"EF5CBA7A43482800FEFAFD06B8CFCCAB7550D0C2022EAEBD438697AD2EBA9168",
INIT_14 => X"AC00A8BBFC8B501CF7A0FED9A548FA19752C4A4EADAE42FCBC38C3B7BEBF42CF",
INIT_15 => X"0000000000000000000000000026E100002F382DBD9ECFE117805F20CFDAAB00",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"09EDCC4052E917114F981800C000000000000000000000000000000000000000",
INIT_19 => X"EBA69AEBA69A69AEBA69AEBA69A69A69A69A69A68698686981D75D7443720030",
INIT_1A => X"46A351A8D068341A0D068341A0D068341A0D46A341A0D46A341A69AEBA69A69A",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000000000046A351A8D46A351A8D46A351A8D",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFEFF7FBEAB450804001EFAAD57FEAA0000000000000000000000",
INIT_22 => X"51401EF087FD74AA087FFFFEFF7D168B55AAD17FFFF552EBFE00007FC00AA087",
INIT_23 => X"82A954BA00003DFEF085155400F78428BEFAAD168A000004020AA5D7BE8B4500",
INIT_24 => X"552A821FF5D00020BA552A82000552A821555D7FEAB55FF80175EFFF80000100",
INIT_25 => X"FAAFBC01EF5D0015555557BFDEBA5D2E975EFF7D568BFFFF80175EF0004000BA",
INIT_26 => X"BAA2FBE8B55A2AE80000F7D5555555D2AAAABAAAD1420BAFFFFFDF45AAD17FFF",
INIT_27 => X"F45555540000082EAABFF00516AA10552E820BA007FEABEF005555555A2D1554",
INIT_28 => X"00000000000000000000000000000000000000000000020AA5D00154005D043F",
INIT_29 => X"B8E38087FC2092147FFFFFFFFFBFDFC7EBF5E8B550000071EFB6DF7AE9200000",
INIT_2A => X"A07082497FEFB6D1451471EF007BD04920871F8FC7E3D56AB6DBEDB7FFEF552A",
INIT_2B => X"8E175FFE38E070280024904AA1C0438FD7005150438F78A2DBFFBED16AA381C0",
INIT_2C => X"38E175EF1400000BA412E871FF550A00092492A850105D2A80155417BEFB6DEB",
INIT_2D => X"FFF5FFF6DAADF7FFD7B6F1C71EF55001756D5D7BFAEBA4920925EFF7D16ABFFE",
INIT_2E => X"700515556DA2DF50492A2FFEDB55B6A080038E3DB50555412AA8ABAAADB40092",
INIT_2F => X"BA410A1240055003FF6D5551420101C2EAFBD7145B6AA28492487082007FEDBD",
INIT_30 => X"5EFFFFBEAA000000000000000000000000000000000000000000000000804050",
INIT_31 => X"ABEFFFFBFDFFF552AAAAAA007BC0000557FFDFEFF7FBFFF55A2D16AB55000017",
INIT_32 => X"BDFEFF7D568AAA5D2A97410007BFFFFF5551555EF087FC200008516AB55A2D16",
INIT_33 => X"A82155087FFFFEFAAAA975EFAAAA974AA0800020BA550028B550855400AAF7AE",
INIT_34 => X"00021EFF7D568BFFA2AA955FF5D04020AA002A955EF5D2E80010002A954005D2",
INIT_35 => X"02AA8AAAAAFFC2000FFD57DFFFAAFFFDF55FFD1575FF5504175EF5D7FEAAAA00",
INIT_36 => X"000415410007BFFF450051555EFA2FBC0000A2FBFFF55FF84000AAAAFBC01450",
INIT_37 => X"00000000000800174BA002E820105D003DFEF5D51420005D2ABFF45557FE8AAA",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000CFFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(2),               -- Port A write enable input
DIA(0)   => data_write_a(17),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(17),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(2),               -- Port B write enable input
DIB(0)   => data_write_b(17),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(17),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_18_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"69844019080000A21A611406840014122A641074155FC28A2024001001801003",
INIT_01 => X"01067920034004180005E9E3C90360C0041C0181002001602025800008440084",
INIT_02 => X"40AC3CAA22D605200000856E2481902400344A20F802C22054001000021E2379",
INIT_03 => X"A54C23B34C81EB2076471000800981140C010101750D1007E58040102B0E0100",
INIT_04 => X"22660C1C0065003C04040013236E105016A028402D618803EB092B9201490B2A",
INIT_05 => X"B8E080000000005889AC41E04508A99070200E010001C1CA11803850C8000100",
INIT_06 => X"800A4CE301545001F40050216C09950004C2047BCF1C8090C02800C0120886B3",
INIT_07 => X"814A0080064C1F300020080182001A9E02C03400082002700000217294007101",
INIT_08 => X"000117088080990419002D86184A01018030430700802541420440022030041A",
INIT_09 => X"7030C30B885200D274004008080003C32A10A19090C02010E102294406168800",
INIT_0A => X"00602A01880980037109700C04C44C92A88DCC2211E44174112840880000060D",
INIT_0B => X"11C0D95C20C2030A003080030800308003080030800308003080018400184004",
INIT_0C => X"8304E02809832E6021002020404042000F00008400811824AD4007ECD9436261",
INIT_0D => X"0AFCE5D22A82B20000520100C801F8A07E103000A1285C84000418360C1B060D",
INIT_0E => X"0AFCFD8CB17E5B4F045557575E6EFBE3942C1040A41D660AFCE1CC1040A41E66",
INIT_0F => X"8E7FFBB385661C08D1455ABA91E6FF5FDFCC1040A41D660AFCF9CC1040A41E66",
INIT_10 => X"015F82C006C3AF31E64CB17E5A9655017F1FC73FAF1D61B1040294C58AD1FF5F",
INIT_11 => X"B95454005BAA36DCF8E519001BF80DEB3EE2020EA678189C6EC32881F7F75648",
INIT_12 => X"67D7EDFCA320037E81BD77D728A800B7546DBDFF12904747A351145FC53ABF8D",
INIT_13 => X"92B764225C57C97EBE76E1254F0C0D4514A84F5573FE9DBA4A38E247C522CC0E",
INIT_14 => X"BE84370001B6922070440556B15F7FABBC40151D7C747D8220673C3B9DB84B20",
INIT_15 => X"06C1B06C1B06C1B06C1B06C1B0491069068000004060300A005A01183F240014",
INIT_16 => X"6C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B",
INIT_17 => X"C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B0",
INIT_18 => X"B80EE173C2300F7DF16000000000000000000000000041B06C1B06C1B06C1B06",
INIT_19 => X"AAAAAA28A28A28AAAAAAA28A28A28A28A28A28A2910591505C104104B28BBECE",
INIT_1A => X"128944A25128944A25128944A25128944A2552A954AA5128944AAAA28A28A28A",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000128944A25128944A25128944A25",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFDFEF5D2A974BA082E954000000000000000000000000",
INIT_22 => X"0028B55002E82000087FFFFFFFFFFFFFEFF7FBEAB450804001EFAAD57FEAA087",
INIT_23 => X"7D168B55AAD17FFFF552EBFE00007FC00AA087FFFFFFFFFBFDF45AAD568B5508",
INIT_24 => X"087FD74AAAAFFFDF45A2D16AB55F7FFFFFFF00043DE10AA843DE00087FFFFEFF",
INIT_25 => X"A55042ABEF5D7FD75FFAAD540145AAD168A000004020AA5D7BE8B450051401EF",
INIT_26 => X"45FF8000010082A954BA00003DFEF085155400F78428BEFAA80000000804154B",
INIT_27 => X"1555D7FEAB55FF80175EF5D00020105D2A97400082E95555085168A10557FD75",
INIT_28 => X"00000000000000000000000000000000000000005D00020BA552A82000552A82",
INIT_29 => X"071EFB6DF7AE921C7FFFFFFFFFFFFFFFF7FBFDFFF5D2A954AA082A9242800000",
INIT_2A => X"1FAF55A2DF6DB7D1C002AB7D002A82028147FFFFFFFFFBFDFC7EBF5E8B550000",
INIT_2B => X"8E38E280871F8FC7E3D56AB6DBEDB7FFEF552AB8E38087FC2092087FFDFC7E3F",
INIT_2C => X"97FEFB6D1451471EF007BD0492B6F1F8F55AADF6DB7DE3F5FAFC708003DE28B6",
INIT_2D => X"A28407038140410492550A2ABC7497BD25FFAADF4516DBED16AA381C0A070824",
INIT_2E => X"D1C516FA28417BD5545E38E070280024904AA1C0438FD7005150438F78A2DBFF",
INIT_2F => X"92492A850105D2A80155417BEFB6DEB8E175FF5D0E05000492097428002E9557",
INIT_30 => X"4AA082A820AA000000000000000000000000000000000000000000000550A000",
INIT_31 => X"FF55A2D16AB550000175EFFFFBEAA00557FFFFFFFFFFFDFEFF7FBFFFEF552E97",
INIT_32 => X"C0000087BFDF45AAD568B55AAFBFDFEF55042ABEF002A800AA557FFDFEFF7FBF",
INIT_33 => X"16AB4500043DEAAFFAEAAAAA08516AB55A2D16ABEFFFFBFDFFF552AAAAAA007B",
INIT_34 => X"D568AAA5D2A97410007BFFFFF5551555EF087FC2000FFD56AB45A2FFFDFFFAAD",
INIT_35 => X"855400AAF7AEBDFEFA280154BA550400000552AA8B45087FC01EFA2FFD55EFF7",
INIT_36 => X"0804154BA082A975EF5D517DEAA007BD5545AAAA974AA0800020BA550028B550",
INIT_37 => X"00000000005D2E80010002A954005D2A82155087FFFFEFAAAA975EF5D2E97400",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000400000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(2),               -- Port A write enable input
DIA(0)   => data_write_a(18),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(18),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(2),               -- Port B write enable input
DIB(0)   => data_write_b(18),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(18),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_19_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"042200000000000041088001001AA00000000000000000000000500802000003",
INIT_01 => X"074018000024000000000404000000000A22000800000800004A200000000001",
INIT_02 => X"0000048002C405000000000006A84000000000200893C246A20000000020031A",
INIT_03 => X"082A58E411004B2000071000000981000C000000002045000200000000000000",
INIT_04 => X"200604000000001C0400001320000000162000002C4000026201201200090800",
INIT_05 => X"1020800000000058840200204000099070200E010001C0400000000000000000",
INIT_06 => X"0012048037805421402850001402498820022802400480405008901100A00102",
INIT_07 => X"00000000020C0130481204919200010C82000000000006002A548902A0020109",
INIT_08 => X"0001150800009900000005861840000000004301000B000000000001C1C00000",
INIT_09 => X"001F00002024B20002000000000002C300000000405000103010204000000000",
INIT_0A => X"00000000000000000000000000000040002000044000000000000000000002F0",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000420003B00000000000000000040012C80000000",
INIT_0D => X"45001A03C0825A0D20800000000018A006001000000000000000000000000000",
INIT_0E => X"450002131E01A1F6EA0A0020211146E069C2ACC01AE80045001D82ACC01AE800",
INIT_0F => X"1188340C3E1CFAD27CC2E004481020892282ACC01AE80045000582ACC01AE800",
INIT_10 => X"DEA03228D810007019931E01A1E5BA02802008C06F029D4C7B76639CEC0A0020",
INIT_11 => X"428AA3592000000206C2A4DAC00000008113C246A181C03FE4662A84575768DF",
INIT_12 => X"08201090549B5800000000261546B24000000000C53807E7CC06618018C51210",
INIT_13 => X"13F6A185A0A0168128411ACB800C0E108A0720288C011046B5986247C5452291",
INIT_14 => X"0000C220010808C10D9A92A74CD7CF4A080031B1515B212143D841431046B58A",
INIT_15 => X"00000000000000000000000000000000000000000000000000000118030004E0",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"3F0C7010C660C744192000000000000000000000000000000000000000000000",
INIT_19 => X"1861861861869A61861861861861861861861861A8208C4C1534D34C07208BBA",
INIT_1A => X"0984C26130984C26130984C26130984D26930984C26130984C261861861869A6",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE000000000000000000984C26130984C26130984C2613",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF552A974AA0004174BA0000000000000000000000",
INIT_22 => X"2E974BAA2FFFFE10087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974BA082E95400F7F",
INIT_23 => X"FFFFFFEFF7FBEAB450804001EFAAD57FEAAF7FFFFFFFFFFFFFFFFF7FBFDFFF55",
INIT_24 => X"002E82000F7FFFFFFFFFFFFDFEFA2D568B550004001EFAAAEA8ABA087FFFFFFF",
INIT_25 => X"5AAD16ABEF5D2ABFF55080402010087FFFFFFFFFBFDF45AAD568B55080028B55",
INIT_26 => X"BA087FFFFEFF7D168B55AAD17FFFF552EBFE00007FC00AAF7FFFFFFFF7FBE8B5",
INIT_27 => X"FFF00043DE10AA843DE00557FFDFEFA2D16AB55A2FFFDFEF5D2EBFE00AAFFFFE",
INIT_28 => X"0000000000000000000000000000000000000000AAFFFDF45A2D16AB55F7FFFF",
INIT_29 => X"954AA082A92428E3FFFFFFFFFFFFFFFFFFFFFFFEF552A974AA0000104AA00000",
INIT_2A => X"FFDFEFF7F5FAFC7492A974AAB6F5F8E101C7FFFFFFFFFFFFFFFF7FBFDFFF5D2A",
INIT_2B => X"A4A8AAA147FFFFFFFFFBFDFC7EBF5E8B550000071EFB6DF7AE92EBFFFFFFFFFF",
INIT_2C => X"2DF6DB7D1C002AB7D002A82028FFFFFFFEFF7F1F8FD7AAD16AB450000001FFBE",
INIT_2D => X"F7FBF8FC7E3F5EAB45B6DF6FBEF5D2AB8F7D000000010087FFDFC7E3F1FAF55A",
INIT_2E => X"7412ABFE28B6F5F8E820871F8FC7E3D56AB6DBEDB7FFEF552AB8E38087FC2092",
INIT_2F => X"55AADF6DB7DE3F5FAFC708003DE28B68E38E284971F8FC7AAD56DB6DBEF5F8FD",
INIT_30 => X"4AA0004000AA000000000000000000000000000000000000000000000B6F1F8F",
INIT_31 => X"DFEFF7FBFFFEF552E974AA082A820AAA2FFFFFFFFFFFFFFFFFFFFFDFEF552E95",
INIT_32 => X"EAA00A2FFFFFFFF7FBFDFFFFFD568B55002A954AAF7D568A00557FFFFFFFFFFF",
INIT_33 => X"56AB450004001EFFF842AAAA557FFDFEFF7FBFFF55A2D16AB550000175EFFFFB",
INIT_34 => X"7BFDF45AAD568B55AAFBFDFEF55042ABEF002A800AAF7FBFDFEFF7D56AB45AAD",
INIT_35 => X"52AAAAAA007BC0000FFFBE8B55AAD168B55F7FFFFFFF552AA8BEF08040200008",
INIT_36 => X"A2D57FFFFF7D568B45002ABDEAAFFD16AA0008516AB55A2D16ABEFFFFBFDFFF5",
INIT_37 => X"0000000000FFD56AB45A2FFFDFFFAAD16AB4500043DEAAFFAEAAAAA08556AB55",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000800000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(2),               -- Port A write enable input
DIA(0)   => data_write_a(19),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(19),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(2),               -- Port B write enable input
DIB(0)   => data_write_b(19),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(19),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_20_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000003",
INIT_01 => X"A65FF80000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000048002CC070000000000000000000000002FF86100200000000220002362",
INIT_03 => X"0000000000080F6000977060009B87A03C000000000000000000000000000000",
INIT_04 => X"3F2EFC040388137C3E20C477600142019E6000003CC0000A6601601A000B0000",
INIT_05 => X"102F91D10802ABFB80000021C8010FB0F0F43E1FE867DFC04400390210000220",
INIT_06 => X"90492261000080003400000010008000004203FE400580000000803000200006",
INIT_07 => X"401000004FFDFF28C4300C0010200100004000002AA001F00000000014000000",
INIT_08 => X"0801F5780259FB00000007BEFBC010002008FF7F00000000010018A81000041C",
INIT_09 => X"00000000020000000000000000000ADF00000020000000800000802830011023",
INIT_0A => X"0000000000000200020000000000000000000000000000000200200290000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"08120000B9090A700000200000004000000400000080002000407FED80000000",
INIT_0D => X"000079804000F00000000000C01FF8A7FE003000000004008100000000000000",
INIT_0E => X"0000798201000000100000000135386000401000010000000079801000010000",
INIT_0F => X"0185C300020004000010000000000252C7801000010000000079801000010000",
INIT_10 => X"00000010C1F30F300002010000080000000000CD8A0000400400000010000000",
INIT_11 => X"008040000000000292C0080000000000A5604000000284000818505200080000",
INIT_12 => X"0015E1B00100000000001496008000000000052B000048080000000000FC3600",
INIT_13 => X"80000000000002BA280000800830300000000000B8B400000401881010000000",
INIT_14 => X"00000000020020020001000040283024E6FB8604020080000383383B00000400",
INIT_15 => X"000000000000000000000004010201001003020200000000000127DBFF004000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"038200010089120104D204002000000000000000000000000000000000000000",
INIT_19 => X"B2CB2CB2CB2CB2CB2CB2CB2CB2C30C30C30C30C306982121A1E79E79A0700030",
INIT_1A => X"432190C86432190C86432190C86432190C86432190C86432190CB2CB2CB2CB2C",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000432190C86432190C86432190C86",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA0804020100000000000000000000000",
INIT_22 => X"2E954AA000400000F7FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0004174BAFFF",
INIT_23 => X"FFFFFFFFFFFFFDFEF5D2A974BA082E95400007FFFFFFFFFFFFFFFFFFFFFFEF55",
INIT_24 => X"A2FFFFE10FFFFFFFFFFFFFFFFFFFFFBFDFFF5D2E954BA007FC00BA087FFFFFFF",
INIT_25 => X"FF7FBFFF550800020BAAAD56AAAAF7FFFFFFFFFFFFFFFFF7FBFDFFF552E974BA",
INIT_26 => X"10087FFFFFFFFFFFFFEFF7FBEAB450804001EFAAD57FEAA007FFFFFFFFFFFFFE",
INIT_27 => X"B550004001EFAAAEA8ABA5D7FFFFFFFFFFFDFEFF7D56AB450000021EFA2D57DE",
INIT_28 => X"0000000000000000000000000000000000000000F7FFFFFFFFFFFFDFEFA2D568",
INIT_29 => X"974AA0000104AAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA08000500000000",
INIT_2A => X"FFFFFFFFFBFDFEF5D2E974AA000A07000E3FFFFFFFFFFFFFFFFFFFFFFFEF552A",
INIT_2B => X"71C50BA1C7FFFFFFFFFFFFFFFF7FBFDFFF5D2A954AA082A92428087FFFFFFFFF",
INIT_2C => X"7F5FAFC7492A974AAB6F5F8E10E3FFFFFFFFFFFFFFEFF7FBFFFFF552E974AA00",
INIT_2D => X"1C7FFFFFFFFFBFDFEFE3F5F8F450004050AABEDF6FABAEBFFFFFFFFFFFFDFEFF",
INIT_2E => X"50804021FFB6D57DE28147FFFFFFFFFBFDFC7EBF5E8B550000071EFB6DF7AE92",
INIT_2F => X"EFF7F1F8FD7AAD16AB450000001FFBEA4A8AAA497FFFFFFF7FBF8FC7EBD168B4",
INIT_30 => X"4AA080017410000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFDFEF552E954AA0004000AAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A95",
INIT_32 => X"820AA087FFFFFFFFFFFFFEFF7FBFDFFF5D2A974AA002E95410A2FFFFFFFFFFFF",
INIT_33 => X"FFDFEF5D2E954AA0051554BA557FFFFFFFFFFFDFEFF7FBFFFEF552E974AA082A",
INIT_34 => X"FFFFFFFF7FBFDFFFFFD568B55002A954AAF7D568A00AAFFFFFFFFFFBFDFEFFFF",
INIT_35 => X"000175EFFFFBEAA005D7FFFFEFF7FBFDFFFAAD16AB450804174AAFFFFFFEBAA2",
INIT_36 => X"F7FFEAB45A2D568B550804001EFF7D57DEBA557FFDFEFF7FBFFF55A2D16AB550",
INIT_37 => X"0000000000F7FBFDFEFF7D56AB45AAD56AB450004001EFFF842AAAA087BFDFEF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000000FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(2),               -- Port A write enable input
DIA(0)   => data_write_a(20),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(20),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(2),               -- Port B write enable input
DIB(0)   => data_write_b(20),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(20),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_21_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"4A302428B824900A128C090A5C1800261500213C005FE812D10420054085A202",
INIT_01 => X"081FFE3440B609703B0427F801A40B8115BC4F655300340288A40D30040E4DD8",
INIT_02 => X"04CA478082CC1740002019824E0203100640303FF8C0B31061096E21A1840814",
INIT_03 => X"8C329E9204020FE002577800405B87047D5042129D8D0248903200013290C800",
INIT_04 => X"3E7FFE02482553FC3C020277E128080A1E6000003CC0000A6601E03A8B0F0008",
INIT_05 => X"F43F8140000203FFC806C8A1C1048FF0F0E07E1F00F7FFC00024010000468310",
INIT_06 => X"08710C10015E083D01A24404786BE0014114C3FE4187A009A663A680100B3096",
INIT_07 => X"200800008FDFFF00290000100211019812E210488228000000900260026C6058",
INIT_08 => X"0EF1F5FA0041FF080AC707FEFBC110008420F7FF388B70A20389346FE8000580",
INIT_09 => X"917FC30010107688862A28C54518DBFF00020004C0A6044901112A0908AA0A30",
INIT_0A => X"006309044081A001B188300E20806520398C6021569249C4B3007127080806FF",
INIT_0B => X"904595123203040D9228D9228D9228D9228D9228D9228D9228D99146C9146C84",
INIT_0C => X"88042090068008003120000806001402504110C48002403601887FEF80022A51",
INIT_0D => X"26C0AC404E43032CA0C205880A7FFAB7FE01409400400C0594A4002200110008",
INIT_0E => X"26C0AC086A170250454004C6012280129B034A080C0B0016A0D20346080C0A80",
INIT_0F => X"0B064092D85938C0112144050224120C500346080C0B0016A0D2034A080C0A80",
INIT_10 => X"40702E058355458967E86A170220D1800093414B0414782E4B5000D81480809A",
INIT_11 => X"081B1545104135443306C35901024F88A88049062A747512B76783C5D040E080",
INIT_12 => X"40160040D86B202049B22198362A8A208279854400A036801480031401900800",
INIT_13 => X"0DD001C002D38334000914028354008301008C0CF1480245108C7640A0604032",
INIT_14 => X"AC0496022300233104662848808E191526205018030060540284FA0C0044022C",
INIT_15 => X"004010040100401004010040102090010008000001C0E010020007DFFFC06E60",
INIT_16 => X"0401004010040100401004010040100401004010040100401004010040100401",
INIT_17 => X"4010040100401004010040100401004010040100401004010040100401004010",
INIT_18 => X"FF7FFDF7FF3E3DFDF7E000000000000000000000000040100401004010040100",
INIT_19 => X"FBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBFFDFDFFFCF3CF3FFFEF9FEE",
INIT_1A => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFEFF7FBFDFEFF7FBFDFEFBEFBEFBEFBE",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0004000100000000000000000000000",
INIT_22 => X"2A954BA0004154BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080402010FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF552A974AA0004174BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"000400000007FFFFFFFFFFFFFFFFFFFFFFEF552E974BA0804000AAF7FFFFFFFF",
INIT_25 => X"FFFFFFDFEF5D2E974BA002E97400007FFFFFFFFFFFFFFFFFFFFFFEF552E954AA",
INIT_26 => X"BA087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974BA082E95400007FFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2E954BA007FC00BA5D7FFFFFFFFFFFFFFFFFFBFDFEF5D2A954AA002E974",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFBFD",
INIT_29 => X"954AA080005000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA00000200000000",
INIT_2A => X"FFFFFFFFFFFFFFF552A974BA0000174AAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0A000AAE3FFFFFFFFFFFFFFFFFFFFFFFEF552A974AA0000104AAF7FFFFFFFFFF",
INIT_2C => X"FFBFDFEF5D2E974AA000A07000007FFFFFFFFFFFFFFFFFFFFDFEF552E954BA08",
INIT_2D => X"1C7FFFFFFFFFFFFFFFFFFBFDFEF5D2A974BA002A95400087FFFFFFFFFFFFFFFF",
INIT_2E => X"F552E974BA0020924BA1C7FFFFFFFFFFFFFFFF7FBFDFFF5D2A954AA082A92428",
INIT_2F => X"FFFFFFFFFEFF7FBFFFFF552E974AA0071C50BA557FFFFFFFFFFFFFFFF7FBFDFF",
INIT_30 => X"4BA000002000000000000000000000000000000000000000000000000E3FFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2A954AA080017410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"000AAF7FFFFFFFFFFFFFFFFFFFFFFFEF552A974BA0000174BAFFFFFFFFFFFFFF",
INIT_33 => X"BFDFEF5D2A954BA082E800AAA2FFFFFFFFFFFFFFFFFFFFFDFEF552E954AA0004",
INIT_34 => X"7FFFFFFFFFFFFFEFF7FBFDFFF5D2A974AA002E95410087FFFFFFFFFFFFFFFF7F",
INIT_35 => X"52E974AA082A820AA557FFFFFFFFFFFFFEFF7FBFFFFF552E954BA002E9741008",
INIT_36 => X"FFFBFDFEFF7FFFFFEF5D2A974BA0000020AA557FFFFFFFFFFFDFEFF7FBFFFEF5",
INIT_37 => X"0000000000AAFFFFFFFFFFBFDFEFFFFFFDFEF5D2E954AA0051554BA5D7FFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(2),               -- Port A write enable input
DIA(0)   => data_write_a(21),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(21),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(2),               -- Port B write enable input
DIB(0)   => data_write_b(21),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(21),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_22_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"5290F4CDE914905A14A43D33F488243E17122300F55FEB189B343A1140548380",
INIT_01 => X"A94007B259F6A975386262000C344BA9573C6FF57B18A5FB0ABFCD3C2C5F4F0C",
INIT_02 => X"D56B4302AC01005111011BD506AA5205274056900596A539584E2E6DFE4B2418",
INIT_03 => X"6B03F2F6151A2081F24001E8400008F401CB10C6594423C8923AD6B55AD0EB5A",
INIT_04 => X"8001023D37E50880436200808BC8492A0089249600101100008087248B64426E",
INIT_05 => X"A51035B41C0A88046CAEE8C23C08E040011C0020F8882001102D620A06D68301",
INIT_06 => X"B93FF975CF7889D085E997A2144E8FC2060B880081A26DCD4047EFF9EF018980",
INIT_07 => X"283800AA500200E8024AD03546A3262FB5AA5542A882040C7A64CBD64065F028",
INIT_08 => X"141008801018040E48D500400015805060040080A2A0F4A82381B4000A0905A0",
INIT_09 => X"4D0000002126F30C902A29C54539C020E11810098D4067EFF9FF284D483E2AB4",
INIT_0A => X"1400006100003202D040050220103D2A512C6A8C4F0008AA800470370000A000",
INIT_0B => X"013456520CA09281C2A81C2A81C2A81C2A81C2A81C2A81C2A81C9540E1540E00",
INIT_0C => X"A1402A13C0A10A893165281A1C2A7283516344C594A85536B1AD800214202C50",
INIT_0D => X"3C70FC20515808A0100820112300011000287B071105034406950A0285014280",
INIT_0E => X"3C70FC48E11CFC48400184CE0D6783139B0959A41606003C70FA0958AC160480",
INIT_0F => X"0D87E8B3B811B52048B10E0402AE1606D80958AC1606003C70FA0959A4160480",
INIT_10 => X"80F84E0185594581E088E11CFC38414020DD42CF909D7E0A551C02180300C0DD",
INIT_11 => X"441154C258012D86F3044A3133004A99BD8455300654458A1D588C4061403000",
INIT_12 => X"A096A240894626600953379822A984B0025B0DEC0345C9200680027181B44887",
INIT_13 => X"E2404160035482BE521C2C04A90783C18000D610B9D8070B12B1A2A62040202A",
INIT_14 => X"304244A91102C93A2D608D2A258DF8034284200C050070E40C80620C870B02C4",
INIT_15 => X"4411044110441104411044110466C440446CA06951D4EA801000980400646002",
INIT_16 => X"0100441104411044110441104411044110441104411044110441104411044110",
INIT_17 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_18 => X"FE8FF1F7DEBDDF7DF7D05122890000000003FFFFFFFF90040100401004010040",
INIT_19 => X"79E79E79E79E79E79E79E79E79E79E79E79E79E7BFFDFD7DDDF7DF7DF7DFBFDE",
INIT_1A => X"3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE79E79E79E79E",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE000000000000000003F9FCFE7F3F9FCFE7F3F9FCFE7F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0800000000000000000000000000000",
INIT_22 => X"2E974AA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000400010FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E954AA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"0004154BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA000015400FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF552A974AA0800154AAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA",
INIT_26 => X"BAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0004174BAFFFFFFFFFFFFFFFFF",
INIT_27 => X"FEF552E974BA0804000AAA2FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0000174",
INIT_28 => X"0000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040001000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E954AA000402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0417410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080005000FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF552A974BA0000174AAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA00",
INIT_2D => X"E3FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0804154BAF7FFFFFFFFFFFFFFFFF",
INIT_2E => X"F552E954BA000E124BAE3FFFFFFFFFFFFFFFFFFFFFFFEF552A974AA0000104AA",
INIT_2F => X"FFFFFFFFFFFFFFFFDFEF552E954BA080A000AAA2FFFFFFFFFFFFFFFFFFFFFFFE",
INIT_30 => X"4BA080400010000000000000000000000000000000000000000000000007FFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"17410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000400010FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF552A954BA000415400FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954AA0800",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFEF552A974BA0000174BAF7FFFFFFFFFFFFFFFFFFF",
INIT_35 => X"52E954AA0004000AAA2FFFFFFFFFFFFFFFFFFFFFDFEF552E974AA0804174AAF7",
INIT_36 => X"FFFFFFFFFFFFBFDFEF5D2E954BA002A820BAA2FFFFFFFFFFFFFFFFFFFFFDFEF5",
INIT_37 => X"0000000000087FFFFFFFFFFFFFFFF7FBFDFEF5D2A954BA082E800AAAAFFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000000FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(2),               -- Port A write enable input
DIA(0)   => data_write_a(22),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(22),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(2),               -- Port B write enable input
DIB(0)   => data_write_b(22),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(22),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_23_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"EF20906D902424807BC8241BC81801B97D38AD3C0800103362A6741C80A12A02",
INIT_01 => X"001FFF8409F089003B4422000D80C80106804A7951C5B9D1C828043EA28838F9",
INIT_02 => X"028406A002DC176444683862400003111001303FFC00F240D50146013B300500",
INIT_03 => X"001B243004080FE000177003145F87017D584B10D804034800200200A1008008",
INIT_04 => X"BEFFFC0248005FFC3C18A2FFE12222425E600000BDC0800AEE01E81A100F0A00",
INIT_05 => X"D03F8000000003FF810640A1C0008FF2F0E17E1F02FFFFC80100004044800080",
INIT_06 => X"800264B4854650040123428C204BF40F439647FF4807E189A477EF81DF0AF116",
INIT_07 => X"01000000FFDFFFE800401005C0A0008F86C60840AAAA100C68D1810C9F4A0020",
INIT_08 => X"1BE1F5F80003FF0002021FFEFBC80000000077FF184B03010004002FE1F29002",
INIT_09 => X"907FC308181204800600000000001BFFA800808189A657EF81DD0C00079CC800",
INIT_0A => X"0063090442A18001B188300C48907120AC810033149249C433200180082A06FF",
INIT_0B => X"9A41C1443243050C1010C1010C1010C1010C1010C1010C1010C1008608086084",
INIT_0C => X"000082A00600200080000500C000400800601200000254A000007FEFC1030221",
INIT_0D => X"0A9080400E0BF30C20CA858E087FFABFFE01409780214EE49620001000080004",
INIT_0E => X"0A908044294700701641005218521210150E5789F90A000A90800E5F81F90880",
INIT_0F => X"0E0220036864A7DCA190440301E2105C000E5F81F90A000A90800E5789F90880",
INIT_10 => X"C1400500C6CE5400032429470068924010164302048156305D66F8701681000E",
INIT_11 => X"2E0CCB0500013440600339C800004D8018000857A82920CE8CB220C81400A180",
INIT_12 => X"220344406739000009B0030019960A00026880C0422C52B01700044901488822",
INIT_13 => X"85C811A010428104128996465ADA020180804A040108A2658217C4008060300C",
INIT_14 => X"BE0692020328CA0028042054A92771C50FC070109000C1C819078280A265920E",
INIT_15 => X"020080200802008020080200800800200200000000000008004807DFFF000470",
INIT_16 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_17 => X"0080200802008020080200802008020080200802008020080200802008020080",
INIT_18 => X"0000000000000000000000000000000000000000000000802008020080200802",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000",
INIT_22 => X"2E974BA080002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E974BA000400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000400000FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF5D2E954AA080000010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA",
INIT_26 => X"10FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080402010FFFFFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2A954BA000015400FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA0804000",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E974BA080002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF5D2E954AA000402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA00",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080002010FFFFFFFFFFFFFFFFFFF",
INIT_2E => X"F5D2A954BA080407000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080005000",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF5D2A954BA000417410FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA080402000000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"02000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000010FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF5D2E974AA000402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0000",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000400010FFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"D2A954AA080017410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954AA080002000FF",
INIT_36 => X"FFFFFFFFFFFFFFFFFF552A954BA080015410FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_37 => X"0000000000F7FFFFFFFFFFFFFFFFFFFFFFFFF552A954BA000415400F7FFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000000FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(2),               -- Port A write enable input
DIA(0)   => data_write_a(23),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(23),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(2),               -- Port B write enable input
DIB(0)   => data_write_b(23),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(23),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_24_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100600007FFF000080108004000800020000840041000080808",
INIT_02 => X"0000068002CC07400000090C080002000000103FF811F150231000520ABE4404",
INIT_03 => X"8428180000080FE000177000001B87003D4000000E8B84010020000000008000",
INIT_04 => X"3E2FFC024800137C3C000077E00000001E6000003CC0000A6601E01A000F0200",
INIT_05 => X"103F8000000003FF80000021C0000FF0F0E03E1F0067FFC00000000000000000",
INIT_06 => X"00132412079001AD00810005E8000001401643FE4007E5501AA00000DC8C3006",
INIT_07 => X"000000000FDFFF62695A5685C094831D966000008002100C2040A178B600C240",
INIT_08 => X"08E1F5F80001FF00000007FEFBC00000000077FF000B00000000002FE0000000",
INIT_09 => X"107FC300000000000600000000001BFFA0000005501AA00000CE200000940000",
INIT_0A => X"00630104408180012188300C00814080008000010012414433000100080806FD",
INIT_0B => X"904181003003000C1000C1000C1000C1000C1000C1000C1000C1000608006084",
INIT_0C => X"00000080060000000000000012002C00000000000000000000007FEF80020201",
INIT_0D => X"440082404E0B332CA2C20188087FFAB7FE000082000000008220000000000000",
INIT_0E => X"4400824903210308074084210002460402009280010D80440084009280010F00",
INIT_0F => X"800A2400401A0C82183248060010280C20009280010D80440084009280010F00",
INIT_10 => X"C0A078160000404A0469032102981380202080026420020D06C002A08481C020",
INIT_11 => X"00164F400860000824059AD01802000208104817B00011306B2D9B0DD5082080",
INIT_12 => X"41021800B35A0300400041202C9E8010C0001040C5836CC01780018601030088",
INIT_13 => X"DB1011E000A140058220004AEFFC8101810021084301880030A8B77400603011",
INIT_14 => X"8C063C0220002201490418082010A57263E010000201033016085A40880030A1",
INIT_15 => X"000000000000000000000000000000000000000000000000000007DFFF0006E0",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"F6E7CC1132CDB444199000000000000000000000000000000000000000000000",
INIT_19 => X"79E79E79E79EFBEFBEFBEFBEFBEF9EF9EF9EF9EFA69861219575D75FF2D0AEEA",
INIT_1A => X"0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1EFBEFBEFBE79E",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE000000000000000000783C1E0F0783C1E0F0783C1E0F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020100000000000000000000000",
INIT_22 => X"2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"080002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_26 => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000400010FFFFFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2E974AA000400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0004000",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040201000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF5D2E974BA080002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFF",
INIT_2E => X"F5D2E974AA000400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF5D2E974AA000400000FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA080402010000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"00010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000010FFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002010FF",
INIT_36 => X"FFFFFFFFFFFFFFFFFF5D2E974AA000002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_37 => X"0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000402010FFFFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(3),               -- Port A write enable input
DIA(0)   => data_write_a(24),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(24),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(3),               -- Port B write enable input
DIB(0)   => data_write_b(24),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(24),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_25_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100200002000000080100004000000020000800041000080808",
INIT_02 => X"0000068002CC474000000800000002000000103FFCE302008000000880844A04",
INIT_03 => X"00000101C0200FF004177800081B87003D400000080000000020000000008000",
INIT_04 => X"3E2FFE024820137C3C004077F01000001E7249213CC1264A660DF05A000F9000",
INIT_05 => X"103F81C1002203FF80000021C1140FF8F0E03E1F0067FFE04800258280010052",
INIT_06 => X"80480AE20000000100000001C8608001401643FE4007C00000000000CC083006",
INIT_07 => X"280800000FDFFFEA4050140540B00100840000080002A00C2040810000000010",
INIT_08 => X"C8E1F5FA21C9FF80040007FEFBE031018C31F7FFBAEBC0020008086FE0000100",
INIT_09 => X"107FC301800000000600000000001BFFE00301000000000000CC020000140000",
INIT_0A => X"0077330C4889CC292588300C0080400000800001001243443B000100880806FD",
INIT_0B => X"904189003003000C1000C1000C1000C1000C1000C1000C1000C1000608006084",
INIT_0C => X"8B04228026824100000000000000000000000000000004A000007FEF80020201",
INIT_0D => X"400000400E03C30C20C2818C087FFAB7FE01409700C10007962418220C110608",
INIT_0E => X"4000000001010000004000000000400400001200000800400000001200000800",
INIT_0F => X"0008000000000480000040000000200000001200000800400000001200000800",
INIT_10 => X"0000001001000002000001010000100000000000202000000440000000800000",
INIT_11 => X"0000410000000008000008400000000200000806300400000820000020004880",
INIT_12 => X"0000080001080000000040000082000000001000000040800800000000020008",
INIT_13 => X"8100000000000000802000000840000200040000020008000000840000804000",
INIT_14 => X"8C04100200000200000610000000210000000018140000000008000008000000",
INIT_15 => X"04411044110441104411044510629041040D180400000010028047DFFF800C60",
INIT_16 => X"4411044110441104411044110441104411044110441104411044110441104411",
INIT_17 => X"4110441104411044110441104411044110441104411044110441104411044110",
INIT_18 => X"196A8C5A2932EC15DA080800002FFFFFFFFFFFFFFFFFC1104411044110441104",
INIT_19 => X"92492492492410410410410410410492410492412000531215A69A6BFBA2894A",
INIT_1A => X"B158AC562B158AC562B158AC562B1588C46231188C46231188C4924924924924",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000B158AC562B158AC562B158AC562",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000",
INIT_22 => X"2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF5D2E974BA080400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_26 => X"10FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0800000",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400000FFFFFFFFFFFFFFFFFFF",
INIT_2E => X"F5D2E974BA080000010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA080402000000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"02000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400000FF",
INIT_36 => X"FFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_37 => X"0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000000FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(3),               -- Port A write enable input
DIA(0)   => data_write_a(25),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(25),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(3),               -- Port B write enable input
DIB(0)   => data_write_b(25),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(25),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_26_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"E9264EAB20190CA3BA4997AA9002AE9C001006B0778015CFA17E0811039879C7",
INIT_01 => X"F1FFF9BB1F773C7F9BB07DFFFDD863FC5FFF3FEFFBBF9FFB22FFFBC7B9F30686",
INIT_02 => X"9B3184F8AFDEAF300029E4E300FC78A6258548EFFA71C00172082400003A2161",
INIT_03 => X"0213C3FDFFFC7F74FFBF737A603B87FEBE1A5294F65628A0001B9CE6CC606E73",
INIT_04 => X"7E2EFEBF6FFEB37C3FF3017776FFCDA43E7B6DFD7DEBFD8E6F5F78DF0BFBD644",
INIT_05 => X"902F87C74E8CCFFBB6FF70E1FE61FFBDF0FEBE1FFD67DFFEFFBDA7F7FED50870",
INIT_06 => X"213246200BCC8920360C1831CD7DF60A244B9BFEE00589DDBCEFEDC1DFA08957",
INIT_07 => X"B1D4223B4FFDFF21CC721C85DCE1458E8782484020A2C1FCA3468D77E0000300",
INIT_08 => X"2C05FD7BC471FBD13D980FBEFBEBF30B8D79FF7F451F33CFD60FE8FFFDF54003",
INIT_09 => X"19FFC71FEFED7B251E35768E8ED6BFDF3EB3EBF9DDBCE7FDC1DF8A760F3EACC0",
INIT_0A => X"56F7730ECCDBDF152199F51EDDCDEBCFF589807B7096CD4CF73AC1FC98884FFF",
INIT_0B => X"B867D3683A03A40F78C0D78C0D78C0D78C0D78C0D78C0D78C0D7A606BC606B8C",
INIT_0C => X"DFBFF5EB36DFE51FC3A80D73D840303983EE7F0EA03BDA680137FFFDFFD7E681",
INIT_0D => X"3F0080425E6BFF8DB0DAE19C09FFFFE7FE3EBEA8EB7AFEE5C9AEBD7F5EBFAF5F",
INIT_0E => X"3F00800DEC010280004000F808020290100FA2F60008003F00800FA2F6000800",
INIT_0F => X"00023002007BC0A14E00400003B8000D000FA2F60008003F00800FA2F6000800",
INIT_10 => X"01E0320007204008040DEC010300100000F600020581003F604D0700008000EE",
INIT_11 => X"201F21A2C40039006807C46426040E101A0259DFE82011A311AA042016040080",
INIT_12 => X"80020048F88C84C101C203403E434588007200D047F00090200007E0010009B0",
INIT_13 => X"0109000003E2000416C0804FE04140E80000F808010AB02033AC048A2A00003D",
INIT_14 => X"FFAFD082003B032FB987E04021D481D4000419060201E1A000044300B02033E8",
INIT_15 => X"AFEBFAFEBFAFEBFAFEBFAFEFFBFBFBFBBFCFBB0FFDFEFFEF2DFFFFFBFF802FFD",
INIT_16 => X"FEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBF",
INIT_17 => X"EBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFA",
INIT_18 => X"F491E166CC8553F86EDB5C88646FFFFFFFFFFFFFFFFFEBFAFEBFAFEBFAFEBFAF",
INIT_19 => X"1861861861861861861861861861869A69A61861AFBD54D5F871C71D475B15BC",
INIT_1A => X"0984C26130984C26130984C26130984C26130984C26130984C26186186186186",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE000000000000000000984C26130984C26130984C2613",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000",
INIT_22 => X"2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_26 => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFF",
INIT_2E => X"F5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA080402000000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"02010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_36 => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_37 => X"0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(3),               -- Port A write enable input
DIA(0)   => data_write_a(26),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(26),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(3),               -- Port B write enable input
DIB(0)   => data_write_b(26),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(26),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_27_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"00080A40000A41248002029000050A088000008242A0004404480002000A1155",
INIT_01 => X"F1FFF1C11F781C129C107DFFFE0860941E81258CA2B71C2220EC1B86E1A00002",
INIT_02 => X"183080988B2EAE00002BE001117C78C6848140CFFA0000800042008000011081",
INIT_03 => X"000003FDF3E47C74F7BCF36A203A47F6B8184210B6160820001318C60C204C63",
INIT_04 => X"7E28FEBF6FEEB3723F71017476DFC524397B6DF572EB6C8E175E70D90F539600",
INIT_05 => X"000F86064C8DDFE3B6FF50D1FC61DE39C8FCB91FF9671FE6B68984B5BCE40834",
INIT_06 => X"0000000800000042020C18300520620A80231BFE200181092CE7ED80DFC00147",
INIT_07 => X"8AC4AA3B0FD1FF201044110560884000840200520002080C23468D0300000282",
INIT_08 => X"2005F0784411E390A4880E3DF7E2FB0B8E717C7F411F3BC6D60B60FFDDE44001",
INIT_09 => X"18FFD757E7ED7A211E81C09818109E1F16B16B71092CE7ED81CF403601228C40",
INIT_0A => X"46FF730E5CCBCD55219AB55F0DEFABC7054880693016DD4C755AC16C1A884FFE",
INIT_0B => X"BC63F1683803C00E3440C3440C3440C3440C3440C3440C3440C3C2061A2061AD",
INIT_0C => X"56BF55CB165EC51D41880FA3F040202883B475062033186801137FF1BAD6F281",
INIT_0D => X"3B0000421E2B0F2E2AE215C808FFFA47FE62BAA86B1AB268E92AB56D5AB6AD5B",
INIT_0E => X"3B000025EC010080004000F808000098100F22520008003B00002F2252000800",
INIT_0F => X"00001042006BC0810600400003B80001002F22520008003B00002F2252000800",
INIT_10 => X"01E032000620000C0405EC010100100000F6000001C1003760410500008000EE",
INIT_11 => X"201D2120840039000817444404040E10020218DE282010A311AA002002040080",
INIT_12 => X"8000000AE888808101C20040BA4241080072001027F00080200007E0000001F0",
INIT_13 => X"0101000003E2000007C0800FE04040280000F8080002F02023AC04080A00003D",
INIT_14 => X"DDAFD082001B03249887E04001D481D4000009020201E1A000040100F02023E8",
INIT_15 => X"ADAB6ADAB6ADAB6ADAB6ADAB6BF1EBDABD8E270BF84A25C6ACB777E3FF800C6D",
INIT_16 => X"DAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6",
INIT_17 => X"AB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6A",
INIT_18 => X"100481CA860402104A471688747FFFFFFFFFFFFFFFFFAB6ADAB6ADAB6ADAB6AD",
INIT_19 => X"0000000000000000000000000008200000000000200072F210000001490E2168",
INIT_1A => X"A05028140A05028140A05028140A050080402010080402010080000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000A05028140A05028140A05028140",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000",
INIT_22 => X"2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_26 => X"10FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFF",
INIT_2E => X"F5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA080402000000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"02000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FF",
INIT_36 => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_37 => X"0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000000FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(3),               -- Port A write enable input
DIA(0)   => data_write_a(27),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(27),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(3),               -- Port B write enable input
DIB(0)   => data_write_b(27),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(27),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_28_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"02200AA400180030808802A900002A08001280A08A801044104A1000001818C3",
INIT_01 => X"50A00011460214428114180000882214413D0A71592A01D92213D28005210202",
INIT_02 => X"8A54800A210200111100C2110054289220810440030404010844000444410001",
INIT_03 => X"4200040822D4500001E0000028000002000211842010092000018C6295200631",
INIT_04 => X"00400000000B8000000140000005840C00000040002008808100048100100044",
INIT_05 => X"0000222200244400135110000135100000000000000000024CA0A01018000320",
INIT_06 => X"A004912008208040024489121144080400081000200008104000000020000041",
INIT_07 => X"A85800994000000A0200802004204420210001022AA8A0001122448142491008",
INIT_08 => X"0414000201800004080A000000124058200408000880004440004080160C4100",
INIT_09 => X"0080000206CB0821082B694D4D29400002002038104000000020003204000440",
INIT_0A => X"12000843066021001400040024440245400082D022040000400800081022C000",
INIT_0B => X"0002002C004001036050160501605016050160501605016050160280B0280B00",
INIT_0C => X"0012400810080414C0A800310840102182C62302A0194C08001680100E4040A0",
INIT_0D => X"05000002003004208208841401800040000A0000200814004198000400020001",
INIT_0E => X"0500000004000080000000000000028000002052000000050000002052000000",
INIT_0F => X"0000300000004001060000000000000900002052000000050000002052000000",
INIT_10 => X"0000000001200000000004000100000000000000050000002001050000000000",
INIT_11 => X"00002020840000004800040404040000120200A9000000010000002002040000",
INIT_12 => X"0000004800808081000002400040410800000090001000002000000000000910",
INIT_13 => X"0001000000000000144000010000402800000000000A1000010000080A000000",
INIT_14 => X"0080000000110006B08140000040000000000902000000000000410010000100",
INIT_15 => X"0080200802008020080200802101210810C39A66A90A85420413A82000000204",
INIT_16 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_17 => X"8020080200802008020080200802008020080200802008020080200802008020",
INIT_18 => X"110A00246972BD89A40A0C22E100000000000000000000200802008020080200",
INIT_19 => X"82082082082082082082082082082082082082080D35050758C30C31DE21102C",
INIT_1A => X"B0582C160B0582C160B0582C160B0580C06030180C06030180C0820820820820",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000B0582C160B0582C160B0582C160",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000",
INIT_22 => X"2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_26 => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFF",
INIT_2E => X"F5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA080402000000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"02000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_36 => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_37 => X"0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000000FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(3),               -- Port A write enable input
DIA(0)   => data_write_a(28),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(28),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(3),               -- Port B write enable input
DIB(0)   => data_write_b(28),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(28),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_29_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"79964E4BA01DACAB9E659792D00AAE160002829C7FDFEFCEE97C2815039D70C3",
INIT_01 => X"50BFF9AB0775343F9AB01DF80D5821FC0FFF3FEFD1AF9FF1207FFBC7B9720586",
INIT_02 => X"0D15846807D207200021C4E200D428A2018408600271C000720A0000003A2161",
INIT_03 => X"0002C009EEFC5F10F9B70178681B80FA3E000100765029A00019084345606421",
INIT_04 => X"3E6E023D27DA937C03E3407712E5CDA41E0924DC3D20B98AE905189F0BF8C000",
INIT_05 => X"902003C30E0447F877F930203E213F8CF01E3E00FC67C03A4D9C87525E510160",
INIT_06 => X"0012460003CC002036040811D919F402244293FEE00400CCB46BA4C164A08857",
INIT_07 => X"914800110FFC0001CC320C81D841418E82800100000041FCA1428575A0001108",
INIT_08 => X"0805FD0180E1F8C1111A0782082B50080508FF00048B124D4005C8AFF4154102",
INIT_09 => X"0180000ABFEF89250815568A8AD6ABC02A02A0B0CCB463B4C0748A720B1EA4C0",
INIT_0A => X"021410028450530014014002D445624DB481806A62840800C22800B8900042FF",
INIT_0B => X"0806522C0A40A50268D0068D0068D0068D0068D0068D0068D006A68034680300",
INIT_0C => X"8912E0A83289641F42A80561D040203182AC3D0AA0118A080036FFFC4F4164A0",
INIT_0D => X"050080424069F5A51250648801BFFFE0003E3E00A0685A85410C0816040B0205",
INIT_0E => X"050080080400028000000000000202900000A0F600000005008000A0F6000000",
INIT_0F => X"00023000001040214E0000000000000D0000A0F600000005008000A0F6000000",
INIT_10 => X"000000000120400800080400030000000000000205800008200D070000000000",
INIT_11 => X"000220A2C400000068008424260400001A0241DAC80001010000042016040000",
INIT_12 => X"00020048108484C10000034004414588000000D04010001020000000010009B0",
INIT_13 => X"000900000000000416C00041000140E800000000010AB0001100008A2A000000",
INIT_14 => X"A282C0000033010FB181E00020400000000419060000000000004300B0001100",
INIT_15 => X"02C0B02C0B02C0B02C0B02C4B12B312912831A27FCFE7FFB175B6FF800802594",
INIT_16 => X"2C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B",
INIT_17 => X"C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B0",
INIT_18 => X"EE7FFDF7FE783FFDFFEA0C00602FFFFFFFFFFFFFFFFFC0B02C0B02C0B02C0B02",
INIT_19 => X"BEFBEFBEFBEFBEFBEFBEFBEFBEEBAEBAEBAEBAEBBFFDF9FBEFFFFFFEBBCF9F96",
INIT_1A => X"FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFBEFBEFBEFBEF",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000FBFDFEFF7FBFDFEFF7FBFDFEFF7",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000",
INIT_22 => X"2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_26 => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFF",
INIT_2E => X"F5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA080402000000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"02000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_36 => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_37 => X"0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(3),               -- Port A write enable input
DIA(0)   => data_write_a(29),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(29),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(3),               -- Port B write enable input
DIB(0)   => data_write_b(29),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(29),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_30_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"FF9FE1F7FFBFFFFDFFD000000000000000000000000000000000000000000000",
INIT_19 => X"79E79E79E79E79E79E79E79E79E79E79E79E79E7AFBD75F5FDF7DF7FF7FFBFFE",
INIT_1A => X"3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE79E79E79E79E",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE000000000000000003F9FCFE7F3F9FCFE7F3F9FCFE7F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000",
INIT_22 => X"2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_26 => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFF",
INIT_2E => X"F5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA080402000000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"02000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_36 => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_37 => X"0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(3),               -- Port A write enable input
DIA(0)   => data_write_a(30),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(30),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(3),               -- Port B write enable input
DIB(0)   => data_write_b(30),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(30),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_31_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"129000008004A00804A40000400800020000000C005FEA005800200400050100",
INIT_01 => X"A15FF18019700810180065FFFC0040801E80258CA2951C2200EC0906A0804140",
INIT_02 => X"146000808A0C060444692000402850040400408FF80000000010000000004000",
INIT_03 => X"000003F5D1202C70F654716A001A07F438184210960600000012108518004842",
INIT_04 => X"3E28FE3F6FE513703F70007472DA4128187B6DB530C1240A060C70580B439200",
INIT_05 => X"000F84040C088BE3E4AE40C1FD04CE38C0FC381FF8671FE01009048084C40010",
INIT_06 => X"0000000000000008000810200420620E00030BFE000181092CE7ED80DF800106",
INIT_07 => X"000000220FD1FF200040100540800000840200408002000C2244890200000200",
INIT_08 => X"0011F0780011E38004800E3CF3E0B1118C31747F000B33820209206FC9E80000",
INIT_09 => X"187FC301B124F2001600000000001A1F00110101092CE7ED81CF000401228800",
INIT_0A => X"0477330C4889CC012188310E08812982050800A91012494C31004124080886FE",
INIT_0B => X"9861D1403803800C1000C1000C1000C1000C1000C1000C1000C1800608006084",
INIT_0C => X"020400830602410901000D02D0002008012054040022102001017FE190022201",
INIT_0D => X"3A0000401E030B0C20C20188087FFA07FE203A80010002608030102008100408",
INIT_0E => X"3A000005E8010000004000F808000010100F02000008003A00000F0200000800",
INIT_0F => X"00000002006B80800000400003B80000000F02000008003A00000F0200000800",
INIT_10 => X"01E03200060000080405E8010000100000F600000081003740400000008000EE",
INIT_11 => X"201D0100000039000007404000000E1000001846282010A211AA000000000080",
INIT_12 => X"80000000E808000001C200003A0200000072000007E00080000007E0000000A0",
INIT_13 => X"0100000003E200000280800EE04000000000F8080000A02022AC04000000003D",
INIT_14 => X"9C06D082000A03200806A040019481D4000000000201E1A000040000A02022E8",
INIT_15 => X"0401004010040100401004010060C040040C200950402090128057C3FF800C60",
INIT_16 => X"4010040100401004010040100401004010040100401004010040100401004010",
INIT_17 => X"0100401004010040100401004010040100401004010040100401004010040100",
INIT_18 => X"000000000000000000001000802FFFFFFFFFFFFFFFFF81004010040100401004",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000",
INIT_22 => X"2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_26 => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFF",
INIT_2E => X"F5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA080402000000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"02000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_36 => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_37 => X"0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_512_2,               -- Port A enable input
WEA      => wbe_a_lo_512_2(3),               -- Port A write enable input
DIA(0)   => data_write_a(31),        -- Port A data input
DOA(0)   => data_read_a_lo_512_2(31),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_512_2,               -- Port B enable input
WEB      => wbe_b_lo_512_2(3),               -- Port B write enable input
DIB(0)   => data_write_b(31),        -- Port B data input
DOB(0)   => data_read_b_lo_512_2(31),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_0_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"ED39BA795990D275FB4A6E96ACC4731DEA4598B0AFB54867F6EE4618C3749803",
INIT_01 => X"58A0047C8607844847CA180001E4A2404042106208408208C2002069161734B3",
INIT_02 => X"8B1EC9562121F8051500147A0E5629A302CF28400615F5787B09FBF999BB1EFD",
INIT_03 => X"404EFC0A2AD6100F01A88E851CE47803C280110521898F6996088862C7B22221",
INIT_04 => X"C0D001C0100AEC83C008E7880D01A64661800002C21A52C590D2012194804844",
INIT_05 => X"650002C3F08754001B51981E007910070F01C1E003980015A204C22F32328BAF",
INIT_06 => X"BCDA4677CAEE7CF5BB870E1DDB9889C5FBFC440129A0604442180238203F70C1",
INIT_07 => X"7AAE0088B02000C2EC3A0E829836E0AF3325372E2AA8FDF3C18306758B24197A",
INIT_08 => X"D7E40002F7AE005FFB4730010411400A61080000F7F4C464B58294901606D5A5",
INIT_09 => X"C4801C40469B0CA9881A28C141118000C5A85A60444210123820B43B40804274",
INIT_0A => X"400800219010107ED453C041B13216656074EA560F0092A24856B05312226900",
INIT_0B => X"27122C3E04E03383E2781EA781E2781EA781E2781EA781E2781C33C0613C0E29",
INIT_0C => X"74EB1F50D0758A9650E520610A6A57A5529E2B439499CF96B086000000B09870",
INIT_0D => X"04F07E024108F4E28638EC57250004480155C1375A97A9121F8BA749D3A4E9D2",
INIT_0E => X"04F07E42177EFDF8570184071575970F8FC07D5BFF078004F07E007D5BFF0780",
INIT_0F => X"8F85ECB1FE047F5FB7B30E0700461E5AF8007D5BFF078004F07E007D5BFF0780",
INIT_10 => X"C0184D07C1DF15C7E3E2177EFDF8C3C03009C3CDD47C7F403FB3FDF89701C011",
INIT_11 => X"4F80FE659C6104C6D7103F9D1D064189B5924418D65FE45DEE55BBEDE34CF900",
INIT_12 => X"6395F64207F3A3A1483136B881FCCB38C2098DACA01FFF603F80001F80FDC81F",
INIT_13 => X"FED151E01015C3BB507D3F811FBEC32B81840714F8D91F4FC513F37C8AE07002",
INIT_14 => X"61692F293185D8D724E15D3FCC6B7C236FE0691A9500125C1F83F8CC1F4FC507",
INIT_15 => X"E93A4E93A4E93A4E93A4E93A4F942F90E9628540052090650525A0000066A00B",
INIT_16 => X"93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4",
INIT_17 => X"3A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E93A4E",
INIT_18 => X"09B56C74DAB15D1CF13501AA495000000000000000003A4E93A4E93A4E93A4E9",
INIT_19 => X"2082082082082082082082082082082082082082082084E41DC71C7155F3898E",
INIT_1A => X"3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F8208208208208",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE5294A5294A52800003E1F0F87C3E1F0F87C3E1F0F87C",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000030FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"A975EFFFAABDE00FFAEBDFFF5D2EAAAAAF7AEBDEBA0000000000000000000000",
INIT_22 => X"8000155087FC0155F7D168B55007BFDF45085168ABA002E82145085155545F7A",
INIT_23 => X"FFFD7545AA8028A00A2802AABAFF8028BEF5D7FFFE10005542145557FD5545FF",
INIT_24 => X"F7AEAAAAAA2FFFDF4500043FE105D2E954BAF7FFC0010080017555555568AAAF",
INIT_25 => X"A5D5168A00A2D142155005142010FFAE820AAFF842AABAA2AE95545FFD168ABA",
INIT_26 => X"FF5D2A821550000000BA007FD55FF5D7FC0145007FD7400550415410002E974B",
INIT_27 => X"F455D5142000082E82145FFD17DFEFFFD168BFFF780000BA007FE8AAAFF803FF",
INIT_28 => X"0000000000000000000000000000000000000000AAFBEAA00007BFDFFF082EBD",
INIT_29 => X"AABEA495FC716F002A975FFE3AA95E00EBAEBDFD75D2AA8A80EA8E2FE3F00000",
INIT_2A => X"56A16D557BC257D415E0216FA3F1E8FC0145B68B551475FAF6D1C556F0AA1C24",
INIT_2B => X"7FD24AFE3D02DAAAE12BD5545A2803AA0000542A0070071C50BAFEF1FAE0016D",
INIT_2C => X"A8B50F55A2F150005A3A438BD04AFAB8F550A8010E004924874825D7FEAA8548",
INIT_2D => X"A2A5504001C74BA42A1571E8028E3DB7816D0120155EA568E870BAEB8A05A2AE",
INIT_2E => X"2FFAFD2A82485FD2415A105C21451ED42A002545E055FFBE81D0BE8EA8A3AA05",
INIT_2F => X"100AA1D0F6F480B6A555A2A57A002A3D5FDB6A5C7E3DFFFE90B45B47ABA497A8",
INIT_30 => X"A0AFE80A8B0A000000000000000000000000000000000000000000000B55EAAA",
INIT_31 => X"ABEF5D557FEBA55022A3F70C6B405F4D2AE975EFAAAAB5E1AF3AABFF45592E88",
INIT_32 => X"411A8DED57CE1055555E5F58EFFC01FE2CACB65F520EBE9EF67D7BEA1FD5D556",
INIT_33 => X"A4AD0079C75D6070CC5CBB0280C029ABAA3EBC114728007521170821CE0FDE69",
INIT_34 => X"2A95E02A2AAB5EB0F280800EFAEE9F5D18F3142341D5DEEBEF55080034E0A592",
INIT_35 => X"B69C30E02116220415A9540AA854140A0A2047F353AAF6C77F7F20D968BF5781",
INIT_36 => X"ABEBE1B4D792A4AD1183454180DD3FDCAAAB7C91565455C141E41887D58AC448",
INIT_37 => X"F0000001FF01EABC4B8014174FF7DA80F52FEDE6BE93172D7D625B556EEAB157",
INIT_38 => X"FF0000001FF0000001FF0000001FF0000001FF0000001FF0000001FF0000001F",
INIT_39 => X"0000000000000000000000000001FF0000001FF0000001FF0000001FF0000001",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000100000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(0),               -- Port A write enable input
DIA(0)   => data_write_a(0),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(0),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(0),               -- Port B write enable input
DIB(0)   => data_write_b(0),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(0),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_1_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"212C001411984004084D000508C53810A03D1450E839B003342114428A000803",
INIT_01 => X"08000011400A100A81160000008C005400400002000000000000028001340000",
INIT_02 => X"C084484000002014400205851002007030450E0000A606C8C44CB4C6666C00E0",
INIT_03 => X"33DF380008164004000002000C80400002031943000101091608463061120118",
INIT_04 => X"4140008000000002000064000400004201000000000210458010070080100433",
INIT_05 => X"8500101040200000010009100000000508000100000000002010600100208D04",
INIT_06 => X"B5EDFDE24618AD433060C182BA860044204C000008A004100008000820280020",
INIT_07 => X"581E02100020000A81244890AA20263030517F122AA801F0983060AC564BF808",
INIT_08 => X"00820800C7A00045B103200000140A02234808000584000004808400020011A4",
INIT_09 => X"0000104000020082800808111008400000200204100000100820800144000414",
INIT_0A => X"12804062945211441E13C051156E800008402802060C94000040901102800000",
INIT_0B => X"24002006406401918C191AC191A4191A4191AC191AC191A4191A00C8560C8D29",
INIT_0C => X"0408010040050880383820080F105F05800302E0E08842422006000000041032",
INIT_0D => X"05000600000090C1841808172580000000008008020084082080204010200810",
INIT_0E => X"0500066210000178470184000000878402C000001E07800500062000001E0780",
INIT_0F => X"00003C404600000011A30E0700000009382000001E07800500062000001E0780",
INIT_10 => X"C0180000012010C20022100000F0C3C03000000055200340000000F88701C000",
INIT_11 => X"05800241186100004D100098190240001290002050068000001010486140F900",
INIT_12 => X"0000164A001303204800026880048230C2000094A0000F601F8000000001C908",
INIT_13 => X"12D051E01000000154200580003C030381840000004B08014401025480E07000",
INIT_14 => X"40082300218450C2800010094000482142E0601895001000000041C408014400",
INIT_15 => X"0802008020080200802008020080008208600500A82A15008000000000468000",
INIT_16 => X"8020080200802008020080200802008020080200802008020080200802008020",
INIT_17 => X"0200802008020080200802008020080200802008020080200802008020080200",
INIT_18 => X"BABEFC54A0810C7452B5420A1000000000000000000002008020080200802008",
INIT_19 => X"AAAAAAAAAAAAAAAAAAAAAAAAAAA28A28A28A28A2A8218D2C0C92492581328A46",
INIT_1A => X"2E974BA5D2E974BA5D2E974BA5D2E975BADD6EB75BADD6EB75BAAAAAAAAAAAAA",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFF6318C6318C63000002E974BA5D2E974BA5D2E974BA5D",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"00000000000000000000000C0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"002155557FFFFFF007FC21EFA2FFD74AAAAD5555550000000000000000000000",
INIT_22 => X"7FD75FFAAAA800AAF7AA974BAFFFBE8B45F7AEBDF455D2EAABEFF7FFE8BFF5D0",
INIT_23 => X"0557DF45AAD1400BAA2AE801550051555EFF7AA95400552AAAABAFFD1574105D",
INIT_24 => X"FFFBEAB55F780020AAAA80020AA082EAAB5500517DF555D2EAAA105500001550",
INIT_25 => X"AF7AE820AA0851574BAA2D1574AA5D7BFDEBAFFD540155557FD5400F78028BFF",
INIT_26 => X"FFFFD56AAAAFFFFD7555AAD168B45AAAEAAABAFF842ABEF5D517DF55552A974A",
INIT_27 => X"4BAF7AE80010082A97410557FEABFFAAFBE8BEFAAD1575EF557FFFE10557FFFF",
INIT_28 => X"00000000000000000000000000000000000000005D7FFDF4500043FE105D2E95",
INIT_29 => X"A8BC2EBDFEAF7F1F840017D4975D2FEF147FC51C7A2FBD5490BFD1C056A00000",
INIT_2A => X"AA8AAAE3D145410F7F1D55D71C002DABAEBAA974BAF7FFEFB45FFAABDF55492A",
INIT_2B => X"0E2AE85028B40155145F7AF6DBED5450AA1C2080BEF495FC71D54124924385FA",
INIT_2C => X"571D2E28E38E0216FA2D1E8E80140F45082B4002D082082AB8B6DBEDB7DF7F54",
INIT_2D => X"A97F7AF6D417E92482BF84020BA495557E3FF78E021FF1471FDEAAFFD56F16D5",
INIT_2E => X"7002FD74951D71EDFFABFD16FAAAE92BD5545A2DA3FB7DAAD4AAAAF487BC70BF",
INIT_2F => X"550A8010E00492487482FFFE82A85EBAE2FFC55554ADBD7A2FFC7BEFF6FFD7FC",
INIT_30 => X"400FBF9424F7000000000000000000000000000000000000000000000547AB8F",
INIT_31 => X"DF55F7AABFF55082CA8B4DF6C1E8F5E5400021EF005162BEF047FD5545AAFBF7",
INIT_32 => X"404547184164AA5D2EBEEB0A2D555410D3555714F8338AAAA1D0AE974AAF7FFF",
INIT_33 => X"AEABFFDF79DCBF755962010BDCBBC21455D7FEABEF75550ACBB7582225FF5843",
INIT_34 => X"D57D412F7D55F5E50C7F401BAAE8403CF5A3FFEAAEB083BC1000FF8409000512",
INIT_35 => X"2AA9FEAFDF7F431A9F7FFE81FF013A8001AFF801F8BA0C57740BDAA0688E5405",
INIT_36 => X"A2FBF7FED2C7F955445079E280A00C56145EF5D16BABAA3EBC3157ABD5FFE55F",
INIT_37 => X"0000000000596EBEF55080034E0A592A4AD00FB863550229BCABEB7DA403FFFD",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000100000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(0),               -- Port A write enable input
DIA(0)   => data_write_a(1),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(1),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(0),               -- Port B write enable input
DIB(0)   => data_write_b(1),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(1),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_2_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10E006600180111284380310006289800480032283E000A34301002001A0817",
INIT_01 => X"A14AC00A1079284D04A044A54E504368404000720885800802000006ECD10200",
INIT_02 => X"92250052A0348C310102048800A8507000040C8550200000480E0080001321E0",
INIT_03 => X"020204E4593C0824400C2220483042809292430400440180000890A4C9400242",
INIT_04 => X"486854B141002252142241502460480031B94420634850069A42241009610A04",
INIT_05 => X"800504244080892105AA6010A44882144840910A21220A8C820025E4A0000B00",
INIT_06 => X"A000442802280000340810209C444804206000AC800088096A0EA8C022208012",
INIT_07 => X"309820A848E0AA09826489A5CC49002001020112028201F8A20488260000108A",
INIT_08 => X"2400582881E0C1419D12041455509341A539C42A0D8208099002801700D10103",
INIT_09 => X"110D525861263100009200151409130A3C80C8C8096A06B8C12088400A9C2080",
INIT_0A => X"0451394CD0391A441583C04B580040089581001342801044877200D002A00DE0",
INIT_0B => X"144423040240450114901149013C9011C9013C9011C90134901144801A4808A5",
INIT_0C => X"D8A5345206D2C10082080A90C00000188150100C202A4640000E2B4081969420",
INIT_0D => X"050080400A0391A51240C480000AA902AA009028C83220008086952B4285A54A",
INIT_0E => X"05008021C00000000040000000020288000500000008000500802A0000000800",
INIT_0F => X"0002300000428000000040000000000D002A0000000800050080250000000800",
INIT_10 => X"0000000001204004000508000000100000000002054000130000000000800000",
INIT_11 => X"000C00000000000068144000000000001A000106200010021002000000000080",
INIT_12 => X"0002004A880000000000034098000000000000D024A000000000000001000900",
INIT_13 => X"00000000000000041400000A8000000000000000010A00000284000000000000",
INIT_14 => X"012100000002000280000000011080C000000000000000000000430000000260",
INIT_15 => X"A769DA769DA769DA368DA36CDA3A9A13A14801404134DA84A024024155000399",
INIT_16 => X"168DA769DA769DA769DA368DA368DA368DA769DA769DA769DA368DA368DA368D",
INIT_17 => X"68DA168DA169DA569DA569DA568DA168DA168DA169DA569DA569DA568DA168DA",
INIT_18 => X"138D70C030B51C50C7D000A2012F81F81F83F03F03F069DA569DA569DA568DA1",
INIT_19 => X"1041041041041041041041041041041041041041024860208165965975960040",
INIT_1A => X"25128944A25128944A25128944A25128944A25128944A2512894104104104104",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFF8421084210840703F25128944A25128944A25128944A",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"00000000000000000000000F0FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"415555087BFFF55A2AA800BAFFAE9540008002AA000000000000000000000000",
INIT_22 => X"7FE8B555551421455D0002145552EBFEBA007FC21EFA2FFD75EFAA8415410AA8",
INIT_23 => X"FFFE8B45552EBDF45FFAEAABFFF7FFE8B55F784155EFA2AEBDEAAA2FBEAABA5D",
INIT_24 => X"5D2AAAAAA5D2E820BAA2FBEAB5555557DF55A2AEBDF555D2E954BAA2AA974BAF",
INIT_25 => X"A5D04021EF557FC21FFAA8428BFFAAAA954AAAAAAAAAAAFFD1574105D7FFFF55",
INIT_26 => X"EFF7800215500557DF55AA80001FFAA80001550055575EFFF84021555D043DEA",
INIT_27 => X"B5500517DF555D042AA10A284154005D0015410085568A00FF80175FFA2D17DF",
INIT_28 => X"00000000000000000000000000000000000000005D00020AAAA80020AA082EAA",
INIT_29 => X"D55D2BE800042AFE8E1557D0075D2F45BEAA800AAFFAA9543A080038A2A00000",
INIT_2A => X"0BDEAAA2FBF8AAA557BE8B6D5D5FFABEF49040017D5D20B8EAA007FC51C7A2FB",
INIT_2B => X"0E174BFA02A974BAF7F5EFB455D2ABDF55492AA8BC7EBDFEAFEFFD00105FFBC2",
INIT_2C => X"3D155E105571D55D71C002DABA5524820BAB6FFEFB6D555578F7DB6A0BDF7D48",
INIT_2D => X"092A071555D5E3AE821D00001FF0871C016DBED1FDE90E3A497492B6AAADAAAE",
INIT_2E => X"0E3DA3DFD5E3DFFFBD5A38A021551C5F7AF6DBE8F401D7B6A0001470155C51D0",
INIT_2F => X"82B4002D082082AB8B6D1C5B7DF7FF78E075C5BE8555400550A38428007FED00",
INIT_30 => X"4AA00042AAA2000000000000000000000000000000000000000000000410F450",
INIT_31 => X"AAAA007FD5555AAFBD7545FBB8020A3F7AE975EF005560B55F7AA800AAF7AA95",
INIT_32 => X"E8F5EFF84165EFF7802BAB0A2FFEAABA557BEABEF057D68F5F5A00021EF55042",
INIT_33 => X"52ABFFFF841FFE75CA882108202E974AAF7D57DF55D7AABFF5428ACA8F45A6C1",
INIT_34 => X"84174A8FFAEBFEB0A2D55541051555694F002CA8AA80800020AAF7FBFFFEF045",
INIT_35 => X"7AAA155F595542455512A975455D3AA8A005500151FF0C57401E5F3D1E00A1A8",
INIT_36 => X"5D2A8A0B882FFFFE10AAAAAB755A66B6AF56A2AA801455D7FE8BFFF680800FFF",
INIT_37 => X"00000000000C3BC1000FF8409000512AEABFF5D79FCAF774AE005BE789555400",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000200000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(0),               -- Port A write enable input
DIA(0)   => data_write_a(2),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(2),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(0),               -- Port B write enable input
DIB(0)   => data_write_b(2),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(2),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_3_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"210C44A20020248B08431120001604B8156023104C4077133420400A02380202",
INIT_01 => X"015A2A424080216D3C2462C99E104B49404040028804A0080A000C16A0D90A0C",
INIT_02 => X"C0A4065000F0A95011000D1501005270B4045AB330860281CC08008222170060",
INIT_03 => X"AD22014098340394A4021320080841C40B411B4298042180002846B06900811A",
INIT_04 => X"244B32A86D20014A0D20403194904900071A24110F0BF400F85F92420E0C946E",
INIT_05 => X"80331030442898B4812840D0500008C528280B063006A64CA30004E5A4E40304",
INIT_06 => X"90016CA00E380042302040A0BC47160424428198C0038C89904E640023600816",
INIT_07 => X"1288020843A66620816049908AA0061011CA0142000009F0A810292E7402F088",
INIT_08 => X"20003C9984A0AC411102014D34EC2200214D5099048823019603A01A49410103",
INIT_09 => X"001CD74C4826220010A8891451284B661CA24A4C899046740121824004100080",
INIT_0A => X"44C9516DC0135C45159BE45F112B48804DC10203021290400772C0F402820D4C",
INIT_0B => X"B400624402404501A49018490184901A4901A4901849018C901A648056480C2D",
INIT_0C => X"D7A9B54000D7C10820680D08C420180381211081A022160000266723E1909021",
INIT_0D => X"400080200E199A4A2CA2994C0399981666409800CA52E4890806BD6B56BDAB52",
INIT_0E => X"40008008E00000000000000000024008000C8000000000400080028000000000",
INIT_0F => X"000A000000588000000000000000200400088000000000400080078000000000",
INIT_10 => X"0000001000004004000D800000000000000000022040000B4000000000000000",
INIT_11 => X"001A0000000000082006C000000000020804087220000122000A000000000000",
INIT_12 => X"00020800B8000000000041002E00000000001040466000000000000001020080",
INIT_13 => X"00000000000000048200004A600000000000000003008000320C000000000000",
INIT_14 => X"432900000222200871028000210400C4000000000000000000080200800030E0",
INIT_15 => X"AF6A5AF6A5AF6A5AF6A5AF6E5AFADA91AB68000101B4D20C08EC461733804A19",
INIT_16 => X"B6B5AF6A5AF6A5AF6A5AF6A5AF6A5AF6A5AB6B5AB6B5AB6B5AB6B5AB6B5AB6B5",
INIT_17 => X"6BDAB6B5A96ADAF6A5AD6ADAF6A5AD6ADAF6A5AD6BDAB6B5A96BDAB6B5A96BDA",
INIT_18 => X"C78C706428A14C586290008A044D54AAB556AA9556AAEBDAB6B5A96BDAB6B5A9",
INIT_19 => X"92492492492492492492492492410410410410412821600001249249015303C0",
INIT_1A => X"351A8D46A351A8D46A351A8D46A351A9D4EA753A9D4EA753A9D4924924924924",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000001543B351A8D46A351A8D46A351A8D46A",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"43DF55FFAA955EFA2D168B55557BEAA000055420000000000000000000000000",
INIT_22 => X"7BE8BFFA2D155410AA8415555087BFFF55A2AA800BAFFAE9554508002AA00AA8",
INIT_23 => X"52ABFEBA007FC21EF007FD75FFAA841541008002AB55AAAA955EF005568A0008",
INIT_24 => X"005168B455D042AB45F7FFD741000042AA10AAAABFF5508003FF555D00021455",
INIT_25 => X"0A2D1575FFF7AA975555D2E80145F78415545082EBDEAAA2FBEAABA5D7FC0155",
INIT_26 => X"55552A954BAFFFFE8B55552EBDE00F7AEAABFFF7FBEAB55F7AABDEBA5D7FC201",
INIT_27 => X"F55A2AEBDF555D2E954BA002EAAABA002A821EF5555554AA087BC01FFFFAAAAB",
INIT_28 => X"0000000000000000000000000000000000000000082E820BAA2FBEAB5555557D",
INIT_29 => X"95578080038A2AA28E3AF55E3A0BA5D7AADB6FB7D5D7FEAA3808554203A00000",
INIT_2A => X"0925D7085F6AA10087FEABD7AAD57AEBAB68E1557D1475FAF45BEAA800AAFFAA",
INIT_2B => X"04AAFFA41040017D5D20B8EAA007FC51C7A2FBD55D7BE80004AA1E8E2AB55B6A",
INIT_2C => X"2FBE80AA557BE8B6D5D5FFABEF49002FB55FFF5D0438140E2FA38B6AEBFF6D1D",
INIT_2D => X"AB8ABAE925D21C7010EADB525D7FFAE975C75D0A901FFFF801557D1C20B8EAAA",
INIT_2E => X"20875C21D5EB8AA8FFF012A954BAFFF5EFB455D20BDE00EBAAA8BC7EBDFEAFEF",
INIT_2F => X"BAB6FFEFB6D555578F7DB6A0BDF7DEB8E125FF002EADA921420871D74971D248",
INIT_30 => X"ABA0051400A20000000000000000000000000000000000000000000001C24820",
INIT_31 => X"8B55F7AA800BAF7AA955EF00042AAA2A2AEAAB55A28408145AAFFFFFFF5D7FEA",
INIT_32 => X"020A35D2ABEF55F7800015F087FEAA00007FEAB55FAD568AA2AFAE975EF55516",
INIT_33 => X"ABFEAAF7AE9DFF759A82AEF70800021EF55042AAAA007FD55558A7BD7145FBB8",
INIT_34 => X"84175EF55002AAB0A2FFEAABA557BEA3EF057968F575D003FF55F7D5420BA5D2",
INIT_35 => X"A8429F45A7D5EAF5FFBAEAAA10554155400AAFFD5145FBAC9755F05040255FFD",
INIT_36 => X"550415557085540000005156155FE90A8F5C082E974AAF7D57DF45552A3FF10A",
INIT_37 => X"00000000005500020AAF7FBFFFEF04552ABFFFF843FFE77C80825BC052ABFE10",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000100000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(0),               -- Port A write enable input
DIA(0)   => data_write_a(3),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(3),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(0),               -- Port B write enable input
DIB(0)   => data_write_b(3),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(3),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_4_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A108400020612C80284210081034849800A000303100048B3432C82904204002",
INIT_01 => X"21066802000820491C00650E1E004360403008418984014902030906A8D10200",
INIT_02 => X"120404E00E4C0600000206100008402005040C00F104008040080080001310E0",
INIT_03 => X"DCA201514D1C0D706C5CF010083A0708BA0841945004010000080084C1000002",
INIT_04 => X"5C4CF21C48B133483C80417570D000083A62488074C1350EA60D785C0A6B0619",
INIT_05 => X"000F0400028083B381A60001E5546EB5C0E2B81E4166DE000139200004E50940",
INIT_06 => X"80004408020800023000102098000204A040038600018019004B800123208806",
INIT_07 => X"120C20204665E1008024188488800000001A01520000A1F08044892400001088",
INIT_08 => X"0801007AC0A1EB413102063CF3E0B3028D29F407059B0B000205A801C2200102",
INIT_09 => X"106052400922D00406BE1002C6150F41200280001900439001FD8A0004142000",
INIT_0A => X"047F2201D899BA503583504B58AB80804540001202805544314041B48A888EC5",
INIT_0B => X"1441E3443043410C5010C3010C1010C3010C1010C1010C3010C14086980861A5",
INIT_0C => X"020000A02600000805400502C0A0004A00625015000A12000026E1E180011220",
INIT_0D => X"400000000E43930C20C20188120782861E4004A800600401A030001008080400",
INIT_0E => X"40000021A8800000000000000000400800170024000000400000310024000000",
INIT_0F => X"0008000000AA80200800000000002000003400240000004000003B0024000000",
INIT_10 => X"00000010000000040004A080000000000000000020400006C008020000000000",
INIT_11 => X"002C008200000008001B4020200000020000090760000200110A040010000000",
INIT_12 => X"00000803E004040000004000E801040000001000086000000000000000020040",
INIT_13 => X"0000000000000000810000164001008000000000020040002240008020000000",
INIT_14 => X"04001040026026004000000002940040000410000000000000080000400000B8",
INIT_15 => X"040080201004008060000001806AC000004890015124D880100886D8F0014420",
INIT_16 => X"4010000180600000018020100400802010000080601000008020000401802000",
INIT_17 => X"0100000004008020180600000000000180600802010000000401802018020000",
INIT_18 => X"3807E05000140634504048820064B261934D964C326980004010000080600806",
INIT_19 => X"AAAAAAAAAAAAAAAAAAAAAAAAAAA28A28A28A28A2934C8D0CCD145144C0A28A06",
INIT_1A => X"068341A0D068341A0D068341A0D068351A8D46A351A8D46A351AAAAAAAAAAAAA",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000000173F068341A0D068341A0D068341A0D",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"57FE10FFFBEAA10007FD7410FFAA97555082A800AA0000000000000000000000",
INIT_22 => X"7FEAA00007BE8AAAAA843DF55FFAA955EFA2D168B55557BEAB45005542000005",
INIT_23 => X"87BFFF55A2AA800BAFFAE9555508002AA000055574105D2A800AA00043FEBA5D",
INIT_24 => X"A2D17DE1000517FE10AAAAA8AAA002E97545557BC00AAA2FFEAAAAAA84155550",
INIT_25 => X"0A2D157400AAAE974AAAAAA974BA08002AB55A2AA955EF005568A00087BE8BFF",
INIT_26 => X"BA080002145552ABFEAA007FC21EF007FD75FFAA8417410A2D140000F7FBC201",
INIT_27 => X"A10AAAABFF5508003FF55F7D568A00552EA8BEFA2AABDEAA087BEAAAAA2FBD54",
INIT_28 => X"000000000000000000000000000000000000000055042AB45F7FFD741000042A",
INIT_29 => X"EAB7808554203A145178E00FFFBE8A101475D5400F7A49057D0824850B800000",
INIT_2A => X"E8008200043FE925571EFA380871C7028A28E3AF55F7A0925D7AADB6FB7D5D7F",
INIT_2B => X"F5FDA38BE8E1557D1475FAF45BEAA800AAFFAA9557D080038AAA145157428492",
INIT_2C => X"85F6AA10087FEABD7AAD57AEBA08517DE00AAAEA8A9200249056D4175C5092AA",
INIT_2D => X"FEDB42028EBFBC2028BED152438AAA092492AAA4954281C0E2FB55B6A0925D70",
INIT_2E => X"A0875EDA80BEF1C743840040017D5520B8EAA007FC51C7007BD55D7BE80004AA",
INIT_2F => X"55FFF5D0438140E2FA38B6AEBFF6DBE84AAEBAF7DF6AA00412EAABFFAA803DEB",
INIT_30 => X"1EF0800154B200000000000000000000000000000000000000000000041002FB",
INIT_31 => X"0145AAFFFFFEF5D7FEABFF0051400A25D5568A00FFFFEAA105D5155410FF8402",
INIT_32 => X"2AAA25555410BA082E8201000043FE005D517DEBA0851574B2AAAEAAB55F7840",
INIT_33 => X"4001FF005575408AA557FEB2FFAE975EF555168B55F7AA800BAF7AA955EF0004",
INIT_34 => X"2ABFF55F7800015F087FEAA00007FEAB55FAD568AA200557DE00AAAAAAA00080",
INIT_35 => X"87BD6145FAAC000A2A6FBC00BAAAFBC00BAF7D1550AAAA8002010F2AC154B25F",
INIT_36 => X"082EA8BFFAA843FEBA08517DE00F3F9574B30800021EF55042AAAA007FD55550",
INIT_37 => X"000000000008003FF55F7D5420BA5D2ABFEAAF7AEBDFF779A82AA43F7FBE8A00",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000200000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(0),               -- Port A write enable input
DIA(0)   => data_write_a(4),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(4),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(0),               -- Port B write enable input
DIB(0)   => data_write_b(4),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(4),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_5_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50DF4A0791B3FCB694379283C81FD996A091832102004A337A20E07C0C1E006",
INIT_01 => X"294014468000A04D5C6A60000C34C24841280A00084000C8C212892EEAD53235",
INIT_02 => X"50AE41540CA1D9100002171C1F0A5171134E2A200D8633F8CD09DBFBBB970E7C",
INIT_03 => X"214E3C521D16021B64430CC51C45B8154689094241898749920842946B90010A",
INIT_04 => X"A2F20F7D7A314CB5C208E28A1BF0224A448920028A185340D0C20B2690000C22",
INIT_05 => X"7520B430B20B984809A8886E230C6106371146E1829941C58310402C600381CF",
INIT_06 => X"9CC96CD7C63A7495B9A356ACBC4601C57FD44F8549A46490261C4B39203F7080",
INIT_07 => X"12A88800B029E0C0A12C4B92AA36A2111167357C220095F3C8952A2E5D26F078",
INIT_08 => X"F3F00503B4AE105B534711820C0C0A1043080300F7E0E728B1829C2FEA0A95A1",
INIT_09 => X"C5184F084136848C9298A8560688F480C58858449026145B3830F40944906234",
INIT_0A => X"50EB4124D2B3902BF5C9700C1199DCA84DF46A974F92C7E28F1630D38088A438",
INIT_0B => X"B3144E5636E3178C86B8CC6B8CA6B8CE6B8C86B8CE6B8CA6B8CC15C6435C670C",
INIT_0C => X"79E51E70E070AA8132252008360A7E91504104C8948047D6B0AE1FE440B28A71",
INIT_0D => X"05F0FE40014090400400080329FF8089FF49611F589765923E139F09C78CE7C6",
INIT_0E => X"05F0FE64037FFD7857418407157797878F005F0DFF0F8005F0FE205F0DFF0F80",
INIT_0F => X"8F87FCB1F8053FDEB9B34E0700461E5FF8205F29FF0F8005F0FE205F29FF0F80",
INIT_10 => X"C0184D07C1FF55C3E3E0037FFCF8D3C03009C3CFD53C7E001FF2FAF89781C011",
INIT_11 => X"4E0CDF47186104C6FF177BD939024189BF900401165D645CEEF5BBCDF148F980",
INIT_12 => X"6397F64AEF7F2320483137F8A9BF8A30C2098DFCA06FFFE01F80001F81FDC94F",
INIT_13 => X"FFD051E01015C3BF553D3E0E5FFE838381840714F9DB4F4FA213F774A0E07002",
INIT_14 => X"8B652E2B3120C81284641D3E8DBF7D636FE070189500125C1F83FBCC4F4F80EF",
INIT_15 => X"E7394E339CE138CE5394E33D4E1E0E30E1208C251134921C12A44103F064014B",
INIT_16 => X"7384E3394E338CE538CE1394E3384E738CE139CE1394E7384E339CE139CE5384",
INIT_17 => X"38CE139CE1384E7384E7394E3384E738CE539CE139CE538CE5384E3394E7384E",
INIT_18 => X"7F7B9DB7FF3A1B6DB7ED438A9C3124B2DA6924965B4D384E7384E339CE138CE5",
INIT_19 => X"FBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEF9F7CFDFDDCF3CF3DF5E5BB4E",
INIT_1A => X"7BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEFBEFBEFBEFBE",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE000000000000118D27BBDDEEF77BBDDEEF77BBDDEEF7",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"E955450055421FFFFFBC0010AAD5574BA557FFDFFF0000000000000000000000",
INIT_22 => X"D5575EF55517FF5500557FE10FFFBEAA10007FD7410FFAA97410082A800AAAAA",
INIT_23 => X"FAA955EFA2D168B55557BEAB55005542000007FD74000055574BA5D7FD7555A2",
INIT_24 => X"007BC00AAAAAEBDF45A28428B45FFD168BFF00002AABA5D2ABFFFFAA843DF55F",
INIT_25 => X"AFF80174BAAAD1555EF5555555550055574105D2A800AA00043FEBA5D7FEAA00",
INIT_26 => X"FFAA8415555087BFFF55A2AA800BAFFAE95555080028A00A2FFFDE00F7D57FEB",
INIT_27 => X"545557BC00AAA2FFEAAAA082A97545F7D5420BA5D2E821FFA2D5554BA557BD75",
INIT_28 => X"000000000000000000000000000000000000000000517FE10AAAAA8AAA002E97",
INIT_29 => X"9043D0824850B8A2AE9756D145B401FFFFFFC7010BEDF524AA5571FDFEF00000",
INIT_2A => X"1524BA5571D757DB6D5525EF555178F6D145178E00EBFBE8A101475D5400F7A4",
INIT_2B => X"24BFFFFA28E3AF55F7A0925D7AADB6FB7D5D7FEAB7D0855420BA1471D7438085",
INIT_2C => X"0043FE925571EFA380871C7028B6AEBDF45B68A28B6DEBDF6DBEF1C0A28AAA55",
INIT_2D => X"A2FBF8E10EBD578EAAFF8415482BED1555EF55555057D145152428492E800820",
INIT_2E => X"FB6DF574A85575C55EFBE8E1557D1475FAF45BEAA800AAFFAA9557D080038AAA",
INIT_2F => X"00AAAEA8A9200249056D4175C50920875FDA381C209256DFFDF420BA552A821F",
INIT_30 => X"0BA55557DFF700000000000000000000000000000000000000000000008517DE",
INIT_31 => X"AA105D5155410FF84020AA0800154B2AAAA975FF5D7BC21EFF7FBD7400F7FBC0",
INIT_32 => X"400A25551554BA0051400BA5551575EFF7D1401FF5D5568BE7555568A00AAFFE",
INIT_33 => X"FFDFFF552EA8AAA55043DFF7AAAEAAB55F78400145AAFFFFFEF5D7FEABFF0051",
INIT_34 => X"55400BA082E8201000043FE005D517DEBA0851574B2FFAABFF45FFAAAABFFAAF",
INIT_35 => X"7AA955EF00002AAA2A2FBE8A00A2D16AAAAFF8002410FFD5575EF5555421E755",
INIT_36 => X"FFFFC00BA552A821EFFFFFD74BA5D51575F7FFAE975EF555168B55F7AA800BAF",
INIT_37 => X"000000000000557DE00AAAAAAA000804001FF0055554088A557FEB25D00021FF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000C00000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(0),               -- Port A write enable input
DIA(0)   => data_write_a(5),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(5),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(0),               -- Port B write enable input
DIB(0)   => data_write_b(5),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(5),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_6_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10800B0061A01002840002C03002818000402322520070B313301C4389B2082",
INIT_01 => X"274008482009404C18A160000C52424841000000090800090210000008510200",
INIT_02 => X"102430600C800110000006100009D070012408000000000648080000001210E0",
INIT_03 => X"000200501D1D02140C420200480140040608010040400104681A0084490C4802",
INIT_04 => X"404402820021000A00824002141000980500000808001114C000080624600600",
INIT_05 => X"120024204209981001A806500304610528000500000080000000300000012940",
INIT_06 => X"2000440832280002300010209C4400142061207A024008900008000220600220",
INIT_07 => X"130C8A220FF41F00902008808800182001020150000001F0800408264000100A",
INIT_08 => X"001BF002C4A01041B1120101000010128568837F04842B080020890008080342",
INIT_09 => X"011847140126805432A62A1596C8B5DF10000008900000100220C00084000008",
INIT_0A => X"44EB4104D09392053589F11C59898888454010830212C54081000410A0088C00",
INIT_0B => X"B0044245B25B456C0096C0096C4096C4096C2096C2096C6096C444B6004B600C",
INIT_0C => X"09040020280010000B3002820110101D0012402CC00802410C26800860070621",
INIT_0D => X"0500819D0000900208201040C4007920004884080000448C281018100C000200",
INIT_0E => X"05008182100000000000000000022AE800C00004000000050081A00004000000",
INIT_0F => X"0002330006000000080000000000000D07A00020000000050081A00020000000",
INIT_10 => X"0000000001204A340002100000000000000000020F4001400000020000000000",
INIT_11 => X"019300020000000068D08000200000001A692121000280000000000010000000",
INIT_12 => X"000201FA100400000000034696010000000000D3478000000000000001003F00",
INIT_13 => X"00000000000000043C0001C0A000008000000000012E000054AC000020000000",
INIT_14 => X"0200000040A410C2810800016000809400001000000000000000433300007600",
INIT_15 => X"060180400000008060180404002AC0200208940041309210B28048180F028000",
INIT_16 => X"2008000100601802000000100601800000000180600800000020180600000000",
INIT_17 => X"0180600000008040100200800000060100000802010040180200002018040100",
INIT_18 => X"7F8FF0F4FA955F7CF7F40A80907638C31C71C718638E00006018040080200004",
INIT_19 => X"38E38E38E38E38E38E38E38E38E38E38E38E38E39B6CEDECDDF7DF7DF5F78BCE",
INIT_1A => X"3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE38E38E38E38E",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFF000000000000196A03F9FCFE7F3F9FCFE7F3F9FCFE7F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"00000000000000000000000C0FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"BFDF45F7AA974AAAAAA97555F784174BAF7D5555FF0000000000000000000000",
INIT_22 => X"FBD7410AA8428AAAAAAE955450055421FFFFFBC0010AAD5574BA557FFDFFF087",
INIT_23 => X"FFBEAA10007FD7410FFAA97400082A800AA08515555508043FE00F7AA97555A2",
INIT_24 => X"55517FF55A2AA97400552AAAB45082E80155F7D1575EFFFAA9555500557FE10F",
INIT_25 => X"FF7AAA8A10082EAAB45A2FFC2000007FD74000055574BA5D7FD7555A2D5575EF",
INIT_26 => X"FFAA843DF55FFAA955EFA2D168B55557BEAB5500554200000003DE10FFD5401F",
INIT_27 => X"BFF00002AABA5D2ABFFFF087BD5545007BFDE10AA803FE105D516AABAFF843FF",
INIT_28 => X"0000000000000000000000000000000000000000AAAEBDF45A28428B45FFD168",
INIT_29 => X"524AA5571FDFEF1C7BFFF55FFA095482B6A49256DEB84104BAFFD1525FF00000",
INIT_2A => X"03DE28F7A49057DAAF5D2428A2842AAAAA2AE9756D145B401FFFFFFC7010BEDF",
INIT_2B => X"A49756D145178E00EBFBE8A101475D5400F7A4904380824850381C5B5057D1C0",
INIT_2C => X"571D757DB6D5525EF555178F6DAAA495428412AAFB451C2A8017DE3DF525FFFF",
INIT_2D => X"1C0E3FE00E3DB471EFE3AAAAA00082EA8B6DA2F1C50381471D74380851524BA5",
INIT_2E => X"049516AAB8FF8428FEFA28E3AF55F7A0925D7AADB6FB7D5D7FEAB7D0855420BA",
INIT_2F => X"45B68A28B6DEBDF6DBEF1C0A28AAA5524BFFFF1C7BD057D1C71FFE10A28038E1",
INIT_30 => X"0AAFFD1401E7000000000000000000000000000000000000000000000B6AEBDF",
INIT_31 => X"21EFF7FBD7400F7FBC00BA55557DFF7557BFDF55F78017400F780001FFAA8400",
INIT_32 => X"154B2557FC01EF55043FEAAFF80021EFA2D1420BAAA8428AA2AAAA975FF5D7BC",
INIT_33 => X"A821EFAAFBC01FFF780155F7555568A00AAFFEAA105D5155410FF84020AA0800",
INIT_34 => X"51554BA0051400BA5551575EFF7D1401FF5D5568BE7AA80174AA082ABDF555D2",
INIT_35 => X"D7FEABFF0051400A25D2EBFE10AAFFD55EFA2AEA8A10082EA8BEFAAD5554B255",
INIT_36 => X"55557DE00AA842AA0000516AABAFF8428BE7AAAEAAB55F78400145AAFFFFFEF5",
INIT_37 => X"0000000000FFAABFF45FFAAAABFFAAFFFDFFF552EA8AAA55043DFF7557BC01EF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000900000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(0),               -- Port A write enable input
DIA(0)   => data_write_a(6),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(6),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(0),               -- Port B write enable input
DIB(0)   => data_write_b(6),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(6),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_7_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10844B00482258A2842112C02450418800002300500030B313300C418992002",
INIT_01 => X"234008422008604D1C20E0000E11426840000000080000080200090000110204",
INIT_02 => X"1025207000B08910000206101188D03080144880010400044808000000122160",
INIT_03 => X"000200401914821004420000CA01000C0600010000605114291A008449484802",
INIT_04 => X"40440200002100080006500210101019040000000B085024D842080244000000",
INIT_05 => X"1A8024200009981001A8224001040104200204000000800CC2092CE4A0004900",
INIT_06 => X"A000440822280002340010209C040014A061200052500810000C490323208E28",
INIT_07 => X"128802020028000890240980A809102001020140000009F0800408264000100A",
INIT_08 => X"001A0602C4A01051B13281010408881203480200448423199046821008082351",
INIT_09 => X"336784144126811054809C1040140A001C8648481000045903318B80A400310A",
INIT_0A => X"000800009010100014114110312388984502148282A08415B032095048008100",
INIT_0B => X"20CDC1C483484D201192011920119201192051920519205192074C9018C90188",
INIT_0C => X"D8A5B44001D2C12901228F82F005310D293054048A2212004466000DA1908528",
INIT_0D => X"800F8108A0D09802082010408580008000000008C85264010816851B428DA146",
INIT_0E => X"800F81321000020000261900E28A204040E000A0000007800F814000A0000007",
INIT_0F => X"7072024807000020400000581C01C1A406400084000007800F81400084000007",
INIT_10 => X"060180E83800E820101210000200000CC3003C32080201C0000C000000160700",
INIT_11 => X"81DD00804086423120B74020023090644840A34000828800000004000420020B",
INIT_12 => X"1C6A0186E8000446120C8905BA0004810C84624237E00010001878007F0030C0",
INIT_13 => X"00080208E4083C44230201AEE0010040261900E30520C0806EAC0082000984C0",
INIT_14 => X"0121011088A600C032128201519480D40005802448160403E0700622C0806EE8",
INIT_15 => X"A1685A1685A168DA368DA36CDA30DA13A108810111349A943AA4401000928A19",
INIT_16 => X"368DA768DA1685A1685A5685A368DA368DA7685A1685A1685A768DA368DA368D",
INIT_17 => X"685A1685A169DA368DA1685A1695A368DA3685A1685A168DA368DA1685A1685A",
INIT_18 => X"00000000000000000000400A8448410400020820800069DA1685A168DA369DA3",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000003667B000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"0155EFAAAEA8ABAAAFBFDE0055556AA005D04155550000000000000000000000",
INIT_22 => X"556AA00FFAE95555087BFDF45F7AA974AAAAAA97555F784174BAF7D5555FFF78",
INIT_23 => X"055421FFFFFBC0010AAD5574BA557FFDFFF5555555EFAAFFFDFEFAAAAAAB455D",
INIT_24 => X"AA8428AAA557BFDFFF55003DFFFF7FBEAA00002EAAAAA082EA8A00AAAE955450",
INIT_25 => X"0552EBDE00007BEAAAAA2D14000008515555508043FE00F7AA97555A2FBD7410",
INIT_26 => X"FF00557FE10FFFBEAA10007FD7410FFAA97400082A800AAF7AE975FFA2800001",
INIT_27 => X"155F7D1575EFFFAA955555D51574AAAAFFD5545087FEAB455D516AB55557BD55",
INIT_28 => X"0000000000000000000000000000000000000000A2AA97400552AAAB45082E80",
INIT_29 => X"104BAFFD1525FFFF8E175C7A2AAAAA82A2F1FAE105D556AA10410E1755500000",
INIT_2A => X"1FFFD7AAAAAFB7D495F6AA10E3AE905551C7BFFF55FFA095482B6A49256DEB84",
INIT_2B => X"2EAAA00A2AE9756D145B401FFFFFFC7010BEDF524AA5571FDFEF415B575D7AAF",
INIT_2C => X"7A49057DAAF5D2428A2842AAAA497BFAFFF49003AFEFEBFBEAA001C2EA8A821C",
INIT_2D => X"F7A4905C7A28A070384120BDE100075EAA82BEDB470101C5B5057D1C003DE28F",
INIT_2E => X"D555F6AB57417BC05D7145178E00EBFBE8A101475D5400F7A490438082485038",
INIT_2F => X"28412AAFB451C2A8017DE3DF525FFFFA49756D495150492BEF1D2555087BE8B7",
INIT_30 => X"A10002E9754D000000000000000000000000000000000000000000000AAA4954",
INIT_31 => X"7400F780001FFAA84000AAFFD1401E7FFAA97555A2AEA8A10AAD568A00555168",
INIT_32 => X"7DFF7007BD5555AAD57DF55AAAEBDFEF007BE8A10AAAE8215D557BFDF55F7801",
INIT_33 => X"FEAA105D2EAAA005D2AAAA18AAAA975FF5D7BC21EFF7FBD7400F7FBC00BA5555",
INIT_34 => X"7FC01EF55043FEAAFF80021EFA2D1420BAAA8428AA2007FE8BFF080028BFFAAF",
INIT_35 => X"F84020AA0800154B2FF8402145A2AA954AA00043DE0000516AA10F7FBD740855",
INIT_36 => X"FFD140145007FE8BEF557BEAB55087FC215D555568A00AAFFEAA105D5155410F",
INIT_37 => X"0000000000AA80174AA082ABDF555D2A821EFAAFBC01FFF780155F7005140000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000000FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(0),               -- Port A write enable input
DIA(0)   => data_write_a(7),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(7),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(0),               -- Port B write enable input
DIB(0)   => data_write_b(7),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(7),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_8_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00000648E2840112C00000418000002700500030B3132000400812086",
INIT_01 => X"214009C21838284D042100000212026840000000180800080200080040510204",
INIT_02 => X"1021004000900110000006100088503000240800014400004808000000122160",
INIT_03 => X"0002004019110214044A82000121400C86000000000000860188008448400002",
INIT_04 => X"000402800031200A0000090214100889A5000000490090104800000224000400",
INIT_05 => X"10C025204289981000A820500344010428008500010080080909304040202004",
INIT_06 => X"8000440003280000340010208C04003420600000C6180810000C490703200010",
INIT_07 => X"130002000028000890240980A809012001020050000009F08004082640000082",
INIT_08 => X"20100402C4201041310041010008801201480200051023090024811008090A1A",
INIT_09 => X"0100001001248100308214528148A48008000008100004590711C04034000083",
INIT_0A => X"10804000801210140001C0103001088845010482004000008420041020008900",
INIT_0B => X"0004404002004400448000480004800048000480004800048000440022400200",
INIT_0C => X"880420000880204909004502D100A10C04205424010216010C26800805000004",
INIT_0D => X"8000801100509802082010400400018000488428800004082014000200010000",
INIT_0E => X"8000800A00000207A8BE7B00000200082040808000F07F80008000808000F07F",
INIT_0F => X"0002000402100000404CB1F8FC0000040000808000F07F80008000808000F07F",
INIT_10 => X"3E07800000004004080A000002072C3FCF0000020040804800040007687E3F00",
INIT_11 => X"10800018639EC00020100002C2F9B0000801016001008100000040120CB3067F",
INIT_12 => X"000200020000585EB6000100800030C73D8000402000001FC07FF80001000080",
INIT_13 => X"002EAE1FEC0000040200408000003C547E7B00000100801004000803551F8FC0",
INIT_14 => X"00000000440610C8000A808040000208901B86E568FE0C000000020080100400",
INIT_15 => X"0040100401004090240902449028D0230249850101349A98BAC0481000888810",
INIT_16 => X"0401004010040100401004010240902409024090240902409004010040100401",
INIT_17 => X"4010040100409024090240902409004010040100401004090240902409024090",
INIT_18 => X"543EBC57A10A1E75D6440A889050000000000000000040902409024010040100",
INIT_19 => X"79E79E79E79E79E79E79E79E79E79E79E79E79E7BF3CCD8DF5B2DB2CA4028A0A",
INIT_1A => X"4F87D3E1F4F87D3E1F4F87D3E1F4F87C3E1F0F87C3E1F0F87C3E79E79E79E79E",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000000D3E94F87D3E1F4F87D3E1F4F87D3E1F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"000000087BEAA10F7803DE00FFAEBFFFF0800155FF0000000000000000000000",
INIT_22 => X"7FC2145005155555F780155EFAAAEA8ABAAAFBFDE0055556AA005D0415555080",
INIT_23 => X"7AA974AAAAAA97555F784174BAF7D5555FF552AA8AAA557FC0010F780154105D",
INIT_24 => X"FFAE95555AAFFE8A00552EBFE00F7D17FF45F7FFFFF55AA80155FF087BFDF45F",
INIT_25 => X"5F7D140010552E821EFAAAABDF555555555EFAAFFFDFEFAAAAAAB455D556AA00",
INIT_26 => X"00AAAE955450055421FFFFFBC0010AAD5574BA557FFDFFF5504000AAAAAAA8B5",
INIT_27 => X"A00002EAAAAA082EA8A00002AA8A10F78402155AA8028A00A2D57FF45557BE8A",
INIT_28 => X"0000000000000000000000000000000000000000557BFDFFF55003DFFFF7FBEA",
INIT_29 => X"6AA10410E17555080E000280071E8A00EB8E3FE10F7AEBAFFF080A175D700000",
INIT_2A => X"1C2000FF8A17400557FC015514555757DFF8E175C7A2AAAAA82A2F1FAE105D55",
INIT_2B => X"8A105D71C7BFFF55FFA095482B6A49256DEB84104BAFFD1525FF492EA8AAA557",
INIT_2C => X"AAAAFB7D495F6AA10E3AE90555A2FBE8A38492ABDE10EBDF7AF6DE3FFF8F7DB6",
INIT_2D => X"550E00082B6A0AFB55F7D1420104124821D7AAA0BDF6D415B575D7AAF1FFFD7A",
INIT_2E => X"0B6D578F6D557FFDA00A2AE9756D145B401FFFFFFC7010BEDF524AA5571FDFEF",
INIT_2F => X"FF49003AFEFEBFBEAA001C2EA8A821C2EAAA001C2EA8A00F7800017DA2842FA0",
INIT_30 => X"BEF082E95545000000000000000000000000000000000000000000000497BFAF",
INIT_31 => X"8A10AAD568A00555168A10002E9754D082E820BA08556AA00AAAABFE00F7AEAA",
INIT_32 => X"401E7082EAAABA5D5140010F7AE974105D7BC21555D51575EFFFAA97555A2AEA",
INIT_33 => X"BEABFFAAFBEABFFF7AA80145557BFDF55F78017400F780001FFAA84000AAFFD1",
INIT_34 => X"7BD5555AAD57DF55AAAEBDFEF007BE8A10AAAE8215DA2FFE8ABA082ABFE00AAF",
INIT_35 => X"7FBC00BA55557DFF75D2E82010F7843DF45FFD540000000402145AA843FFFF00",
INIT_36 => X"F780021FFA2803DE10FFD16ABFF5D7BFDE10AAAA975FF5D7BC21EFF7FBD7400F",
INIT_37 => X"0000000000007FE8BFF080028BFFAAFFEAA105D2EAAA005D2AAAA185D2AAAA10",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000400000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(1),               -- Port A write enable input
DIA(0)   => data_write_a(8),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(8),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(1),               -- Port B write enable input
DIB(0)   => data_write_b(8),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(8),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_9_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000B0001800002840002C0000281800000030000000033022000000000002",
INIT_01 => X"8000098218302849180060000C004240413C0A61590001D90213C90008510200",
INIT_02 => X"000008700CB089100002061031200074810448800104008048080080001210E2",
INIT_03 => X"000200140C1822000A028010408100000628000140402080041A100040024840",
INIT_04 => X"41040000000400080002040200080800040000000B08D1055842080604600700",
INIT_05 => X"10002024000020102400010000026104200004000400800C8B0024E4E0010C40",
INIT_06 => X"8000440802280002700800008A840004A0610000C0000810000C590103600810",
INIT_07 => X"538600220028001890240980A80800200102025000000BF08200002440000883",
INIT_08 => X"00000402C220104131102101040810028528820005100003900E884000010007",
INIT_09 => X"00000005E000000600BCA284140200800C834948100004590111824404012080",
INIT_0A => X"04080000901012100A1141005922000245410002008880000032005080000800",
INIT_0B => X"2000020040044010440104401004010440100401044010040104400802008208",
INIT_0C => X"D1A1344420D2E100000808000000000481000000202002400006800825908402",
INIT_0D => X"0500000000109000000000000580008000080000C852240100068D0B4685A342",
INIT_0E => X"0500000A00000000000000000000028000408020000000050000208020000000",
INIT_0F => X"0000304002100020000000000000000900208004000000050000208004000000",
INIT_10 => X"0000000001200000000A00000000000000000000050000480008000000000000",
INIT_11 => X"009F0080000000004807C0200000000012000020000081000000040000000000",
INIT_12 => X"00000048F8000400000002403E0004000000009067E000000000000000000900",
INIT_13 => X"0000000000000000140000CEE001000000000000000A000036AC008000000000",
INIT_14 => X"03210000000400CA81000000619480D4000400000000000000004100000036E8",
INIT_15 => X"A368DA368DA3685A1685A1685A121A11A1419001512490040024001000008019",
INIT_16 => X"1685A1685A1685A1685A1685A368DA368DA368DA368DA368DA368DA368DA368D",
INIT_17 => X"685A1685A168DA368DA368DA368DA368DA368DA368DA3685A1685A1685A1685A",
INIT_18 => X"CCF48DE68A895C38E250080000000000000000000000685A1685A1685A1685A1",
INIT_19 => X"514514514514514514514514514D34D34D34D34D28E10040392482090157344C",
INIT_1A => X"4D268341A0D069349A0D069349A0D068341A0D068341A0D06834514514514514",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000001654D0D069349A0D068341A4D268341A",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"BE8B45002A974AAAA803DFFFAA843DF45FFFFEAABA0000000000000000000000",
INIT_22 => X"AEBDE00AAFBEAABA080000000087BEAA10F7803DE00FFAEBFFFF0800155FFAAF",
INIT_23 => X"AAEA8ABAAAFBFDE0055556AA005D0415555087BFDE00A2FBD7400F7FBFDFFFA2",
INIT_24 => X"005155555557BE8BEF007FFDEAAAAD1555EF0055401FFF7AEAAA10F780155EFA",
INIT_25 => X"0F7AA974AA082E80010A2AAAAA10552AA8AAA557FC0010F780154105D7FC2145",
INIT_26 => X"BA087BFDF45F7AA974AAAAAA97555F784174BAF7D5555FFF780154AA5D2AA8A1",
INIT_27 => X"F45F7FFFFF55AA80155FF080400145FFFBEAABAF7D17FEBAA2AEBDF45002EAAA",
INIT_28 => X"0000000000000000000000000000000000000000AAFFE8A00552EBFE00F7D17F",
INIT_29 => X"BAFFF080A175D7BEF1E8B6D002090482B68E38FC7BE8A3DF7DF7F5E8A9200000",
INIT_2A => X"BD0400FFF5FDFC7B6A0BDE38B6F5E8A92080E000280071E8A00EB8E3FE10F7AE",
INIT_2B => X"AAA8A38FF8E175C7A2AAAAA82A2F1FAE105D556AA10410E175550871FFE00A2F",
INIT_2C => X"F8A17400557FC015514555757D5D71E8BEF147BFAE82A2DB555C71C5B451D7FF",
INIT_2D => X"FF84174BA5D20AAA00E3AA904BA142A87010A2AEADA38492EA8AAA5571C2000F",
INIT_2E => X"AAAA0BFF7D0024ADA921C7BFFF55FFA095482B6A49256DEB84104BAFFD1525FF",
INIT_2F => X"38492ABDE10EBDF7AF6DE3FFF8F7DB68A105D7000400155FFFBEDA82FFD57DEB",
INIT_30 => X"FEFF7D16AA00000000000000000000000000000000000000000000000A2FBE8A",
INIT_31 => X"AA00AAAABFE00F7AEAABEF082E95545F7D568BEF080402000F7AAA8B55FFAABD",
INIT_32 => X"9754D00517DE00A2FFC2000F7D17FF55FF803FEAAFFD16AA00082E820BA08556",
INIT_33 => X"FD55555D7FD5555FFAAA8AAAFFAA97555A2AEA8A10AAD568A00555168A10002E",
INIT_34 => X"2EAAABA5D5140010F7AE974105D7BC21555D51575EF555568BEF5D7FE8A10AAF",
INIT_35 => X"A84000AAFFD1401E7FF80174AA5D0028A00AAAE800AA552A97400A2AEBDEAA08",
INIT_36 => X"F7FBFFE00FFD17FEAAA2803DFEF08043FE00557BFDF55F78017400F780001FFA",
INIT_37 => X"0000000000A2FFE8ABA082ABFE00AAFBEABFFAAFBEABFFF7AA80145080002145",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000800000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(1),               -- Port A write enable input
DIA(0)   => data_write_a(9),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(9),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(1),               -- Port B write enable input
DIB(0)   => data_write_b(9),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(9),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_10_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000B0001800002840002C0000281800020030000000033022000000180006",
INIT_01 => X"000008000000004C002000000010026840000000080000080200000000110200",
INIT_02 => X"0000004000800110000006100000003000040800010400004808000000120060",
INIT_03 => X"000200000810020000020000400100000600000000400000001A000040004800",
INIT_04 => X"0004000000000008000200020000000004000000080010004000000200000000",
INIT_05 => X"1000202000011010000000000000010520000400000080000000200000200004",
INIT_06 => X"80004408022800023000000088040004A061000040000810000C490103600000",
INIT_07 => X"120420020028000890240980A808002001020050000009F08000002440000082",
INIT_08 => X"00000402C0201051311001000000020201080200440400000000800000000000",
INIT_09 => X"0000105808000000000000000000008000008088100004590111800004000000",
INIT_0A => X"00804000801210440003C1411008800045000002000014000040009002800000",
INIT_0B => X"0400200000000000000004000040000000000000040000400000000000000221",
INIT_0C => X"0100802000000000000002802000000400100000000002000026000840011400",
INIT_0D => X"0500000000409002082010400400008000400008002044082000081004080204",
INIT_0E => X"0500000200000000000000000000028000400000000000050000200000000000",
INIT_0F => X"0000304002000000000000000000000900200000000000050000200000000000",
INIT_10 => X"0000000001200000000200000000000000000000050000400000000000000000",
INIT_11 => X"0082000000000000480080000000000012000101000080000000000000000000",
INIT_12 => X"0000004810000000000002400400000000000090400000000000000000000940",
INIT_13 => X"0000000000000000150000C00000000000000000000A40001400000000000000",
INIT_14 => X"02000000002400C2810000006000000000000000000000000000410040001400",
INIT_15 => X"020080200802008020080200800800220200840001309A08A848001000008000",
INIT_16 => X"0000000000000000000000000200802008020080200802008020080200802008",
INIT_17 => X"0080200802000000000000000000000000000000000000000000000000000000",
INIT_18 => X"940FE0D397124355520542821010000000000000000000802008020080200802",
INIT_19 => X"28A28A28A28A28A28A28A28A28A28A28A28A28A29554199854514514F546890A",
INIT_1A => X"32994CA6532995CAE572B94CA6532994CA6532994CA6532994CA28A28A28A28A",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000001867172B94CA6532994CA6572B95CAE5",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FC2155F7D155545AA80001EFAAFBEAB45557FFDE100000000000000000000000",
INIT_22 => X"FBE8BFFF78402155AAFBE8B45002A974AAAA803DFFFAA843DF45FFFFEAABA007",
INIT_23 => X"87BEAA10F7803DE00FFAEBFFFF0800155FF00042AB55FFD168B55AA8000010FF",
INIT_24 => X"AAFBEAABAA2FFD741055003DFEFF7AA801FFAAD16AABA002ABDE100800000000",
INIT_25 => X"FF7FBC0145F78028A00A2D142155087BFDE00A2FBD7400F7FBFDFFFA2AEBDE00",
INIT_26 => X"BAF780155EFAAAEA8ABAAAFBFDE0055556AA005D0415555007FD74105555555E",
INIT_27 => X"5EF0055401FFF7AEAAA105D042ABFF5D556AB55AAD168ABA002A975FFF7AEBDE",
INIT_28 => X"0000000000000000000000000000000000000000557BE8BEF007FFDEAAAAD155",
INIT_29 => X"3DF7DF7F5E8A92007BC217DEBDB55555AA8E071D7AAFBEFB455D71F8E0000000",
INIT_2A => X"B6DB55BE8E05000EBFFE8BC7E38E07145BEF1E8B6D002090482B68E38FC7BE8A",
INIT_2B => X"2EB8E00080E000280071E8A00EB8E3FE10F7AEBAFFF080A175D700042AB7DEBD",
INIT_2C => X"FF5FDFC7B6A0BDE38B6F5E8A92B6FBD5410490A3DFD7F7A4821D7A2D16FA8214",
INIT_2D => X"0071D54104951555D7EBF5C5155E3842AA00BED1421450871FFE00A2FBD0400F",
INIT_2E => X"20820955EFE3AEBDEAAFF8E175C7A2AAAAA82A2F1FAE105D556AA10410E17555",
INIT_2F => X"EF147BFAE82A2DB555C71C5B451D7FFAAA8A38410E2ABD749516FB55BED16FA8",
INIT_30 => X"F455D556AA000000000000000000000000000000000000000000000005D71E8B",
INIT_31 => X"2000F7AAA8B55FFAABDFEFF7D16AA00087FC01EFA2FFD7545AAAE97555A2FBFD",
INIT_32 => X"9554500042ABFFA2FFFFF45F7AE97400AAFFE8B45AAAA95545F7D568BEF08040",
INIT_33 => X"400155A2D57FE00552EA8A00082E820BA08556AA00AAAABFE00F7AEAABEF082E",
INIT_34 => X"517DE00A2FFC2000F7D17FF55FF803FEAAFFD16AA00FFFBD5400082EBFF45F78",
INIT_35 => X"55168A10002E9754D085155410085557555AAD557555A2802AA10FFD54214500",
INIT_36 => X"08557DF55F7D17FE000804155FFAAAABDEAAFFAA97555A2AEA8A10AAD568A005",
INIT_37 => X"0000000000555568BEF5D7FE8A10AAFFD55555D7FD5555FFAAA8AAA002AAAB45",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000008FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(1),               -- Port A write enable input
DIA(0)   => data_write_a(10),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(10),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(1),               -- Port B write enable input
DIB(0)   => data_write_b(10),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(10),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_11_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10180B05A0010402840602C2D001019000000300000000330A20080EC180002",
INIT_01 => X"AB400986B830284D1820E0000C3642484000000008000008820009080A512220",
INIT_02 => X"102A68440080011000000618062AD03502640800010410424908136019920868",
INIT_03 => X"004A0846191B22120642000442C110044600000101E9225CDC9A10844A9A4842",
INIT_04 => X"0094024000250808800216021138000B848000000800100040000102A0600200",
INIT_05 => X"7E4024242008A8102CA88A44010401042200444000888000000028000002A002",
INIT_06 => X"8088445712280000B18812288E0400253855200045C86810000C5B0503286A28",
INIT_07 => X"10008822A028004880200A80880208200122006C000015F0C20408264902C840",
INIT_08 => X"9390040280241041D1754100000018108728820024002B3A01A89540080824C8",
INIT_09 => X"A1001C41A1348498B080801010000080D00301081000045B0511D28D94012339",
INIT_0A => X"44080000901012428003414158230CBA4576708241C010908040341322008000",
INIT_0B => X"040464D280144050C72A0872A0C72A0872A0C72A0C72A0872A0C595043950421",
INIT_0C => X"0804001400000820110A42822204880CD81040442900021704E6000800001D54",
INIT_0D => X"80C62D0500409002082010404580018000404012004004192C10000000000000",
INIT_0E => X"80C62D5803161C526DB40506C120A806ABB0D808CC334A80A54B70D408CC32D2",
INIT_0F => X"2B5144D0DD903C54916D15458C0513005570D408CC334A80A54B70D808CC32D2",
INIT_10 => X"52148C4DB05621E363F813961C20EDA944016558C2347A080B10D8DD6422AA10",
INIT_11 => X"1880144D3345C65593800319C18BD1ECA1C9010112566F10AC4183C340DAE02D",
INIT_12 => X"5810503000633830DE3C2C9C00289A66AA8DE50E0800360614AC281430890600",
INIT_13 => X"0CD2A9CEA8199B6B082B55900314140365320485C4F00AD544407241C175C402",
INIT_14 => X"0000074044C4801832701A89D20A38093631425969020855A281844E00540404",
INIT_15 => X"0000000000000000000000000020C00200088101513492101280401000400200",
INIT_16 => X"2008020080200802008020080000000000000000000000000000000000000000",
INIT_17 => X"0080200802008020080200802008020080200802008020080200802008020080",
INIT_18 => X"804180C0B10A4210420140028400000000000000000000802008020080200802",
INIT_19 => X"000000000000000000000000000820820820820801C414947000000055062608",
INIT_1A => X"0000000004020000000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000001F87E000000000000010080000000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"ABDF5508557DF45002ABDFFFF7803DE10AA80000AA0000000000000000000000",
INIT_22 => X"FFE8A10A28000000007FC2155F7D155545AA80001EFAAFBEAB45557FFDE10082",
INIT_23 => X"02A974AAAA803DFFFAA843DF45FFFFEAABAA2AEBFF45FFAEBFEAA002A801FFF7",
INIT_24 => X"F78402155AAD155555A28428BFF002ABDE00A2AABFE10082ABFFEFAAFBE8B450",
INIT_25 => X"0002A80010A2842AAAA007BFFF4500042AB55FFD168B55AA8000010FFFBE8BFF",
INIT_26 => X"00080000000087BEAA10F7803DE00FFAEBFFFF0800155FF00557FF45557FC201",
INIT_27 => X"1FFAAD16AABA002ABDE10A2D168A10A284021FF5D00154BAF7FBE8BEFFFD5400",
INIT_28 => X"0000000000000000000000000000000000000000A2FFD741055003DFEFF7AA80",
INIT_29 => X"EFB455D71F8E00002EBDF6D005B78F7D142ABDFC7F78E3FE28B684070AA00000",
INIT_2A => X"0BDEAA1C2A801C7E3FFEFA10B68407038007BC217DEBDB55555AA8E071D7AAFB",
INIT_2B => X"20B8FEFBEF1E8B6D002090482B68E38FC7BE8A3DF7DF7F5E8A92BEAEBFF7DEBA",
INIT_2C => X"E8E05000EBFFE8BC7E38E07145B6D15756DA28A28BFF082ABAE10B6AAB8E2808",
INIT_2D => X"08517DF7D497BC5028142A87000A28A2AA92007FF8F7D00042AB7DEBDB6DB55B",
INIT_2E => X"2FFFFEFBC7E3DF42028080E000280071E8A00EB8E3FE10F7AEBAFFF080A175D7",
INIT_2F => X"10490A3DFD7F7A4821D7A2D16FA82142EB8E00B6DB6AA28A280001FF5D0A1048",
INIT_30 => X"EAAF784154BA000000000000000000000000000000000000000000000B6FBD54",
INIT_31 => X"7545AAAE97555A2FBFDF455D556AA00082EBFFEF007BE8BFF5D2ABDF55F7AABD",
INIT_32 => X"6AA00FFAEBFFEFAA803DEBA5D2E82155A2FBFDE00FF84154BA087FC01EFA2FFD",
INIT_33 => X"AAAA00FFAAA8AAA080028BFFF7D568BEF080402000F7AAA8B55FFAABDFEFF7D1",
INIT_34 => X"042ABFFA2FFFFF45F7AE97400AAFFE8B45AAAA95545F7D5555FFAAAAA8BFF002",
INIT_35 => X"7AEAABEF082E9554508557DFFF007BD54BA5D2E95400A2AEA8A00007FEABFF00",
INIT_36 => X"AA80001FF5D2E82000F7FFFFF45AAFFC20BA082E820BA08556AA00AAAABFE00F",
INIT_37 => X"0000000000FFFBD5400082EBFF45F78400155A2D57FE00552EA8A00FFFFE8AAA",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000800000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(1),               -- Port A write enable input
DIA(0)   => data_write_a(11),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(11),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(1),               -- Port B write enable input
DIB(0)   => data_write_b(11),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(11),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_12_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A500C4B01BC0268A6940312C0DE045196A831A300500032B333287E4FC812006",
INIT_01 => X"AF400D869830E84D5823E0000C1742484000000008000008820009280A553235",
INIT_02 => X"502A7144008001100000171C022BD13412762A000586235ECC09C8423B960866",
INIT_03 => X"31863846191BA218064204000281200406A10843010022DEDF0852944A9C014A",
INIT_04 => X"0014030000250409000014821038080B840000400800102040000302F0600233",
INIT_05 => X"7FC034348008A8102CA88F48010601042400048000188000000938000002E088",
INIT_06 => X"9CC96CC6F63A5001F12B56A0AC8601F47AC06400D1F80C10020C493F03343A38",
INIT_07 => X"1020002030280098A12048908A16BA311177124C000003F08A94282E5C262861",
INIT_08 => X"827A0602902A10491165E10000049010C52882008600A73A01E8974008092CF8",
INIT_09 => X"47000001A1248008F000000000000080000F010C100204593F11A6CDF48023BF",
INIT_0A => X"040000208010120ACA01400058010CBA4D277C86CCE802B380003C1360008000",
INIT_0B => X"011C46D3C7BC1EF083AF0C3AF083AF083AF0C3AF083AF083AF0C1D7861D78400",
INIT_0C => X"08040014C9001AE91D17E50AD79FEFC87C2154745F82131FFCCE00080000095E",
INIT_0D => X"807BF7118180984004000803D40001880001001400C005031010000000000000",
INIT_0E => X"807BF76A109C944B5891BF06C5EEB14FCBF0D90076D61C807BF7D0D80876D49C",
INIT_0F => X"6DE38EB9FB10350C00A99F7CA80757365E50D80876D61C807BF7D0D90076D49C",
INIT_10 => X"841BCC69A0D8C6F7F0AA001C943A65756A0976EB5A7E7FC8951018186334F311",
INIT_11 => X"D5A014481991C6A737D80211912970CDCDD1864116D6C7080651CB4661F33615",
INIT_12 => X"349E929300423224AE19B9BEC0289033238D4E6EA805892946A9B011A7B152CF",
INIT_13 => X"6244CD7AC01CAAA56B3E6D9001068715D64006D2A961CF9B44512A2504532182",
INIT_14 => X"00000439FDC25C58067A9FAB46095A0B5289A0282D2E1444ACB12A17CF9B4414",
INIT_15 => X"0000000000000000000000040026C00000288401513492909280401000F70A00",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"088881360A95090CB05442029010000000000000000000000000000000000000",
INIT_19 => X"1041041041041041041041041049249249249249200100002D4514510051B946",
INIT_1A => X"592C964B2592C964B2592C964B2592C86432190C86432190C864104104104104",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000002007F592C964B2592C964B2592C964B2",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"43FE0008557DFFF0800020105D557FEAA00557DE100000000000000000000000",
INIT_22 => X"557DFFFF7AA80000082ABDF5508557DF45002ABDFFFF7803DE10AA80000AAAA8",
INIT_23 => X"7D155545AA80001EFAAFBEAB45557FFDE10AAD5420000051555FFA2AA8200000",
INIT_24 => X"A28000000A2D155410F7FFFFEBA08003FE00082AA8AAAAAFFC00BA007FC2155F",
INIT_25 => X"0A2AABFE1055516ABEF5D517DEAAA2AEBFF45FFAEBFEAA002A801FFF7FFE8A10",
INIT_26 => X"55AAFBE8B45002A974AAAA803DFFFAA843DF45FFFFEAABA000028A105D2ABFE1",
INIT_27 => X"E00A2AABFE10082ABFFEF085542000000417555002A820AA08557DFFFF7AA821",
INIT_28 => X"0000000000000000000000000000000000000000AAD155555A28428BFF002ABD",
INIT_29 => X"3FE28B684070AABE803AE38145B78FD7000005010495B7AE921C517DE1000000",
INIT_2A => X"B505FFB6A487000005F7AFD7F7A482038002EBDF6D005B78F7D142ABDFC7F78E",
INIT_2B => X"F5C2082007BC217DEBDB55555AA8E071D7AAFBEFB455D71F8E00BED547038145",
INIT_2C => X"C2A801C7E3FFEFA10B68407038B6D550428FFF1FDE821C003FE001C2EAAAAAB6",
INIT_2D => X"00002FA285D20BDE28A2A4B8E10555B68BEF5D517DEAABEAEBFF7DEBA0BDEAA1",
INIT_2E => X"2005F7DFD7F7A482155BEF1E8B6D002090482B68E38FC7BE8A3DF7DF7F5E8A92",
INIT_2F => X"6DA28A28BFF082ABAE10B6AAB8E280820B8FEF085F4703814001055514208208",
INIT_30 => X"A0055517DE00000000000000000000000000000000000000000000000B6D1575",
INIT_31 => X"8BFF5D2ABDF55F7AABDEAAF784154BAF7802AABA5D7FEAB45080015410007FEA",
INIT_32 => X"6AA00F7D1554BA5D7BC01FFFF8015410007FEAB45F780020BA082EBFFEF007BE",
INIT_33 => X"43FE10552EAAAAAFFD140000087FC01EFA2FFD7545AAAE97555A2FBFDF455D55",
INIT_34 => X"AEBFFEFAA803DEBA5D2E82155A2FBFDE00FF84154BAF7D1400BAFFD57FE005D0",
INIT_35 => X"FAABDFEFF7D16AA0008003FEBA55003DEBAA28428A105D7FEABEF55557DEBAFF",
INIT_36 => X"550402145550000010087FFFF45F78402145F7D568BEF080402000F7AAA8B55F",
INIT_37 => X"0000000000F7D5555FFAAAAA8BFF002AAAA00FFAAA8AAA080028BFF087BD54AA",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000000FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(1),               -- Port A write enable input
DIA(0)   => data_write_a(12),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(12),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(1),               -- Port B write enable input
DIB(0)   => data_write_b(12),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(12),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_13_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10110A0441812402840402822007818000E00700000000330A3000000008042",
INIT_01 => X"A1400984B830C848180260000C0042604001000008220008A200100802110200",
INIT_02 => X"10A00860009141100000C6180C285035000E0800010431004908135980120C60",
INIT_03 => X"004E20441910221B06420C85D5013804060000000040324C441A108468024842",
INIT_04 => X"0184034010250089C00EA8021938325B04800002091090014880080200000900",
INIT_05 => X"18002424B008881024A8004E01040104270004E0000080090500604840000481",
INIT_06 => X"80004414022A2490B00A142C8C840005794540015E006810001C4B01032C7E20",
INIT_07 => X"510200028028004880280A808816002101022468000011F082040A264006C000",
INIT_08 => X"D2B00402B220104B531001000008001041080200B660E30B200C8040080A9206",
INIT_09 => X"A1000809A93484D21000000000000080C90391881000145B0111A30404015000",
INIT_0A => X"000000008010102A82014100101118BA4510008241480290882400900000A000",
INIT_0B => X"0284484000000000400000000040000000000000040000000000000020000000",
INIT_0C => X"A944AA2000A02000212800020000000D80004084A0000390002E001843210400",
INIT_0D => X"859C1881A04090000000000021800180010341179065441356150A1285094284",
INIT_0E => X"859C188810C65A72A617520252781EA02520D589B9A260859C1840DD81B9A0E0",
INIT_0F => X"0E71F1052D942748C19484E39442D15961C0DD81B9A260859C1840D589B9A0E0",
INIT_10 => X"E60605C0C12CBD400B0810C65A61AA459D0047398500D5889D26907356533C00",
INIT_11 => X"8F60CA1562094650CA28398A42C051E0332181010109294C8E1160CB8C80A561",
INIT_12 => X"2645056D073148580A3C065141942AC4128CA199180C5232575138094450AD0A",
INIT_13 => X"84CA93A2FC008962142B17301A9A1A5196A80245208E0AC5C853C8028163B8C0",
INIT_14 => X"0240034000E4DC8A84000014982372011FC1E475F0F0084A3961F5A80AC5C816",
INIT_15 => X"4250942509425094250942509428D421420882020120981812C8403000088212",
INIT_16 => X"2509425094250942509425094250942509425094250942509425094250942509",
INIT_17 => X"5094250942509425094250942509425094250942509425094250942509425094",
INIT_18 => X"FF3F7DF7FF3E9F7DF7E24502A800000000000000000050942509425094250942",
INIT_19 => X"EBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBF7DFDFDDD555555F7EFBBEE",
INIT_1A => X"7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAEBAEBAEBAEBA",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000000007F7EBF5FAFD7EBF5FAFD7EBF5FAFD",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5554BA087FFFF55557BD54AAF7FBC01FFA2802ABEF0000000000000000000000",
INIT_22 => X"2E80155AA802AB45AA843FE0008557DFFF0800020105D557FEAA00557DE10AAD",
INIT_23 => X"8557DF45002ABDFFFF7803DE10AA80000AA087BD75EF087FFFFEF557BEAB4555",
INIT_24 => X"F7AA80000AAD1420AA087BD7555FFD168AAAFFAE820AA5D5557555082ABDF550",
INIT_25 => X"5FFD157555085140010F7AEAABFFAAD5420000051555FFA2AA8200000557DFFF",
INIT_26 => X"45007FC2155F7D155545AA80001EFAAFBEAB45557FFDE10AAAEA8BFFA2FBD754",
INIT_27 => X"E00082AA8AAAAAFFC00BA00002AAAAF7D5574BA557BE8A10A284154BAFFAAAAB",
INIT_28 => X"0000000000000000000000000000000000000000A2D155410F7FFFFEBA08003F",
INIT_29 => X"7AE921C517DE10A2DB50482147FFAF554971D0492E3F1C71C7BE8A2ABD700000",
INIT_2A => X"FFAFD7497BE8B5555208217DBE8A2AB45BE803AE38145B78FD7000005010495B",
INIT_2B => X"5F5056D002EBDF6D005B78F7D142ABDFC7F78E3FE28B684070AA1C71D25D7007",
INIT_2C => X"6A487000005F7AFD7F7A482038AADF47092147FD257DFFD568A82FFA4870BA55",
INIT_2D => X"A2A0ADBC7A2FFD257DE3DF52555085142000FFAAAFBFFBED547038145B505FFB",
INIT_2E => X"0B680124BAFFAAAFB45007BC217DEBDB55555AA8E071D7AAFBEFB455D71F8E00",
INIT_2F => X"28FFF1FDE821C003FE001C2EAAAAAB6F5C20821C002AA92FFDF574824171EAA1",
INIT_30 => X"545F7AEA8B55000000000000000000000000000000000000000000000B6D5504",
INIT_31 => X"AB45080015410007FEAA0055517DE00A2FFC00105D7BE8B55085142010AAD157",
INIT_32 => X"154BA5D5140145007BE8B55087BEAB555D04001EFF7AAA8B55F7802AABA5D7FE",
INIT_33 => X"16AA10FF80174AA557FC21EF082EBFFEF007BE8BFF5D2ABDF55F7AABDEAAF784",
INIT_34 => X"D1554BA5D7BC01FFFF8015410007FEAB45F780020BAA2FFD54105D7FC21EFFFD",
INIT_35 => X"2FBFDF455D556AA00A2803FF45AAFFC21EFAAFBC0155085540000FFAEBFFEFF7",
INIT_36 => X"F7FBD5410085568A10FF80020AAFFAABFF55087FC01EFA2FFD7545AAAE97555A",
INIT_37 => X"0000000000F7D1400BAFFD57FE005D043FE10552EAAAAAFFD1400005D042AA00",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000CFFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(1),               -- Port A write enable input
DIA(0)   => data_write_a(13),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(13),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(1),               -- Port B write enable input
DIB(0)   => data_write_b(13),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(13),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_14_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10020A000180000284008280000281800000030000000033022000000580002",
INIT_01 => X"A140098018300848184860000C20C24040000000084000084200000000110200",
INIT_02 => X"1020006000900110000006102028503400040800010400204908012018120E64",
INIT_03 => X"000200441910221006420000400100040600000000E9E401209A108448004842",
INIT_04 => X"0004020000250008000200021038000804000000090090004800080200000000",
INIT_05 => X"500024240008881024A800400104010420000400000080080100204040000000",
INIT_06 => X"8000440102282015B10A10288E0400042345400040006810000C5901033D7880",
INIT_07 => X"1100000200280048802008828812002001220064000005F1C2850A2649204070",
INIT_08 => X"00B00402802010411110010000080010010802000400230B000C804008080002",
INIT_09 => X"01000009A92480001000000000000080C8038188100004590111B68404010000",
INIT_0A => X"0000000080101000000141001001088A45000082400000008020009000008000",
INIT_0B => X"0004404000000000400004000000000000004000000000000004000000000000",
INIT_0C => X"8904A0200080200001080002000000088000400420000200002E000841010400",
INIT_0D => X"0500000C80409000000000000000018000000000806044010014081204090204",
INIT_0E => X"0500005813A0210D072E8D012001028402908004000587050000108004000707",
INIT_0F => X"9004300044900812386A280E5800088980108020000587050000108020000707",
INIT_10 => X"DE00482E19E30002007813A02096038AE200880405200308828062A68C0BC700",
INIT_11 => X"00000E5A08E6000048001292B83280001208A1011004011060049A1C59192055",
INIT_12 => X"492060480256530650000240001DB011CC00009000032C4C979E3806180C0900",
INIT_13 => X"5A3433EDE00154181400000007BCBD858F120120541A0000000033757465B2C0",
INIT_14 => X"02002C000024008A84001A0902000422E3E99681004802115652594000000001",
INIT_15 => X"0240902409024090240902409028D021020880000120901812C8401000000210",
INIT_16 => X"2409024090240902409024090240902409024090240902409024090240902409",
INIT_17 => X"4090240902409024090240902409024090240902409024090240902409024090",
INIT_18 => X"5C8FF0F7BE9D5F7DF65040028000000000000000000040902409024090240902",
INIT_19 => X"79E79E79E79E79E79E79E79E79E79E79E79E79E7BF7DDDDDFCF3CF3DF5579B4E",
INIT_1A => X"3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE79E79E79E79E",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000003FF803F9FCFE7F3F9FCFE7F3F9FCFE7F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"BE8B55A2AE80000F7D5555555D2AAAABAAAD1420BA0000000000000000000000",
INIT_22 => X"00155EF0804155EFAAD5554BA087FFFF55557BD54AAF7FBC01FFA2802ABEFA2F",
INIT_23 => X"8557DFFF0800020105D557FEAA00557DE10A2AA801FFA28402000AAAE9554555",
INIT_24 => X"AA802AB4500516AA00A2AE800BAFFFFC20BAF7AEA8B45080417400AA843FE000",
INIT_25 => X"0A2843FEBAFFFBD7410A2D168BFF087BD75EF087FFFFEF557BEAB45552E80155",
INIT_26 => X"AA082ABDF5508557DF45002ABDFFFF7803DE10AA80000AA005568ABAA2840201",
INIT_27 => X"AAAFFAE820AA5D5557555002E80155A280000005D7FFDF4555517DFEF00043FE",
INIT_28 => X"0000000000000000000000000000000000000000AAD1420AA087BD7555FFD168",
INIT_29 => X"C71C7BE8A2ABD7A2FFEDB55B6A080038E3DB50555412AA8ABAAADB4009200000",
INIT_2A => X"402038AAAA955554900105FF0800175D7A2DB50482147FFAF554971D0492E3F1",
INIT_2B => X"0A12410BE803AE38145B78FD7000005010495B7AE921C517DE10A2AE851FFB68",
INIT_2C => X"97BE8B5555208217DBE8A2AB451C556FA00A2A0800BAE3F1C0092EBAAADB6D08",
INIT_2D => X"00516DABAA28402038B6803DE82F7F5D5410A2D568BC71C71D25D7007FFAFD74",
INIT_2E => X"55D5F78FD7000E3FEAA002EBDF6D005B78F7D142ABDFC7F78E3FE28B684070AA",
INIT_2F => X"92147FD257DFFD568A82FFA4870BA555F5056D002A80155B680000105D7FF8F4",
INIT_30 => X"AAAAAFFC2000000000000000000000000000000000000000000000000AADF470",
INIT_31 => X"8B55085142010AAD157545F7AEA8B55A2FBFFF55FF84000AAAAFBC0145002AA8",
INIT_32 => X"7DE00A2AA955FFFF80020BAAAAA975450800001EF080417555A2FFC00105D7BE",
INIT_33 => X"140000A2AEBFFEF082A82010F7802AABA5D7FEAB45080015410007FEAA005551",
INIT_34 => X"5140145007BE8B55087BEAB555D04001EFF7AAA8B555D557FE00A280020BAAAD",
INIT_35 => X"7AABDEAAF784154BA08557FEAAA284000AAFF803DE00FFD557400AAD56AB455D",
INIT_36 => X"F780020105D7BEAB45557BE8B45082EBFEBA082EBFFEF007BE8BFF5D2ABDF55F",
INIT_37 => X"0000000000A2FFD54105D7FC21EFFFD16AA10FF80174AA557FC21EF082A80145",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000000FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(1),               -- Port A write enable input
DIA(0)   => data_write_a(14),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(14),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(1),               -- Port B write enable input
DIB(0)   => data_write_b(14),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(14),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_15_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000A000000000284000280000001800020030000000033022000000180002",
INIT_01 => X"A140098018300848180060000C00424040000000080000080200000000110200",
INIT_02 => X"102100400C8011100000061000A8503401044880010430004808000180122378",
INIT_03 => X"000200541D102210064200000045000546080000400020000008108448400042",
INIT_04 => X"8094020000254C880000028A1018000844000000880013504000002600000000",
INIT_05 => X"10002424000AA81024A82040010C61062001440002988000000024808001004B",
INIT_06 => X"80004400022A00003C8912248E0400042854400040006810000C4901032B1800",
INIT_07 => X"50200000B0280048A0280A828801002101020040000005F38204082640000000",
INIT_08 => X"01F00402802610411100110000000010010802000400230A0008884008080004",
INIT_09 => X"01000001A12481041000000000000080C0030108100004590111820404000000",
INIT_0A => X"0000000080101000004140001001088A45000082000000008000001080008000",
INIT_0B => X"0004404000000000400004000040000400000000000000000004000020000200",
INIT_0C => X"0804000020024100012808020000000981004004A0200310000C000800000000",
INIT_0D => X"0000001180009000000000002100018000000000004004010010000000000000",
INIT_0E => X"00000008000002000000000000000000000080A40000000000000080A4000000",
INIT_0F => X"00000000001000204800000000000000000080A40000000000000080A4000000",
INIT_10 => X"000000000000000000080000020000000000000000000008000C020000000000",
INIT_11 => X"000000824000000000000020220000000001800100020300000004003420480A",
INIT_12 => X"0000000000040440000000000001048000000000000000100800400000000000",
INIT_13 => X"000800000000000000000000000100C220050000000000000000008220884400",
INIT_14 => X"000000000000000830000000000000000016101C5C1400000000000000000000",
INIT_15 => X"0000000000000000000000000020C00000088000012090101280401000000200",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000040028000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"000010082A954BA00003DFEF085155400F78428BEF0000000000000000000000",
INIT_22 => X"8015400FF84001EFA2FBE8B55A2AE80000F7D5555555D2AAAABAAAD1420BAFF8",
INIT_23 => X"87FFFF55557BD54AAF7FBC01FFA2802ABEFF7AE95555A2FBE8BEFA2843DE00AA",
INIT_24 => X"0804155EFFFFBE8BFF0800174AA557BFDE10A2FBEAB45F7D56AABAAAD5554BA0",
INIT_25 => X"5FFD568BEF087FE8A1055003FE00A2AA801FFA28402000AAAE955455500155EF",
INIT_26 => X"45AA843FE0008557DFFF0800020105D557FEAA00557DE10F7D1574AAA2D16AB5",
INIT_27 => X"0BAF7AEA8B45080417400FFFFC2145080015400AA802AA00AAAE800BA5D00155",
INIT_28 => X"000000000000000000000000000000000000000000516AA00A2AE800BAFFFFC2",
INIT_29 => X"A8ABAAADB40092E38E070280024904AA1C0438FD7005150438F78A2DBFF00000",
INIT_2A => X"FE8BC7BE8E38E10A28017400E38A051FFA2FFEDB55B6A080038E3DB50555412A",
INIT_2B => X"D16AABAA2DB50482147FFAF554971D0492E3F1C71C7BE8A2ABD7E3AA9257DA2F",
INIT_2C => X"AAA955554900105FF0800175D7E3FFEFBD70000124AA557FFDE10A2FBEDB6DF7",
INIT_2D => X"FFDF50482A2DB6AB45FFD56DBD7087BEAA38410038E38A2AE851FFB68402038A",
INIT_2E => X"0AAA085082550A1057DBE803AE38145B78FD7000005010495B7AE921C517DE10",
INIT_2F => X"00A2A0800BAE3F1C0092EBAAADB6D080A12410FFF1C017D140410400BE8E28A1",
INIT_30 => X"0AAF7AEBDFEF0000000000000000000000000000000000000000000001C556FA",
INIT_31 => X"00AAAAFBC0145002AA8AAAAAFFC2000AAAA974AA0800020BA550028B55085540",
INIT_32 => X"A8B55AAAE821EFAAFBEAB55F7AAA8A00AA8417400AAAE975EFA2FBFFF55FF840",
INIT_33 => X"BFFE10A2FFFFFEFF7D568ABAA2FFC00105D7BE8B55085142010AAD157545F7AE",
INIT_34 => X"AA955FFFF80020BAAAAA975450800001EF080417555AAFFFDF450804020AA557",
INIT_35 => X"07FEAA0055517DE00FFFBC2000AAFBE8B55F7D17DF45007FE8AAA08002AAAAA2",
INIT_36 => X"5D0000010F7AAA8A10AA8017400552A801EFF7802AABA5D7FEAB450800154100",
INIT_37 => X"00000000005D557FE00A280020BAAAD140000A2AEBFFEF082A82010FFD5421EF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000C00000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(1),               -- Port A write enable input
DIA(0)   => data_write_a(15),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(15),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(1),               -- Port B write enable input
DIB(0)   => data_write_b(15),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(15),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_16_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"DA22C618B1000482B688B186588884862A400438255FC38381441205BA803003",
INIT_01 => X"264AC80028404C211203A952A90341080B173340412000E1005D628000820484",
INIT_02 => X"400034C206C405000001A48202084004003008255040826EE008B440200E2042",
INIT_03 => X"A459C1240181AB20AD27315B7F1983CA1C900040422A005762010010000C0400",
INIT_04 => X"296E542B6E3A825C15FB385321B4ADFE16AB45FD2C400002E205231201290A28",
INIT_05 => X"B9E5815006028179808C00A0D2152B90707A1E0BD423CAC0000D610000000710",
INIT_06 => X"81F104A1415C292164280081C6AB88742086ACACDE240000A80090CE82A803B9",
INIT_07 => X"400800000ACCAA280940580400A37B8896CA4D000A80C1102A00001C14028009",
INIT_08 => X"0015452880C8D90409A02D965965200100104F2B00822512000000231520A024",
INIT_09 => X"A5AA80018120E00066000000000012C9000A0000D0A80000BF8028E87C1B9927",
INIT_0A => X"00520228080108039501200848002912300208092B940192D1000000000000A8",
INIT_0B => X"03561180063DB4F6110001100011000110001100011000110001080008800080",
INIT_0C => X"080200854409418B02ED0000502A02972000040BB401100010012B4C90000100",
INIT_0D => X"6D061A1F8D60D80820500101244AA8A2AA242E80000009200120000000000000",
INIT_0E => X"6D066210E5001DB4A5B400C7D553847165A99000C6564CDD051DC99000C65555",
INIT_0F => X"21D0C48F254946148107354292673D1F72C99000C6564CDD0565C99000C65555",
INIT_10 => X"952D2058F33225787810F5001D6121A9559224D1FF97D0272F04D89441A56D8A",
INIT_11 => X"6C1C74485B81E31306C71D1093AB8A64811BADC00992180D58033B1172F2A025",
INIT_12 => X"7B86DED8E3A212748F0E0CA638E890B7A8546120C0AFF5B548AC431FB1C7DB07",
INIT_13 => X"EFCE9B26DECA1AD36A2E4F40DF6AAAF260AF88899E8B8B93D12A877178DD0032",
INIT_14 => X"A8009F8B108C80A1021B9A8BB8056662CA1951596800FC01A38D4D4B072B922F",
INIT_15 => X"00000000000000000000000000044000102A0001148442A1108103595580A840",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"4C690DA64C1C4F68A36040000000000000000000000000000000000000000000",
INIT_19 => X"D14D14D14D14D14D14D14D14D14514514514514529E5F87869E79E78558D1154",
INIT_1A => X"3D1E8F47A7D3E9F4FA7D3E9F4FA7D3E9F47A7D1E9F47A7D1E9F4D14D14D14D14",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE000000000000000007D3E9F4FA7D3E8F47A3D1E8F47A",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFEFF7D168B55AAD17FFFF552EBFE00007FC00AA0000000000000000000000",
INIT_22 => X"04000BA552A821FFFF8000010082A954BA00003DFEF085155400F78428BEF087",
INIT_23 => X"2AE80000F7D5555555D2AAAABAAAD1420BA5D2E975EFF7D568BFFFF80175EF00",
INIT_24 => X"FF84001EF0000020AA5D00154005D043FF45555540000082EAABFFA2FBE8B55A",
INIT_25 => X"0087FD74BAAAAEBFFEF557FC00AAF7AE95555A2FBE8BEFA2843DE00AA8015400",
INIT_26 => X"FFAAD5554BA087FFFF55557BD54AAF7FBC01FFA2802ABEF557BEABEF5D041541",
INIT_27 => X"E10A2FBEAB45F7D56AABA082A97545F7D16ABFFFFAABFEAAFF84001FF002A821",
INIT_28 => X"0000000000000000000000000000000000000000FFFBE8BFF0800174AA557BFD",
INIT_29 => X"50438F78A2DBFF0871F8FC7E3D56AB6DBEDB7FFEF552AB8E38087FC209200000",
INIT_2A => X"16ABFFE38E175EF1400000BA412E871FFE38E070280024904AA1C0438FD70051",
INIT_2B => X"2EAFBD7A2FFEDB55B6A080038E3DB50555412AA8ABAAADB400924920925EFF7D",
INIT_2C => X"E8E38E10A28017400E38A051FF0804050BA410A1240055003FF6D5551420101C",
INIT_2D => X"4975EDBC7550E12410087FD74AAB6AABFFC7557FC00BAE3AA9257DA2FFE8BC7B",
INIT_2E => X"AF780051C70824851D7A2DB50482147FFAF554971D0492E3F1C71C7BE8A2ABD7",
INIT_2F => X"D70000124AA557FFDE10A2FBEDB6DF7D16AABA08249756DF7D168BC7F7AABAEA",
INIT_30 => X"AAA007BC0000000000000000000000000000000000000000000000000E3FFEFB",
INIT_31 => X"20BA550028B550855400AAF7AEBDFEF08516AB55A2D16ABEFFFFBFDFFF552AAA",
INIT_32 => X"C20000000021EFF7D568BFFA2AA955FF5D04020AA002A955EFAAAA974AA08000",
INIT_33 => X"03DFEF5D51420005D2ABFF45A2FBFFF55FF84000AAAAFBC0145002AA8AAAAAFF",
INIT_34 => X"AE821EFAAFBEAB55F7AAA8A00AA8417400AAAE975EF0800174BA002E820105D0",
INIT_35 => X"AD157545F7AEA8B5500557DF45552A82000007BD74AAF7AEBDF455D7BC20BAAA",
INIT_36 => X"F7D568B55FFAAAAABAFF8415545000015555A2FFC00105D7BE8B55085142010A",
INIT_37 => X"0000000000AAFFFDF450804020AA557BFFE10A2FFFFFEFF7D568ABA0804155FF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000400000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(2),               -- Port A write enable input
DIA(0)   => data_write_a(16),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(16),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(2),               -- Port B write enable input
DIB(0)   => data_write_b(16),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(16),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_17_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"5284CE4FB7BD2C8994A13392DBD02E14006B82AC7E800D44D3DD2FD5F9B961C0",
INIT_01 => X"F9BA301F7E03FC6793F2199B39FC233C11D93AE6F3BB92B32091DBC339B24542",
INIT_02 => X"1D5FC0C08F040404446965C0607FB8A217C400C33A908078551BD04222186338",
INIT_03 => X"8504930A37F65820CB24111B7F08014A0AB84A52B6D2AFF97C1B5AC757F06D6B",
INIT_04 => X"250834336D1E81500FDB38302292ADFE103B6DBD204037F202042075E2B1D00A",
INIT_05 => X"8F039786062C6CE092F5FE005236781C402A0807B4070670083DC68206D7E6D0",
INIT_06 => X"0CD26803C3582408962C58B183F8AEF42045919B30E085DD2ED57D4EED08CA6A",
INIT_07 => X"700000B30380670B8142500448E3E01E94EF1340A28AC1AC8156044D1400AA00",
INIT_08 => X"009F3A1B0120A1C51DFFC40C30E5F0182D0950190C0810BE00E9A76E4C6FFBE4",
INIT_09 => X"8FCCC200A59BDD2FFE3F3EC7C7DEF207000F00059D2ED56D7EED2ED3C9A867DC",
INIT_0A => X"0617112E46F05D02DD814102F800633F1D0A7CC9AE7A08BFF0001D35682AC0CE",
INIT_0B => X"8A3F06ABD73DBCF4FBCF4FBCF4FBCF4FBCF4FBCF4FBCF4FBCF4FBE7A7DE7A780",
INIT_0C => X"001000974F08518F5AFFC94B533FADA7FDE97D6BFF329E1B50FF99F086000D9E",
INIT_0D => X"F50B018F95EA3DED1652EC0B27E67F419E2E1E8000C0036340B8000000000000",
INIT_0E => X"F50B01C8DF7F96197DB4AFC8C8886AF672A1537F759299F50B03C1537F759199",
INIT_0F => X"6068331C5103E7EF0FBEED6BB6A9412007C1537F759299F50B03C1537F759199",
INIT_10 => X"21F2CD7F252CDABB3CE8CF7F963AB9FD6AD434201AA68B837FFD1F7B7125B68C",
INIT_11 => X"BD055EB6D555CB2949C15BA7270FF256526BBFD55BBE71D79F73C7AC6DB9BF37",
INIT_12 => X"94080BF82B74E4E1FE4ACA4E0ABD6DAAAB965293036FF6B652A99A6026027FBE",
INIT_13 => X"EF5CBA7A43482800FEFAFD06B8CFCCAB7550D0C2022EAEBD438697AD2EBA9168",
INIT_14 => X"AC00A8BBFC8B501CF7A0FED9A548FA19752C4A4EADAE42FCBC38C3B7BEBF42CF",
INIT_15 => X"0000000000000000000000000026E100002F382DBD9ECFE117805F20CFDAAB00",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"09EDCC4052E917114F981800C000000000000000000000000000000000000000",
INIT_19 => X"EBA69AEBA69A69AEBA69AEBA69A69A69A69A69A68698686981D75D7443720030",
INIT_1A => X"46A351A8D068341A0D068341A0D068341A0D46A341A0D46A341A69AEBA69A69A",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE0000000000000000046A351A8D46A351A8D46A351A8D",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFEFF7FBEAB450804001EFAAD57FEAA0000000000000000000000",
INIT_22 => X"51401EF087FD74AA087FFFFEFF7D168B55AAD17FFFF552EBFE00007FC00AA087",
INIT_23 => X"82A954BA00003DFEF085155400F78428BEFAAD168A000004020AA5D7BE8B4500",
INIT_24 => X"552A821FF5D00020BA552A82000552A821555D7FEAB55FF80175EFFF80000100",
INIT_25 => X"FAAFBC01EF5D0015555557BFDEBA5D2E975EFF7D568BFFFF80175EF0004000BA",
INIT_26 => X"BAA2FBE8B55A2AE80000F7D5555555D2AAAABAAAD1420BAFFFFFDF45AAD17FFF",
INIT_27 => X"F45555540000082EAABFF00516AA10552E820BA007FEABEF005555555A2D1554",
INIT_28 => X"00000000000000000000000000000000000000000000020AA5D00154005D043F",
INIT_29 => X"B8E38087FC2092147FFFFFFFFFBFDFC7EBF5E8B550000071EFB6DF7AE9200000",
INIT_2A => X"A07082497FEFB6D1451471EF007BD04920871F8FC7E3D56AB6DBEDB7FFEF552A",
INIT_2B => X"8E175FFE38E070280024904AA1C0438FD7005150438F78A2DBFFBED16AA381C0",
INIT_2C => X"38E175EF1400000BA412E871FF550A00092492A850105D2A80155417BEFB6DEB",
INIT_2D => X"FFF5FFF6DAADF7FFD7B6F1C71EF55001756D5D7BFAEBA4920925EFF7D16ABFFE",
INIT_2E => X"700515556DA2DF50492A2FFEDB55B6A080038E3DB50555412AA8ABAAADB40092",
INIT_2F => X"BA410A1240055003FF6D5551420101C2EAFBD7145B6AA28492487082007FEDBD",
INIT_30 => X"5EFFFFBEAA000000000000000000000000000000000000000000000000804050",
INIT_31 => X"ABEFFFFBFDFFF552AAAAAA007BC0000557FFDFEFF7FBFFF55A2D16AB55000017",
INIT_32 => X"BDFEFF7D568AAA5D2A97410007BFFFFF5551555EF087FC200008516AB55A2D16",
INIT_33 => X"A82155087FFFFEFAAAA975EFAAAA974AA0800020BA550028B550855400AAF7AE",
INIT_34 => X"00021EFF7D568BFFA2AA955FF5D04020AA002A955EF5D2E80010002A954005D2",
INIT_35 => X"02AA8AAAAAFFC2000FFD57DFFFAAFFFDF55FFD1575FF5504175EF5D7FEAAAA00",
INIT_36 => X"000415410007BFFF450051555EFA2FBC0000A2FBFFF55FF84000AAAAFBC01450",
INIT_37 => X"00000000000800174BA002E820105D003DFEF5D51420005D2ABFF45557FE8AAA",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000CFFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(2),               -- Port A write enable input
DIA(0)   => data_write_a(17),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(17),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(2),               -- Port B write enable input
DIB(0)   => data_write_b(17),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(17),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_18_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"69844019080000A21A611406840014122A641074155FC28A2024001001801003",
INIT_01 => X"01067920034004180005E9E3C90360C0041C0181002001602025800008440084",
INIT_02 => X"40AC3CAA22D605200000856E2481902400344A20F802C22054001000021E2379",
INIT_03 => X"A54C23B34C81EB2076471000800981140C010101750D1007E58040102B0E0100",
INIT_04 => X"22660C1C0065003C04040013236E105016A028402D618803EB092B9201490B2A",
INIT_05 => X"B8E080000000005889AC41E04508A99070200E010001C1CA11803850C8000100",
INIT_06 => X"800A4CE301545001F40050216C09950004C2047BCF1C8090C02800C0120886B3",
INIT_07 => X"814A0080064C1F300020080182001A9E02C03400082002700000217294007101",
INIT_08 => X"000117088080990419002D86184A01018030430700802541420440022030041A",
INIT_09 => X"7030C30B885200D274004008080003C32A10A19090C02010E102294406168800",
INIT_0A => X"00602A01880980037109700C04C44C92A88DCC2211E44174112840880000060D",
INIT_0B => X"11C0D95C20C2030A003080030800308003080030800308003080018400184004",
INIT_0C => X"8304E02809832E6021002020404042000F00008400811824AD4007ECD9436261",
INIT_0D => X"0AFCE5D22A82B20000520100C801F8A07E103000A1285C84000418360C1B060D",
INIT_0E => X"0AFCFD8CB17E5B4F045557575E6EFBE3942C1040A41D660AFCE1CC1040A41E66",
INIT_0F => X"8E7FFBB385661C08D1455ABA91E6FF5FDFCC1040A41D660AFCF9CC1040A41E66",
INIT_10 => X"015F82C006C3AF31E64CB17E5A9655017F1FC73FAF1D61B1040294C58AD1FF5F",
INIT_11 => X"B95454005BAA36DCF8E519001BF80DEB3EE2020EA678189C6EC32881F7F75648",
INIT_12 => X"67D7EDFCA320037E81BD77D728A800B7546DBDFF12904747A351145FC53ABF8D",
INIT_13 => X"92B764225C57C97EBE76E1254F0C0D4514A84F5573FE9DBA4A38E247C522CC0E",
INIT_14 => X"BE84370001B6922070440556B15F7FABBC40151D7C747D8220673C3B9DB84B20",
INIT_15 => X"06C1B06C1B06C1B06C1B06C1B0491069068000004060300A005A01183F240014",
INIT_16 => X"6C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B",
INIT_17 => X"C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B0",
INIT_18 => X"B80EE173C2300F7DF16000000000000000000000000041B06C1B06C1B06C1B06",
INIT_19 => X"AAAAAA28A28A28AAAAAAA28A28A28A28A28A28A2910591505C104104B28BBECE",
INIT_1A => X"128944A25128944A25128944A25128944A2552A954AA5128944AAAA28A28A28A",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000128944A25128944A25128944A25",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFDFEF5D2A974BA082E954000000000000000000000000",
INIT_22 => X"0028B55002E82000087FFFFFFFFFFFFFEFF7FBEAB450804001EFAAD57FEAA087",
INIT_23 => X"7D168B55AAD17FFFF552EBFE00007FC00AA087FFFFFFFFFBFDF45AAD568B5508",
INIT_24 => X"087FD74AAAAFFFDF45A2D16AB55F7FFFFFFF00043DE10AA843DE00087FFFFEFF",
INIT_25 => X"A55042ABEF5D7FD75FFAAD540145AAD168A000004020AA5D7BE8B450051401EF",
INIT_26 => X"45FF8000010082A954BA00003DFEF085155400F78428BEFAA80000000804154B",
INIT_27 => X"1555D7FEAB55FF80175EF5D00020105D2A97400082E95555085168A10557FD75",
INIT_28 => X"00000000000000000000000000000000000000005D00020BA552A82000552A82",
INIT_29 => X"071EFB6DF7AE921C7FFFFFFFFFFFFFFFF7FBFDFFF5D2A954AA082A9242800000",
INIT_2A => X"1FAF55A2DF6DB7D1C002AB7D002A82028147FFFFFFFFFBFDFC7EBF5E8B550000",
INIT_2B => X"8E38E280871F8FC7E3D56AB6DBEDB7FFEF552AB8E38087FC2092087FFDFC7E3F",
INIT_2C => X"97FEFB6D1451471EF007BD0492B6F1F8F55AADF6DB7DE3F5FAFC708003DE28B6",
INIT_2D => X"A28407038140410492550A2ABC7497BD25FFAADF4516DBED16AA381C0A070824",
INIT_2E => X"D1C516FA28417BD5545E38E070280024904AA1C0438FD7005150438F78A2DBFF",
INIT_2F => X"92492A850105D2A80155417BEFB6DEB8E175FF5D0E05000492097428002E9557",
INIT_30 => X"4AA082A820AA000000000000000000000000000000000000000000000550A000",
INIT_31 => X"FF55A2D16AB550000175EFFFFBEAA00557FFFFFFFFFFFDFEFF7FBFFFEF552E97",
INIT_32 => X"C0000087BFDF45AAD568B55AAFBFDFEF55042ABEF002A800AA557FFDFEFF7FBF",
INIT_33 => X"16AB4500043DEAAFFAEAAAAA08516AB55A2D16ABEFFFFBFDFFF552AAAAAA007B",
INIT_34 => X"D568AAA5D2A97410007BFFFFF5551555EF087FC2000FFD56AB45A2FFFDFFFAAD",
INIT_35 => X"855400AAF7AEBDFEFA280154BA550400000552AA8B45087FC01EFA2FFD55EFF7",
INIT_36 => X"0804154BA082A975EF5D517DEAA007BD5545AAAA974AA0800020BA550028B550",
INIT_37 => X"00000000005D2E80010002A954005D2A82155087FFFFEFAAAA975EF5D2E97400",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000400000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(2),               -- Port A write enable input
DIA(0)   => data_write_a(18),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(18),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(2),               -- Port B write enable input
DIB(0)   => data_write_b(18),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(18),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_19_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"042200000000000041088001001AA00000000000000000000000500802000003",
INIT_01 => X"074018000024000000000404000000000A22000800000800004A200000000001",
INIT_02 => X"0000048002C405000000000006A84000000000200893C246A20000000020031A",
INIT_03 => X"082A58E411004B2000071000000981000C000000002045000200000000000000",
INIT_04 => X"200604000000001C0400001320000000162000002C4000026201201200090800",
INIT_05 => X"1020800000000058840200204000099070200E010001C0400000000000000000",
INIT_06 => X"0012048037805421402850001402498820022802400480405008901100A00102",
INIT_07 => X"00000000020C0130481204919200010C82000000000006002A548902A0020109",
INIT_08 => X"0001150800009900000005861840000000004301000B000000000001C1C00000",
INIT_09 => X"001F00002024B20002000000000002C300000000405000103010204000000000",
INIT_0A => X"00000000000000000000000000000040002000044000000000000000000002F0",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000420003B00000000000000000040012C80000000",
INIT_0D => X"45001A03C0825A0D20800000000018A006001000000000000000000000000000",
INIT_0E => X"450002131E01A1F6EA0A0020211146E069C2ACC01AE80045001D82ACC01AE800",
INIT_0F => X"1188340C3E1CFAD27CC2E004481020892282ACC01AE80045000582ACC01AE800",
INIT_10 => X"DEA03228D810007019931E01A1E5BA02802008C06F029D4C7B76639CEC0A0020",
INIT_11 => X"428AA3592000000206C2A4DAC00000008113C246A181C03FE4662A84575768DF",
INIT_12 => X"08201090549B5800000000261546B24000000000C53807E7CC06618018C51210",
INIT_13 => X"13F6A185A0A0168128411ACB800C0E108A0720288C011046B5986247C5452291",
INIT_14 => X"0000C220010808C10D9A92A74CD7CF4A080031B1515B212143D841431046B58A",
INIT_15 => X"00000000000000000000000000000000000000000000000000000118030004E0",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"3F0C7010C660C744192000000000000000000000000000000000000000000000",
INIT_19 => X"1861861861869A61861861861861861861861861A8208C4C1534D34C07208BBA",
INIT_1A => X"0984C26130984C26130984C26130984D26930984C26130984C261861861869A6",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE000000000000000000984C26130984C26130984C2613",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF552A974AA0004174BA0000000000000000000000",
INIT_22 => X"2E974BAA2FFFFE10087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974BA082E95400F7F",
INIT_23 => X"FFFFFFEFF7FBEAB450804001EFAAD57FEAAF7FFFFFFFFFFFFFFFFF7FBFDFFF55",
INIT_24 => X"002E82000F7FFFFFFFFFFFFDFEFA2D568B550004001EFAAAEA8ABA087FFFFFFF",
INIT_25 => X"5AAD16ABEF5D2ABFF55080402010087FFFFFFFFFBFDF45AAD568B55080028B55",
INIT_26 => X"BA087FFFFEFF7D168B55AAD17FFFF552EBFE00007FC00AAF7FFFFFFFF7FBE8B5",
INIT_27 => X"FFF00043DE10AA843DE00557FFDFEFA2D16AB55A2FFFDFEF5D2EBFE00AAFFFFE",
INIT_28 => X"0000000000000000000000000000000000000000AAFFFDF45A2D16AB55F7FFFF",
INIT_29 => X"954AA082A92428E3FFFFFFFFFFFFFFFFFFFFFFFEF552A974AA0000104AA00000",
INIT_2A => X"FFDFEFF7F5FAFC7492A974AAB6F5F8E101C7FFFFFFFFFFFFFFFF7FBFDFFF5D2A",
INIT_2B => X"A4A8AAA147FFFFFFFFFBFDFC7EBF5E8B550000071EFB6DF7AE92EBFFFFFFFFFF",
INIT_2C => X"2DF6DB7D1C002AB7D002A82028FFFFFFFEFF7F1F8FD7AAD16AB450000001FFBE",
INIT_2D => X"F7FBF8FC7E3F5EAB45B6DF6FBEF5D2AB8F7D000000010087FFDFC7E3F1FAF55A",
INIT_2E => X"7412ABFE28B6F5F8E820871F8FC7E3D56AB6DBEDB7FFEF552AB8E38087FC2092",
INIT_2F => X"55AADF6DB7DE3F5FAFC708003DE28B68E38E284971F8FC7AAD56DB6DBEF5F8FD",
INIT_30 => X"4AA0004000AA000000000000000000000000000000000000000000000B6F1F8F",
INIT_31 => X"DFEFF7FBFFFEF552E974AA082A820AAA2FFFFFFFFFFFFFFFFFFFFFDFEF552E95",
INIT_32 => X"EAA00A2FFFFFFFF7FBFDFFFFFD568B55002A954AAF7D568A00557FFFFFFFFFFF",
INIT_33 => X"56AB450004001EFFF842AAAA557FFDFEFF7FBFFF55A2D16AB550000175EFFFFB",
INIT_34 => X"7BFDF45AAD568B55AAFBFDFEF55042ABEF002A800AAF7FBFDFEFF7D56AB45AAD",
INIT_35 => X"52AAAAAA007BC0000FFFBE8B55AAD168B55F7FFFFFFF552AA8BEF08040200008",
INIT_36 => X"A2D57FFFFF7D568B45002ABDEAAFFD16AA0008516AB55A2D16ABEFFFFBFDFFF5",
INIT_37 => X"0000000000FFD56AB45A2FFFDFFFAAD16AB4500043DEAAFFAEAAAAA08556AB55",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000800000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(2),               -- Port A write enable input
DIA(0)   => data_write_a(19),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(19),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(2),               -- Port B write enable input
DIB(0)   => data_write_b(19),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(19),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_20_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000003",
INIT_01 => X"A65FF80000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000048002CC070000000000000000000000002FF86100200000000220002362",
INIT_03 => X"0000000000080F6000977060009B87A03C000000000000000000000000000000",
INIT_04 => X"3F2EFC040388137C3E20C477600142019E6000003CC0000A6601601A000B0000",
INIT_05 => X"102F91D10802ABFB80000021C8010FB0F0F43E1FE867DFC04400390210000220",
INIT_06 => X"90492261000080003400000010008000004203FE400580000000803000200006",
INIT_07 => X"401000004FFDFF28C4300C0010200100004000002AA001F00000000014000000",
INIT_08 => X"0801F5780259FB00000007BEFBC010002008FF7F00000000010018A81000041C",
INIT_09 => X"00000000020000000000000000000ADF00000020000000800000802830011023",
INIT_0A => X"0000000000000200020000000000000000000000000000000200200290000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"08120000B9090A700000200000004000000400000080002000407FED80000000",
INIT_0D => X"000079804000F00000000000C01FF8A7FE003000000004008100000000000000",
INIT_0E => X"0000798201000000100000000135386000401000010000000079801000010000",
INIT_0F => X"0185C300020004000010000000000252C7801000010000000079801000010000",
INIT_10 => X"00000010C1F30F300002010000080000000000CD8A0000400400000010000000",
INIT_11 => X"008040000000000292C0080000000000A5604000000284000818505200080000",
INIT_12 => X"0015E1B00100000000001496008000000000052B000048080000000000FC3600",
INIT_13 => X"80000000000002BA280000800830300000000000B8B400000401881010000000",
INIT_14 => X"00000000020020020001000040283024E6FB8604020080000383383B00000400",
INIT_15 => X"000000000000000000000004010201001003020200000000000127DBFF004000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"038200010089120104D204002000000000000000000000000000000000000000",
INIT_19 => X"B2CB2CB2CB2CB2CB2CB2CB2CB2C30C30C30C30C306982121A1E79E79A0700030",
INIT_1A => X"432190C86432190C86432190C86432190C86432190C86432190CB2CB2CB2CB2C",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000432190C86432190C86432190C86",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA0804020100000000000000000000000",
INIT_22 => X"2E954AA000400000F7FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0004174BAFFF",
INIT_23 => X"FFFFFFFFFFFFFDFEF5D2A974BA082E95400007FFFFFFFFFFFFFFFFFFFFFFEF55",
INIT_24 => X"A2FFFFE10FFFFFFFFFFFFFFFFFFFFFBFDFFF5D2E954BA007FC00BA087FFFFFFF",
INIT_25 => X"FF7FBFFF550800020BAAAD56AAAAF7FFFFFFFFFFFFFFFFF7FBFDFFF552E974BA",
INIT_26 => X"10087FFFFFFFFFFFFFEFF7FBEAB450804001EFAAD57FEAA007FFFFFFFFFFFFFE",
INIT_27 => X"B550004001EFAAAEA8ABA5D7FFFFFFFFFFFDFEFF7D56AB450000021EFA2D57DE",
INIT_28 => X"0000000000000000000000000000000000000000F7FFFFFFFFFFFFDFEFA2D568",
INIT_29 => X"974AA0000104AAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA08000500000000",
INIT_2A => X"FFFFFFFFFBFDFEF5D2E974AA000A07000E3FFFFFFFFFFFFFFFFFFFFFFFEF552A",
INIT_2B => X"71C50BA1C7FFFFFFFFFFFFFFFF7FBFDFFF5D2A954AA082A92428087FFFFFFFFF",
INIT_2C => X"7F5FAFC7492A974AAB6F5F8E10E3FFFFFFFFFFFFFFEFF7FBFFFFF552E974AA00",
INIT_2D => X"1C7FFFFFFFFFBFDFEFE3F5F8F450004050AABEDF6FABAEBFFFFFFFFFFFFDFEFF",
INIT_2E => X"50804021FFB6D57DE28147FFFFFFFFFBFDFC7EBF5E8B550000071EFB6DF7AE92",
INIT_2F => X"EFF7F1F8FD7AAD16AB450000001FFBEA4A8AAA497FFFFFFF7FBF8FC7EBD168B4",
INIT_30 => X"4AA080017410000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFDFEF552E954AA0004000AAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A95",
INIT_32 => X"820AA087FFFFFFFFFFFFFEFF7FBFDFFF5D2A974AA002E95410A2FFFFFFFFFFFF",
INIT_33 => X"FFDFEF5D2E954AA0051554BA557FFFFFFFFFFFDFEFF7FBFFFEF552E974AA082A",
INIT_34 => X"FFFFFFFF7FBFDFFFFFD568B55002A954AAF7D568A00AAFFFFFFFFFFBFDFEFFFF",
INIT_35 => X"000175EFFFFBEAA005D7FFFFEFF7FBFDFFFAAD16AB450804174AAFFFFFFEBAA2",
INIT_36 => X"F7FFEAB45A2D568B550804001EFF7D57DEBA557FFDFEFF7FBFFF55A2D16AB550",
INIT_37 => X"0000000000F7FBFDFEFF7D56AB45AAD56AB450004001EFFF842AAAA087BFDFEF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000000FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(2),               -- Port A write enable input
DIA(0)   => data_write_a(20),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(20),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(2),               -- Port B write enable input
DIB(0)   => data_write_b(20),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(20),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_21_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"4A302428B824900A128C090A5C1800261500213C005FE812D10420054085A202",
INIT_01 => X"081FFE3440B609703B0427F801A40B8115BC4F655300340288A40D30040E4DD8",
INIT_02 => X"04CA478082CC1740002019824E0203100640303FF8C0B31061096E21A1840814",
INIT_03 => X"8C329E9204020FE002577800405B87047D5042129D8D0248903200013290C800",
INIT_04 => X"3E7FFE02482553FC3C020277E128080A1E6000003CC0000A6601E03A8B0F0008",
INIT_05 => X"F43F8140000203FFC806C8A1C1048FF0F0E07E1F00F7FFC00024010000468310",
INIT_06 => X"08710C10015E083D01A24404786BE0014114C3FE4187A009A663A680100B3096",
INIT_07 => X"200800008FDFFF00290000100211019812E210488228000000900260026C6058",
INIT_08 => X"0EF1F5FA0041FF080AC707FEFBC110008420F7FF388B70A20389346FE8000580",
INIT_09 => X"917FC30010107688862A28C54518DBFF00020004C0A6044901112A0908AA0A30",
INIT_0A => X"006309044081A001B188300E20806520398C6021569249C4B3007127080806FF",
INIT_0B => X"904595123203040D9228D9228D9228D9228D9228D9228D9228D99146C9146C84",
INIT_0C => X"88042090068008003120000806001402504110C48002403601887FEF80022A51",
INIT_0D => X"26C0AC404E43032CA0C205880A7FFAB7FE01409400400C0594A4002200110008",
INIT_0E => X"26C0AC086A170250454004C6012280129B034A080C0B0016A0D20346080C0A80",
INIT_0F => X"0B064092D85938C0112144050224120C500346080C0B0016A0D2034A080C0A80",
INIT_10 => X"40702E058355458967E86A170220D1800093414B0414782E4B5000D81480809A",
INIT_11 => X"081B1545104135443306C35901024F88A88049062A747512B76783C5D040E080",
INIT_12 => X"40160040D86B202049B22198362A8A208279854400A036801480031401900800",
INIT_13 => X"0DD001C002D38334000914028354008301008C0CF1480245108C7640A0604032",
INIT_14 => X"AC0496022300233104662848808E191526205018030060540284FA0C0044022C",
INIT_15 => X"004010040100401004010040102090010008000001C0E010020007DFFFC06E60",
INIT_16 => X"0401004010040100401004010040100401004010040100401004010040100401",
INIT_17 => X"4010040100401004010040100401004010040100401004010040100401004010",
INIT_18 => X"FF7FFDF7FF3E3DFDF7E000000000000000000000000040100401004010040100",
INIT_19 => X"FBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBFFDFDFFFCF3CF3FFFEF9FEE",
INIT_1A => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFEFF7FBFDFEFF7FBFDFEFBEFBEFBEFBE",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0004000100000000000000000000000",
INIT_22 => X"2A954BA0004154BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080402010FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF552A974AA0004174BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"000400000007FFFFFFFFFFFFFFFFFFFFFFEF552E974BA0804000AAF7FFFFFFFF",
INIT_25 => X"FFFFFFDFEF5D2E974BA002E97400007FFFFFFFFFFFFFFFFFFFFFFEF552E954AA",
INIT_26 => X"BA087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974BA082E95400007FFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2E954BA007FC00BA5D7FFFFFFFFFFFFFFFFFFBFDFEF5D2A954AA002E974",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFBFD",
INIT_29 => X"954AA080005000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA00000200000000",
INIT_2A => X"FFFFFFFFFFFFFFF552A974BA0000174AAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0A000AAE3FFFFFFFFFFFFFFFFFFFFFFFEF552A974AA0000104AAF7FFFFFFFFFF",
INIT_2C => X"FFBFDFEF5D2E974AA000A07000007FFFFFFFFFFFFFFFFFFFFDFEF552E954BA08",
INIT_2D => X"1C7FFFFFFFFFFFFFFFFFFBFDFEF5D2A974BA002A95400087FFFFFFFFFFFFFFFF",
INIT_2E => X"F552E974BA0020924BA1C7FFFFFFFFFFFFFFFF7FBFDFFF5D2A954AA082A92428",
INIT_2F => X"FFFFFFFFFEFF7FBFFFFF552E974AA0071C50BA557FFFFFFFFFFFFFFFF7FBFDFF",
INIT_30 => X"4BA000002000000000000000000000000000000000000000000000000E3FFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2A954AA080017410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"000AAF7FFFFFFFFFFFFFFFFFFFFFFFEF552A974BA0000174BAFFFFFFFFFFFFFF",
INIT_33 => X"BFDFEF5D2A954BA082E800AAA2FFFFFFFFFFFFFFFFFFFFFDFEF552E954AA0004",
INIT_34 => X"7FFFFFFFFFFFFFEFF7FBFDFFF5D2A974AA002E95410087FFFFFFFFFFFFFFFF7F",
INIT_35 => X"52E974AA082A820AA557FFFFFFFFFFFFFEFF7FBFFFFF552E954BA002E9741008",
INIT_36 => X"FFFBFDFEFF7FFFFFEF5D2A974BA0000020AA557FFFFFFFFFFFDFEFF7FBFFFEF5",
INIT_37 => X"0000000000AAFFFFFFFFFFBFDFEFFFFFFDFEF5D2E954AA0051554BA5D7FFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(2),               -- Port A write enable input
DIA(0)   => data_write_a(21),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(21),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(2),               -- Port B write enable input
DIB(0)   => data_write_b(21),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(21),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_22_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"5290F4CDE914905A14A43D33F488243E17122300F55FEB189B343A1140548380",
INIT_01 => X"A94007B259F6A975386262000C344BA9573C6FF57B18A5FB0ABFCD3C2C5F4F0C",
INIT_02 => X"D56B4302AC01005111011BD506AA5205274056900596A539584E2E6DFE4B2418",
INIT_03 => X"6B03F2F6151A2081F24001E8400008F401CB10C6594423C8923AD6B55AD0EB5A",
INIT_04 => X"8001023D37E50880436200808BC8492A0089249600101100008087248B64426E",
INIT_05 => X"A51035B41C0A88046CAEE8C23C08E040011C0020F8882001102D620A06D68301",
INIT_06 => X"B93FF975CF7889D085E997A2144E8FC2060B880081A26DCD4047EFF9EF018980",
INIT_07 => X"283800AA500200E8024AD03546A3262FB5AA5542A882040C7A64CBD64065F028",
INIT_08 => X"141008801018040E48D500400015805060040080A2A0F4A82381B4000A0905A0",
INIT_09 => X"4D0000002126F30C902A29C54539C020E11810098D4067EFF9FF284D483E2AB4",
INIT_0A => X"1400006100003202D040050220103D2A512C6A8C4F0008AA800470370000A000",
INIT_0B => X"013456520CA09281C2A81C2A81C2A81C2A81C2A81C2A81C2A81C9540E1540E00",
INIT_0C => X"A1402A13C0A10A893165281A1C2A7283516344C594A85536B1AD800214202C50",
INIT_0D => X"3C70FC20515808A0100820112300011000287B071105034406950A0285014280",
INIT_0E => X"3C70FC48E11CFC48400184CE0D6783139B0959A41606003C70FA0958AC160480",
INIT_0F => X"0D87E8B3B811B52048B10E0402AE1606D80958AC1606003C70FA0959A4160480",
INIT_10 => X"80F84E0185594581E088E11CFC38414020DD42CF909D7E0A551C02180300C0DD",
INIT_11 => X"441154C258012D86F3044A3133004A99BD8455300654458A1D588C4061403000",
INIT_12 => X"A096A240894626600953379822A984B0025B0DEC0345C9200680027181B44887",
INIT_13 => X"E2404160035482BE521C2C04A90783C18000D610B9D8070B12B1A2A62040202A",
INIT_14 => X"304244A91102C93A2D608D2A258DF8034284200C050070E40C80620C870B02C4",
INIT_15 => X"4411044110441104411044110466C440446CA06951D4EA801000980400646002",
INIT_16 => X"0100441104411044110441104411044110441104411044110441104411044110",
INIT_17 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_18 => X"FE8FF1F7DEBDDF7DF7D05122890000000003FFFFFFFF90040100401004010040",
INIT_19 => X"79E79E79E79E79E79E79E79E79E79E79E79E79E7BFFDFD7DDDF7DF7DF7DFBFDE",
INIT_1A => X"3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE79E79E79E79E",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE000000000000000003F9FCFE7F3F9FCFE7F3F9FCFE7F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0800000000000000000000000000000",
INIT_22 => X"2E974AA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000400010FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E954AA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"0004154BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA000015400FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF552A974AA0800154AAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA",
INIT_26 => X"BAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0004174BAFFFFFFFFFFFFFFFFF",
INIT_27 => X"FEF552E974BA0804000AAA2FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0000174",
INIT_28 => X"0000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040001000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E954AA000402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0417410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080005000FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF552A974BA0000174AAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA00",
INIT_2D => X"E3FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0804154BAF7FFFFFFFFFFFFFFFFF",
INIT_2E => X"F552E954BA000E124BAE3FFFFFFFFFFFFFFFFFFFFFFFEF552A974AA0000104AA",
INIT_2F => X"FFFFFFFFFFFFFFFFDFEF552E954BA080A000AAA2FFFFFFFFFFFFFFFFFFFFFFFE",
INIT_30 => X"4BA080400010000000000000000000000000000000000000000000000007FFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"17410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000400010FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF552A954BA000415400FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954AA0800",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFEF552A974BA0000174BAF7FFFFFFFFFFFFFFFFFFF",
INIT_35 => X"52E954AA0004000AAA2FFFFFFFFFFFFFFFFFFFFFDFEF552E974AA0804174AAF7",
INIT_36 => X"FFFFFFFFFFFFBFDFEF5D2E954BA002A820BAA2FFFFFFFFFFFFFFFFFFFFFDFEF5",
INIT_37 => X"0000000000087FFFFFFFFFFFFFFFF7FBFDFEF5D2A954BA082E800AAAAFFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000000FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(2),               -- Port A write enable input
DIA(0)   => data_write_a(22),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(22),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(2),               -- Port B write enable input
DIB(0)   => data_write_b(22),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(22),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_23_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"EF20906D902424807BC8241BC81801B97D38AD3C0800103362A6741C80A12A02",
INIT_01 => X"001FFF8409F089003B4422000D80C80106804A7951C5B9D1C828043EA28838F9",
INIT_02 => X"028406A002DC176444683862400003111001303FFC00F240D50146013B300500",
INIT_03 => X"001B243004080FE000177003145F87017D584B10D804034800200200A1008008",
INIT_04 => X"BEFFFC0248005FFC3C18A2FFE12222425E600000BDC0800AEE01E81A100F0A00",
INIT_05 => X"D03F8000000003FF810640A1C0008FF2F0E17E1F02FFFFC80100004044800080",
INIT_06 => X"800264B4854650040123428C204BF40F439647FF4807E189A477EF81DF0AF116",
INIT_07 => X"01000000FFDFFFE800401005C0A0008F86C60840AAAA100C68D1810C9F4A0020",
INIT_08 => X"1BE1F5F80003FF0002021FFEFBC80000000077FF184B03010004002FE1F29002",
INIT_09 => X"907FC308181204800600000000001BFFA800808189A657EF81DD0C00079CC800",
INIT_0A => X"0063090442A18001B188300C48907120AC810033149249C433200180082A06FF",
INIT_0B => X"9A41C1443243050C1010C1010C1010C1010C1010C1010C1010C1008608086084",
INIT_0C => X"000082A00600200080000500C000400800601200000254A000007FEFC1030221",
INIT_0D => X"0A9080400E0BF30C20CA858E087FFABFFE01409780214EE49620001000080004",
INIT_0E => X"0A908044294700701641005218521210150E5789F90A000A90800E5F81F90880",
INIT_0F => X"0E0220036864A7DCA190440301E2105C000E5F81F90A000A90800E5789F90880",
INIT_10 => X"C1400500C6CE5400032429470068924010164302048156305D66F8701681000E",
INIT_11 => X"2E0CCB0500013440600339C800004D8018000857A82920CE8CB220C81400A180",
INIT_12 => X"220344406739000009B0030019960A00026880C0422C52B01700044901488822",
INIT_13 => X"85C811A010428104128996465ADA020180804A040108A2658217C4008060300C",
INIT_14 => X"BE0692020328CA0028042054A92771C50FC070109000C1C819078280A265920E",
INIT_15 => X"020080200802008020080200800800200200000000000008004807DFFF000470",
INIT_16 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_17 => X"0080200802008020080200802008020080200802008020080200802008020080",
INIT_18 => X"0000000000000000000000000000000000000000000000802008020080200802",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000",
INIT_22 => X"2E974BA080002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E974BA000400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000400000FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF5D2E954AA080000010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA",
INIT_26 => X"10FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080402010FFFFFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2A954BA000015400FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA0804000",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E974BA080002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF5D2E954AA000402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA00",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080002010FFFFFFFFFFFFFFFFFFF",
INIT_2E => X"F5D2A954BA080407000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080005000",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF5D2A954BA000417410FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA080402000000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"02000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000010FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF5D2E974AA000402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0000",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000400010FFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"D2A954AA080017410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954AA080002000FF",
INIT_36 => X"FFFFFFFFFFFFFFFFFF552A954BA080015410FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_37 => X"0000000000F7FFFFFFFFFFFFFFFFFFFFFFFFF552A954BA000415400F7FFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000000FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(2),               -- Port A write enable input
DIA(0)   => data_write_a(23),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(23),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(2),               -- Port B write enable input
DIB(0)   => data_write_b(23),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(23),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_24_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100600007FFF000080108004000800020000840041000080808",
INIT_02 => X"0000068002CC07400000090C080002000000103FF811F150231000520ABE4404",
INIT_03 => X"8428180000080FE000177000001B87003D4000000E8B84010020000000008000",
INIT_04 => X"3E2FFC024800137C3C000077E00000001E6000003CC0000A6601E01A000F0200",
INIT_05 => X"103F8000000003FF80000021C0000FF0F0E03E1F0067FFC00000000000000000",
INIT_06 => X"00132412079001AD00810005E8000001401643FE4007E5501AA00000DC8C3006",
INIT_07 => X"000000000FDFFF62695A5685C094831D966000008002100C2040A178B600C240",
INIT_08 => X"08E1F5F80001FF00000007FEFBC00000000077FF000B00000000002FE0000000",
INIT_09 => X"107FC300000000000600000000001BFFA0000005501AA00000CE200000940000",
INIT_0A => X"00630104408180012188300C00814080008000010012414433000100080806FD",
INIT_0B => X"904181003003000C1000C1000C1000C1000C1000C1000C1000C1000608006084",
INIT_0C => X"00000080060000000000000012002C00000000000000000000007FEF80020201",
INIT_0D => X"440082404E0B332CA2C20188087FFAB7FE000082000000008220000000000000",
INIT_0E => X"4400824903210308074084210002460402009280010D80440084009280010F00",
INIT_0F => X"800A2400401A0C82183248060010280C20009280010D80440084009280010F00",
INIT_10 => X"C0A078160000404A0469032102981380202080026420020D06C002A08481C020",
INIT_11 => X"00164F400860000824059AD01802000208104817B00011306B2D9B0DD5082080",
INIT_12 => X"41021800B35A0300400041202C9E8010C0001040C5836CC01780018601030088",
INIT_13 => X"DB1011E000A140058220004AEFFC8101810021084301880030A8B77400603011",
INIT_14 => X"8C063C0220002201490418082010A57263E010000201033016085A40880030A1",
INIT_15 => X"000000000000000000000000000000000000000000000000000007DFFF0006E0",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"F6E7CC1132CDB444199000000000000000000000000000000000000000000000",
INIT_19 => X"79E79E79E79EFBEFBEFBEFBEFBEF9EF9EF9EF9EFA69861219575D75FF2D0AEEA",
INIT_1A => X"0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1EFBEFBEFBE79E",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE000000000000000000783C1E0F0783C1E0F0783C1E0F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020100000000000000000000000",
INIT_22 => X"2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"080002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_26 => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000400010FFFFFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2E974AA000400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0004000",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040201000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF5D2E974BA080002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFF",
INIT_2E => X"F5D2E974AA000400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF5D2E974AA000400000FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA080402010000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"00010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000010FFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002010FF",
INIT_36 => X"FFFFFFFFFFFFFFFFFF5D2E974AA000002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_37 => X"0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000402010FFFFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(3),               -- Port A write enable input
DIA(0)   => data_write_a(24),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(24),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(3),               -- Port B write enable input
DIB(0)   => data_write_b(24),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(24),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_25_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100200002000000080100004000000020000800041000080808",
INIT_02 => X"0000068002CC474000000800000002000000103FFCE302008000000880844A04",
INIT_03 => X"00000101C0200FF004177800081B87003D400000080000000020000000008000",
INIT_04 => X"3E2FFE024820137C3C004077F01000001E7249213CC1264A660DF05A000F9000",
INIT_05 => X"103F81C1002203FF80000021C1140FF8F0E03E1F0067FFE04800258280010052",
INIT_06 => X"80480AE20000000100000001C8608001401643FE4007C00000000000CC083006",
INIT_07 => X"280800000FDFFFEA4050140540B00100840000080002A00C2040810000000010",
INIT_08 => X"C8E1F5FA21C9FF80040007FEFBE031018C31F7FFBAEBC0020008086FE0000100",
INIT_09 => X"107FC301800000000600000000001BFFE00301000000000000CC020000140000",
INIT_0A => X"0077330C4889CC292588300C0080400000800001001243443B000100880806FD",
INIT_0B => X"904189003003000C1000C1000C1000C1000C1000C1000C1000C1000608006084",
INIT_0C => X"8B04228026824100000000000000000000000000000004A000007FEF80020201",
INIT_0D => X"400000400E03C30C20C2818C087FFAB7FE01409700C10007962418220C110608",
INIT_0E => X"4000000001010000004000000000400400001200000800400000001200000800",
INIT_0F => X"0008000000000480000040000000200000001200000800400000001200000800",
INIT_10 => X"0000001001000002000001010000100000000000202000000440000000800000",
INIT_11 => X"0000410000000008000008400000000200000806300400000820000020004880",
INIT_12 => X"0000080001080000000040000082000000001000000040800800000000020008",
INIT_13 => X"8100000000000000802000000840000200040000020008000000840000804000",
INIT_14 => X"8C04100200000200000610000000210000000018140000000008000008000000",
INIT_15 => X"04411044110441104411044510629041040D180400000010028047DFFF800C60",
INIT_16 => X"4411044110441104411044110441104411044110441104411044110441104411",
INIT_17 => X"4110441104411044110441104411044110441104411044110441104411044110",
INIT_18 => X"196A8C5A2932EC15DA080800002FFFFFFFFFFFFFFFFFC1104411044110441104",
INIT_19 => X"92492492492410410410410410410492410492412000531215A69A6BFBA2894A",
INIT_1A => X"B158AC562B158AC562B158AC562B1588C46231188C46231188C4924924924924",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000B158AC562B158AC562B158AC562",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000",
INIT_22 => X"2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF5D2E974BA080400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_26 => X"10FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0800000",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400000FFFFFFFFFFFFFFFFFFF",
INIT_2E => X"F5D2E974BA080000010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA080402000000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"02000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400000FF",
INIT_36 => X"FFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_37 => X"0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000000FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(3),               -- Port A write enable input
DIA(0)   => data_write_a(25),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(25),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(3),               -- Port B write enable input
DIB(0)   => data_write_b(25),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(25),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_26_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"E9264EAB20190CA3BA4997AA9002AE9C001006B0778015CFA17E0811039879C7",
INIT_01 => X"F1FFF9BB1F773C7F9BB07DFFFDD863FC5FFF3FEFFBBF9FFB22FFFBC7B9F30686",
INIT_02 => X"9B3184F8AFDEAF300029E4E300FC78A6258548EFFA71C00172082400003A2161",
INIT_03 => X"0213C3FDFFFC7F74FFBF737A603B87FEBE1A5294F65628A0001B9CE6CC606E73",
INIT_04 => X"7E2EFEBF6FFEB37C3FF3017776FFCDA43E7B6DFD7DEBFD8E6F5F78DF0BFBD644",
INIT_05 => X"902F87C74E8CCFFBB6FF70E1FE61FFBDF0FEBE1FFD67DFFEFFBDA7F7FED50870",
INIT_06 => X"213246200BCC8920360C1831CD7DF60A244B9BFEE00589DDBCEFEDC1DFA08957",
INIT_07 => X"B1D4223B4FFDFF21CC721C85DCE1458E8782484020A2C1FCA3468D77E0000300",
INIT_08 => X"2C05FD7BC471FBD13D980FBEFBEBF30B8D79FF7F451F33CFD60FE8FFFDF54003",
INIT_09 => X"19FFC71FEFED7B251E35768E8ED6BFDF3EB3EBF9DDBCE7FDC1DF8A760F3EACC0",
INIT_0A => X"56F7730ECCDBDF152199F51EDDCDEBCFF589807B7096CD4CF73AC1FC98884FFF",
INIT_0B => X"B867D3683A03A40F78C0D78C0D78C0D78C0D78C0D78C0D78C0D7A606BC606B8C",
INIT_0C => X"DFBFF5EB36DFE51FC3A80D73D840303983EE7F0EA03BDA680137FFFDFFD7E681",
INIT_0D => X"3F0080425E6BFF8DB0DAE19C09FFFFE7FE3EBEA8EB7AFEE5C9AEBD7F5EBFAF5F",
INIT_0E => X"3F00800DEC010280004000F808020290100FA2F60008003F00800FA2F6000800",
INIT_0F => X"00023002007BC0A14E00400003B8000D000FA2F60008003F00800FA2F6000800",
INIT_10 => X"01E0320007204008040DEC010300100000F600020581003F604D0700008000EE",
INIT_11 => X"201F21A2C40039006807C46426040E101A0259DFE82011A311AA042016040080",
INIT_12 => X"80020048F88C84C101C203403E434588007200D047F00090200007E0010009B0",
INIT_13 => X"0109000003E2000416C0804FE04140E80000F808010AB02033AC048A2A00003D",
INIT_14 => X"FFAFD082003B032FB987E04021D481D4000419060201E1A000044300B02033E8",
INIT_15 => X"AFEBFAFEBFAFEBFAFEBFAFEFFBFBFBFBBFCFBB0FFDFEFFEF2DFFFFFBFF802FFD",
INIT_16 => X"FEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBF",
INIT_17 => X"EBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFA",
INIT_18 => X"F491E166CC8553F86EDB5C88646FFFFFFFFFFFFFFFFFEBFAFEBFAFEBFAFEBFAF",
INIT_19 => X"1861861861861861861861861861869A69A61861AFBD54D5F871C71D475B15BC",
INIT_1A => X"0984C26130984C26130984C26130984C26130984C26130984C26186186186186",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE000000000000000000984C26130984C26130984C2613",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000",
INIT_22 => X"2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_26 => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFF",
INIT_2E => X"F5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA080402000000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"02010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_36 => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_37 => X"0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(3),               -- Port A write enable input
DIA(0)   => data_write_a(26),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(26),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(3),               -- Port B write enable input
DIB(0)   => data_write_b(26),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(26),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_27_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"00080A40000A41248002029000050A088000008242A0004404480002000A1155",
INIT_01 => X"F1FFF1C11F781C129C107DFFFE0860941E81258CA2B71C2220EC1B86E1A00002",
INIT_02 => X"183080988B2EAE00002BE001117C78C6848140CFFA0000800042008000011081",
INIT_03 => X"000003FDF3E47C74F7BCF36A203A47F6B8184210B6160820001318C60C204C63",
INIT_04 => X"7E28FEBF6FEEB3723F71017476DFC524397B6DF572EB6C8E175E70D90F539600",
INIT_05 => X"000F86064C8DDFE3B6FF50D1FC61DE39C8FCB91FF9671FE6B68984B5BCE40834",
INIT_06 => X"0000000800000042020C18300520620A80231BFE200181092CE7ED80DFC00147",
INIT_07 => X"8AC4AA3B0FD1FF201044110560884000840200520002080C23468D0300000282",
INIT_08 => X"2005F0784411E390A4880E3DF7E2FB0B8E717C7F411F3BC6D60B60FFDDE44001",
INIT_09 => X"18FFD757E7ED7A211E81C09818109E1F16B16B71092CE7ED81CF403601228C40",
INIT_0A => X"46FF730E5CCBCD55219AB55F0DEFABC7054880693016DD4C755AC16C1A884FFE",
INIT_0B => X"BC63F1683803C00E3440C3440C3440C3440C3440C3440C3440C3C2061A2061AD",
INIT_0C => X"56BF55CB165EC51D41880FA3F040202883B475062033186801137FF1BAD6F281",
INIT_0D => X"3B0000421E2B0F2E2AE215C808FFFA47FE62BAA86B1AB268E92AB56D5AB6AD5B",
INIT_0E => X"3B000025EC010080004000F808000098100F22520008003B00002F2252000800",
INIT_0F => X"00001042006BC0810600400003B80001002F22520008003B00002F2252000800",
INIT_10 => X"01E032000620000C0405EC010100100000F6000001C1003760410500008000EE",
INIT_11 => X"201D2120840039000817444404040E10020218DE282010A311AA002002040080",
INIT_12 => X"8000000AE888808101C20040BA4241080072001027F00080200007E0000001F0",
INIT_13 => X"0101000003E2000007C0800FE04040280000F8080002F02023AC04080A00003D",
INIT_14 => X"DDAFD082001B03249887E04001D481D4000009020201E1A000040100F02023E8",
INIT_15 => X"ADAB6ADAB6ADAB6ADAB6ADAB6BF1EBDABD8E270BF84A25C6ACB777E3FF800C6D",
INIT_16 => X"DAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6",
INIT_17 => X"AB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6A",
INIT_18 => X"100481CA860402104A471688747FFFFFFFFFFFFFFFFFAB6ADAB6ADAB6ADAB6AD",
INIT_19 => X"0000000000000000000000000008200000000000200072F210000001490E2168",
INIT_1A => X"A05028140A05028140A05028140A050080402010080402010080000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000A05028140A05028140A05028140",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000",
INIT_22 => X"2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_26 => X"10FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFF",
INIT_2E => X"F5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA080402000000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"02000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FF",
INIT_36 => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_37 => X"0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000000FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(3),               -- Port A write enable input
DIA(0)   => data_write_a(27),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(27),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(3),               -- Port B write enable input
DIB(0)   => data_write_b(27),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(27),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_28_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"02200AA400180030808802A900002A08001280A08A801044104A1000001818C3",
INIT_01 => X"50A00011460214428114180000882214413D0A71592A01D92213D28005210202",
INIT_02 => X"8A54800A210200111100C2110054289220810440030404010844000444410001",
INIT_03 => X"4200040822D4500001E0000028000002000211842010092000018C6295200631",
INIT_04 => X"00400000000B8000000140000005840C00000040002008808100048100100044",
INIT_05 => X"0000222200244400135110000135100000000000000000024CA0A01018000320",
INIT_06 => X"A004912008208040024489121144080400081000200008104000000020000041",
INIT_07 => X"A85800994000000A0200802004204420210001022AA8A0001122448142491008",
INIT_08 => X"0414000201800004080A000000124058200408000880004440004080160C4100",
INIT_09 => X"0080000206CB0821082B694D4D29400002002038104000000020003204000440",
INIT_0A => X"12000843066021001400040024440245400082D022040000400800081022C000",
INIT_0B => X"0002002C004001036050160501605016050160501605016050160280B0280B00",
INIT_0C => X"0012400810080414C0A800310840102182C62302A0194C08001680100E4040A0",
INIT_0D => X"05000002003004208208841401800040000A0000200814004198000400020001",
INIT_0E => X"0500000004000080000000000000028000002052000000050000002052000000",
INIT_0F => X"0000300000004001060000000000000900002052000000050000002052000000",
INIT_10 => X"0000000001200000000004000100000000000000050000002001050000000000",
INIT_11 => X"00002020840000004800040404040000120200A9000000010000002002040000",
INIT_12 => X"0000004800808081000002400040410800000090001000002000000000000910",
INIT_13 => X"0001000000000000144000010000402800000000000A1000010000080A000000",
INIT_14 => X"0080000000110006B08140000040000000000902000000000000410010000100",
INIT_15 => X"0080200802008020080200802101210810C39A66A90A85420413A82000000204",
INIT_16 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_17 => X"8020080200802008020080200802008020080200802008020080200802008020",
INIT_18 => X"110A00246972BD89A40A0C22E100000000000000000000200802008020080200",
INIT_19 => X"82082082082082082082082082082082082082080D35050758C30C31DE21102C",
INIT_1A => X"B0582C160B0582C160B0582C160B0580C06030180C06030180C0820820820820",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000B0582C160B0582C160B0582C160",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000",
INIT_22 => X"2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_26 => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFF",
INIT_2E => X"F5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA080402000000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"02000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_36 => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_37 => X"0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"00000000000000000000000000000000000FFFFFFFFF00000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(3),               -- Port A write enable input
DIA(0)   => data_write_a(28),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(28),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(3),               -- Port B write enable input
DIB(0)   => data_write_b(28),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(28),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_29_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"79964E4BA01DACAB9E659792D00AAE160002829C7FDFEFCEE97C2815039D70C3",
INIT_01 => X"50BFF9AB0775343F9AB01DF80D5821FC0FFF3FEFD1AF9FF1207FFBC7B9720586",
INIT_02 => X"0D15846807D207200021C4E200D428A2018408600271C000720A0000003A2161",
INIT_03 => X"0002C009EEFC5F10F9B70178681B80FA3E000100765029A00019084345606421",
INIT_04 => X"3E6E023D27DA937C03E3407712E5CDA41E0924DC3D20B98AE905189F0BF8C000",
INIT_05 => X"902003C30E0447F877F930203E213F8CF01E3E00FC67C03A4D9C87525E510160",
INIT_06 => X"0012460003CC002036040811D919F402244293FEE00400CCB46BA4C164A08857",
INIT_07 => X"914800110FFC0001CC320C81D841418E82800100000041FCA1428575A0001108",
INIT_08 => X"0805FD0180E1F8C1111A0782082B50080508FF00048B124D4005C8AFF4154102",
INIT_09 => X"0180000ABFEF89250815568A8AD6ABC02A02A0B0CCB463B4C0748A720B1EA4C0",
INIT_0A => X"021410028450530014014002D445624DB481806A62840800C22800B8900042FF",
INIT_0B => X"0806522C0A40A50268D0068D0068D0068D0068D0068D0068D006A68034680300",
INIT_0C => X"8912E0A83289641F42A80561D040203182AC3D0AA0118A080036FFFC4F4164A0",
INIT_0D => X"050080424069F5A51250648801BFFFE0003E3E00A0685A85410C0816040B0205",
INIT_0E => X"050080080400028000000000000202900000A0F600000005008000A0F6000000",
INIT_0F => X"00023000001040214E0000000000000D0000A0F600000005008000A0F6000000",
INIT_10 => X"000000000120400800080400030000000000000205800008200D070000000000",
INIT_11 => X"000220A2C400000068008424260400001A0241DAC80001010000042016040000",
INIT_12 => X"00020048108484C10000034004414588000000D04010001020000000010009B0",
INIT_13 => X"000900000000000416C00041000140E800000000010AB0001100008A2A000000",
INIT_14 => X"A282C0000033010FB181E00020400000000419060000000000004300B0001100",
INIT_15 => X"02C0B02C0B02C0B02C0B02C4B12B312912831A27FCFE7FFB175B6FF800802594",
INIT_16 => X"2C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B",
INIT_17 => X"C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B0",
INIT_18 => X"EE7FFDF7FE783FFDFFEA0C00602FFFFFFFFFFFFFFFFFC0B02C0B02C0B02C0B02",
INIT_19 => X"BEFBEFBEFBEFBEFBEFBEFBEFBEEBAEBAEBAEBAEBBFFDF9FBEFFFFFFEBBCF9F96",
INIT_1A => X"FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFBEFBEFBEFBEF",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000FBFDFEFF7FBFDFEFF7FBFDFEFF7",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000",
INIT_22 => X"2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_26 => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFF",
INIT_2E => X"F5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA080402000000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"02000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_36 => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_37 => X"0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(3),               -- Port A write enable input
DIA(0)   => data_write_a(29),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(29),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(3),               -- Port B write enable input
DIB(0)   => data_write_b(29),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(29),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_30_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"FF9FE1F7FFBFFFFDFFD000000000000000000000000000000000000000000000",
INIT_19 => X"79E79E79E79E79E79E79E79E79E79E79E79E79E7AFBD75F5FDF7DF7FF7FFBFFE",
INIT_1A => X"3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE79E79E79E79E",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE000000000000000003F9FCFE7F3F9FCFE7F3F9FCFE7F",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000",
INIT_22 => X"2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_26 => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFF",
INIT_2E => X"F5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA080402000000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"02000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_36 => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_37 => X"0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(3),               -- Port A write enable input
DIA(0)   => data_write_a(30),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(30),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(3),               -- Port B write enable input
DIB(0)   => data_write_b(30),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(30),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_31_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"129000008004A00804A40000400800020000000C005FEA005800200400050100",
INIT_01 => X"A15FF18019700810180065FFFC0040801E80258CA2951C2200EC0906A0804140",
INIT_02 => X"146000808A0C060444692000402850040400408FF80000000010000000004000",
INIT_03 => X"000003F5D1202C70F654716A001A07F438184210960600000012108518004842",
INIT_04 => X"3E28FE3F6FE513703F70007472DA4128187B6DB530C1240A060C70580B439200",
INIT_05 => X"000F84040C088BE3E4AE40C1FD04CE38C0FC381FF8671FE01009048084C40010",
INIT_06 => X"0000000000000008000810200420620E00030BFE000181092CE7ED80DF800106",
INIT_07 => X"000000220FD1FF200040100540800000840200408002000C2244890200000200",
INIT_08 => X"0011F0780011E38004800E3CF3E0B1118C31747F000B33820209206FC9E80000",
INIT_09 => X"187FC301B124F2001600000000001A1F00110101092CE7ED81CF000401228800",
INIT_0A => X"0477330C4889CC012188310E08812982050800A91012494C31004124080886FE",
INIT_0B => X"9861D1403803800C1000C1000C1000C1000C1000C1000C1000C1800608006084",
INIT_0C => X"020400830602410901000D02D0002008012054040022102001017FE190022201",
INIT_0D => X"3A0000401E030B0C20C20188087FFA07FE203A80010002608030102008100408",
INIT_0E => X"3A000005E8010000004000F808000010100F02000008003A00000F0200000800",
INIT_0F => X"00000002006B80800000400003B80000000F02000008003A00000F0200000800",
INIT_10 => X"01E03200060000080405E8010000100000F600000081003740400000008000EE",
INIT_11 => X"201D0100000039000007404000000E1000001846282010A211AA000000000080",
INIT_12 => X"80000000E808000001C200003A0200000072000007E00080000007E0000000A0",
INIT_13 => X"0100000003E200000280800EE04000000000F8080000A02022AC04000000003D",
INIT_14 => X"9C06D082000A03200806A040019481D4000000000201E1A000040000A02022E8",
INIT_15 => X"0401004010040100401004010060C040040C200950402090128057C3FF800C60",
INIT_16 => X"4010040100401004010040100401004010040100401004010040100401004010",
INIT_17 => X"0100401004010040100401004010040100401004010040100401004010040100",
INIT_18 => X"000000000000000000001000802FFFFFFFFFFFFFFFFF81004010040100401004",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"FFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_20 => X"0000000000000000000000000FFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000000000000",
INIT_22 => X"2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_23 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_24 => X"080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFF",
INIT_25 => X"FFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_26 => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFF",
INIT_27 => X"FFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020",
INIT_28 => X"0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040200000000",
INIT_2A => X"FFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_2B => X"0402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFF",
INIT_2C => X"FFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_2D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFF",
INIT_2E => X"F5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"4BA080402000000000000000000000000000000000000000000000000FFFFFFF",
INIT_31 => X"FFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E97",
INIT_32 => X"02000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFF",
INIT_33 => X"FFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804",
INIT_34 => X"FFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFF",
INIT_35 => X"D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FF",
INIT_36 => X"FFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5",
INIT_37 => X"0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFF",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_512_2,               -- Port A enable input
WEA      => wbe_a_hi_512_2(3),               -- Port A write enable input
DIA(0)   => data_write_a(31),        -- Port A data input
DOA(0)   => data_read_a_hi_512_2(31),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_512_2,               -- Port B enable input
WEB      => wbe_b_hi_512_2(3),               -- Port B write enable input
DIB(0)   => data_write_b(31),        -- Port B data input
DOB(0)   => data_read_b_hi_512_2(31),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


end;